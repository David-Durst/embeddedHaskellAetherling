module FIFO(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0,
  input  [31:0] I_1,
  input  [31:0] I_2,
  input  [31:0] I_3,
  input  [31:0] I_4,
  input  [31:0] I_5,
  input  [31:0] I_6,
  input  [31:0] I_7,
  output [31:0] O_0,
  output [31:0] O_1,
  output [31:0] O_2,
  output [31:0] O_3,
  output [31:0] O_4,
  output [31:0] O_5,
  output [31:0] O_6,
  output [31:0] O_7
);
  reg [31:0] _T__0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_0;
  reg [31:0] _T__1; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_1;
  reg [31:0] _T__2; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_2;
  reg [31:0] _T__3; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_3;
  reg [31:0] _T__4; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_4;
  reg [31:0] _T__5; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_5;
  reg [31:0] _T__6; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_6;
  reg [31:0] _T__7; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_7;
  reg  _T_1; // @[FIFO.scala 15:27]
  reg [31:0] _RAND_8;
  assign valid_down = _T_1; // @[FIFO.scala 16:16]
  assign O_0 = _T__0; // @[FIFO.scala 14:7]
  assign O_1 = _T__1; // @[FIFO.scala 14:7]
  assign O_2 = _T__2; // @[FIFO.scala 14:7]
  assign O_3 = _T__3; // @[FIFO.scala 14:7]
  assign O_4 = _T__4; // @[FIFO.scala 14:7]
  assign O_5 = _T__5; // @[FIFO.scala 14:7]
  assign O_6 = _T__6; // @[FIFO.scala 14:7]
  assign O_7 = _T__7; // @[FIFO.scala 14:7]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T__0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T__1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T__2 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T__3 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T__4 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T__5 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T__6 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T__7 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_1 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T__0 <= I_0;
    _T__1 <= I_1;
    _T__2 <= I_2;
    _T__3 <= I_3;
    _T__4 <= I_4;
    _T__5 <= I_5;
    _T__6 <= I_6;
    _T__7 <= I_7;
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      _T_1 <= valid_up;
    end
  end
endmodule
module NestedCounters(
  input   CE,
  output  valid
);
  assign valid = CE; // @[NestedCounters.scala 65:13]
endmodule
module NestedCounters_1(
  input   CE,
  output  valid
);
  wire  NestedCounters_CE; // @[NestedCounters.scala 53:31]
  wire  NestedCounters_valid; // @[NestedCounters.scala 53:31]
  NestedCounters NestedCounters ( // @[NestedCounters.scala 53:31]
    .CE(NestedCounters_CE),
    .valid(NestedCounters_valid)
  );
  assign valid = NestedCounters_valid; // @[NestedCounters.scala 56:11]
  assign NestedCounters_CE = CE; // @[NestedCounters.scala 57:22]
endmodule
module NestedCountersWithNumValid(
  input   CE,
  output  valid
);
  wire  NestedCounters_CE; // @[NestedCounters.scala 20:44]
  wire  NestedCounters_valid; // @[NestedCounters.scala 20:44]
  NestedCounters_1 NestedCounters ( // @[NestedCounters.scala 20:44]
    .CE(NestedCounters_CE),
    .valid(NestedCounters_valid)
  );
  assign valid = NestedCounters_valid; // @[NestedCounters.scala 22:9]
  assign NestedCounters_CE = CE; // @[NestedCounters.scala 21:27]
endmodule
module RAM_ST(
  input         clock,
  input         RE,
  input  [7:0]  RADDR,
  output [31:0] RDATA_0,
  output [31:0] RDATA_1,
  output [31:0] RDATA_2,
  output [31:0] RDATA_3,
  output [31:0] RDATA_4,
  output [31:0] RDATA_5,
  output [31:0] RDATA_6,
  output [31:0] RDATA_7,
  input         WE,
  input  [7:0]  WADDR,
  input  [31:0] WDATA_0,
  input  [31:0] WDATA_1,
  input  [31:0] WDATA_2,
  input  [31:0] WDATA_3,
  input  [31:0] WDATA_4,
  input  [31:0] WDATA_5,
  input  [31:0] WDATA_6,
  input  [31:0] WDATA_7
);
  wire  write_elem_counter_CE; // @[RAM_ST.scala 20:34]
  wire  write_elem_counter_valid; // @[RAM_ST.scala 20:34]
  wire  read_elem_counter_CE; // @[RAM_ST.scala 21:33]
  wire  read_elem_counter_valid; // @[RAM_ST.scala 21:33]
  reg [255:0] ram [0:239]; // @[RAM_ST.scala 29:24]
  reg [255:0] _RAND_0;
  wire [255:0] ram__T_15_data; // @[RAM_ST.scala 29:24]
  wire [7:0] ram__T_15_addr; // @[RAM_ST.scala 29:24]
  reg [255:0] _RAND_1;
  wire [255:0] ram__T_9_data; // @[RAM_ST.scala 29:24]
  wire [7:0] ram__T_9_addr; // @[RAM_ST.scala 29:24]
  wire  ram__T_9_mask; // @[RAM_ST.scala 29:24]
  wire  ram__T_9_en; // @[RAM_ST.scala 29:24]
  reg  ram__T_15_en_pipe_0;
  reg [31:0] _RAND_2;
  reg [7:0] ram__T_15_addr_pipe_0;
  reg [31:0] _RAND_3;
  wire [7:0] _GEN_1; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_2; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_3; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_4; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_5; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_6; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_7; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_8; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_9; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_10; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_11; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_12; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_13; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_14; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_15; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_16; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_17; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_18; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_19; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_20; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_21; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_22; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_23; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_24; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_25; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_26; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_27; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_28; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_29; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_30; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_31; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_32; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_33; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_34; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_35; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_36; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_37; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_38; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_39; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_40; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_41; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_42; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_43; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_44; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_45; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_46; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_47; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_48; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_49; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_50; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_51; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_52; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_53; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_54; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_55; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_56; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_57; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_58; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_59; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_60; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_61; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_62; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_63; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_64; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_65; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_66; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_67; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_68; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_69; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_70; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_71; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_72; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_73; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_74; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_75; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_76; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_77; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_78; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_79; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_80; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_81; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_82; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_83; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_84; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_85; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_86; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_87; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_88; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_89; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_90; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_91; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_92; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_93; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_94; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_95; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_96; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_97; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_98; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_99; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_100; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_101; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_102; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_103; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_104; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_105; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_106; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_107; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_108; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_109; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_110; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_111; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_112; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_113; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_114; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_115; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_116; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_117; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_118; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_119; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_120; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_121; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_122; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_123; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_124; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_125; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_126; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_127; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_128; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_129; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_130; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_131; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_132; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_133; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_134; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_135; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_136; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_137; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_138; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_139; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_140; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_141; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_142; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_143; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_144; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_145; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_146; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_147; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_148; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_149; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_150; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_151; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_152; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_153; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_154; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_155; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_156; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_157; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_158; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_159; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_160; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_161; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_162; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_163; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_164; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_165; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_166; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_167; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_168; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_169; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_170; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_171; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_172; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_173; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_174; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_175; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_176; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_177; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_178; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_179; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_180; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_181; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_182; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_183; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_184; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_185; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_186; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_187; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_188; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_189; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_190; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_191; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_192; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_193; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_194; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_195; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_196; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_197; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_198; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_199; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_200; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_201; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_202; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_203; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_204; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_205; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_206; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_207; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_208; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_209; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_210; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_211; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_212; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_213; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_214; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_215; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_216; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_217; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_218; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_219; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_220; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_221; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_222; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_223; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_224; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_225; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_226; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_227; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_228; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_229; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_230; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_231; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_232; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_233; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_234; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_235; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_236; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_237; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_238; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_239; // @[RAM_ST.scala 31:71]
  wire [8:0] _T; // @[RAM_ST.scala 31:71]
  wire [127:0] _T_4; // @[RAM_ST.scala 31:115]
  wire [127:0] _T_7; // @[RAM_ST.scala 31:115]
  wire [7:0] _GEN_246; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_247; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_248; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_249; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_250; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_251; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_252; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_253; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_254; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_255; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_256; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_257; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_258; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_259; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_260; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_261; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_262; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_263; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_264; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_265; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_266; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_267; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_268; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_269; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_270; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_271; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_272; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_273; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_274; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_275; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_276; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_277; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_278; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_279; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_280; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_281; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_282; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_283; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_284; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_285; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_286; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_287; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_288; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_289; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_290; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_291; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_292; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_293; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_294; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_295; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_296; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_297; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_298; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_299; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_300; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_301; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_302; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_303; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_304; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_305; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_306; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_307; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_308; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_309; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_310; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_311; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_312; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_313; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_314; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_315; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_316; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_317; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_318; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_319; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_320; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_321; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_322; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_323; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_324; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_325; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_326; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_327; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_328; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_329; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_330; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_331; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_332; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_333; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_334; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_335; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_336; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_337; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_338; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_339; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_340; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_341; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_342; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_343; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_344; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_345; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_346; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_347; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_348; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_349; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_350; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_351; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_352; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_353; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_354; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_355; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_356; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_357; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_358; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_359; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_360; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_361; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_362; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_363; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_364; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_365; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_366; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_367; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_368; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_369; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_370; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_371; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_372; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_373; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_374; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_375; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_376; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_377; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_378; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_379; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_380; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_381; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_382; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_383; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_384; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_385; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_386; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_387; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_388; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_389; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_390; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_391; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_392; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_393; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_394; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_395; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_396; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_397; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_398; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_399; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_400; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_401; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_402; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_403; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_404; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_405; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_406; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_407; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_408; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_409; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_410; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_411; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_412; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_413; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_414; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_415; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_416; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_417; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_418; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_419; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_420; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_421; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_422; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_423; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_424; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_425; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_426; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_427; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_428; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_429; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_430; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_431; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_432; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_433; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_434; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_435; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_436; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_437; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_438; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_439; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_440; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_441; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_442; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_443; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_444; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_445; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_446; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_447; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_448; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_449; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_450; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_451; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_452; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_453; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_454; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_455; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_456; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_457; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_458; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_459; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_460; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_461; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_462; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_463; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_464; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_465; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_466; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_467; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_468; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_469; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_470; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_471; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_472; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_473; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_474; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_475; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_476; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_477; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_478; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_479; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_480; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_481; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_482; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_483; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_484; // @[RAM_ST.scala 32:46]
  wire [8:0] _T_10; // @[RAM_ST.scala 32:46]
  wire [255:0] _T_17;
  NestedCountersWithNumValid write_elem_counter ( // @[RAM_ST.scala 20:34]
    .CE(write_elem_counter_CE),
    .valid(write_elem_counter_valid)
  );
  NestedCountersWithNumValid read_elem_counter ( // @[RAM_ST.scala 21:33]
    .CE(read_elem_counter_CE),
    .valid(read_elem_counter_valid)
  );
  assign ram__T_15_addr = ram__T_15_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram__T_15_data = ram[ram__T_15_addr]; // @[RAM_ST.scala 29:24]
  `else
  assign ram__T_15_data = ram__T_15_addr >= 8'hf0 ? _RAND_1[255:0] : ram[ram__T_15_addr]; // @[RAM_ST.scala 29:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram__T_9_data = {_T_7,_T_4};
  assign ram__T_9_addr = _T[7:0];
  assign ram__T_9_mask = 1'h1;
  assign ram__T_9_en = write_elem_counter_valid;
  assign _GEN_1 = 8'h1 == WADDR ? 8'h1 : 8'h0; // @[RAM_ST.scala 31:71]
  assign _GEN_2 = 8'h2 == WADDR ? 8'h2 : _GEN_1; // @[RAM_ST.scala 31:71]
  assign _GEN_3 = 8'h3 == WADDR ? 8'h3 : _GEN_2; // @[RAM_ST.scala 31:71]
  assign _GEN_4 = 8'h4 == WADDR ? 8'h4 : _GEN_3; // @[RAM_ST.scala 31:71]
  assign _GEN_5 = 8'h5 == WADDR ? 8'h5 : _GEN_4; // @[RAM_ST.scala 31:71]
  assign _GEN_6 = 8'h6 == WADDR ? 8'h6 : _GEN_5; // @[RAM_ST.scala 31:71]
  assign _GEN_7 = 8'h7 == WADDR ? 8'h7 : _GEN_6; // @[RAM_ST.scala 31:71]
  assign _GEN_8 = 8'h8 == WADDR ? 8'h8 : _GEN_7; // @[RAM_ST.scala 31:71]
  assign _GEN_9 = 8'h9 == WADDR ? 8'h9 : _GEN_8; // @[RAM_ST.scala 31:71]
  assign _GEN_10 = 8'ha == WADDR ? 8'ha : _GEN_9; // @[RAM_ST.scala 31:71]
  assign _GEN_11 = 8'hb == WADDR ? 8'hb : _GEN_10; // @[RAM_ST.scala 31:71]
  assign _GEN_12 = 8'hc == WADDR ? 8'hc : _GEN_11; // @[RAM_ST.scala 31:71]
  assign _GEN_13 = 8'hd == WADDR ? 8'hd : _GEN_12; // @[RAM_ST.scala 31:71]
  assign _GEN_14 = 8'he == WADDR ? 8'he : _GEN_13; // @[RAM_ST.scala 31:71]
  assign _GEN_15 = 8'hf == WADDR ? 8'hf : _GEN_14; // @[RAM_ST.scala 31:71]
  assign _GEN_16 = 8'h10 == WADDR ? 8'h10 : _GEN_15; // @[RAM_ST.scala 31:71]
  assign _GEN_17 = 8'h11 == WADDR ? 8'h11 : _GEN_16; // @[RAM_ST.scala 31:71]
  assign _GEN_18 = 8'h12 == WADDR ? 8'h12 : _GEN_17; // @[RAM_ST.scala 31:71]
  assign _GEN_19 = 8'h13 == WADDR ? 8'h13 : _GEN_18; // @[RAM_ST.scala 31:71]
  assign _GEN_20 = 8'h14 == WADDR ? 8'h14 : _GEN_19; // @[RAM_ST.scala 31:71]
  assign _GEN_21 = 8'h15 == WADDR ? 8'h15 : _GEN_20; // @[RAM_ST.scala 31:71]
  assign _GEN_22 = 8'h16 == WADDR ? 8'h16 : _GEN_21; // @[RAM_ST.scala 31:71]
  assign _GEN_23 = 8'h17 == WADDR ? 8'h17 : _GEN_22; // @[RAM_ST.scala 31:71]
  assign _GEN_24 = 8'h18 == WADDR ? 8'h18 : _GEN_23; // @[RAM_ST.scala 31:71]
  assign _GEN_25 = 8'h19 == WADDR ? 8'h19 : _GEN_24; // @[RAM_ST.scala 31:71]
  assign _GEN_26 = 8'h1a == WADDR ? 8'h1a : _GEN_25; // @[RAM_ST.scala 31:71]
  assign _GEN_27 = 8'h1b == WADDR ? 8'h1b : _GEN_26; // @[RAM_ST.scala 31:71]
  assign _GEN_28 = 8'h1c == WADDR ? 8'h1c : _GEN_27; // @[RAM_ST.scala 31:71]
  assign _GEN_29 = 8'h1d == WADDR ? 8'h1d : _GEN_28; // @[RAM_ST.scala 31:71]
  assign _GEN_30 = 8'h1e == WADDR ? 8'h1e : _GEN_29; // @[RAM_ST.scala 31:71]
  assign _GEN_31 = 8'h1f == WADDR ? 8'h1f : _GEN_30; // @[RAM_ST.scala 31:71]
  assign _GEN_32 = 8'h20 == WADDR ? 8'h20 : _GEN_31; // @[RAM_ST.scala 31:71]
  assign _GEN_33 = 8'h21 == WADDR ? 8'h21 : _GEN_32; // @[RAM_ST.scala 31:71]
  assign _GEN_34 = 8'h22 == WADDR ? 8'h22 : _GEN_33; // @[RAM_ST.scala 31:71]
  assign _GEN_35 = 8'h23 == WADDR ? 8'h23 : _GEN_34; // @[RAM_ST.scala 31:71]
  assign _GEN_36 = 8'h24 == WADDR ? 8'h24 : _GEN_35; // @[RAM_ST.scala 31:71]
  assign _GEN_37 = 8'h25 == WADDR ? 8'h25 : _GEN_36; // @[RAM_ST.scala 31:71]
  assign _GEN_38 = 8'h26 == WADDR ? 8'h26 : _GEN_37; // @[RAM_ST.scala 31:71]
  assign _GEN_39 = 8'h27 == WADDR ? 8'h27 : _GEN_38; // @[RAM_ST.scala 31:71]
  assign _GEN_40 = 8'h28 == WADDR ? 8'h28 : _GEN_39; // @[RAM_ST.scala 31:71]
  assign _GEN_41 = 8'h29 == WADDR ? 8'h29 : _GEN_40; // @[RAM_ST.scala 31:71]
  assign _GEN_42 = 8'h2a == WADDR ? 8'h2a : _GEN_41; // @[RAM_ST.scala 31:71]
  assign _GEN_43 = 8'h2b == WADDR ? 8'h2b : _GEN_42; // @[RAM_ST.scala 31:71]
  assign _GEN_44 = 8'h2c == WADDR ? 8'h2c : _GEN_43; // @[RAM_ST.scala 31:71]
  assign _GEN_45 = 8'h2d == WADDR ? 8'h2d : _GEN_44; // @[RAM_ST.scala 31:71]
  assign _GEN_46 = 8'h2e == WADDR ? 8'h2e : _GEN_45; // @[RAM_ST.scala 31:71]
  assign _GEN_47 = 8'h2f == WADDR ? 8'h2f : _GEN_46; // @[RAM_ST.scala 31:71]
  assign _GEN_48 = 8'h30 == WADDR ? 8'h30 : _GEN_47; // @[RAM_ST.scala 31:71]
  assign _GEN_49 = 8'h31 == WADDR ? 8'h31 : _GEN_48; // @[RAM_ST.scala 31:71]
  assign _GEN_50 = 8'h32 == WADDR ? 8'h32 : _GEN_49; // @[RAM_ST.scala 31:71]
  assign _GEN_51 = 8'h33 == WADDR ? 8'h33 : _GEN_50; // @[RAM_ST.scala 31:71]
  assign _GEN_52 = 8'h34 == WADDR ? 8'h34 : _GEN_51; // @[RAM_ST.scala 31:71]
  assign _GEN_53 = 8'h35 == WADDR ? 8'h35 : _GEN_52; // @[RAM_ST.scala 31:71]
  assign _GEN_54 = 8'h36 == WADDR ? 8'h36 : _GEN_53; // @[RAM_ST.scala 31:71]
  assign _GEN_55 = 8'h37 == WADDR ? 8'h37 : _GEN_54; // @[RAM_ST.scala 31:71]
  assign _GEN_56 = 8'h38 == WADDR ? 8'h38 : _GEN_55; // @[RAM_ST.scala 31:71]
  assign _GEN_57 = 8'h39 == WADDR ? 8'h39 : _GEN_56; // @[RAM_ST.scala 31:71]
  assign _GEN_58 = 8'h3a == WADDR ? 8'h3a : _GEN_57; // @[RAM_ST.scala 31:71]
  assign _GEN_59 = 8'h3b == WADDR ? 8'h3b : _GEN_58; // @[RAM_ST.scala 31:71]
  assign _GEN_60 = 8'h3c == WADDR ? 8'h3c : _GEN_59; // @[RAM_ST.scala 31:71]
  assign _GEN_61 = 8'h3d == WADDR ? 8'h3d : _GEN_60; // @[RAM_ST.scala 31:71]
  assign _GEN_62 = 8'h3e == WADDR ? 8'h3e : _GEN_61; // @[RAM_ST.scala 31:71]
  assign _GEN_63 = 8'h3f == WADDR ? 8'h3f : _GEN_62; // @[RAM_ST.scala 31:71]
  assign _GEN_64 = 8'h40 == WADDR ? 8'h40 : _GEN_63; // @[RAM_ST.scala 31:71]
  assign _GEN_65 = 8'h41 == WADDR ? 8'h41 : _GEN_64; // @[RAM_ST.scala 31:71]
  assign _GEN_66 = 8'h42 == WADDR ? 8'h42 : _GEN_65; // @[RAM_ST.scala 31:71]
  assign _GEN_67 = 8'h43 == WADDR ? 8'h43 : _GEN_66; // @[RAM_ST.scala 31:71]
  assign _GEN_68 = 8'h44 == WADDR ? 8'h44 : _GEN_67; // @[RAM_ST.scala 31:71]
  assign _GEN_69 = 8'h45 == WADDR ? 8'h45 : _GEN_68; // @[RAM_ST.scala 31:71]
  assign _GEN_70 = 8'h46 == WADDR ? 8'h46 : _GEN_69; // @[RAM_ST.scala 31:71]
  assign _GEN_71 = 8'h47 == WADDR ? 8'h47 : _GEN_70; // @[RAM_ST.scala 31:71]
  assign _GEN_72 = 8'h48 == WADDR ? 8'h48 : _GEN_71; // @[RAM_ST.scala 31:71]
  assign _GEN_73 = 8'h49 == WADDR ? 8'h49 : _GEN_72; // @[RAM_ST.scala 31:71]
  assign _GEN_74 = 8'h4a == WADDR ? 8'h4a : _GEN_73; // @[RAM_ST.scala 31:71]
  assign _GEN_75 = 8'h4b == WADDR ? 8'h4b : _GEN_74; // @[RAM_ST.scala 31:71]
  assign _GEN_76 = 8'h4c == WADDR ? 8'h4c : _GEN_75; // @[RAM_ST.scala 31:71]
  assign _GEN_77 = 8'h4d == WADDR ? 8'h4d : _GEN_76; // @[RAM_ST.scala 31:71]
  assign _GEN_78 = 8'h4e == WADDR ? 8'h4e : _GEN_77; // @[RAM_ST.scala 31:71]
  assign _GEN_79 = 8'h4f == WADDR ? 8'h4f : _GEN_78; // @[RAM_ST.scala 31:71]
  assign _GEN_80 = 8'h50 == WADDR ? 8'h50 : _GEN_79; // @[RAM_ST.scala 31:71]
  assign _GEN_81 = 8'h51 == WADDR ? 8'h51 : _GEN_80; // @[RAM_ST.scala 31:71]
  assign _GEN_82 = 8'h52 == WADDR ? 8'h52 : _GEN_81; // @[RAM_ST.scala 31:71]
  assign _GEN_83 = 8'h53 == WADDR ? 8'h53 : _GEN_82; // @[RAM_ST.scala 31:71]
  assign _GEN_84 = 8'h54 == WADDR ? 8'h54 : _GEN_83; // @[RAM_ST.scala 31:71]
  assign _GEN_85 = 8'h55 == WADDR ? 8'h55 : _GEN_84; // @[RAM_ST.scala 31:71]
  assign _GEN_86 = 8'h56 == WADDR ? 8'h56 : _GEN_85; // @[RAM_ST.scala 31:71]
  assign _GEN_87 = 8'h57 == WADDR ? 8'h57 : _GEN_86; // @[RAM_ST.scala 31:71]
  assign _GEN_88 = 8'h58 == WADDR ? 8'h58 : _GEN_87; // @[RAM_ST.scala 31:71]
  assign _GEN_89 = 8'h59 == WADDR ? 8'h59 : _GEN_88; // @[RAM_ST.scala 31:71]
  assign _GEN_90 = 8'h5a == WADDR ? 8'h5a : _GEN_89; // @[RAM_ST.scala 31:71]
  assign _GEN_91 = 8'h5b == WADDR ? 8'h5b : _GEN_90; // @[RAM_ST.scala 31:71]
  assign _GEN_92 = 8'h5c == WADDR ? 8'h5c : _GEN_91; // @[RAM_ST.scala 31:71]
  assign _GEN_93 = 8'h5d == WADDR ? 8'h5d : _GEN_92; // @[RAM_ST.scala 31:71]
  assign _GEN_94 = 8'h5e == WADDR ? 8'h5e : _GEN_93; // @[RAM_ST.scala 31:71]
  assign _GEN_95 = 8'h5f == WADDR ? 8'h5f : _GEN_94; // @[RAM_ST.scala 31:71]
  assign _GEN_96 = 8'h60 == WADDR ? 8'h60 : _GEN_95; // @[RAM_ST.scala 31:71]
  assign _GEN_97 = 8'h61 == WADDR ? 8'h61 : _GEN_96; // @[RAM_ST.scala 31:71]
  assign _GEN_98 = 8'h62 == WADDR ? 8'h62 : _GEN_97; // @[RAM_ST.scala 31:71]
  assign _GEN_99 = 8'h63 == WADDR ? 8'h63 : _GEN_98; // @[RAM_ST.scala 31:71]
  assign _GEN_100 = 8'h64 == WADDR ? 8'h64 : _GEN_99; // @[RAM_ST.scala 31:71]
  assign _GEN_101 = 8'h65 == WADDR ? 8'h65 : _GEN_100; // @[RAM_ST.scala 31:71]
  assign _GEN_102 = 8'h66 == WADDR ? 8'h66 : _GEN_101; // @[RAM_ST.scala 31:71]
  assign _GEN_103 = 8'h67 == WADDR ? 8'h67 : _GEN_102; // @[RAM_ST.scala 31:71]
  assign _GEN_104 = 8'h68 == WADDR ? 8'h68 : _GEN_103; // @[RAM_ST.scala 31:71]
  assign _GEN_105 = 8'h69 == WADDR ? 8'h69 : _GEN_104; // @[RAM_ST.scala 31:71]
  assign _GEN_106 = 8'h6a == WADDR ? 8'h6a : _GEN_105; // @[RAM_ST.scala 31:71]
  assign _GEN_107 = 8'h6b == WADDR ? 8'h6b : _GEN_106; // @[RAM_ST.scala 31:71]
  assign _GEN_108 = 8'h6c == WADDR ? 8'h6c : _GEN_107; // @[RAM_ST.scala 31:71]
  assign _GEN_109 = 8'h6d == WADDR ? 8'h6d : _GEN_108; // @[RAM_ST.scala 31:71]
  assign _GEN_110 = 8'h6e == WADDR ? 8'h6e : _GEN_109; // @[RAM_ST.scala 31:71]
  assign _GEN_111 = 8'h6f == WADDR ? 8'h6f : _GEN_110; // @[RAM_ST.scala 31:71]
  assign _GEN_112 = 8'h70 == WADDR ? 8'h70 : _GEN_111; // @[RAM_ST.scala 31:71]
  assign _GEN_113 = 8'h71 == WADDR ? 8'h71 : _GEN_112; // @[RAM_ST.scala 31:71]
  assign _GEN_114 = 8'h72 == WADDR ? 8'h72 : _GEN_113; // @[RAM_ST.scala 31:71]
  assign _GEN_115 = 8'h73 == WADDR ? 8'h73 : _GEN_114; // @[RAM_ST.scala 31:71]
  assign _GEN_116 = 8'h74 == WADDR ? 8'h74 : _GEN_115; // @[RAM_ST.scala 31:71]
  assign _GEN_117 = 8'h75 == WADDR ? 8'h75 : _GEN_116; // @[RAM_ST.scala 31:71]
  assign _GEN_118 = 8'h76 == WADDR ? 8'h76 : _GEN_117; // @[RAM_ST.scala 31:71]
  assign _GEN_119 = 8'h77 == WADDR ? 8'h77 : _GEN_118; // @[RAM_ST.scala 31:71]
  assign _GEN_120 = 8'h78 == WADDR ? 8'h78 : _GEN_119; // @[RAM_ST.scala 31:71]
  assign _GEN_121 = 8'h79 == WADDR ? 8'h79 : _GEN_120; // @[RAM_ST.scala 31:71]
  assign _GEN_122 = 8'h7a == WADDR ? 8'h7a : _GEN_121; // @[RAM_ST.scala 31:71]
  assign _GEN_123 = 8'h7b == WADDR ? 8'h7b : _GEN_122; // @[RAM_ST.scala 31:71]
  assign _GEN_124 = 8'h7c == WADDR ? 8'h7c : _GEN_123; // @[RAM_ST.scala 31:71]
  assign _GEN_125 = 8'h7d == WADDR ? 8'h7d : _GEN_124; // @[RAM_ST.scala 31:71]
  assign _GEN_126 = 8'h7e == WADDR ? 8'h7e : _GEN_125; // @[RAM_ST.scala 31:71]
  assign _GEN_127 = 8'h7f == WADDR ? 8'h7f : _GEN_126; // @[RAM_ST.scala 31:71]
  assign _GEN_128 = 8'h80 == WADDR ? 8'h80 : _GEN_127; // @[RAM_ST.scala 31:71]
  assign _GEN_129 = 8'h81 == WADDR ? 8'h81 : _GEN_128; // @[RAM_ST.scala 31:71]
  assign _GEN_130 = 8'h82 == WADDR ? 8'h82 : _GEN_129; // @[RAM_ST.scala 31:71]
  assign _GEN_131 = 8'h83 == WADDR ? 8'h83 : _GEN_130; // @[RAM_ST.scala 31:71]
  assign _GEN_132 = 8'h84 == WADDR ? 8'h84 : _GEN_131; // @[RAM_ST.scala 31:71]
  assign _GEN_133 = 8'h85 == WADDR ? 8'h85 : _GEN_132; // @[RAM_ST.scala 31:71]
  assign _GEN_134 = 8'h86 == WADDR ? 8'h86 : _GEN_133; // @[RAM_ST.scala 31:71]
  assign _GEN_135 = 8'h87 == WADDR ? 8'h87 : _GEN_134; // @[RAM_ST.scala 31:71]
  assign _GEN_136 = 8'h88 == WADDR ? 8'h88 : _GEN_135; // @[RAM_ST.scala 31:71]
  assign _GEN_137 = 8'h89 == WADDR ? 8'h89 : _GEN_136; // @[RAM_ST.scala 31:71]
  assign _GEN_138 = 8'h8a == WADDR ? 8'h8a : _GEN_137; // @[RAM_ST.scala 31:71]
  assign _GEN_139 = 8'h8b == WADDR ? 8'h8b : _GEN_138; // @[RAM_ST.scala 31:71]
  assign _GEN_140 = 8'h8c == WADDR ? 8'h8c : _GEN_139; // @[RAM_ST.scala 31:71]
  assign _GEN_141 = 8'h8d == WADDR ? 8'h8d : _GEN_140; // @[RAM_ST.scala 31:71]
  assign _GEN_142 = 8'h8e == WADDR ? 8'h8e : _GEN_141; // @[RAM_ST.scala 31:71]
  assign _GEN_143 = 8'h8f == WADDR ? 8'h8f : _GEN_142; // @[RAM_ST.scala 31:71]
  assign _GEN_144 = 8'h90 == WADDR ? 8'h90 : _GEN_143; // @[RAM_ST.scala 31:71]
  assign _GEN_145 = 8'h91 == WADDR ? 8'h91 : _GEN_144; // @[RAM_ST.scala 31:71]
  assign _GEN_146 = 8'h92 == WADDR ? 8'h92 : _GEN_145; // @[RAM_ST.scala 31:71]
  assign _GEN_147 = 8'h93 == WADDR ? 8'h93 : _GEN_146; // @[RAM_ST.scala 31:71]
  assign _GEN_148 = 8'h94 == WADDR ? 8'h94 : _GEN_147; // @[RAM_ST.scala 31:71]
  assign _GEN_149 = 8'h95 == WADDR ? 8'h95 : _GEN_148; // @[RAM_ST.scala 31:71]
  assign _GEN_150 = 8'h96 == WADDR ? 8'h96 : _GEN_149; // @[RAM_ST.scala 31:71]
  assign _GEN_151 = 8'h97 == WADDR ? 8'h97 : _GEN_150; // @[RAM_ST.scala 31:71]
  assign _GEN_152 = 8'h98 == WADDR ? 8'h98 : _GEN_151; // @[RAM_ST.scala 31:71]
  assign _GEN_153 = 8'h99 == WADDR ? 8'h99 : _GEN_152; // @[RAM_ST.scala 31:71]
  assign _GEN_154 = 8'h9a == WADDR ? 8'h9a : _GEN_153; // @[RAM_ST.scala 31:71]
  assign _GEN_155 = 8'h9b == WADDR ? 8'h9b : _GEN_154; // @[RAM_ST.scala 31:71]
  assign _GEN_156 = 8'h9c == WADDR ? 8'h9c : _GEN_155; // @[RAM_ST.scala 31:71]
  assign _GEN_157 = 8'h9d == WADDR ? 8'h9d : _GEN_156; // @[RAM_ST.scala 31:71]
  assign _GEN_158 = 8'h9e == WADDR ? 8'h9e : _GEN_157; // @[RAM_ST.scala 31:71]
  assign _GEN_159 = 8'h9f == WADDR ? 8'h9f : _GEN_158; // @[RAM_ST.scala 31:71]
  assign _GEN_160 = 8'ha0 == WADDR ? 8'ha0 : _GEN_159; // @[RAM_ST.scala 31:71]
  assign _GEN_161 = 8'ha1 == WADDR ? 8'ha1 : _GEN_160; // @[RAM_ST.scala 31:71]
  assign _GEN_162 = 8'ha2 == WADDR ? 8'ha2 : _GEN_161; // @[RAM_ST.scala 31:71]
  assign _GEN_163 = 8'ha3 == WADDR ? 8'ha3 : _GEN_162; // @[RAM_ST.scala 31:71]
  assign _GEN_164 = 8'ha4 == WADDR ? 8'ha4 : _GEN_163; // @[RAM_ST.scala 31:71]
  assign _GEN_165 = 8'ha5 == WADDR ? 8'ha5 : _GEN_164; // @[RAM_ST.scala 31:71]
  assign _GEN_166 = 8'ha6 == WADDR ? 8'ha6 : _GEN_165; // @[RAM_ST.scala 31:71]
  assign _GEN_167 = 8'ha7 == WADDR ? 8'ha7 : _GEN_166; // @[RAM_ST.scala 31:71]
  assign _GEN_168 = 8'ha8 == WADDR ? 8'ha8 : _GEN_167; // @[RAM_ST.scala 31:71]
  assign _GEN_169 = 8'ha9 == WADDR ? 8'ha9 : _GEN_168; // @[RAM_ST.scala 31:71]
  assign _GEN_170 = 8'haa == WADDR ? 8'haa : _GEN_169; // @[RAM_ST.scala 31:71]
  assign _GEN_171 = 8'hab == WADDR ? 8'hab : _GEN_170; // @[RAM_ST.scala 31:71]
  assign _GEN_172 = 8'hac == WADDR ? 8'hac : _GEN_171; // @[RAM_ST.scala 31:71]
  assign _GEN_173 = 8'had == WADDR ? 8'had : _GEN_172; // @[RAM_ST.scala 31:71]
  assign _GEN_174 = 8'hae == WADDR ? 8'hae : _GEN_173; // @[RAM_ST.scala 31:71]
  assign _GEN_175 = 8'haf == WADDR ? 8'haf : _GEN_174; // @[RAM_ST.scala 31:71]
  assign _GEN_176 = 8'hb0 == WADDR ? 8'hb0 : _GEN_175; // @[RAM_ST.scala 31:71]
  assign _GEN_177 = 8'hb1 == WADDR ? 8'hb1 : _GEN_176; // @[RAM_ST.scala 31:71]
  assign _GEN_178 = 8'hb2 == WADDR ? 8'hb2 : _GEN_177; // @[RAM_ST.scala 31:71]
  assign _GEN_179 = 8'hb3 == WADDR ? 8'hb3 : _GEN_178; // @[RAM_ST.scala 31:71]
  assign _GEN_180 = 8'hb4 == WADDR ? 8'hb4 : _GEN_179; // @[RAM_ST.scala 31:71]
  assign _GEN_181 = 8'hb5 == WADDR ? 8'hb5 : _GEN_180; // @[RAM_ST.scala 31:71]
  assign _GEN_182 = 8'hb6 == WADDR ? 8'hb6 : _GEN_181; // @[RAM_ST.scala 31:71]
  assign _GEN_183 = 8'hb7 == WADDR ? 8'hb7 : _GEN_182; // @[RAM_ST.scala 31:71]
  assign _GEN_184 = 8'hb8 == WADDR ? 8'hb8 : _GEN_183; // @[RAM_ST.scala 31:71]
  assign _GEN_185 = 8'hb9 == WADDR ? 8'hb9 : _GEN_184; // @[RAM_ST.scala 31:71]
  assign _GEN_186 = 8'hba == WADDR ? 8'hba : _GEN_185; // @[RAM_ST.scala 31:71]
  assign _GEN_187 = 8'hbb == WADDR ? 8'hbb : _GEN_186; // @[RAM_ST.scala 31:71]
  assign _GEN_188 = 8'hbc == WADDR ? 8'hbc : _GEN_187; // @[RAM_ST.scala 31:71]
  assign _GEN_189 = 8'hbd == WADDR ? 8'hbd : _GEN_188; // @[RAM_ST.scala 31:71]
  assign _GEN_190 = 8'hbe == WADDR ? 8'hbe : _GEN_189; // @[RAM_ST.scala 31:71]
  assign _GEN_191 = 8'hbf == WADDR ? 8'hbf : _GEN_190; // @[RAM_ST.scala 31:71]
  assign _GEN_192 = 8'hc0 == WADDR ? 8'hc0 : _GEN_191; // @[RAM_ST.scala 31:71]
  assign _GEN_193 = 8'hc1 == WADDR ? 8'hc1 : _GEN_192; // @[RAM_ST.scala 31:71]
  assign _GEN_194 = 8'hc2 == WADDR ? 8'hc2 : _GEN_193; // @[RAM_ST.scala 31:71]
  assign _GEN_195 = 8'hc3 == WADDR ? 8'hc3 : _GEN_194; // @[RAM_ST.scala 31:71]
  assign _GEN_196 = 8'hc4 == WADDR ? 8'hc4 : _GEN_195; // @[RAM_ST.scala 31:71]
  assign _GEN_197 = 8'hc5 == WADDR ? 8'hc5 : _GEN_196; // @[RAM_ST.scala 31:71]
  assign _GEN_198 = 8'hc6 == WADDR ? 8'hc6 : _GEN_197; // @[RAM_ST.scala 31:71]
  assign _GEN_199 = 8'hc7 == WADDR ? 8'hc7 : _GEN_198; // @[RAM_ST.scala 31:71]
  assign _GEN_200 = 8'hc8 == WADDR ? 8'hc8 : _GEN_199; // @[RAM_ST.scala 31:71]
  assign _GEN_201 = 8'hc9 == WADDR ? 8'hc9 : _GEN_200; // @[RAM_ST.scala 31:71]
  assign _GEN_202 = 8'hca == WADDR ? 8'hca : _GEN_201; // @[RAM_ST.scala 31:71]
  assign _GEN_203 = 8'hcb == WADDR ? 8'hcb : _GEN_202; // @[RAM_ST.scala 31:71]
  assign _GEN_204 = 8'hcc == WADDR ? 8'hcc : _GEN_203; // @[RAM_ST.scala 31:71]
  assign _GEN_205 = 8'hcd == WADDR ? 8'hcd : _GEN_204; // @[RAM_ST.scala 31:71]
  assign _GEN_206 = 8'hce == WADDR ? 8'hce : _GEN_205; // @[RAM_ST.scala 31:71]
  assign _GEN_207 = 8'hcf == WADDR ? 8'hcf : _GEN_206; // @[RAM_ST.scala 31:71]
  assign _GEN_208 = 8'hd0 == WADDR ? 8'hd0 : _GEN_207; // @[RAM_ST.scala 31:71]
  assign _GEN_209 = 8'hd1 == WADDR ? 8'hd1 : _GEN_208; // @[RAM_ST.scala 31:71]
  assign _GEN_210 = 8'hd2 == WADDR ? 8'hd2 : _GEN_209; // @[RAM_ST.scala 31:71]
  assign _GEN_211 = 8'hd3 == WADDR ? 8'hd3 : _GEN_210; // @[RAM_ST.scala 31:71]
  assign _GEN_212 = 8'hd4 == WADDR ? 8'hd4 : _GEN_211; // @[RAM_ST.scala 31:71]
  assign _GEN_213 = 8'hd5 == WADDR ? 8'hd5 : _GEN_212; // @[RAM_ST.scala 31:71]
  assign _GEN_214 = 8'hd6 == WADDR ? 8'hd6 : _GEN_213; // @[RAM_ST.scala 31:71]
  assign _GEN_215 = 8'hd7 == WADDR ? 8'hd7 : _GEN_214; // @[RAM_ST.scala 31:71]
  assign _GEN_216 = 8'hd8 == WADDR ? 8'hd8 : _GEN_215; // @[RAM_ST.scala 31:71]
  assign _GEN_217 = 8'hd9 == WADDR ? 8'hd9 : _GEN_216; // @[RAM_ST.scala 31:71]
  assign _GEN_218 = 8'hda == WADDR ? 8'hda : _GEN_217; // @[RAM_ST.scala 31:71]
  assign _GEN_219 = 8'hdb == WADDR ? 8'hdb : _GEN_218; // @[RAM_ST.scala 31:71]
  assign _GEN_220 = 8'hdc == WADDR ? 8'hdc : _GEN_219; // @[RAM_ST.scala 31:71]
  assign _GEN_221 = 8'hdd == WADDR ? 8'hdd : _GEN_220; // @[RAM_ST.scala 31:71]
  assign _GEN_222 = 8'hde == WADDR ? 8'hde : _GEN_221; // @[RAM_ST.scala 31:71]
  assign _GEN_223 = 8'hdf == WADDR ? 8'hdf : _GEN_222; // @[RAM_ST.scala 31:71]
  assign _GEN_224 = 8'he0 == WADDR ? 8'he0 : _GEN_223; // @[RAM_ST.scala 31:71]
  assign _GEN_225 = 8'he1 == WADDR ? 8'he1 : _GEN_224; // @[RAM_ST.scala 31:71]
  assign _GEN_226 = 8'he2 == WADDR ? 8'he2 : _GEN_225; // @[RAM_ST.scala 31:71]
  assign _GEN_227 = 8'he3 == WADDR ? 8'he3 : _GEN_226; // @[RAM_ST.scala 31:71]
  assign _GEN_228 = 8'he4 == WADDR ? 8'he4 : _GEN_227; // @[RAM_ST.scala 31:71]
  assign _GEN_229 = 8'he5 == WADDR ? 8'he5 : _GEN_228; // @[RAM_ST.scala 31:71]
  assign _GEN_230 = 8'he6 == WADDR ? 8'he6 : _GEN_229; // @[RAM_ST.scala 31:71]
  assign _GEN_231 = 8'he7 == WADDR ? 8'he7 : _GEN_230; // @[RAM_ST.scala 31:71]
  assign _GEN_232 = 8'he8 == WADDR ? 8'he8 : _GEN_231; // @[RAM_ST.scala 31:71]
  assign _GEN_233 = 8'he9 == WADDR ? 8'he9 : _GEN_232; // @[RAM_ST.scala 31:71]
  assign _GEN_234 = 8'hea == WADDR ? 8'hea : _GEN_233; // @[RAM_ST.scala 31:71]
  assign _GEN_235 = 8'heb == WADDR ? 8'heb : _GEN_234; // @[RAM_ST.scala 31:71]
  assign _GEN_236 = 8'hec == WADDR ? 8'hec : _GEN_235; // @[RAM_ST.scala 31:71]
  assign _GEN_237 = 8'hed == WADDR ? 8'hed : _GEN_236; // @[RAM_ST.scala 31:71]
  assign _GEN_238 = 8'hee == WADDR ? 8'hee : _GEN_237; // @[RAM_ST.scala 31:71]
  assign _GEN_239 = 8'hef == WADDR ? 8'hef : _GEN_238; // @[RAM_ST.scala 31:71]
  assign _T = {{1'd0}, _GEN_239}; // @[RAM_ST.scala 31:71]
  assign _T_4 = {WDATA_3,WDATA_2,WDATA_1,WDATA_0}; // @[RAM_ST.scala 31:115]
  assign _T_7 = {WDATA_7,WDATA_6,WDATA_5,WDATA_4}; // @[RAM_ST.scala 31:115]
  assign _GEN_246 = 8'h1 == RADDR ? 8'h1 : 8'h0; // @[RAM_ST.scala 32:46]
  assign _GEN_247 = 8'h2 == RADDR ? 8'h2 : _GEN_246; // @[RAM_ST.scala 32:46]
  assign _GEN_248 = 8'h3 == RADDR ? 8'h3 : _GEN_247; // @[RAM_ST.scala 32:46]
  assign _GEN_249 = 8'h4 == RADDR ? 8'h4 : _GEN_248; // @[RAM_ST.scala 32:46]
  assign _GEN_250 = 8'h5 == RADDR ? 8'h5 : _GEN_249; // @[RAM_ST.scala 32:46]
  assign _GEN_251 = 8'h6 == RADDR ? 8'h6 : _GEN_250; // @[RAM_ST.scala 32:46]
  assign _GEN_252 = 8'h7 == RADDR ? 8'h7 : _GEN_251; // @[RAM_ST.scala 32:46]
  assign _GEN_253 = 8'h8 == RADDR ? 8'h8 : _GEN_252; // @[RAM_ST.scala 32:46]
  assign _GEN_254 = 8'h9 == RADDR ? 8'h9 : _GEN_253; // @[RAM_ST.scala 32:46]
  assign _GEN_255 = 8'ha == RADDR ? 8'ha : _GEN_254; // @[RAM_ST.scala 32:46]
  assign _GEN_256 = 8'hb == RADDR ? 8'hb : _GEN_255; // @[RAM_ST.scala 32:46]
  assign _GEN_257 = 8'hc == RADDR ? 8'hc : _GEN_256; // @[RAM_ST.scala 32:46]
  assign _GEN_258 = 8'hd == RADDR ? 8'hd : _GEN_257; // @[RAM_ST.scala 32:46]
  assign _GEN_259 = 8'he == RADDR ? 8'he : _GEN_258; // @[RAM_ST.scala 32:46]
  assign _GEN_260 = 8'hf == RADDR ? 8'hf : _GEN_259; // @[RAM_ST.scala 32:46]
  assign _GEN_261 = 8'h10 == RADDR ? 8'h10 : _GEN_260; // @[RAM_ST.scala 32:46]
  assign _GEN_262 = 8'h11 == RADDR ? 8'h11 : _GEN_261; // @[RAM_ST.scala 32:46]
  assign _GEN_263 = 8'h12 == RADDR ? 8'h12 : _GEN_262; // @[RAM_ST.scala 32:46]
  assign _GEN_264 = 8'h13 == RADDR ? 8'h13 : _GEN_263; // @[RAM_ST.scala 32:46]
  assign _GEN_265 = 8'h14 == RADDR ? 8'h14 : _GEN_264; // @[RAM_ST.scala 32:46]
  assign _GEN_266 = 8'h15 == RADDR ? 8'h15 : _GEN_265; // @[RAM_ST.scala 32:46]
  assign _GEN_267 = 8'h16 == RADDR ? 8'h16 : _GEN_266; // @[RAM_ST.scala 32:46]
  assign _GEN_268 = 8'h17 == RADDR ? 8'h17 : _GEN_267; // @[RAM_ST.scala 32:46]
  assign _GEN_269 = 8'h18 == RADDR ? 8'h18 : _GEN_268; // @[RAM_ST.scala 32:46]
  assign _GEN_270 = 8'h19 == RADDR ? 8'h19 : _GEN_269; // @[RAM_ST.scala 32:46]
  assign _GEN_271 = 8'h1a == RADDR ? 8'h1a : _GEN_270; // @[RAM_ST.scala 32:46]
  assign _GEN_272 = 8'h1b == RADDR ? 8'h1b : _GEN_271; // @[RAM_ST.scala 32:46]
  assign _GEN_273 = 8'h1c == RADDR ? 8'h1c : _GEN_272; // @[RAM_ST.scala 32:46]
  assign _GEN_274 = 8'h1d == RADDR ? 8'h1d : _GEN_273; // @[RAM_ST.scala 32:46]
  assign _GEN_275 = 8'h1e == RADDR ? 8'h1e : _GEN_274; // @[RAM_ST.scala 32:46]
  assign _GEN_276 = 8'h1f == RADDR ? 8'h1f : _GEN_275; // @[RAM_ST.scala 32:46]
  assign _GEN_277 = 8'h20 == RADDR ? 8'h20 : _GEN_276; // @[RAM_ST.scala 32:46]
  assign _GEN_278 = 8'h21 == RADDR ? 8'h21 : _GEN_277; // @[RAM_ST.scala 32:46]
  assign _GEN_279 = 8'h22 == RADDR ? 8'h22 : _GEN_278; // @[RAM_ST.scala 32:46]
  assign _GEN_280 = 8'h23 == RADDR ? 8'h23 : _GEN_279; // @[RAM_ST.scala 32:46]
  assign _GEN_281 = 8'h24 == RADDR ? 8'h24 : _GEN_280; // @[RAM_ST.scala 32:46]
  assign _GEN_282 = 8'h25 == RADDR ? 8'h25 : _GEN_281; // @[RAM_ST.scala 32:46]
  assign _GEN_283 = 8'h26 == RADDR ? 8'h26 : _GEN_282; // @[RAM_ST.scala 32:46]
  assign _GEN_284 = 8'h27 == RADDR ? 8'h27 : _GEN_283; // @[RAM_ST.scala 32:46]
  assign _GEN_285 = 8'h28 == RADDR ? 8'h28 : _GEN_284; // @[RAM_ST.scala 32:46]
  assign _GEN_286 = 8'h29 == RADDR ? 8'h29 : _GEN_285; // @[RAM_ST.scala 32:46]
  assign _GEN_287 = 8'h2a == RADDR ? 8'h2a : _GEN_286; // @[RAM_ST.scala 32:46]
  assign _GEN_288 = 8'h2b == RADDR ? 8'h2b : _GEN_287; // @[RAM_ST.scala 32:46]
  assign _GEN_289 = 8'h2c == RADDR ? 8'h2c : _GEN_288; // @[RAM_ST.scala 32:46]
  assign _GEN_290 = 8'h2d == RADDR ? 8'h2d : _GEN_289; // @[RAM_ST.scala 32:46]
  assign _GEN_291 = 8'h2e == RADDR ? 8'h2e : _GEN_290; // @[RAM_ST.scala 32:46]
  assign _GEN_292 = 8'h2f == RADDR ? 8'h2f : _GEN_291; // @[RAM_ST.scala 32:46]
  assign _GEN_293 = 8'h30 == RADDR ? 8'h30 : _GEN_292; // @[RAM_ST.scala 32:46]
  assign _GEN_294 = 8'h31 == RADDR ? 8'h31 : _GEN_293; // @[RAM_ST.scala 32:46]
  assign _GEN_295 = 8'h32 == RADDR ? 8'h32 : _GEN_294; // @[RAM_ST.scala 32:46]
  assign _GEN_296 = 8'h33 == RADDR ? 8'h33 : _GEN_295; // @[RAM_ST.scala 32:46]
  assign _GEN_297 = 8'h34 == RADDR ? 8'h34 : _GEN_296; // @[RAM_ST.scala 32:46]
  assign _GEN_298 = 8'h35 == RADDR ? 8'h35 : _GEN_297; // @[RAM_ST.scala 32:46]
  assign _GEN_299 = 8'h36 == RADDR ? 8'h36 : _GEN_298; // @[RAM_ST.scala 32:46]
  assign _GEN_300 = 8'h37 == RADDR ? 8'h37 : _GEN_299; // @[RAM_ST.scala 32:46]
  assign _GEN_301 = 8'h38 == RADDR ? 8'h38 : _GEN_300; // @[RAM_ST.scala 32:46]
  assign _GEN_302 = 8'h39 == RADDR ? 8'h39 : _GEN_301; // @[RAM_ST.scala 32:46]
  assign _GEN_303 = 8'h3a == RADDR ? 8'h3a : _GEN_302; // @[RAM_ST.scala 32:46]
  assign _GEN_304 = 8'h3b == RADDR ? 8'h3b : _GEN_303; // @[RAM_ST.scala 32:46]
  assign _GEN_305 = 8'h3c == RADDR ? 8'h3c : _GEN_304; // @[RAM_ST.scala 32:46]
  assign _GEN_306 = 8'h3d == RADDR ? 8'h3d : _GEN_305; // @[RAM_ST.scala 32:46]
  assign _GEN_307 = 8'h3e == RADDR ? 8'h3e : _GEN_306; // @[RAM_ST.scala 32:46]
  assign _GEN_308 = 8'h3f == RADDR ? 8'h3f : _GEN_307; // @[RAM_ST.scala 32:46]
  assign _GEN_309 = 8'h40 == RADDR ? 8'h40 : _GEN_308; // @[RAM_ST.scala 32:46]
  assign _GEN_310 = 8'h41 == RADDR ? 8'h41 : _GEN_309; // @[RAM_ST.scala 32:46]
  assign _GEN_311 = 8'h42 == RADDR ? 8'h42 : _GEN_310; // @[RAM_ST.scala 32:46]
  assign _GEN_312 = 8'h43 == RADDR ? 8'h43 : _GEN_311; // @[RAM_ST.scala 32:46]
  assign _GEN_313 = 8'h44 == RADDR ? 8'h44 : _GEN_312; // @[RAM_ST.scala 32:46]
  assign _GEN_314 = 8'h45 == RADDR ? 8'h45 : _GEN_313; // @[RAM_ST.scala 32:46]
  assign _GEN_315 = 8'h46 == RADDR ? 8'h46 : _GEN_314; // @[RAM_ST.scala 32:46]
  assign _GEN_316 = 8'h47 == RADDR ? 8'h47 : _GEN_315; // @[RAM_ST.scala 32:46]
  assign _GEN_317 = 8'h48 == RADDR ? 8'h48 : _GEN_316; // @[RAM_ST.scala 32:46]
  assign _GEN_318 = 8'h49 == RADDR ? 8'h49 : _GEN_317; // @[RAM_ST.scala 32:46]
  assign _GEN_319 = 8'h4a == RADDR ? 8'h4a : _GEN_318; // @[RAM_ST.scala 32:46]
  assign _GEN_320 = 8'h4b == RADDR ? 8'h4b : _GEN_319; // @[RAM_ST.scala 32:46]
  assign _GEN_321 = 8'h4c == RADDR ? 8'h4c : _GEN_320; // @[RAM_ST.scala 32:46]
  assign _GEN_322 = 8'h4d == RADDR ? 8'h4d : _GEN_321; // @[RAM_ST.scala 32:46]
  assign _GEN_323 = 8'h4e == RADDR ? 8'h4e : _GEN_322; // @[RAM_ST.scala 32:46]
  assign _GEN_324 = 8'h4f == RADDR ? 8'h4f : _GEN_323; // @[RAM_ST.scala 32:46]
  assign _GEN_325 = 8'h50 == RADDR ? 8'h50 : _GEN_324; // @[RAM_ST.scala 32:46]
  assign _GEN_326 = 8'h51 == RADDR ? 8'h51 : _GEN_325; // @[RAM_ST.scala 32:46]
  assign _GEN_327 = 8'h52 == RADDR ? 8'h52 : _GEN_326; // @[RAM_ST.scala 32:46]
  assign _GEN_328 = 8'h53 == RADDR ? 8'h53 : _GEN_327; // @[RAM_ST.scala 32:46]
  assign _GEN_329 = 8'h54 == RADDR ? 8'h54 : _GEN_328; // @[RAM_ST.scala 32:46]
  assign _GEN_330 = 8'h55 == RADDR ? 8'h55 : _GEN_329; // @[RAM_ST.scala 32:46]
  assign _GEN_331 = 8'h56 == RADDR ? 8'h56 : _GEN_330; // @[RAM_ST.scala 32:46]
  assign _GEN_332 = 8'h57 == RADDR ? 8'h57 : _GEN_331; // @[RAM_ST.scala 32:46]
  assign _GEN_333 = 8'h58 == RADDR ? 8'h58 : _GEN_332; // @[RAM_ST.scala 32:46]
  assign _GEN_334 = 8'h59 == RADDR ? 8'h59 : _GEN_333; // @[RAM_ST.scala 32:46]
  assign _GEN_335 = 8'h5a == RADDR ? 8'h5a : _GEN_334; // @[RAM_ST.scala 32:46]
  assign _GEN_336 = 8'h5b == RADDR ? 8'h5b : _GEN_335; // @[RAM_ST.scala 32:46]
  assign _GEN_337 = 8'h5c == RADDR ? 8'h5c : _GEN_336; // @[RAM_ST.scala 32:46]
  assign _GEN_338 = 8'h5d == RADDR ? 8'h5d : _GEN_337; // @[RAM_ST.scala 32:46]
  assign _GEN_339 = 8'h5e == RADDR ? 8'h5e : _GEN_338; // @[RAM_ST.scala 32:46]
  assign _GEN_340 = 8'h5f == RADDR ? 8'h5f : _GEN_339; // @[RAM_ST.scala 32:46]
  assign _GEN_341 = 8'h60 == RADDR ? 8'h60 : _GEN_340; // @[RAM_ST.scala 32:46]
  assign _GEN_342 = 8'h61 == RADDR ? 8'h61 : _GEN_341; // @[RAM_ST.scala 32:46]
  assign _GEN_343 = 8'h62 == RADDR ? 8'h62 : _GEN_342; // @[RAM_ST.scala 32:46]
  assign _GEN_344 = 8'h63 == RADDR ? 8'h63 : _GEN_343; // @[RAM_ST.scala 32:46]
  assign _GEN_345 = 8'h64 == RADDR ? 8'h64 : _GEN_344; // @[RAM_ST.scala 32:46]
  assign _GEN_346 = 8'h65 == RADDR ? 8'h65 : _GEN_345; // @[RAM_ST.scala 32:46]
  assign _GEN_347 = 8'h66 == RADDR ? 8'h66 : _GEN_346; // @[RAM_ST.scala 32:46]
  assign _GEN_348 = 8'h67 == RADDR ? 8'h67 : _GEN_347; // @[RAM_ST.scala 32:46]
  assign _GEN_349 = 8'h68 == RADDR ? 8'h68 : _GEN_348; // @[RAM_ST.scala 32:46]
  assign _GEN_350 = 8'h69 == RADDR ? 8'h69 : _GEN_349; // @[RAM_ST.scala 32:46]
  assign _GEN_351 = 8'h6a == RADDR ? 8'h6a : _GEN_350; // @[RAM_ST.scala 32:46]
  assign _GEN_352 = 8'h6b == RADDR ? 8'h6b : _GEN_351; // @[RAM_ST.scala 32:46]
  assign _GEN_353 = 8'h6c == RADDR ? 8'h6c : _GEN_352; // @[RAM_ST.scala 32:46]
  assign _GEN_354 = 8'h6d == RADDR ? 8'h6d : _GEN_353; // @[RAM_ST.scala 32:46]
  assign _GEN_355 = 8'h6e == RADDR ? 8'h6e : _GEN_354; // @[RAM_ST.scala 32:46]
  assign _GEN_356 = 8'h6f == RADDR ? 8'h6f : _GEN_355; // @[RAM_ST.scala 32:46]
  assign _GEN_357 = 8'h70 == RADDR ? 8'h70 : _GEN_356; // @[RAM_ST.scala 32:46]
  assign _GEN_358 = 8'h71 == RADDR ? 8'h71 : _GEN_357; // @[RAM_ST.scala 32:46]
  assign _GEN_359 = 8'h72 == RADDR ? 8'h72 : _GEN_358; // @[RAM_ST.scala 32:46]
  assign _GEN_360 = 8'h73 == RADDR ? 8'h73 : _GEN_359; // @[RAM_ST.scala 32:46]
  assign _GEN_361 = 8'h74 == RADDR ? 8'h74 : _GEN_360; // @[RAM_ST.scala 32:46]
  assign _GEN_362 = 8'h75 == RADDR ? 8'h75 : _GEN_361; // @[RAM_ST.scala 32:46]
  assign _GEN_363 = 8'h76 == RADDR ? 8'h76 : _GEN_362; // @[RAM_ST.scala 32:46]
  assign _GEN_364 = 8'h77 == RADDR ? 8'h77 : _GEN_363; // @[RAM_ST.scala 32:46]
  assign _GEN_365 = 8'h78 == RADDR ? 8'h78 : _GEN_364; // @[RAM_ST.scala 32:46]
  assign _GEN_366 = 8'h79 == RADDR ? 8'h79 : _GEN_365; // @[RAM_ST.scala 32:46]
  assign _GEN_367 = 8'h7a == RADDR ? 8'h7a : _GEN_366; // @[RAM_ST.scala 32:46]
  assign _GEN_368 = 8'h7b == RADDR ? 8'h7b : _GEN_367; // @[RAM_ST.scala 32:46]
  assign _GEN_369 = 8'h7c == RADDR ? 8'h7c : _GEN_368; // @[RAM_ST.scala 32:46]
  assign _GEN_370 = 8'h7d == RADDR ? 8'h7d : _GEN_369; // @[RAM_ST.scala 32:46]
  assign _GEN_371 = 8'h7e == RADDR ? 8'h7e : _GEN_370; // @[RAM_ST.scala 32:46]
  assign _GEN_372 = 8'h7f == RADDR ? 8'h7f : _GEN_371; // @[RAM_ST.scala 32:46]
  assign _GEN_373 = 8'h80 == RADDR ? 8'h80 : _GEN_372; // @[RAM_ST.scala 32:46]
  assign _GEN_374 = 8'h81 == RADDR ? 8'h81 : _GEN_373; // @[RAM_ST.scala 32:46]
  assign _GEN_375 = 8'h82 == RADDR ? 8'h82 : _GEN_374; // @[RAM_ST.scala 32:46]
  assign _GEN_376 = 8'h83 == RADDR ? 8'h83 : _GEN_375; // @[RAM_ST.scala 32:46]
  assign _GEN_377 = 8'h84 == RADDR ? 8'h84 : _GEN_376; // @[RAM_ST.scala 32:46]
  assign _GEN_378 = 8'h85 == RADDR ? 8'h85 : _GEN_377; // @[RAM_ST.scala 32:46]
  assign _GEN_379 = 8'h86 == RADDR ? 8'h86 : _GEN_378; // @[RAM_ST.scala 32:46]
  assign _GEN_380 = 8'h87 == RADDR ? 8'h87 : _GEN_379; // @[RAM_ST.scala 32:46]
  assign _GEN_381 = 8'h88 == RADDR ? 8'h88 : _GEN_380; // @[RAM_ST.scala 32:46]
  assign _GEN_382 = 8'h89 == RADDR ? 8'h89 : _GEN_381; // @[RAM_ST.scala 32:46]
  assign _GEN_383 = 8'h8a == RADDR ? 8'h8a : _GEN_382; // @[RAM_ST.scala 32:46]
  assign _GEN_384 = 8'h8b == RADDR ? 8'h8b : _GEN_383; // @[RAM_ST.scala 32:46]
  assign _GEN_385 = 8'h8c == RADDR ? 8'h8c : _GEN_384; // @[RAM_ST.scala 32:46]
  assign _GEN_386 = 8'h8d == RADDR ? 8'h8d : _GEN_385; // @[RAM_ST.scala 32:46]
  assign _GEN_387 = 8'h8e == RADDR ? 8'h8e : _GEN_386; // @[RAM_ST.scala 32:46]
  assign _GEN_388 = 8'h8f == RADDR ? 8'h8f : _GEN_387; // @[RAM_ST.scala 32:46]
  assign _GEN_389 = 8'h90 == RADDR ? 8'h90 : _GEN_388; // @[RAM_ST.scala 32:46]
  assign _GEN_390 = 8'h91 == RADDR ? 8'h91 : _GEN_389; // @[RAM_ST.scala 32:46]
  assign _GEN_391 = 8'h92 == RADDR ? 8'h92 : _GEN_390; // @[RAM_ST.scala 32:46]
  assign _GEN_392 = 8'h93 == RADDR ? 8'h93 : _GEN_391; // @[RAM_ST.scala 32:46]
  assign _GEN_393 = 8'h94 == RADDR ? 8'h94 : _GEN_392; // @[RAM_ST.scala 32:46]
  assign _GEN_394 = 8'h95 == RADDR ? 8'h95 : _GEN_393; // @[RAM_ST.scala 32:46]
  assign _GEN_395 = 8'h96 == RADDR ? 8'h96 : _GEN_394; // @[RAM_ST.scala 32:46]
  assign _GEN_396 = 8'h97 == RADDR ? 8'h97 : _GEN_395; // @[RAM_ST.scala 32:46]
  assign _GEN_397 = 8'h98 == RADDR ? 8'h98 : _GEN_396; // @[RAM_ST.scala 32:46]
  assign _GEN_398 = 8'h99 == RADDR ? 8'h99 : _GEN_397; // @[RAM_ST.scala 32:46]
  assign _GEN_399 = 8'h9a == RADDR ? 8'h9a : _GEN_398; // @[RAM_ST.scala 32:46]
  assign _GEN_400 = 8'h9b == RADDR ? 8'h9b : _GEN_399; // @[RAM_ST.scala 32:46]
  assign _GEN_401 = 8'h9c == RADDR ? 8'h9c : _GEN_400; // @[RAM_ST.scala 32:46]
  assign _GEN_402 = 8'h9d == RADDR ? 8'h9d : _GEN_401; // @[RAM_ST.scala 32:46]
  assign _GEN_403 = 8'h9e == RADDR ? 8'h9e : _GEN_402; // @[RAM_ST.scala 32:46]
  assign _GEN_404 = 8'h9f == RADDR ? 8'h9f : _GEN_403; // @[RAM_ST.scala 32:46]
  assign _GEN_405 = 8'ha0 == RADDR ? 8'ha0 : _GEN_404; // @[RAM_ST.scala 32:46]
  assign _GEN_406 = 8'ha1 == RADDR ? 8'ha1 : _GEN_405; // @[RAM_ST.scala 32:46]
  assign _GEN_407 = 8'ha2 == RADDR ? 8'ha2 : _GEN_406; // @[RAM_ST.scala 32:46]
  assign _GEN_408 = 8'ha3 == RADDR ? 8'ha3 : _GEN_407; // @[RAM_ST.scala 32:46]
  assign _GEN_409 = 8'ha4 == RADDR ? 8'ha4 : _GEN_408; // @[RAM_ST.scala 32:46]
  assign _GEN_410 = 8'ha5 == RADDR ? 8'ha5 : _GEN_409; // @[RAM_ST.scala 32:46]
  assign _GEN_411 = 8'ha6 == RADDR ? 8'ha6 : _GEN_410; // @[RAM_ST.scala 32:46]
  assign _GEN_412 = 8'ha7 == RADDR ? 8'ha7 : _GEN_411; // @[RAM_ST.scala 32:46]
  assign _GEN_413 = 8'ha8 == RADDR ? 8'ha8 : _GEN_412; // @[RAM_ST.scala 32:46]
  assign _GEN_414 = 8'ha9 == RADDR ? 8'ha9 : _GEN_413; // @[RAM_ST.scala 32:46]
  assign _GEN_415 = 8'haa == RADDR ? 8'haa : _GEN_414; // @[RAM_ST.scala 32:46]
  assign _GEN_416 = 8'hab == RADDR ? 8'hab : _GEN_415; // @[RAM_ST.scala 32:46]
  assign _GEN_417 = 8'hac == RADDR ? 8'hac : _GEN_416; // @[RAM_ST.scala 32:46]
  assign _GEN_418 = 8'had == RADDR ? 8'had : _GEN_417; // @[RAM_ST.scala 32:46]
  assign _GEN_419 = 8'hae == RADDR ? 8'hae : _GEN_418; // @[RAM_ST.scala 32:46]
  assign _GEN_420 = 8'haf == RADDR ? 8'haf : _GEN_419; // @[RAM_ST.scala 32:46]
  assign _GEN_421 = 8'hb0 == RADDR ? 8'hb0 : _GEN_420; // @[RAM_ST.scala 32:46]
  assign _GEN_422 = 8'hb1 == RADDR ? 8'hb1 : _GEN_421; // @[RAM_ST.scala 32:46]
  assign _GEN_423 = 8'hb2 == RADDR ? 8'hb2 : _GEN_422; // @[RAM_ST.scala 32:46]
  assign _GEN_424 = 8'hb3 == RADDR ? 8'hb3 : _GEN_423; // @[RAM_ST.scala 32:46]
  assign _GEN_425 = 8'hb4 == RADDR ? 8'hb4 : _GEN_424; // @[RAM_ST.scala 32:46]
  assign _GEN_426 = 8'hb5 == RADDR ? 8'hb5 : _GEN_425; // @[RAM_ST.scala 32:46]
  assign _GEN_427 = 8'hb6 == RADDR ? 8'hb6 : _GEN_426; // @[RAM_ST.scala 32:46]
  assign _GEN_428 = 8'hb7 == RADDR ? 8'hb7 : _GEN_427; // @[RAM_ST.scala 32:46]
  assign _GEN_429 = 8'hb8 == RADDR ? 8'hb8 : _GEN_428; // @[RAM_ST.scala 32:46]
  assign _GEN_430 = 8'hb9 == RADDR ? 8'hb9 : _GEN_429; // @[RAM_ST.scala 32:46]
  assign _GEN_431 = 8'hba == RADDR ? 8'hba : _GEN_430; // @[RAM_ST.scala 32:46]
  assign _GEN_432 = 8'hbb == RADDR ? 8'hbb : _GEN_431; // @[RAM_ST.scala 32:46]
  assign _GEN_433 = 8'hbc == RADDR ? 8'hbc : _GEN_432; // @[RAM_ST.scala 32:46]
  assign _GEN_434 = 8'hbd == RADDR ? 8'hbd : _GEN_433; // @[RAM_ST.scala 32:46]
  assign _GEN_435 = 8'hbe == RADDR ? 8'hbe : _GEN_434; // @[RAM_ST.scala 32:46]
  assign _GEN_436 = 8'hbf == RADDR ? 8'hbf : _GEN_435; // @[RAM_ST.scala 32:46]
  assign _GEN_437 = 8'hc0 == RADDR ? 8'hc0 : _GEN_436; // @[RAM_ST.scala 32:46]
  assign _GEN_438 = 8'hc1 == RADDR ? 8'hc1 : _GEN_437; // @[RAM_ST.scala 32:46]
  assign _GEN_439 = 8'hc2 == RADDR ? 8'hc2 : _GEN_438; // @[RAM_ST.scala 32:46]
  assign _GEN_440 = 8'hc3 == RADDR ? 8'hc3 : _GEN_439; // @[RAM_ST.scala 32:46]
  assign _GEN_441 = 8'hc4 == RADDR ? 8'hc4 : _GEN_440; // @[RAM_ST.scala 32:46]
  assign _GEN_442 = 8'hc5 == RADDR ? 8'hc5 : _GEN_441; // @[RAM_ST.scala 32:46]
  assign _GEN_443 = 8'hc6 == RADDR ? 8'hc6 : _GEN_442; // @[RAM_ST.scala 32:46]
  assign _GEN_444 = 8'hc7 == RADDR ? 8'hc7 : _GEN_443; // @[RAM_ST.scala 32:46]
  assign _GEN_445 = 8'hc8 == RADDR ? 8'hc8 : _GEN_444; // @[RAM_ST.scala 32:46]
  assign _GEN_446 = 8'hc9 == RADDR ? 8'hc9 : _GEN_445; // @[RAM_ST.scala 32:46]
  assign _GEN_447 = 8'hca == RADDR ? 8'hca : _GEN_446; // @[RAM_ST.scala 32:46]
  assign _GEN_448 = 8'hcb == RADDR ? 8'hcb : _GEN_447; // @[RAM_ST.scala 32:46]
  assign _GEN_449 = 8'hcc == RADDR ? 8'hcc : _GEN_448; // @[RAM_ST.scala 32:46]
  assign _GEN_450 = 8'hcd == RADDR ? 8'hcd : _GEN_449; // @[RAM_ST.scala 32:46]
  assign _GEN_451 = 8'hce == RADDR ? 8'hce : _GEN_450; // @[RAM_ST.scala 32:46]
  assign _GEN_452 = 8'hcf == RADDR ? 8'hcf : _GEN_451; // @[RAM_ST.scala 32:46]
  assign _GEN_453 = 8'hd0 == RADDR ? 8'hd0 : _GEN_452; // @[RAM_ST.scala 32:46]
  assign _GEN_454 = 8'hd1 == RADDR ? 8'hd1 : _GEN_453; // @[RAM_ST.scala 32:46]
  assign _GEN_455 = 8'hd2 == RADDR ? 8'hd2 : _GEN_454; // @[RAM_ST.scala 32:46]
  assign _GEN_456 = 8'hd3 == RADDR ? 8'hd3 : _GEN_455; // @[RAM_ST.scala 32:46]
  assign _GEN_457 = 8'hd4 == RADDR ? 8'hd4 : _GEN_456; // @[RAM_ST.scala 32:46]
  assign _GEN_458 = 8'hd5 == RADDR ? 8'hd5 : _GEN_457; // @[RAM_ST.scala 32:46]
  assign _GEN_459 = 8'hd6 == RADDR ? 8'hd6 : _GEN_458; // @[RAM_ST.scala 32:46]
  assign _GEN_460 = 8'hd7 == RADDR ? 8'hd7 : _GEN_459; // @[RAM_ST.scala 32:46]
  assign _GEN_461 = 8'hd8 == RADDR ? 8'hd8 : _GEN_460; // @[RAM_ST.scala 32:46]
  assign _GEN_462 = 8'hd9 == RADDR ? 8'hd9 : _GEN_461; // @[RAM_ST.scala 32:46]
  assign _GEN_463 = 8'hda == RADDR ? 8'hda : _GEN_462; // @[RAM_ST.scala 32:46]
  assign _GEN_464 = 8'hdb == RADDR ? 8'hdb : _GEN_463; // @[RAM_ST.scala 32:46]
  assign _GEN_465 = 8'hdc == RADDR ? 8'hdc : _GEN_464; // @[RAM_ST.scala 32:46]
  assign _GEN_466 = 8'hdd == RADDR ? 8'hdd : _GEN_465; // @[RAM_ST.scala 32:46]
  assign _GEN_467 = 8'hde == RADDR ? 8'hde : _GEN_466; // @[RAM_ST.scala 32:46]
  assign _GEN_468 = 8'hdf == RADDR ? 8'hdf : _GEN_467; // @[RAM_ST.scala 32:46]
  assign _GEN_469 = 8'he0 == RADDR ? 8'he0 : _GEN_468; // @[RAM_ST.scala 32:46]
  assign _GEN_470 = 8'he1 == RADDR ? 8'he1 : _GEN_469; // @[RAM_ST.scala 32:46]
  assign _GEN_471 = 8'he2 == RADDR ? 8'he2 : _GEN_470; // @[RAM_ST.scala 32:46]
  assign _GEN_472 = 8'he3 == RADDR ? 8'he3 : _GEN_471; // @[RAM_ST.scala 32:46]
  assign _GEN_473 = 8'he4 == RADDR ? 8'he4 : _GEN_472; // @[RAM_ST.scala 32:46]
  assign _GEN_474 = 8'he5 == RADDR ? 8'he5 : _GEN_473; // @[RAM_ST.scala 32:46]
  assign _GEN_475 = 8'he6 == RADDR ? 8'he6 : _GEN_474; // @[RAM_ST.scala 32:46]
  assign _GEN_476 = 8'he7 == RADDR ? 8'he7 : _GEN_475; // @[RAM_ST.scala 32:46]
  assign _GEN_477 = 8'he8 == RADDR ? 8'he8 : _GEN_476; // @[RAM_ST.scala 32:46]
  assign _GEN_478 = 8'he9 == RADDR ? 8'he9 : _GEN_477; // @[RAM_ST.scala 32:46]
  assign _GEN_479 = 8'hea == RADDR ? 8'hea : _GEN_478; // @[RAM_ST.scala 32:46]
  assign _GEN_480 = 8'heb == RADDR ? 8'heb : _GEN_479; // @[RAM_ST.scala 32:46]
  assign _GEN_481 = 8'hec == RADDR ? 8'hec : _GEN_480; // @[RAM_ST.scala 32:46]
  assign _GEN_482 = 8'hed == RADDR ? 8'hed : _GEN_481; // @[RAM_ST.scala 32:46]
  assign _GEN_483 = 8'hee == RADDR ? 8'hee : _GEN_482; // @[RAM_ST.scala 32:46]
  assign _GEN_484 = 8'hef == RADDR ? 8'hef : _GEN_483; // @[RAM_ST.scala 32:46]
  assign _T_10 = {{1'd0}, _GEN_484}; // @[RAM_ST.scala 32:46]
  assign _T_17 = ram__T_15_data;
  assign RDATA_0 = _T_17[31:0]; // @[RAM_ST.scala 32:9]
  assign RDATA_1 = _T_17[63:32]; // @[RAM_ST.scala 32:9]
  assign RDATA_2 = _T_17[95:64]; // @[RAM_ST.scala 32:9]
  assign RDATA_3 = _T_17[127:96]; // @[RAM_ST.scala 32:9]
  assign RDATA_4 = _T_17[159:128]; // @[RAM_ST.scala 32:9]
  assign RDATA_5 = _T_17[191:160]; // @[RAM_ST.scala 32:9]
  assign RDATA_6 = _T_17[223:192]; // @[RAM_ST.scala 32:9]
  assign RDATA_7 = _T_17[255:224]; // @[RAM_ST.scala 32:9]
  assign write_elem_counter_CE = WE; // @[RAM_ST.scala 23:25]
  assign read_elem_counter_CE = RE; // @[RAM_ST.scala 24:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {8{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 240; initvar = initvar+1)
    ram[initvar] = _RAND_0[255:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {8{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram__T_15_en_pipe_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  ram__T_15_addr_pipe_0 = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram__T_9_en & ram__T_9_mask) begin
      ram[ram__T_9_addr] <= ram__T_9_data; // @[RAM_ST.scala 29:24]
    end
    ram__T_15_en_pipe_0 <= read_elem_counter_valid;
    if (read_elem_counter_valid) begin
      ram__T_15_addr_pipe_0 <= _T_10[7:0];
    end
  end
endmodule
module ShiftT(
  input         clock,
  input         reset,
  input         valid_up,
  input  [31:0] I_0,
  input  [31:0] I_1,
  input  [31:0] I_2,
  input  [31:0] I_3,
  input  [31:0] I_4,
  input  [31:0] I_5,
  input  [31:0] I_6,
  input  [31:0] I_7,
  output [31:0] O_0,
  output [31:0] O_1,
  output [31:0] O_2,
  output [31:0] O_3,
  output [31:0] O_4,
  output [31:0] O_5,
  output [31:0] O_6,
  output [31:0] O_7
);
  wire  RAM_ST_clock; // @[ShiftT.scala 39:29]
  wire  RAM_ST_RE; // @[ShiftT.scala 39:29]
  wire [7:0] RAM_ST_RADDR; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_RDATA_0; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_RDATA_1; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_RDATA_2; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_RDATA_3; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_RDATA_4; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_RDATA_5; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_RDATA_6; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_RDATA_7; // @[ShiftT.scala 39:29]
  wire  RAM_ST_WE; // @[ShiftT.scala 39:29]
  wire [7:0] RAM_ST_WADDR; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_WDATA_0; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_WDATA_1; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_WDATA_2; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_WDATA_3; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_WDATA_4; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_WDATA_5; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_WDATA_6; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_WDATA_7; // @[ShiftT.scala 39:29]
  wire  NestedCounters_CE; // @[ShiftT.scala 41:31]
  wire  NestedCounters_valid; // @[ShiftT.scala 41:31]
  reg [7:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[Counter.scala 37:24]
  wire [7:0] _T_3; // @[Counter.scala 38:22]
  RAM_ST RAM_ST ( // @[ShiftT.scala 39:29]
    .clock(RAM_ST_clock),
    .RE(RAM_ST_RE),
    .RADDR(RAM_ST_RADDR),
    .RDATA_0(RAM_ST_RDATA_0),
    .RDATA_1(RAM_ST_RDATA_1),
    .RDATA_2(RAM_ST_RDATA_2),
    .RDATA_3(RAM_ST_RDATA_3),
    .RDATA_4(RAM_ST_RDATA_4),
    .RDATA_5(RAM_ST_RDATA_5),
    .RDATA_6(RAM_ST_RDATA_6),
    .RDATA_7(RAM_ST_RDATA_7),
    .WE(RAM_ST_WE),
    .WADDR(RAM_ST_WADDR),
    .WDATA_0(RAM_ST_WDATA_0),
    .WDATA_1(RAM_ST_WDATA_1),
    .WDATA_2(RAM_ST_WDATA_2),
    .WDATA_3(RAM_ST_WDATA_3),
    .WDATA_4(RAM_ST_WDATA_4),
    .WDATA_5(RAM_ST_WDATA_5),
    .WDATA_6(RAM_ST_WDATA_6),
    .WDATA_7(RAM_ST_WDATA_7)
  );
  NestedCounters_1 NestedCounters ( // @[ShiftT.scala 41:31]
    .CE(NestedCounters_CE),
    .valid(NestedCounters_valid)
  );
  assign _T_1 = value == 8'hef; // @[Counter.scala 37:24]
  assign _T_3 = value + 8'h1; // @[Counter.scala 38:22]
  assign O_0 = RAM_ST_RDATA_0; // @[ShiftT.scala 51:7]
  assign O_1 = RAM_ST_RDATA_1; // @[ShiftT.scala 51:7]
  assign O_2 = RAM_ST_RDATA_2; // @[ShiftT.scala 51:7]
  assign O_3 = RAM_ST_RDATA_3; // @[ShiftT.scala 51:7]
  assign O_4 = RAM_ST_RDATA_4; // @[ShiftT.scala 51:7]
  assign O_5 = RAM_ST_RDATA_5; // @[ShiftT.scala 51:7]
  assign O_6 = RAM_ST_RDATA_6; // @[ShiftT.scala 51:7]
  assign O_7 = RAM_ST_RDATA_7; // @[ShiftT.scala 51:7]
  assign RAM_ST_clock = clock;
  assign RAM_ST_RE = valid_up; // @[ShiftT.scala 49:20]
  assign RAM_ST_RADDR = _T_1 ? 8'h0 : _T_3; // @[ShiftT.scala 46:76 ShiftT.scala 47:38]
  assign RAM_ST_WE = valid_up; // @[ShiftT.scala 48:20]
  assign RAM_ST_WADDR = value; // @[ShiftT.scala 45:23]
  assign RAM_ST_WDATA_0 = I_0; // @[ShiftT.scala 50:23]
  assign RAM_ST_WDATA_1 = I_1; // @[ShiftT.scala 50:23]
  assign RAM_ST_WDATA_2 = I_2; // @[ShiftT.scala 50:23]
  assign RAM_ST_WDATA_3 = I_3; // @[ShiftT.scala 50:23]
  assign RAM_ST_WDATA_4 = I_4; // @[ShiftT.scala 50:23]
  assign RAM_ST_WDATA_5 = I_5; // @[ShiftT.scala 50:23]
  assign RAM_ST_WDATA_6 = I_6; // @[ShiftT.scala 50:23]
  assign RAM_ST_WDATA_7 = I_7; // @[ShiftT.scala 50:23]
  assign NestedCounters_CE = valid_up; // @[ShiftT.scala 42:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 8'h0;
    end else if (valid_up) begin
      if (_T_1) begin
        value <= 8'h0;
      end else begin
        value <= _T_3;
      end
    end
  end
endmodule
module ShiftTS(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0,
  input  [31:0] I_1,
  input  [31:0] I_2,
  input  [31:0] I_3,
  input  [31:0] I_4,
  input  [31:0] I_5,
  input  [31:0] I_6,
  input  [31:0] I_7,
  output [31:0] O_0,
  output [31:0] O_1,
  output [31:0] O_2,
  output [31:0] O_3,
  output [31:0] O_4,
  output [31:0] O_5,
  output [31:0] O_6,
  output [31:0] O_7
);
  wire  ShiftT_clock; // @[ShiftTS.scala 32:26]
  wire  ShiftT_reset; // @[ShiftTS.scala 32:26]
  wire  ShiftT_valid_up; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_I_0; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_I_1; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_I_2; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_I_3; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_I_4; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_I_5; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_I_6; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_I_7; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_O_0; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_O_1; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_O_2; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_O_3; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_O_4; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_O_5; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_O_6; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_O_7; // @[ShiftTS.scala 32:26]
  ShiftT ShiftT ( // @[ShiftTS.scala 32:26]
    .clock(ShiftT_clock),
    .reset(ShiftT_reset),
    .valid_up(ShiftT_valid_up),
    .I_0(ShiftT_I_0),
    .I_1(ShiftT_I_1),
    .I_2(ShiftT_I_2),
    .I_3(ShiftT_I_3),
    .I_4(ShiftT_I_4),
    .I_5(ShiftT_I_5),
    .I_6(ShiftT_I_6),
    .I_7(ShiftT_I_7),
    .O_0(ShiftT_O_0),
    .O_1(ShiftT_O_1),
    .O_2(ShiftT_O_2),
    .O_3(ShiftT_O_3),
    .O_4(ShiftT_O_4),
    .O_5(ShiftT_O_5),
    .O_6(ShiftT_O_6),
    .O_7(ShiftT_O_7)
  );
  assign valid_down = valid_up; // @[ShiftTS.scala 58:14]
  assign O_0 = ShiftT_O_0; // @[ShiftTS.scala 51:36]
  assign O_1 = ShiftT_O_1; // @[ShiftTS.scala 51:36]
  assign O_2 = ShiftT_O_2; // @[ShiftTS.scala 51:36]
  assign O_3 = ShiftT_O_3; // @[ShiftTS.scala 51:36]
  assign O_4 = ShiftT_O_4; // @[ShiftTS.scala 51:36]
  assign O_5 = ShiftT_O_5; // @[ShiftTS.scala 51:36]
  assign O_6 = ShiftT_O_6; // @[ShiftTS.scala 51:36]
  assign O_7 = ShiftT_O_7; // @[ShiftTS.scala 51:36]
  assign ShiftT_clock = clock;
  assign ShiftT_reset = reset;
  assign ShiftT_valid_up = valid_up; // @[ShiftTS.scala 53:29]
  assign ShiftT_I_0 = I_0; // @[ShiftTS.scala 50:25]
  assign ShiftT_I_1 = I_1; // @[ShiftTS.scala 50:25]
  assign ShiftT_I_2 = I_2; // @[ShiftTS.scala 50:25]
  assign ShiftT_I_3 = I_3; // @[ShiftTS.scala 50:25]
  assign ShiftT_I_4 = I_4; // @[ShiftTS.scala 50:25]
  assign ShiftT_I_5 = I_5; // @[ShiftTS.scala 50:25]
  assign ShiftT_I_6 = I_6; // @[ShiftTS.scala 50:25]
  assign ShiftT_I_7 = I_7; // @[ShiftTS.scala 50:25]
endmodule
module ShiftT_2(
  input         clock,
  input  [31:0] I_0,
  output [31:0] O_0
);
  reg [31:0] _T_0; // @[ShiftT.scala 24:82]
  reg [31:0] _RAND_0;
  assign O_0 = _T_0; // @[ShiftT.scala 24:7]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_0 <= I_0;
  end
endmodule
module ShiftTS_2(
  input         clock,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0,
  input  [31:0] I_1,
  input  [31:0] I_2,
  input  [31:0] I_3,
  input  [31:0] I_4,
  input  [31:0] I_5,
  input  [31:0] I_6,
  input  [31:0] I_7,
  output [31:0] O_0,
  output [31:0] O_1,
  output [31:0] O_2,
  output [31:0] O_3,
  output [31:0] O_4,
  output [31:0] O_5,
  output [31:0] O_6,
  output [31:0] O_7
);
  wire  ShiftT_clock; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_I_0; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_O_0; // @[ShiftTS.scala 32:26]
  ShiftT_2 ShiftT ( // @[ShiftTS.scala 32:26]
    .clock(ShiftT_clock),
    .I_0(ShiftT_I_0),
    .O_0(ShiftT_O_0)
  );
  assign valid_down = valid_up; // @[ShiftTS.scala 58:14]
  assign O_0 = ShiftT_O_0; // @[ShiftTS.scala 51:36]
  assign O_1 = I_0; // @[ShiftTS.scala 40:36]
  assign O_2 = I_1; // @[ShiftTS.scala 40:36]
  assign O_3 = I_2; // @[ShiftTS.scala 40:36]
  assign O_4 = I_3; // @[ShiftTS.scala 40:36]
  assign O_5 = I_4; // @[ShiftTS.scala 40:36]
  assign O_6 = I_5; // @[ShiftTS.scala 40:36]
  assign O_7 = I_6; // @[ShiftTS.scala 40:36]
  assign ShiftT_clock = clock;
  assign ShiftT_I_0 = I_7; // @[ShiftTS.scala 50:25]
endmodule
module SSeqTupleCreator(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0,
  input  [31:0] I1,
  output [31:0] O_0,
  output [31:0] O_1
);
  assign valid_down = valid_up; // @[Tuple.scala 15:14]
  assign O_0 = I0; // @[Tuple.scala 12:32]
  assign O_1 = I1; // @[Tuple.scala 13:32]
endmodule
module Map2S(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0,
  input  [31:0] I0_1,
  input  [31:0] I0_2,
  input  [31:0] I0_3,
  input  [31:0] I0_4,
  input  [31:0] I0_5,
  input  [31:0] I0_6,
  input  [31:0] I0_7,
  input  [31:0] I1_0,
  input  [31:0] I1_1,
  input  [31:0] I1_2,
  input  [31:0] I1_3,
  input  [31:0] I1_4,
  input  [31:0] I1_5,
  input  [31:0] I1_6,
  input  [31:0] I1_7,
  output [31:0] O_0_0,
  output [31:0] O_0_1,
  output [31:0] O_1_0,
  output [31:0] O_1_1,
  output [31:0] O_2_0,
  output [31:0] O_2_1,
  output [31:0] O_3_0,
  output [31:0] O_3_1,
  output [31:0] O_4_0,
  output [31:0] O_4_1,
  output [31:0] O_5_0,
  output [31:0] O_5_1,
  output [31:0] O_6_0,
  output [31:0] O_6_1,
  output [31:0] O_7_0,
  output [31:0] O_7_1
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_1; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_1; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  wire  _T_2; // @[Map2S.scala 26:83]
  wire  _T_3; // @[Map2S.scala 26:83]
  wire  _T_4; // @[Map2S.scala 26:83]
  wire  _T_5; // @[Map2S.scala 26:83]
  SSeqTupleCreator fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1(fst_op_I1),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1)
  );
  SSeqTupleCreator other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0(other_ops_0_I0),
    .I1(other_ops_0_I1),
    .O_0(other_ops_0_O_0),
    .O_1(other_ops_0_O_1)
  );
  SSeqTupleCreator other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0(other_ops_1_I0),
    .I1(other_ops_1_I1),
    .O_0(other_ops_1_O_0),
    .O_1(other_ops_1_O_1)
  );
  SSeqTupleCreator other_ops_2 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0(other_ops_2_I0),
    .I1(other_ops_2_I1),
    .O_0(other_ops_2_O_0),
    .O_1(other_ops_2_O_1)
  );
  SSeqTupleCreator other_ops_3 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I0(other_ops_3_I0),
    .I1(other_ops_3_I1),
    .O_0(other_ops_3_O_0),
    .O_1(other_ops_3_O_1)
  );
  SSeqTupleCreator other_ops_4 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I0(other_ops_4_I0),
    .I1(other_ops_4_I1),
    .O_0(other_ops_4_O_0),
    .O_1(other_ops_4_O_1)
  );
  SSeqTupleCreator other_ops_5 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I0(other_ops_5_I0),
    .I1(other_ops_5_I1),
    .O_0(other_ops_5_O_0),
    .O_1(other_ops_5_O_1)
  );
  SSeqTupleCreator other_ops_6 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I0(other_ops_6_I0),
    .I1(other_ops_6_I1),
    .O_0(other_ops_6_O_0),
    .O_1(other_ops_6_O_1)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[Map2S.scala 26:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[Map2S.scala 26:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_5 & other_ops_6_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0 = fst_op_O_0; // @[Map2S.scala 19:8]
  assign O_0_1 = fst_op_O_1; // @[Map2S.scala 19:8]
  assign O_1_0 = other_ops_0_O_0; // @[Map2S.scala 24:12]
  assign O_1_1 = other_ops_0_O_1; // @[Map2S.scala 24:12]
  assign O_2_0 = other_ops_1_O_0; // @[Map2S.scala 24:12]
  assign O_2_1 = other_ops_1_O_1; // @[Map2S.scala 24:12]
  assign O_3_0 = other_ops_2_O_0; // @[Map2S.scala 24:12]
  assign O_3_1 = other_ops_2_O_1; // @[Map2S.scala 24:12]
  assign O_4_0 = other_ops_3_O_0; // @[Map2S.scala 24:12]
  assign O_4_1 = other_ops_3_O_1; // @[Map2S.scala 24:12]
  assign O_5_0 = other_ops_4_O_0; // @[Map2S.scala 24:12]
  assign O_5_1 = other_ops_4_O_1; // @[Map2S.scala 24:12]
  assign O_6_0 = other_ops_5_O_0; // @[Map2S.scala 24:12]
  assign O_6_1 = other_ops_5_O_1; // @[Map2S.scala 24:12]
  assign O_7_0 = other_ops_6_O_0; // @[Map2S.scala 24:12]
  assign O_7_1 = other_ops_6_O_1; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0 = I0_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I1 = I1_1; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0 = I0_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1 = I1_2; // @[Map2S.scala 23:43]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0 = I0_3; // @[Map2S.scala 22:43]
  assign other_ops_2_I1 = I1_3; // @[Map2S.scala 23:43]
  assign other_ops_3_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_3_I0 = I0_4; // @[Map2S.scala 22:43]
  assign other_ops_3_I1 = I1_4; // @[Map2S.scala 23:43]
  assign other_ops_4_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_4_I0 = I0_5; // @[Map2S.scala 22:43]
  assign other_ops_4_I1 = I1_5; // @[Map2S.scala 23:43]
  assign other_ops_5_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_5_I0 = I0_6; // @[Map2S.scala 22:43]
  assign other_ops_5_I1 = I1_6; // @[Map2S.scala 23:43]
  assign other_ops_6_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_6_I0 = I0_7; // @[Map2S.scala 22:43]
  assign other_ops_6_I1 = I1_7; // @[Map2S.scala 23:43]
endmodule
module Map2T(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0,
  input  [31:0] I0_1,
  input  [31:0] I0_2,
  input  [31:0] I0_3,
  input  [31:0] I0_4,
  input  [31:0] I0_5,
  input  [31:0] I0_6,
  input  [31:0] I0_7,
  input  [31:0] I1_0,
  input  [31:0] I1_1,
  input  [31:0] I1_2,
  input  [31:0] I1_3,
  input  [31:0] I1_4,
  input  [31:0] I1_5,
  input  [31:0] I1_6,
  input  [31:0] I1_7,
  output [31:0] O_0_0,
  output [31:0] O_0_1,
  output [31:0] O_1_0,
  output [31:0] O_1_1,
  output [31:0] O_2_0,
  output [31:0] O_2_1,
  output [31:0] O_3_0,
  output [31:0] O_3_1,
  output [31:0] O_4_0,
  output [31:0] O_4_1,
  output [31:0] O_5_0,
  output [31:0] O_5_1,
  output [31:0] O_6_0,
  output [31:0] O_6_1,
  output [31:0] O_7_0,
  output [31:0] O_7_1
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_3; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_4; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_5; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_6; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_7; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_1; // @[Map2T.scala 8:20]
  Map2S op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0(op_I0_0),
    .I0_1(op_I0_1),
    .I0_2(op_I0_2),
    .I0_3(op_I0_3),
    .I0_4(op_I0_4),
    .I0_5(op_I0_5),
    .I0_6(op_I0_6),
    .I0_7(op_I0_7),
    .I1_0(op_I1_0),
    .I1_1(op_I1_1),
    .I1_2(op_I1_2),
    .I1_3(op_I1_3),
    .I1_4(op_I1_4),
    .I1_5(op_I1_5),
    .I1_6(op_I1_6),
    .I1_7(op_I1_7),
    .O_0_0(op_O_0_0),
    .O_0_1(op_O_0_1),
    .O_1_0(op_O_1_0),
    .O_1_1(op_O_1_1),
    .O_2_0(op_O_2_0),
    .O_2_1(op_O_2_1),
    .O_3_0(op_O_3_0),
    .O_3_1(op_O_3_1),
    .O_4_0(op_O_4_0),
    .O_4_1(op_O_4_1),
    .O_5_0(op_O_5_0),
    .O_5_1(op_O_5_1),
    .O_6_0(op_O_6_0),
    .O_6_1(op_O_6_1),
    .O_7_0(op_O_7_0),
    .O_7_1(op_O_7_1)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_0 = op_O_0_0; // @[Map2T.scala 17:7]
  assign O_0_1 = op_O_0_1; // @[Map2T.scala 17:7]
  assign O_1_0 = op_O_1_0; // @[Map2T.scala 17:7]
  assign O_1_1 = op_O_1_1; // @[Map2T.scala 17:7]
  assign O_2_0 = op_O_2_0; // @[Map2T.scala 17:7]
  assign O_2_1 = op_O_2_1; // @[Map2T.scala 17:7]
  assign O_3_0 = op_O_3_0; // @[Map2T.scala 17:7]
  assign O_3_1 = op_O_3_1; // @[Map2T.scala 17:7]
  assign O_4_0 = op_O_4_0; // @[Map2T.scala 17:7]
  assign O_4_1 = op_O_4_1; // @[Map2T.scala 17:7]
  assign O_5_0 = op_O_5_0; // @[Map2T.scala 17:7]
  assign O_5_1 = op_O_5_1; // @[Map2T.scala 17:7]
  assign O_6_0 = op_O_6_0; // @[Map2T.scala 17:7]
  assign O_6_1 = op_O_6_1; // @[Map2T.scala 17:7]
  assign O_7_0 = op_O_7_0; // @[Map2T.scala 17:7]
  assign O_7_1 = op_O_7_1; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0 = I0_0; // @[Map2T.scala 15:11]
  assign op_I0_1 = I0_1; // @[Map2T.scala 15:11]
  assign op_I0_2 = I0_2; // @[Map2T.scala 15:11]
  assign op_I0_3 = I0_3; // @[Map2T.scala 15:11]
  assign op_I0_4 = I0_4; // @[Map2T.scala 15:11]
  assign op_I0_5 = I0_5; // @[Map2T.scala 15:11]
  assign op_I0_6 = I0_6; // @[Map2T.scala 15:11]
  assign op_I0_7 = I0_7; // @[Map2T.scala 15:11]
  assign op_I1_0 = I1_0; // @[Map2T.scala 16:11]
  assign op_I1_1 = I1_1; // @[Map2T.scala 16:11]
  assign op_I1_2 = I1_2; // @[Map2T.scala 16:11]
  assign op_I1_3 = I1_3; // @[Map2T.scala 16:11]
  assign op_I1_4 = I1_4; // @[Map2T.scala 16:11]
  assign op_I1_5 = I1_5; // @[Map2T.scala 16:11]
  assign op_I1_6 = I1_6; // @[Map2T.scala 16:11]
  assign op_I1_7 = I1_7; // @[Map2T.scala 16:11]
endmodule
module SSeqTupleAppender(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0,
  input  [31:0] I0_1,
  input  [31:0] I1,
  output [31:0] O_0,
  output [31:0] O_1,
  output [31:0] O_2
);
  assign valid_down = valid_up; // @[Tuple.scala 28:14]
  assign O_0 = I0_0; // @[Tuple.scala 24:34]
  assign O_1 = I0_1; // @[Tuple.scala 24:34]
  assign O_2 = I1; // @[Tuple.scala 26:32]
endmodule
module Map2S_1(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0_0,
  input  [31:0] I0_0_1,
  input  [31:0] I0_1_0,
  input  [31:0] I0_1_1,
  input  [31:0] I0_2_0,
  input  [31:0] I0_2_1,
  input  [31:0] I0_3_0,
  input  [31:0] I0_3_1,
  input  [31:0] I0_4_0,
  input  [31:0] I0_4_1,
  input  [31:0] I0_5_0,
  input  [31:0] I0_5_1,
  input  [31:0] I0_6_0,
  input  [31:0] I0_6_1,
  input  [31:0] I0_7_0,
  input  [31:0] I0_7_1,
  input  [31:0] I1_0,
  input  [31:0] I1_1,
  input  [31:0] I1_2,
  input  [31:0] I1_3,
  input  [31:0] I1_4,
  input  [31:0] I1_5,
  input  [31:0] I1_6,
  input  [31:0] I1_7,
  output [31:0] O_0_0,
  output [31:0] O_0_1,
  output [31:0] O_0_2,
  output [31:0] O_1_0,
  output [31:0] O_1_1,
  output [31:0] O_1_2,
  output [31:0] O_2_0,
  output [31:0] O_2_1,
  output [31:0] O_2_2,
  output [31:0] O_3_0,
  output [31:0] O_3_1,
  output [31:0] O_3_2,
  output [31:0] O_4_0,
  output [31:0] O_4_1,
  output [31:0] O_4_2,
  output [31:0] O_5_0,
  output [31:0] O_5_1,
  output [31:0] O_5_2,
  output [31:0] O_6_0,
  output [31:0] O_6_1,
  output [31:0] O_6_2,
  output [31:0] O_7_0,
  output [31:0] O_7_1,
  output [31:0] O_7_2
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_2; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_2; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  wire  _T_2; // @[Map2S.scala 26:83]
  wire  _T_3; // @[Map2S.scala 26:83]
  wire  _T_4; // @[Map2S.scala 26:83]
  wire  _T_5; // @[Map2S.scala 26:83]
  SSeqTupleAppender fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I0_1(fst_op_I0_1),
    .I1(fst_op_I1),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1),
    .O_2(fst_op_O_2)
  );
  SSeqTupleAppender other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0(other_ops_0_I0_0),
    .I0_1(other_ops_0_I0_1),
    .I1(other_ops_0_I1),
    .O_0(other_ops_0_O_0),
    .O_1(other_ops_0_O_1),
    .O_2(other_ops_0_O_2)
  );
  SSeqTupleAppender other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0_0(other_ops_1_I0_0),
    .I0_1(other_ops_1_I0_1),
    .I1(other_ops_1_I1),
    .O_0(other_ops_1_O_0),
    .O_1(other_ops_1_O_1),
    .O_2(other_ops_1_O_2)
  );
  SSeqTupleAppender other_ops_2 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0_0(other_ops_2_I0_0),
    .I0_1(other_ops_2_I0_1),
    .I1(other_ops_2_I1),
    .O_0(other_ops_2_O_0),
    .O_1(other_ops_2_O_1),
    .O_2(other_ops_2_O_2)
  );
  SSeqTupleAppender other_ops_3 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I0_0(other_ops_3_I0_0),
    .I0_1(other_ops_3_I0_1),
    .I1(other_ops_3_I1),
    .O_0(other_ops_3_O_0),
    .O_1(other_ops_3_O_1),
    .O_2(other_ops_3_O_2)
  );
  SSeqTupleAppender other_ops_4 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I0_0(other_ops_4_I0_0),
    .I0_1(other_ops_4_I0_1),
    .I1(other_ops_4_I1),
    .O_0(other_ops_4_O_0),
    .O_1(other_ops_4_O_1),
    .O_2(other_ops_4_O_2)
  );
  SSeqTupleAppender other_ops_5 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I0_0(other_ops_5_I0_0),
    .I0_1(other_ops_5_I0_1),
    .I1(other_ops_5_I1),
    .O_0(other_ops_5_O_0),
    .O_1(other_ops_5_O_1),
    .O_2(other_ops_5_O_2)
  );
  SSeqTupleAppender other_ops_6 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I0_0(other_ops_6_I0_0),
    .I0_1(other_ops_6_I0_1),
    .I1(other_ops_6_I1),
    .O_0(other_ops_6_O_0),
    .O_1(other_ops_6_O_1),
    .O_2(other_ops_6_O_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[Map2S.scala 26:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[Map2S.scala 26:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_5 & other_ops_6_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0 = fst_op_O_0; // @[Map2S.scala 19:8]
  assign O_0_1 = fst_op_O_1; // @[Map2S.scala 19:8]
  assign O_0_2 = fst_op_O_2; // @[Map2S.scala 19:8]
  assign O_1_0 = other_ops_0_O_0; // @[Map2S.scala 24:12]
  assign O_1_1 = other_ops_0_O_1; // @[Map2S.scala 24:12]
  assign O_1_2 = other_ops_0_O_2; // @[Map2S.scala 24:12]
  assign O_2_0 = other_ops_1_O_0; // @[Map2S.scala 24:12]
  assign O_2_1 = other_ops_1_O_1; // @[Map2S.scala 24:12]
  assign O_2_2 = other_ops_1_O_2; // @[Map2S.scala 24:12]
  assign O_3_0 = other_ops_2_O_0; // @[Map2S.scala 24:12]
  assign O_3_1 = other_ops_2_O_1; // @[Map2S.scala 24:12]
  assign O_3_2 = other_ops_2_O_2; // @[Map2S.scala 24:12]
  assign O_4_0 = other_ops_3_O_0; // @[Map2S.scala 24:12]
  assign O_4_1 = other_ops_3_O_1; // @[Map2S.scala 24:12]
  assign O_4_2 = other_ops_3_O_2; // @[Map2S.scala 24:12]
  assign O_5_0 = other_ops_4_O_0; // @[Map2S.scala 24:12]
  assign O_5_1 = other_ops_4_O_1; // @[Map2S.scala 24:12]
  assign O_5_2 = other_ops_4_O_2; // @[Map2S.scala 24:12]
  assign O_6_0 = other_ops_5_O_0; // @[Map2S.scala 24:12]
  assign O_6_1 = other_ops_5_O_1; // @[Map2S.scala 24:12]
  assign O_6_2 = other_ops_5_O_2; // @[Map2S.scala 24:12]
  assign O_7_0 = other_ops_6_O_0; // @[Map2S.scala 24:12]
  assign O_7_1 = other_ops_6_O_1; // @[Map2S.scala 24:12]
  assign O_7_2 = other_ops_6_O_2; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1 = I0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0 = I0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1 = I0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I1 = I1_1; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0_0 = I0_2_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1 = I0_2_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I1 = I1_2; // @[Map2S.scala 23:43]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0_0 = I0_3_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_1 = I0_3_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I1 = I1_3; // @[Map2S.scala 23:43]
  assign other_ops_3_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_3_I0_0 = I0_4_0; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_1 = I0_4_1; // @[Map2S.scala 22:43]
  assign other_ops_3_I1 = I1_4; // @[Map2S.scala 23:43]
  assign other_ops_4_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_4_I0_0 = I0_5_0; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_1 = I0_5_1; // @[Map2S.scala 22:43]
  assign other_ops_4_I1 = I1_5; // @[Map2S.scala 23:43]
  assign other_ops_5_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_5_I0_0 = I0_6_0; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_1 = I0_6_1; // @[Map2S.scala 22:43]
  assign other_ops_5_I1 = I1_6; // @[Map2S.scala 23:43]
  assign other_ops_6_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_6_I0_0 = I0_7_0; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_1 = I0_7_1; // @[Map2S.scala 22:43]
  assign other_ops_6_I1 = I1_7; // @[Map2S.scala 23:43]
endmodule
module Map2T_1(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0_0,
  input  [31:0] I0_0_1,
  input  [31:0] I0_1_0,
  input  [31:0] I0_1_1,
  input  [31:0] I0_2_0,
  input  [31:0] I0_2_1,
  input  [31:0] I0_3_0,
  input  [31:0] I0_3_1,
  input  [31:0] I0_4_0,
  input  [31:0] I0_4_1,
  input  [31:0] I0_5_0,
  input  [31:0] I0_5_1,
  input  [31:0] I0_6_0,
  input  [31:0] I0_6_1,
  input  [31:0] I0_7_0,
  input  [31:0] I0_7_1,
  input  [31:0] I1_0,
  input  [31:0] I1_1,
  input  [31:0] I1_2,
  input  [31:0] I1_3,
  input  [31:0] I1_4,
  input  [31:0] I1_5,
  input  [31:0] I1_6,
  input  [31:0] I1_7,
  output [31:0] O_0_0,
  output [31:0] O_0_1,
  output [31:0] O_0_2,
  output [31:0] O_1_0,
  output [31:0] O_1_1,
  output [31:0] O_1_2,
  output [31:0] O_2_0,
  output [31:0] O_2_1,
  output [31:0] O_2_2,
  output [31:0] O_3_0,
  output [31:0] O_3_1,
  output [31:0] O_3_2,
  output [31:0] O_4_0,
  output [31:0] O_4_1,
  output [31:0] O_4_2,
  output [31:0] O_5_0,
  output [31:0] O_5_1,
  output [31:0] O_5_2,
  output [31:0] O_6_0,
  output [31:0] O_6_1,
  output [31:0] O_6_2,
  output [31:0] O_7_0,
  output [31:0] O_7_1,
  output [31:0] O_7_2
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_3; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_4; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_5; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_6; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_7; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_2; // @[Map2T.scala 8:20]
  Map2S_1 op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0_0(op_I0_0_0),
    .I0_0_1(op_I0_0_1),
    .I0_1_0(op_I0_1_0),
    .I0_1_1(op_I0_1_1),
    .I0_2_0(op_I0_2_0),
    .I0_2_1(op_I0_2_1),
    .I0_3_0(op_I0_3_0),
    .I0_3_1(op_I0_3_1),
    .I0_4_0(op_I0_4_0),
    .I0_4_1(op_I0_4_1),
    .I0_5_0(op_I0_5_0),
    .I0_5_1(op_I0_5_1),
    .I0_6_0(op_I0_6_0),
    .I0_6_1(op_I0_6_1),
    .I0_7_0(op_I0_7_0),
    .I0_7_1(op_I0_7_1),
    .I1_0(op_I1_0),
    .I1_1(op_I1_1),
    .I1_2(op_I1_2),
    .I1_3(op_I1_3),
    .I1_4(op_I1_4),
    .I1_5(op_I1_5),
    .I1_6(op_I1_6),
    .I1_7(op_I1_7),
    .O_0_0(op_O_0_0),
    .O_0_1(op_O_0_1),
    .O_0_2(op_O_0_2),
    .O_1_0(op_O_1_0),
    .O_1_1(op_O_1_1),
    .O_1_2(op_O_1_2),
    .O_2_0(op_O_2_0),
    .O_2_1(op_O_2_1),
    .O_2_2(op_O_2_2),
    .O_3_0(op_O_3_0),
    .O_3_1(op_O_3_1),
    .O_3_2(op_O_3_2),
    .O_4_0(op_O_4_0),
    .O_4_1(op_O_4_1),
    .O_4_2(op_O_4_2),
    .O_5_0(op_O_5_0),
    .O_5_1(op_O_5_1),
    .O_5_2(op_O_5_2),
    .O_6_0(op_O_6_0),
    .O_6_1(op_O_6_1),
    .O_6_2(op_O_6_2),
    .O_7_0(op_O_7_0),
    .O_7_1(op_O_7_1),
    .O_7_2(op_O_7_2)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_0 = op_O_0_0; // @[Map2T.scala 17:7]
  assign O_0_1 = op_O_0_1; // @[Map2T.scala 17:7]
  assign O_0_2 = op_O_0_2; // @[Map2T.scala 17:7]
  assign O_1_0 = op_O_1_0; // @[Map2T.scala 17:7]
  assign O_1_1 = op_O_1_1; // @[Map2T.scala 17:7]
  assign O_1_2 = op_O_1_2; // @[Map2T.scala 17:7]
  assign O_2_0 = op_O_2_0; // @[Map2T.scala 17:7]
  assign O_2_1 = op_O_2_1; // @[Map2T.scala 17:7]
  assign O_2_2 = op_O_2_2; // @[Map2T.scala 17:7]
  assign O_3_0 = op_O_3_0; // @[Map2T.scala 17:7]
  assign O_3_1 = op_O_3_1; // @[Map2T.scala 17:7]
  assign O_3_2 = op_O_3_2; // @[Map2T.scala 17:7]
  assign O_4_0 = op_O_4_0; // @[Map2T.scala 17:7]
  assign O_4_1 = op_O_4_1; // @[Map2T.scala 17:7]
  assign O_4_2 = op_O_4_2; // @[Map2T.scala 17:7]
  assign O_5_0 = op_O_5_0; // @[Map2T.scala 17:7]
  assign O_5_1 = op_O_5_1; // @[Map2T.scala 17:7]
  assign O_5_2 = op_O_5_2; // @[Map2T.scala 17:7]
  assign O_6_0 = op_O_6_0; // @[Map2T.scala 17:7]
  assign O_6_1 = op_O_6_1; // @[Map2T.scala 17:7]
  assign O_6_2 = op_O_6_2; // @[Map2T.scala 17:7]
  assign O_7_0 = op_O_7_0; // @[Map2T.scala 17:7]
  assign O_7_1 = op_O_7_1; // @[Map2T.scala 17:7]
  assign O_7_2 = op_O_7_2; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0_0 = I0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_0_1 = I0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_1_0 = I0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_1_1 = I0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_2_0 = I0_2_0; // @[Map2T.scala 15:11]
  assign op_I0_2_1 = I0_2_1; // @[Map2T.scala 15:11]
  assign op_I0_3_0 = I0_3_0; // @[Map2T.scala 15:11]
  assign op_I0_3_1 = I0_3_1; // @[Map2T.scala 15:11]
  assign op_I0_4_0 = I0_4_0; // @[Map2T.scala 15:11]
  assign op_I0_4_1 = I0_4_1; // @[Map2T.scala 15:11]
  assign op_I0_5_0 = I0_5_0; // @[Map2T.scala 15:11]
  assign op_I0_5_1 = I0_5_1; // @[Map2T.scala 15:11]
  assign op_I0_6_0 = I0_6_0; // @[Map2T.scala 15:11]
  assign op_I0_6_1 = I0_6_1; // @[Map2T.scala 15:11]
  assign op_I0_7_0 = I0_7_0; // @[Map2T.scala 15:11]
  assign op_I0_7_1 = I0_7_1; // @[Map2T.scala 15:11]
  assign op_I1_0 = I1_0; // @[Map2T.scala 16:11]
  assign op_I1_1 = I1_1; // @[Map2T.scala 16:11]
  assign op_I1_2 = I1_2; // @[Map2T.scala 16:11]
  assign op_I1_3 = I1_3; // @[Map2T.scala 16:11]
  assign op_I1_4 = I1_4; // @[Map2T.scala 16:11]
  assign op_I1_5 = I1_5; // @[Map2T.scala 16:11]
  assign op_I1_6 = I1_6; // @[Map2T.scala 16:11]
  assign op_I1_7 = I1_7; // @[Map2T.scala 16:11]
endmodule
module PartitionS(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0,
  input  [31:0] I_0_1,
  input  [31:0] I_0_2,
  input  [31:0] I_1_0,
  input  [31:0] I_1_1,
  input  [31:0] I_1_2,
  input  [31:0] I_2_0,
  input  [31:0] I_2_1,
  input  [31:0] I_2_2,
  input  [31:0] I_3_0,
  input  [31:0] I_3_1,
  input  [31:0] I_3_2,
  input  [31:0] I_4_0,
  input  [31:0] I_4_1,
  input  [31:0] I_4_2,
  input  [31:0] I_5_0,
  input  [31:0] I_5_1,
  input  [31:0] I_5_2,
  input  [31:0] I_6_0,
  input  [31:0] I_6_1,
  input  [31:0] I_6_2,
  input  [31:0] I_7_0,
  input  [31:0] I_7_1,
  input  [31:0] I_7_2,
  output [31:0] O_0_0_0,
  output [31:0] O_0_0_1,
  output [31:0] O_0_0_2,
  output [31:0] O_1_0_0,
  output [31:0] O_1_0_1,
  output [31:0] O_1_0_2,
  output [31:0] O_2_0_0,
  output [31:0] O_2_0_1,
  output [31:0] O_2_0_2,
  output [31:0] O_3_0_0,
  output [31:0] O_3_0_1,
  output [31:0] O_3_0_2,
  output [31:0] O_4_0_0,
  output [31:0] O_4_0_1,
  output [31:0] O_4_0_2,
  output [31:0] O_5_0_0,
  output [31:0] O_5_0_1,
  output [31:0] O_5_0_2,
  output [31:0] O_6_0_0,
  output [31:0] O_6_0_1,
  output [31:0] O_6_0_2,
  output [31:0] O_7_0_0,
  output [31:0] O_7_0_1,
  output [31:0] O_7_0_2
);
  assign valid_down = valid_up; // @[Partition.scala 18:14]
  assign O_0_0_0 = I_0_0; // @[Partition.scala 15:39]
  assign O_0_0_1 = I_0_1; // @[Partition.scala 15:39]
  assign O_0_0_2 = I_0_2; // @[Partition.scala 15:39]
  assign O_1_0_0 = I_1_0; // @[Partition.scala 15:39]
  assign O_1_0_1 = I_1_1; // @[Partition.scala 15:39]
  assign O_1_0_2 = I_1_2; // @[Partition.scala 15:39]
  assign O_2_0_0 = I_2_0; // @[Partition.scala 15:39]
  assign O_2_0_1 = I_2_1; // @[Partition.scala 15:39]
  assign O_2_0_2 = I_2_2; // @[Partition.scala 15:39]
  assign O_3_0_0 = I_3_0; // @[Partition.scala 15:39]
  assign O_3_0_1 = I_3_1; // @[Partition.scala 15:39]
  assign O_3_0_2 = I_3_2; // @[Partition.scala 15:39]
  assign O_4_0_0 = I_4_0; // @[Partition.scala 15:39]
  assign O_4_0_1 = I_4_1; // @[Partition.scala 15:39]
  assign O_4_0_2 = I_4_2; // @[Partition.scala 15:39]
  assign O_5_0_0 = I_5_0; // @[Partition.scala 15:39]
  assign O_5_0_1 = I_5_1; // @[Partition.scala 15:39]
  assign O_5_0_2 = I_5_2; // @[Partition.scala 15:39]
  assign O_6_0_0 = I_6_0; // @[Partition.scala 15:39]
  assign O_6_0_1 = I_6_1; // @[Partition.scala 15:39]
  assign O_6_0_2 = I_6_2; // @[Partition.scala 15:39]
  assign O_7_0_0 = I_7_0; // @[Partition.scala 15:39]
  assign O_7_0_1 = I_7_1; // @[Partition.scala 15:39]
  assign O_7_0_2 = I_7_2; // @[Partition.scala 15:39]
endmodule
module MapT(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0,
  input  [31:0] I_0_1,
  input  [31:0] I_0_2,
  input  [31:0] I_1_0,
  input  [31:0] I_1_1,
  input  [31:0] I_1_2,
  input  [31:0] I_2_0,
  input  [31:0] I_2_1,
  input  [31:0] I_2_2,
  input  [31:0] I_3_0,
  input  [31:0] I_3_1,
  input  [31:0] I_3_2,
  input  [31:0] I_4_0,
  input  [31:0] I_4_1,
  input  [31:0] I_4_2,
  input  [31:0] I_5_0,
  input  [31:0] I_5_1,
  input  [31:0] I_5_2,
  input  [31:0] I_6_0,
  input  [31:0] I_6_1,
  input  [31:0] I_6_2,
  input  [31:0] I_7_0,
  input  [31:0] I_7_1,
  input  [31:0] I_7_2,
  output [31:0] O_0_0_0,
  output [31:0] O_0_0_1,
  output [31:0] O_0_0_2,
  output [31:0] O_1_0_0,
  output [31:0] O_1_0_1,
  output [31:0] O_1_0_2,
  output [31:0] O_2_0_0,
  output [31:0] O_2_0_1,
  output [31:0] O_2_0_2,
  output [31:0] O_3_0_0,
  output [31:0] O_3_0_1,
  output [31:0] O_3_0_2,
  output [31:0] O_4_0_0,
  output [31:0] O_4_0_1,
  output [31:0] O_4_0_2,
  output [31:0] O_5_0_0,
  output [31:0] O_5_0_1,
  output [31:0] O_5_0_2,
  output [31:0] O_6_0_0,
  output [31:0] O_6_0_1,
  output [31:0] O_6_0_2,
  output [31:0] O_7_0_0,
  output [31:0] O_7_0_1,
  output [31:0] O_7_0_2
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_0_2; // @[MapT.scala 8:20]
  PartitionS op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0(op_I_0_0),
    .I_0_1(op_I_0_1),
    .I_0_2(op_I_0_2),
    .I_1_0(op_I_1_0),
    .I_1_1(op_I_1_1),
    .I_1_2(op_I_1_2),
    .I_2_0(op_I_2_0),
    .I_2_1(op_I_2_1),
    .I_2_2(op_I_2_2),
    .I_3_0(op_I_3_0),
    .I_3_1(op_I_3_1),
    .I_3_2(op_I_3_2),
    .I_4_0(op_I_4_0),
    .I_4_1(op_I_4_1),
    .I_4_2(op_I_4_2),
    .I_5_0(op_I_5_0),
    .I_5_1(op_I_5_1),
    .I_5_2(op_I_5_2),
    .I_6_0(op_I_6_0),
    .I_6_1(op_I_6_1),
    .I_6_2(op_I_6_2),
    .I_7_0(op_I_7_0),
    .I_7_1(op_I_7_1),
    .I_7_2(op_I_7_2),
    .O_0_0_0(op_O_0_0_0),
    .O_0_0_1(op_O_0_0_1),
    .O_0_0_2(op_O_0_0_2),
    .O_1_0_0(op_O_1_0_0),
    .O_1_0_1(op_O_1_0_1),
    .O_1_0_2(op_O_1_0_2),
    .O_2_0_0(op_O_2_0_0),
    .O_2_0_1(op_O_2_0_1),
    .O_2_0_2(op_O_2_0_2),
    .O_3_0_0(op_O_3_0_0),
    .O_3_0_1(op_O_3_0_1),
    .O_3_0_2(op_O_3_0_2),
    .O_4_0_0(op_O_4_0_0),
    .O_4_0_1(op_O_4_0_1),
    .O_4_0_2(op_O_4_0_2),
    .O_5_0_0(op_O_5_0_0),
    .O_5_0_1(op_O_5_0_1),
    .O_5_0_2(op_O_5_0_2),
    .O_6_0_0(op_O_6_0_0),
    .O_6_0_1(op_O_6_0_1),
    .O_6_0_2(op_O_6_0_2),
    .O_7_0_0(op_O_7_0_0),
    .O_7_0_1(op_O_7_0_1),
    .O_7_0_2(op_O_7_0_2)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0 = op_O_0_0_0; // @[MapT.scala 15:7]
  assign O_0_0_1 = op_O_0_0_1; // @[MapT.scala 15:7]
  assign O_0_0_2 = op_O_0_0_2; // @[MapT.scala 15:7]
  assign O_1_0_0 = op_O_1_0_0; // @[MapT.scala 15:7]
  assign O_1_0_1 = op_O_1_0_1; // @[MapT.scala 15:7]
  assign O_1_0_2 = op_O_1_0_2; // @[MapT.scala 15:7]
  assign O_2_0_0 = op_O_2_0_0; // @[MapT.scala 15:7]
  assign O_2_0_1 = op_O_2_0_1; // @[MapT.scala 15:7]
  assign O_2_0_2 = op_O_2_0_2; // @[MapT.scala 15:7]
  assign O_3_0_0 = op_O_3_0_0; // @[MapT.scala 15:7]
  assign O_3_0_1 = op_O_3_0_1; // @[MapT.scala 15:7]
  assign O_3_0_2 = op_O_3_0_2; // @[MapT.scala 15:7]
  assign O_4_0_0 = op_O_4_0_0; // @[MapT.scala 15:7]
  assign O_4_0_1 = op_O_4_0_1; // @[MapT.scala 15:7]
  assign O_4_0_2 = op_O_4_0_2; // @[MapT.scala 15:7]
  assign O_5_0_0 = op_O_5_0_0; // @[MapT.scala 15:7]
  assign O_5_0_1 = op_O_5_0_1; // @[MapT.scala 15:7]
  assign O_5_0_2 = op_O_5_0_2; // @[MapT.scala 15:7]
  assign O_6_0_0 = op_O_6_0_0; // @[MapT.scala 15:7]
  assign O_6_0_1 = op_O_6_0_1; // @[MapT.scala 15:7]
  assign O_6_0_2 = op_O_6_0_2; // @[MapT.scala 15:7]
  assign O_7_0_0 = op_O_7_0_0; // @[MapT.scala 15:7]
  assign O_7_0_1 = op_O_7_0_1; // @[MapT.scala 15:7]
  assign O_7_0_2 = op_O_7_0_2; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0 = I_0_0; // @[MapT.scala 14:10]
  assign op_I_0_1 = I_0_1; // @[MapT.scala 14:10]
  assign op_I_0_2 = I_0_2; // @[MapT.scala 14:10]
  assign op_I_1_0 = I_1_0; // @[MapT.scala 14:10]
  assign op_I_1_1 = I_1_1; // @[MapT.scala 14:10]
  assign op_I_1_2 = I_1_2; // @[MapT.scala 14:10]
  assign op_I_2_0 = I_2_0; // @[MapT.scala 14:10]
  assign op_I_2_1 = I_2_1; // @[MapT.scala 14:10]
  assign op_I_2_2 = I_2_2; // @[MapT.scala 14:10]
  assign op_I_3_0 = I_3_0; // @[MapT.scala 14:10]
  assign op_I_3_1 = I_3_1; // @[MapT.scala 14:10]
  assign op_I_3_2 = I_3_2; // @[MapT.scala 14:10]
  assign op_I_4_0 = I_4_0; // @[MapT.scala 14:10]
  assign op_I_4_1 = I_4_1; // @[MapT.scala 14:10]
  assign op_I_4_2 = I_4_2; // @[MapT.scala 14:10]
  assign op_I_5_0 = I_5_0; // @[MapT.scala 14:10]
  assign op_I_5_1 = I_5_1; // @[MapT.scala 14:10]
  assign op_I_5_2 = I_5_2; // @[MapT.scala 14:10]
  assign op_I_6_0 = I_6_0; // @[MapT.scala 14:10]
  assign op_I_6_1 = I_6_1; // @[MapT.scala 14:10]
  assign op_I_6_2 = I_6_2; // @[MapT.scala 14:10]
  assign op_I_7_0 = I_7_0; // @[MapT.scala 14:10]
  assign op_I_7_1 = I_7_1; // @[MapT.scala 14:10]
  assign op_I_7_2 = I_7_2; // @[MapT.scala 14:10]
endmodule
module SSeqTupleToSSeq(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0,
  input  [31:0] I_1,
  input  [31:0] I_2,
  output [31:0] O_0,
  output [31:0] O_1,
  output [31:0] O_2
);
  assign valid_down = valid_up; // @[Tuple.scala 42:14]
  assign O_0 = I_0; // @[Tuple.scala 41:5]
  assign O_1 = I_1; // @[Tuple.scala 41:5]
  assign O_2 = I_2; // @[Tuple.scala 41:5]
endmodule
module Remove1S(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0,
  input  [31:0] I_0_1,
  input  [31:0] I_0_2,
  output [31:0] O_0,
  output [31:0] O_1,
  output [31:0] O_2
);
  wire  op_inst_valid_up; // @[Remove1S.scala 9:23]
  wire  op_inst_valid_down; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_I_0; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_I_1; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_I_2; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_O_0; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_O_1; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_O_2; // @[Remove1S.scala 9:23]
  SSeqTupleToSSeq op_inst ( // @[Remove1S.scala 9:23]
    .valid_up(op_inst_valid_up),
    .valid_down(op_inst_valid_down),
    .I_0(op_inst_I_0),
    .I_1(op_inst_I_1),
    .I_2(op_inst_I_2),
    .O_0(op_inst_O_0),
    .O_1(op_inst_O_1),
    .O_2(op_inst_O_2)
  );
  assign valid_down = op_inst_valid_down; // @[Remove1S.scala 16:14]
  assign O_0 = op_inst_O_0; // @[Remove1S.scala 14:5]
  assign O_1 = op_inst_O_1; // @[Remove1S.scala 14:5]
  assign O_2 = op_inst_O_2; // @[Remove1S.scala 14:5]
  assign op_inst_valid_up = valid_up; // @[Remove1S.scala 15:20]
  assign op_inst_I_0 = I_0_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_1 = I_0_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_2 = I_0_2; // @[Remove1S.scala 13:13]
endmodule
module MapS(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0_0,
  input  [31:0] I_0_0_1,
  input  [31:0] I_0_0_2,
  input  [31:0] I_1_0_0,
  input  [31:0] I_1_0_1,
  input  [31:0] I_1_0_2,
  input  [31:0] I_2_0_0,
  input  [31:0] I_2_0_1,
  input  [31:0] I_2_0_2,
  input  [31:0] I_3_0_0,
  input  [31:0] I_3_0_1,
  input  [31:0] I_3_0_2,
  input  [31:0] I_4_0_0,
  input  [31:0] I_4_0_1,
  input  [31:0] I_4_0_2,
  input  [31:0] I_5_0_0,
  input  [31:0] I_5_0_1,
  input  [31:0] I_5_0_2,
  input  [31:0] I_6_0_0,
  input  [31:0] I_6_0_1,
  input  [31:0] I_6_0_2,
  input  [31:0] I_7_0_0,
  input  [31:0] I_7_0_1,
  input  [31:0] I_7_0_2,
  output [31:0] O_0_0,
  output [31:0] O_0_1,
  output [31:0] O_0_2,
  output [31:0] O_1_0,
  output [31:0] O_1_1,
  output [31:0] O_1_2,
  output [31:0] O_2_0,
  output [31:0] O_2_1,
  output [31:0] O_2_2,
  output [31:0] O_3_0,
  output [31:0] O_3_1,
  output [31:0] O_3_2,
  output [31:0] O_4_0,
  output [31:0] O_4_1,
  output [31:0] O_4_2,
  output [31:0] O_5_0,
  output [31:0] O_5_1,
  output [31:0] O_5_2,
  output [31:0] O_6_0,
  output [31:0] O_6_1,
  output [31:0] O_6_2,
  output [31:0] O_7_0,
  output [31:0] O_7_1,
  output [31:0] O_7_2
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_0; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_1; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_2; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_0; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_1; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_2; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_O_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_O_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_O_2; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_O_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_O_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_O_2; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_O_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_O_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_O_2; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_O_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_O_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_O_2; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_O_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_O_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_O_2; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_O_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_O_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_O_2; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_O_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_O_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_O_2; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  wire  _T_1; // @[MapS.scala 23:83]
  wire  _T_2; // @[MapS.scala 23:83]
  wire  _T_3; // @[MapS.scala 23:83]
  wire  _T_4; // @[MapS.scala 23:83]
  wire  _T_5; // @[MapS.scala 23:83]
  Remove1S fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_0(fst_op_I_0_0),
    .I_0_1(fst_op_I_0_1),
    .I_0_2(fst_op_I_0_2),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1),
    .O_2(fst_op_O_2)
  );
  Remove1S other_ops_0 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_0(other_ops_0_I_0_0),
    .I_0_1(other_ops_0_I_0_1),
    .I_0_2(other_ops_0_I_0_2),
    .O_0(other_ops_0_O_0),
    .O_1(other_ops_0_O_1),
    .O_2(other_ops_0_O_2)
  );
  Remove1S other_ops_1 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0_0(other_ops_1_I_0_0),
    .I_0_1(other_ops_1_I_0_1),
    .I_0_2(other_ops_1_I_0_2),
    .O_0(other_ops_1_O_0),
    .O_1(other_ops_1_O_1),
    .O_2(other_ops_1_O_2)
  );
  Remove1S other_ops_2 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I_0_0(other_ops_2_I_0_0),
    .I_0_1(other_ops_2_I_0_1),
    .I_0_2(other_ops_2_I_0_2),
    .O_0(other_ops_2_O_0),
    .O_1(other_ops_2_O_1),
    .O_2(other_ops_2_O_2)
  );
  Remove1S other_ops_3 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I_0_0(other_ops_3_I_0_0),
    .I_0_1(other_ops_3_I_0_1),
    .I_0_2(other_ops_3_I_0_2),
    .O_0(other_ops_3_O_0),
    .O_1(other_ops_3_O_1),
    .O_2(other_ops_3_O_2)
  );
  Remove1S other_ops_4 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I_0_0(other_ops_4_I_0_0),
    .I_0_1(other_ops_4_I_0_1),
    .I_0_2(other_ops_4_I_0_2),
    .O_0(other_ops_4_O_0),
    .O_1(other_ops_4_O_1),
    .O_2(other_ops_4_O_2)
  );
  Remove1S other_ops_5 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I_0_0(other_ops_5_I_0_0),
    .I_0_1(other_ops_5_I_0_1),
    .I_0_2(other_ops_5_I_0_2),
    .O_0(other_ops_5_O_0),
    .O_1(other_ops_5_O_1),
    .O_2(other_ops_5_O_2)
  );
  Remove1S other_ops_6 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I_0_0(other_ops_6_I_0_0),
    .I_0_1(other_ops_6_I_0_1),
    .I_0_2(other_ops_6_I_0_2),
    .O_0(other_ops_6_O_0),
    .O_1(other_ops_6_O_1),
    .O_2(other_ops_6_O_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[MapS.scala 23:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[MapS.scala 23:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[MapS.scala 23:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[MapS.scala 23:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T_5 & other_ops_6_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign O_0_1 = fst_op_O_1; // @[MapS.scala 17:8]
  assign O_0_2 = fst_op_O_2; // @[MapS.scala 17:8]
  assign O_1_0 = other_ops_0_O_0; // @[MapS.scala 21:12]
  assign O_1_1 = other_ops_0_O_1; // @[MapS.scala 21:12]
  assign O_1_2 = other_ops_0_O_2; // @[MapS.scala 21:12]
  assign O_2_0 = other_ops_1_O_0; // @[MapS.scala 21:12]
  assign O_2_1 = other_ops_1_O_1; // @[MapS.scala 21:12]
  assign O_2_2 = other_ops_1_O_2; // @[MapS.scala 21:12]
  assign O_3_0 = other_ops_2_O_0; // @[MapS.scala 21:12]
  assign O_3_1 = other_ops_2_O_1; // @[MapS.scala 21:12]
  assign O_3_2 = other_ops_2_O_2; // @[MapS.scala 21:12]
  assign O_4_0 = other_ops_3_O_0; // @[MapS.scala 21:12]
  assign O_4_1 = other_ops_3_O_1; // @[MapS.scala 21:12]
  assign O_4_2 = other_ops_3_O_2; // @[MapS.scala 21:12]
  assign O_5_0 = other_ops_4_O_0; // @[MapS.scala 21:12]
  assign O_5_1 = other_ops_4_O_1; // @[MapS.scala 21:12]
  assign O_5_2 = other_ops_4_O_2; // @[MapS.scala 21:12]
  assign O_6_0 = other_ops_5_O_0; // @[MapS.scala 21:12]
  assign O_6_1 = other_ops_5_O_1; // @[MapS.scala 21:12]
  assign O_6_2 = other_ops_5_O_2; // @[MapS.scala 21:12]
  assign O_7_0 = other_ops_6_O_0; // @[MapS.scala 21:12]
  assign O_7_1 = other_ops_6_O_1; // @[MapS.scala 21:12]
  assign O_7_2 = other_ops_6_O_2; // @[MapS.scala 21:12]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_0 = I_0_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_1 = I_0_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_2 = I_0_0_2; // @[MapS.scala 16:12]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_0 = I_1_0_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1 = I_1_0_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2 = I_1_0_2; // @[MapS.scala 20:41]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0_0 = I_2_0_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1 = I_2_0_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2 = I_2_0_2; // @[MapS.scala 20:41]
  assign other_ops_2_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_2_I_0_0 = I_3_0_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1 = I_3_0_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2 = I_3_0_2; // @[MapS.scala 20:41]
  assign other_ops_3_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_3_I_0_0 = I_4_0_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_1 = I_4_0_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_2 = I_4_0_2; // @[MapS.scala 20:41]
  assign other_ops_4_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_4_I_0_0 = I_5_0_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_1 = I_5_0_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_2 = I_5_0_2; // @[MapS.scala 20:41]
  assign other_ops_5_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_5_I_0_0 = I_6_0_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_1 = I_6_0_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_2 = I_6_0_2; // @[MapS.scala 20:41]
  assign other_ops_6_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_6_I_0_0 = I_7_0_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_1 = I_7_0_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_2 = I_7_0_2; // @[MapS.scala 20:41]
endmodule
module MapT_1(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0_0,
  input  [31:0] I_0_0_1,
  input  [31:0] I_0_0_2,
  input  [31:0] I_1_0_0,
  input  [31:0] I_1_0_1,
  input  [31:0] I_1_0_2,
  input  [31:0] I_2_0_0,
  input  [31:0] I_2_0_1,
  input  [31:0] I_2_0_2,
  input  [31:0] I_3_0_0,
  input  [31:0] I_3_0_1,
  input  [31:0] I_3_0_2,
  input  [31:0] I_4_0_0,
  input  [31:0] I_4_0_1,
  input  [31:0] I_4_0_2,
  input  [31:0] I_5_0_0,
  input  [31:0] I_5_0_1,
  input  [31:0] I_5_0_2,
  input  [31:0] I_6_0_0,
  input  [31:0] I_6_0_1,
  input  [31:0] I_6_0_2,
  input  [31:0] I_7_0_0,
  input  [31:0] I_7_0_1,
  input  [31:0] I_7_0_2,
  output [31:0] O_0_0,
  output [31:0] O_0_1,
  output [31:0] O_0_2,
  output [31:0] O_1_0,
  output [31:0] O_1_1,
  output [31:0] O_1_2,
  output [31:0] O_2_0,
  output [31:0] O_2_1,
  output [31:0] O_2_2,
  output [31:0] O_3_0,
  output [31:0] O_3_1,
  output [31:0] O_3_2,
  output [31:0] O_4_0,
  output [31:0] O_4_1,
  output [31:0] O_4_2,
  output [31:0] O_5_0,
  output [31:0] O_5_1,
  output [31:0] O_5_2,
  output [31:0] O_6_0,
  output [31:0] O_6_1,
  output [31:0] O_6_2,
  output [31:0] O_7_0,
  output [31:0] O_7_1,
  output [31:0] O_7_2
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_2; // @[MapT.scala 8:20]
  MapS op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0(op_I_0_0_0),
    .I_0_0_1(op_I_0_0_1),
    .I_0_0_2(op_I_0_0_2),
    .I_1_0_0(op_I_1_0_0),
    .I_1_0_1(op_I_1_0_1),
    .I_1_0_2(op_I_1_0_2),
    .I_2_0_0(op_I_2_0_0),
    .I_2_0_1(op_I_2_0_1),
    .I_2_0_2(op_I_2_0_2),
    .I_3_0_0(op_I_3_0_0),
    .I_3_0_1(op_I_3_0_1),
    .I_3_0_2(op_I_3_0_2),
    .I_4_0_0(op_I_4_0_0),
    .I_4_0_1(op_I_4_0_1),
    .I_4_0_2(op_I_4_0_2),
    .I_5_0_0(op_I_5_0_0),
    .I_5_0_1(op_I_5_0_1),
    .I_5_0_2(op_I_5_0_2),
    .I_6_0_0(op_I_6_0_0),
    .I_6_0_1(op_I_6_0_1),
    .I_6_0_2(op_I_6_0_2),
    .I_7_0_0(op_I_7_0_0),
    .I_7_0_1(op_I_7_0_1),
    .I_7_0_2(op_I_7_0_2),
    .O_0_0(op_O_0_0),
    .O_0_1(op_O_0_1),
    .O_0_2(op_O_0_2),
    .O_1_0(op_O_1_0),
    .O_1_1(op_O_1_1),
    .O_1_2(op_O_1_2),
    .O_2_0(op_O_2_0),
    .O_2_1(op_O_2_1),
    .O_2_2(op_O_2_2),
    .O_3_0(op_O_3_0),
    .O_3_1(op_O_3_1),
    .O_3_2(op_O_3_2),
    .O_4_0(op_O_4_0),
    .O_4_1(op_O_4_1),
    .O_4_2(op_O_4_2),
    .O_5_0(op_O_5_0),
    .O_5_1(op_O_5_1),
    .O_5_2(op_O_5_2),
    .O_6_0(op_O_6_0),
    .O_6_1(op_O_6_1),
    .O_6_2(op_O_6_2),
    .O_7_0(op_O_7_0),
    .O_7_1(op_O_7_1),
    .O_7_2(op_O_7_2)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0 = op_O_0_0; // @[MapT.scala 15:7]
  assign O_0_1 = op_O_0_1; // @[MapT.scala 15:7]
  assign O_0_2 = op_O_0_2; // @[MapT.scala 15:7]
  assign O_1_0 = op_O_1_0; // @[MapT.scala 15:7]
  assign O_1_1 = op_O_1_1; // @[MapT.scala 15:7]
  assign O_1_2 = op_O_1_2; // @[MapT.scala 15:7]
  assign O_2_0 = op_O_2_0; // @[MapT.scala 15:7]
  assign O_2_1 = op_O_2_1; // @[MapT.scala 15:7]
  assign O_2_2 = op_O_2_2; // @[MapT.scala 15:7]
  assign O_3_0 = op_O_3_0; // @[MapT.scala 15:7]
  assign O_3_1 = op_O_3_1; // @[MapT.scala 15:7]
  assign O_3_2 = op_O_3_2; // @[MapT.scala 15:7]
  assign O_4_0 = op_O_4_0; // @[MapT.scala 15:7]
  assign O_4_1 = op_O_4_1; // @[MapT.scala 15:7]
  assign O_4_2 = op_O_4_2; // @[MapT.scala 15:7]
  assign O_5_0 = op_O_5_0; // @[MapT.scala 15:7]
  assign O_5_1 = op_O_5_1; // @[MapT.scala 15:7]
  assign O_5_2 = op_O_5_2; // @[MapT.scala 15:7]
  assign O_6_0 = op_O_6_0; // @[MapT.scala 15:7]
  assign O_6_1 = op_O_6_1; // @[MapT.scala 15:7]
  assign O_6_2 = op_O_6_2; // @[MapT.scala 15:7]
  assign O_7_0 = op_O_7_0; // @[MapT.scala 15:7]
  assign O_7_1 = op_O_7_1; // @[MapT.scala 15:7]
  assign O_7_2 = op_O_7_2; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0 = I_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_1 = I_0_0_1; // @[MapT.scala 14:10]
  assign op_I_0_0_2 = I_0_0_2; // @[MapT.scala 14:10]
  assign op_I_1_0_0 = I_1_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_1 = I_1_0_1; // @[MapT.scala 14:10]
  assign op_I_1_0_2 = I_1_0_2; // @[MapT.scala 14:10]
  assign op_I_2_0_0 = I_2_0_0; // @[MapT.scala 14:10]
  assign op_I_2_0_1 = I_2_0_1; // @[MapT.scala 14:10]
  assign op_I_2_0_2 = I_2_0_2; // @[MapT.scala 14:10]
  assign op_I_3_0_0 = I_3_0_0; // @[MapT.scala 14:10]
  assign op_I_3_0_1 = I_3_0_1; // @[MapT.scala 14:10]
  assign op_I_3_0_2 = I_3_0_2; // @[MapT.scala 14:10]
  assign op_I_4_0_0 = I_4_0_0; // @[MapT.scala 14:10]
  assign op_I_4_0_1 = I_4_0_1; // @[MapT.scala 14:10]
  assign op_I_4_0_2 = I_4_0_2; // @[MapT.scala 14:10]
  assign op_I_5_0_0 = I_5_0_0; // @[MapT.scala 14:10]
  assign op_I_5_0_1 = I_5_0_1; // @[MapT.scala 14:10]
  assign op_I_5_0_2 = I_5_0_2; // @[MapT.scala 14:10]
  assign op_I_6_0_0 = I_6_0_0; // @[MapT.scala 14:10]
  assign op_I_6_0_1 = I_6_0_1; // @[MapT.scala 14:10]
  assign op_I_6_0_2 = I_6_0_2; // @[MapT.scala 14:10]
  assign op_I_7_0_0 = I_7_0_0; // @[MapT.scala 14:10]
  assign op_I_7_0_1 = I_7_0_1; // @[MapT.scala 14:10]
  assign op_I_7_0_2 = I_7_0_2; // @[MapT.scala 14:10]
endmodule
module SSeqTupleCreator_2(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0,
  input  [31:0] I0_1,
  input  [31:0] I0_2,
  input  [31:0] I1_0,
  input  [31:0] I1_1,
  input  [31:0] I1_2,
  output [31:0] O_0_0,
  output [31:0] O_0_1,
  output [31:0] O_0_2,
  output [31:0] O_1_0,
  output [31:0] O_1_1,
  output [31:0] O_1_2
);
  assign valid_down = valid_up; // @[Tuple.scala 15:14]
  assign O_0_0 = I0_0; // @[Tuple.scala 12:32]
  assign O_0_1 = I0_1; // @[Tuple.scala 12:32]
  assign O_0_2 = I0_2; // @[Tuple.scala 12:32]
  assign O_1_0 = I1_0; // @[Tuple.scala 13:32]
  assign O_1_1 = I1_1; // @[Tuple.scala 13:32]
  assign O_1_2 = I1_2; // @[Tuple.scala 13:32]
endmodule
module Map2S_4(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0_0,
  input  [31:0] I0_0_1,
  input  [31:0] I0_0_2,
  input  [31:0] I0_1_0,
  input  [31:0] I0_1_1,
  input  [31:0] I0_1_2,
  input  [31:0] I0_2_0,
  input  [31:0] I0_2_1,
  input  [31:0] I0_2_2,
  input  [31:0] I0_3_0,
  input  [31:0] I0_3_1,
  input  [31:0] I0_3_2,
  input  [31:0] I0_4_0,
  input  [31:0] I0_4_1,
  input  [31:0] I0_4_2,
  input  [31:0] I0_5_0,
  input  [31:0] I0_5_1,
  input  [31:0] I0_5_2,
  input  [31:0] I0_6_0,
  input  [31:0] I0_6_1,
  input  [31:0] I0_6_2,
  input  [31:0] I0_7_0,
  input  [31:0] I0_7_1,
  input  [31:0] I0_7_2,
  input  [31:0] I1_0_0,
  input  [31:0] I1_0_1,
  input  [31:0] I1_0_2,
  input  [31:0] I1_1_0,
  input  [31:0] I1_1_1,
  input  [31:0] I1_1_2,
  input  [31:0] I1_2_0,
  input  [31:0] I1_2_1,
  input  [31:0] I1_2_2,
  input  [31:0] I1_3_0,
  input  [31:0] I1_3_1,
  input  [31:0] I1_3_2,
  input  [31:0] I1_4_0,
  input  [31:0] I1_4_1,
  input  [31:0] I1_4_2,
  input  [31:0] I1_5_0,
  input  [31:0] I1_5_1,
  input  [31:0] I1_5_2,
  input  [31:0] I1_6_0,
  input  [31:0] I1_6_1,
  input  [31:0] I1_6_2,
  input  [31:0] I1_7_0,
  input  [31:0] I1_7_1,
  input  [31:0] I1_7_2,
  output [31:0] O_0_0_0,
  output [31:0] O_0_0_1,
  output [31:0] O_0_0_2,
  output [31:0] O_0_1_0,
  output [31:0] O_0_1_1,
  output [31:0] O_0_1_2,
  output [31:0] O_1_0_0,
  output [31:0] O_1_0_1,
  output [31:0] O_1_0_2,
  output [31:0] O_1_1_0,
  output [31:0] O_1_1_1,
  output [31:0] O_1_1_2,
  output [31:0] O_2_0_0,
  output [31:0] O_2_0_1,
  output [31:0] O_2_0_2,
  output [31:0] O_2_1_0,
  output [31:0] O_2_1_1,
  output [31:0] O_2_1_2,
  output [31:0] O_3_0_0,
  output [31:0] O_3_0_1,
  output [31:0] O_3_0_2,
  output [31:0] O_3_1_0,
  output [31:0] O_3_1_1,
  output [31:0] O_3_1_2,
  output [31:0] O_4_0_0,
  output [31:0] O_4_0_1,
  output [31:0] O_4_0_2,
  output [31:0] O_4_1_0,
  output [31:0] O_4_1_1,
  output [31:0] O_4_1_2,
  output [31:0] O_5_0_0,
  output [31:0] O_5_0_1,
  output [31:0] O_5_0_2,
  output [31:0] O_5_1_0,
  output [31:0] O_5_1_1,
  output [31:0] O_5_1_2,
  output [31:0] O_6_0_0,
  output [31:0] O_6_0_1,
  output [31:0] O_6_0_2,
  output [31:0] O_6_1_0,
  output [31:0] O_6_1_1,
  output [31:0] O_6_1_2,
  output [31:0] O_7_0_0,
  output [31:0] O_7_0_1,
  output [31:0] O_7_0_2,
  output [31:0] O_7_1_0,
  output [31:0] O_7_1_1,
  output [31:0] O_7_1_2
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_2; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_2; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_2; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_1_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_1_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_1_2; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_1_2; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  wire  _T_2; // @[Map2S.scala 26:83]
  wire  _T_3; // @[Map2S.scala 26:83]
  wire  _T_4; // @[Map2S.scala 26:83]
  wire  _T_5; // @[Map2S.scala 26:83]
  SSeqTupleCreator_2 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I0_1(fst_op_I0_1),
    .I0_2(fst_op_I0_2),
    .I1_0(fst_op_I1_0),
    .I1_1(fst_op_I1_1),
    .I1_2(fst_op_I1_2),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1),
    .O_0_2(fst_op_O_0_2),
    .O_1_0(fst_op_O_1_0),
    .O_1_1(fst_op_O_1_1),
    .O_1_2(fst_op_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0(other_ops_0_I0_0),
    .I0_1(other_ops_0_I0_1),
    .I0_2(other_ops_0_I0_2),
    .I1_0(other_ops_0_I1_0),
    .I1_1(other_ops_0_I1_1),
    .I1_2(other_ops_0_I1_2),
    .O_0_0(other_ops_0_O_0_0),
    .O_0_1(other_ops_0_O_0_1),
    .O_0_2(other_ops_0_O_0_2),
    .O_1_0(other_ops_0_O_1_0),
    .O_1_1(other_ops_0_O_1_1),
    .O_1_2(other_ops_0_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0_0(other_ops_1_I0_0),
    .I0_1(other_ops_1_I0_1),
    .I0_2(other_ops_1_I0_2),
    .I1_0(other_ops_1_I1_0),
    .I1_1(other_ops_1_I1_1),
    .I1_2(other_ops_1_I1_2),
    .O_0_0(other_ops_1_O_0_0),
    .O_0_1(other_ops_1_O_0_1),
    .O_0_2(other_ops_1_O_0_2),
    .O_1_0(other_ops_1_O_1_0),
    .O_1_1(other_ops_1_O_1_1),
    .O_1_2(other_ops_1_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_2 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0_0(other_ops_2_I0_0),
    .I0_1(other_ops_2_I0_1),
    .I0_2(other_ops_2_I0_2),
    .I1_0(other_ops_2_I1_0),
    .I1_1(other_ops_2_I1_1),
    .I1_2(other_ops_2_I1_2),
    .O_0_0(other_ops_2_O_0_0),
    .O_0_1(other_ops_2_O_0_1),
    .O_0_2(other_ops_2_O_0_2),
    .O_1_0(other_ops_2_O_1_0),
    .O_1_1(other_ops_2_O_1_1),
    .O_1_2(other_ops_2_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_3 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I0_0(other_ops_3_I0_0),
    .I0_1(other_ops_3_I0_1),
    .I0_2(other_ops_3_I0_2),
    .I1_0(other_ops_3_I1_0),
    .I1_1(other_ops_3_I1_1),
    .I1_2(other_ops_3_I1_2),
    .O_0_0(other_ops_3_O_0_0),
    .O_0_1(other_ops_3_O_0_1),
    .O_0_2(other_ops_3_O_0_2),
    .O_1_0(other_ops_3_O_1_0),
    .O_1_1(other_ops_3_O_1_1),
    .O_1_2(other_ops_3_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_4 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I0_0(other_ops_4_I0_0),
    .I0_1(other_ops_4_I0_1),
    .I0_2(other_ops_4_I0_2),
    .I1_0(other_ops_4_I1_0),
    .I1_1(other_ops_4_I1_1),
    .I1_2(other_ops_4_I1_2),
    .O_0_0(other_ops_4_O_0_0),
    .O_0_1(other_ops_4_O_0_1),
    .O_0_2(other_ops_4_O_0_2),
    .O_1_0(other_ops_4_O_1_0),
    .O_1_1(other_ops_4_O_1_1),
    .O_1_2(other_ops_4_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_5 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I0_0(other_ops_5_I0_0),
    .I0_1(other_ops_5_I0_1),
    .I0_2(other_ops_5_I0_2),
    .I1_0(other_ops_5_I1_0),
    .I1_1(other_ops_5_I1_1),
    .I1_2(other_ops_5_I1_2),
    .O_0_0(other_ops_5_O_0_0),
    .O_0_1(other_ops_5_O_0_1),
    .O_0_2(other_ops_5_O_0_2),
    .O_1_0(other_ops_5_O_1_0),
    .O_1_1(other_ops_5_O_1_1),
    .O_1_2(other_ops_5_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_6 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I0_0(other_ops_6_I0_0),
    .I0_1(other_ops_6_I0_1),
    .I0_2(other_ops_6_I0_2),
    .I1_0(other_ops_6_I1_0),
    .I1_1(other_ops_6_I1_1),
    .I1_2(other_ops_6_I1_2),
    .O_0_0(other_ops_6_O_0_0),
    .O_0_1(other_ops_6_O_0_1),
    .O_0_2(other_ops_6_O_0_2),
    .O_1_0(other_ops_6_O_1_0),
    .O_1_1(other_ops_6_O_1_1),
    .O_1_2(other_ops_6_O_1_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[Map2S.scala 26:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[Map2S.scala 26:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_5 & other_ops_6_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[Map2S.scala 19:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[Map2S.scala 19:8]
  assign O_0_0_2 = fst_op_O_0_2; // @[Map2S.scala 19:8]
  assign O_0_1_0 = fst_op_O_1_0; // @[Map2S.scala 19:8]
  assign O_0_1_1 = fst_op_O_1_1; // @[Map2S.scala 19:8]
  assign O_0_1_2 = fst_op_O_1_2; // @[Map2S.scala 19:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[Map2S.scala 24:12]
  assign O_1_0_1 = other_ops_0_O_0_1; // @[Map2S.scala 24:12]
  assign O_1_0_2 = other_ops_0_O_0_2; // @[Map2S.scala 24:12]
  assign O_1_1_0 = other_ops_0_O_1_0; // @[Map2S.scala 24:12]
  assign O_1_1_1 = other_ops_0_O_1_1; // @[Map2S.scala 24:12]
  assign O_1_1_2 = other_ops_0_O_1_2; // @[Map2S.scala 24:12]
  assign O_2_0_0 = other_ops_1_O_0_0; // @[Map2S.scala 24:12]
  assign O_2_0_1 = other_ops_1_O_0_1; // @[Map2S.scala 24:12]
  assign O_2_0_2 = other_ops_1_O_0_2; // @[Map2S.scala 24:12]
  assign O_2_1_0 = other_ops_1_O_1_0; // @[Map2S.scala 24:12]
  assign O_2_1_1 = other_ops_1_O_1_1; // @[Map2S.scala 24:12]
  assign O_2_1_2 = other_ops_1_O_1_2; // @[Map2S.scala 24:12]
  assign O_3_0_0 = other_ops_2_O_0_0; // @[Map2S.scala 24:12]
  assign O_3_0_1 = other_ops_2_O_0_1; // @[Map2S.scala 24:12]
  assign O_3_0_2 = other_ops_2_O_0_2; // @[Map2S.scala 24:12]
  assign O_3_1_0 = other_ops_2_O_1_0; // @[Map2S.scala 24:12]
  assign O_3_1_1 = other_ops_2_O_1_1; // @[Map2S.scala 24:12]
  assign O_3_1_2 = other_ops_2_O_1_2; // @[Map2S.scala 24:12]
  assign O_4_0_0 = other_ops_3_O_0_0; // @[Map2S.scala 24:12]
  assign O_4_0_1 = other_ops_3_O_0_1; // @[Map2S.scala 24:12]
  assign O_4_0_2 = other_ops_3_O_0_2; // @[Map2S.scala 24:12]
  assign O_4_1_0 = other_ops_3_O_1_0; // @[Map2S.scala 24:12]
  assign O_4_1_1 = other_ops_3_O_1_1; // @[Map2S.scala 24:12]
  assign O_4_1_2 = other_ops_3_O_1_2; // @[Map2S.scala 24:12]
  assign O_5_0_0 = other_ops_4_O_0_0; // @[Map2S.scala 24:12]
  assign O_5_0_1 = other_ops_4_O_0_1; // @[Map2S.scala 24:12]
  assign O_5_0_2 = other_ops_4_O_0_2; // @[Map2S.scala 24:12]
  assign O_5_1_0 = other_ops_4_O_1_0; // @[Map2S.scala 24:12]
  assign O_5_1_1 = other_ops_4_O_1_1; // @[Map2S.scala 24:12]
  assign O_5_1_2 = other_ops_4_O_1_2; // @[Map2S.scala 24:12]
  assign O_6_0_0 = other_ops_5_O_0_0; // @[Map2S.scala 24:12]
  assign O_6_0_1 = other_ops_5_O_0_1; // @[Map2S.scala 24:12]
  assign O_6_0_2 = other_ops_5_O_0_2; // @[Map2S.scala 24:12]
  assign O_6_1_0 = other_ops_5_O_1_0; // @[Map2S.scala 24:12]
  assign O_6_1_1 = other_ops_5_O_1_1; // @[Map2S.scala 24:12]
  assign O_6_1_2 = other_ops_5_O_1_2; // @[Map2S.scala 24:12]
  assign O_7_0_0 = other_ops_6_O_0_0; // @[Map2S.scala 24:12]
  assign O_7_0_1 = other_ops_6_O_0_1; // @[Map2S.scala 24:12]
  assign O_7_0_2 = other_ops_6_O_0_2; // @[Map2S.scala 24:12]
  assign O_7_1_0 = other_ops_6_O_1_0; // @[Map2S.scala 24:12]
  assign O_7_1_1 = other_ops_6_O_1_1; // @[Map2S.scala 24:12]
  assign O_7_1_2 = other_ops_6_O_1_2; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1 = I0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_2 = I0_0_2; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = I1_0_0; // @[Map2S.scala 18:13]
  assign fst_op_I1_1 = I1_0_1; // @[Map2S.scala 18:13]
  assign fst_op_I1_2 = I1_0_2; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0 = I0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1 = I0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_2 = I0_1_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I1_0 = I1_1_0; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_1 = I1_1_1; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_2 = I1_1_2; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0_0 = I0_2_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1 = I0_2_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_2 = I0_2_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1_0 = I1_2_0; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_1 = I1_2_1; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_2 = I1_2_2; // @[Map2S.scala 23:43]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0_0 = I0_3_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_1 = I0_3_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_2 = I0_3_2; // @[Map2S.scala 22:43]
  assign other_ops_2_I1_0 = I1_3_0; // @[Map2S.scala 23:43]
  assign other_ops_2_I1_1 = I1_3_1; // @[Map2S.scala 23:43]
  assign other_ops_2_I1_2 = I1_3_2; // @[Map2S.scala 23:43]
  assign other_ops_3_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_3_I0_0 = I0_4_0; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_1 = I0_4_1; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_2 = I0_4_2; // @[Map2S.scala 22:43]
  assign other_ops_3_I1_0 = I1_4_0; // @[Map2S.scala 23:43]
  assign other_ops_3_I1_1 = I1_4_1; // @[Map2S.scala 23:43]
  assign other_ops_3_I1_2 = I1_4_2; // @[Map2S.scala 23:43]
  assign other_ops_4_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_4_I0_0 = I0_5_0; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_1 = I0_5_1; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_2 = I0_5_2; // @[Map2S.scala 22:43]
  assign other_ops_4_I1_0 = I1_5_0; // @[Map2S.scala 23:43]
  assign other_ops_4_I1_1 = I1_5_1; // @[Map2S.scala 23:43]
  assign other_ops_4_I1_2 = I1_5_2; // @[Map2S.scala 23:43]
  assign other_ops_5_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_5_I0_0 = I0_6_0; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_1 = I0_6_1; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_2 = I0_6_2; // @[Map2S.scala 22:43]
  assign other_ops_5_I1_0 = I1_6_0; // @[Map2S.scala 23:43]
  assign other_ops_5_I1_1 = I1_6_1; // @[Map2S.scala 23:43]
  assign other_ops_5_I1_2 = I1_6_2; // @[Map2S.scala 23:43]
  assign other_ops_6_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_6_I0_0 = I0_7_0; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_1 = I0_7_1; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_2 = I0_7_2; // @[Map2S.scala 22:43]
  assign other_ops_6_I1_0 = I1_7_0; // @[Map2S.scala 23:43]
  assign other_ops_6_I1_1 = I1_7_1; // @[Map2S.scala 23:43]
  assign other_ops_6_I1_2 = I1_7_2; // @[Map2S.scala 23:43]
endmodule
module Map2T_4(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0_0,
  input  [31:0] I0_0_1,
  input  [31:0] I0_0_2,
  input  [31:0] I0_1_0,
  input  [31:0] I0_1_1,
  input  [31:0] I0_1_2,
  input  [31:0] I0_2_0,
  input  [31:0] I0_2_1,
  input  [31:0] I0_2_2,
  input  [31:0] I0_3_0,
  input  [31:0] I0_3_1,
  input  [31:0] I0_3_2,
  input  [31:0] I0_4_0,
  input  [31:0] I0_4_1,
  input  [31:0] I0_4_2,
  input  [31:0] I0_5_0,
  input  [31:0] I0_5_1,
  input  [31:0] I0_5_2,
  input  [31:0] I0_6_0,
  input  [31:0] I0_6_1,
  input  [31:0] I0_6_2,
  input  [31:0] I0_7_0,
  input  [31:0] I0_7_1,
  input  [31:0] I0_7_2,
  input  [31:0] I1_0_0,
  input  [31:0] I1_0_1,
  input  [31:0] I1_0_2,
  input  [31:0] I1_1_0,
  input  [31:0] I1_1_1,
  input  [31:0] I1_1_2,
  input  [31:0] I1_2_0,
  input  [31:0] I1_2_1,
  input  [31:0] I1_2_2,
  input  [31:0] I1_3_0,
  input  [31:0] I1_3_1,
  input  [31:0] I1_3_2,
  input  [31:0] I1_4_0,
  input  [31:0] I1_4_1,
  input  [31:0] I1_4_2,
  input  [31:0] I1_5_0,
  input  [31:0] I1_5_1,
  input  [31:0] I1_5_2,
  input  [31:0] I1_6_0,
  input  [31:0] I1_6_1,
  input  [31:0] I1_6_2,
  input  [31:0] I1_7_0,
  input  [31:0] I1_7_1,
  input  [31:0] I1_7_2,
  output [31:0] O_0_0_0,
  output [31:0] O_0_0_1,
  output [31:0] O_0_0_2,
  output [31:0] O_0_1_0,
  output [31:0] O_0_1_1,
  output [31:0] O_0_1_2,
  output [31:0] O_1_0_0,
  output [31:0] O_1_0_1,
  output [31:0] O_1_0_2,
  output [31:0] O_1_1_0,
  output [31:0] O_1_1_1,
  output [31:0] O_1_1_2,
  output [31:0] O_2_0_0,
  output [31:0] O_2_0_1,
  output [31:0] O_2_0_2,
  output [31:0] O_2_1_0,
  output [31:0] O_2_1_1,
  output [31:0] O_2_1_2,
  output [31:0] O_3_0_0,
  output [31:0] O_3_0_1,
  output [31:0] O_3_0_2,
  output [31:0] O_3_1_0,
  output [31:0] O_3_1_1,
  output [31:0] O_3_1_2,
  output [31:0] O_4_0_0,
  output [31:0] O_4_0_1,
  output [31:0] O_4_0_2,
  output [31:0] O_4_1_0,
  output [31:0] O_4_1_1,
  output [31:0] O_4_1_2,
  output [31:0] O_5_0_0,
  output [31:0] O_5_0_1,
  output [31:0] O_5_0_2,
  output [31:0] O_5_1_0,
  output [31:0] O_5_1_1,
  output [31:0] O_5_1_2,
  output [31:0] O_6_0_0,
  output [31:0] O_6_0_1,
  output [31:0] O_6_0_2,
  output [31:0] O_6_1_0,
  output [31:0] O_6_1_1,
  output [31:0] O_6_1_2,
  output [31:0] O_7_0_0,
  output [31:0] O_7_0_1,
  output [31:0] O_7_0_2,
  output [31:0] O_7_1_0,
  output [31:0] O_7_1_1,
  output [31:0] O_7_1_2
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_3_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_3_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_3_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_4_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_4_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_4_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_5_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_5_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_5_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_6_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_6_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_6_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_7_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_7_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_7_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_1_2; // @[Map2T.scala 8:20]
  Map2S_4 op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0_0(op_I0_0_0),
    .I0_0_1(op_I0_0_1),
    .I0_0_2(op_I0_0_2),
    .I0_1_0(op_I0_1_0),
    .I0_1_1(op_I0_1_1),
    .I0_1_2(op_I0_1_2),
    .I0_2_0(op_I0_2_0),
    .I0_2_1(op_I0_2_1),
    .I0_2_2(op_I0_2_2),
    .I0_3_0(op_I0_3_0),
    .I0_3_1(op_I0_3_1),
    .I0_3_2(op_I0_3_2),
    .I0_4_0(op_I0_4_0),
    .I0_4_1(op_I0_4_1),
    .I0_4_2(op_I0_4_2),
    .I0_5_0(op_I0_5_0),
    .I0_5_1(op_I0_5_1),
    .I0_5_2(op_I0_5_2),
    .I0_6_0(op_I0_6_0),
    .I0_6_1(op_I0_6_1),
    .I0_6_2(op_I0_6_2),
    .I0_7_0(op_I0_7_0),
    .I0_7_1(op_I0_7_1),
    .I0_7_2(op_I0_7_2),
    .I1_0_0(op_I1_0_0),
    .I1_0_1(op_I1_0_1),
    .I1_0_2(op_I1_0_2),
    .I1_1_0(op_I1_1_0),
    .I1_1_1(op_I1_1_1),
    .I1_1_2(op_I1_1_2),
    .I1_2_0(op_I1_2_0),
    .I1_2_1(op_I1_2_1),
    .I1_2_2(op_I1_2_2),
    .I1_3_0(op_I1_3_0),
    .I1_3_1(op_I1_3_1),
    .I1_3_2(op_I1_3_2),
    .I1_4_0(op_I1_4_0),
    .I1_4_1(op_I1_4_1),
    .I1_4_2(op_I1_4_2),
    .I1_5_0(op_I1_5_0),
    .I1_5_1(op_I1_5_1),
    .I1_5_2(op_I1_5_2),
    .I1_6_0(op_I1_6_0),
    .I1_6_1(op_I1_6_1),
    .I1_6_2(op_I1_6_2),
    .I1_7_0(op_I1_7_0),
    .I1_7_1(op_I1_7_1),
    .I1_7_2(op_I1_7_2),
    .O_0_0_0(op_O_0_0_0),
    .O_0_0_1(op_O_0_0_1),
    .O_0_0_2(op_O_0_0_2),
    .O_0_1_0(op_O_0_1_0),
    .O_0_1_1(op_O_0_1_1),
    .O_0_1_2(op_O_0_1_2),
    .O_1_0_0(op_O_1_0_0),
    .O_1_0_1(op_O_1_0_1),
    .O_1_0_2(op_O_1_0_2),
    .O_1_1_0(op_O_1_1_0),
    .O_1_1_1(op_O_1_1_1),
    .O_1_1_2(op_O_1_1_2),
    .O_2_0_0(op_O_2_0_0),
    .O_2_0_1(op_O_2_0_1),
    .O_2_0_2(op_O_2_0_2),
    .O_2_1_0(op_O_2_1_0),
    .O_2_1_1(op_O_2_1_1),
    .O_2_1_2(op_O_2_1_2),
    .O_3_0_0(op_O_3_0_0),
    .O_3_0_1(op_O_3_0_1),
    .O_3_0_2(op_O_3_0_2),
    .O_3_1_0(op_O_3_1_0),
    .O_3_1_1(op_O_3_1_1),
    .O_3_1_2(op_O_3_1_2),
    .O_4_0_0(op_O_4_0_0),
    .O_4_0_1(op_O_4_0_1),
    .O_4_0_2(op_O_4_0_2),
    .O_4_1_0(op_O_4_1_0),
    .O_4_1_1(op_O_4_1_1),
    .O_4_1_2(op_O_4_1_2),
    .O_5_0_0(op_O_5_0_0),
    .O_5_0_1(op_O_5_0_1),
    .O_5_0_2(op_O_5_0_2),
    .O_5_1_0(op_O_5_1_0),
    .O_5_1_1(op_O_5_1_1),
    .O_5_1_2(op_O_5_1_2),
    .O_6_0_0(op_O_6_0_0),
    .O_6_0_1(op_O_6_0_1),
    .O_6_0_2(op_O_6_0_2),
    .O_6_1_0(op_O_6_1_0),
    .O_6_1_1(op_O_6_1_1),
    .O_6_1_2(op_O_6_1_2),
    .O_7_0_0(op_O_7_0_0),
    .O_7_0_1(op_O_7_0_1),
    .O_7_0_2(op_O_7_0_2),
    .O_7_1_0(op_O_7_1_0),
    .O_7_1_1(op_O_7_1_1),
    .O_7_1_2(op_O_7_1_2)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_0_0 = op_O_0_0_0; // @[Map2T.scala 17:7]
  assign O_0_0_1 = op_O_0_0_1; // @[Map2T.scala 17:7]
  assign O_0_0_2 = op_O_0_0_2; // @[Map2T.scala 17:7]
  assign O_0_1_0 = op_O_0_1_0; // @[Map2T.scala 17:7]
  assign O_0_1_1 = op_O_0_1_1; // @[Map2T.scala 17:7]
  assign O_0_1_2 = op_O_0_1_2; // @[Map2T.scala 17:7]
  assign O_1_0_0 = op_O_1_0_0; // @[Map2T.scala 17:7]
  assign O_1_0_1 = op_O_1_0_1; // @[Map2T.scala 17:7]
  assign O_1_0_2 = op_O_1_0_2; // @[Map2T.scala 17:7]
  assign O_1_1_0 = op_O_1_1_0; // @[Map2T.scala 17:7]
  assign O_1_1_1 = op_O_1_1_1; // @[Map2T.scala 17:7]
  assign O_1_1_2 = op_O_1_1_2; // @[Map2T.scala 17:7]
  assign O_2_0_0 = op_O_2_0_0; // @[Map2T.scala 17:7]
  assign O_2_0_1 = op_O_2_0_1; // @[Map2T.scala 17:7]
  assign O_2_0_2 = op_O_2_0_2; // @[Map2T.scala 17:7]
  assign O_2_1_0 = op_O_2_1_0; // @[Map2T.scala 17:7]
  assign O_2_1_1 = op_O_2_1_1; // @[Map2T.scala 17:7]
  assign O_2_1_2 = op_O_2_1_2; // @[Map2T.scala 17:7]
  assign O_3_0_0 = op_O_3_0_0; // @[Map2T.scala 17:7]
  assign O_3_0_1 = op_O_3_0_1; // @[Map2T.scala 17:7]
  assign O_3_0_2 = op_O_3_0_2; // @[Map2T.scala 17:7]
  assign O_3_1_0 = op_O_3_1_0; // @[Map2T.scala 17:7]
  assign O_3_1_1 = op_O_3_1_1; // @[Map2T.scala 17:7]
  assign O_3_1_2 = op_O_3_1_2; // @[Map2T.scala 17:7]
  assign O_4_0_0 = op_O_4_0_0; // @[Map2T.scala 17:7]
  assign O_4_0_1 = op_O_4_0_1; // @[Map2T.scala 17:7]
  assign O_4_0_2 = op_O_4_0_2; // @[Map2T.scala 17:7]
  assign O_4_1_0 = op_O_4_1_0; // @[Map2T.scala 17:7]
  assign O_4_1_1 = op_O_4_1_1; // @[Map2T.scala 17:7]
  assign O_4_1_2 = op_O_4_1_2; // @[Map2T.scala 17:7]
  assign O_5_0_0 = op_O_5_0_0; // @[Map2T.scala 17:7]
  assign O_5_0_1 = op_O_5_0_1; // @[Map2T.scala 17:7]
  assign O_5_0_2 = op_O_5_0_2; // @[Map2T.scala 17:7]
  assign O_5_1_0 = op_O_5_1_0; // @[Map2T.scala 17:7]
  assign O_5_1_1 = op_O_5_1_1; // @[Map2T.scala 17:7]
  assign O_5_1_2 = op_O_5_1_2; // @[Map2T.scala 17:7]
  assign O_6_0_0 = op_O_6_0_0; // @[Map2T.scala 17:7]
  assign O_6_0_1 = op_O_6_0_1; // @[Map2T.scala 17:7]
  assign O_6_0_2 = op_O_6_0_2; // @[Map2T.scala 17:7]
  assign O_6_1_0 = op_O_6_1_0; // @[Map2T.scala 17:7]
  assign O_6_1_1 = op_O_6_1_1; // @[Map2T.scala 17:7]
  assign O_6_1_2 = op_O_6_1_2; // @[Map2T.scala 17:7]
  assign O_7_0_0 = op_O_7_0_0; // @[Map2T.scala 17:7]
  assign O_7_0_1 = op_O_7_0_1; // @[Map2T.scala 17:7]
  assign O_7_0_2 = op_O_7_0_2; // @[Map2T.scala 17:7]
  assign O_7_1_0 = op_O_7_1_0; // @[Map2T.scala 17:7]
  assign O_7_1_1 = op_O_7_1_1; // @[Map2T.scala 17:7]
  assign O_7_1_2 = op_O_7_1_2; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0_0 = I0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_0_1 = I0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_0_2 = I0_0_2; // @[Map2T.scala 15:11]
  assign op_I0_1_0 = I0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_1_1 = I0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_1_2 = I0_1_2; // @[Map2T.scala 15:11]
  assign op_I0_2_0 = I0_2_0; // @[Map2T.scala 15:11]
  assign op_I0_2_1 = I0_2_1; // @[Map2T.scala 15:11]
  assign op_I0_2_2 = I0_2_2; // @[Map2T.scala 15:11]
  assign op_I0_3_0 = I0_3_0; // @[Map2T.scala 15:11]
  assign op_I0_3_1 = I0_3_1; // @[Map2T.scala 15:11]
  assign op_I0_3_2 = I0_3_2; // @[Map2T.scala 15:11]
  assign op_I0_4_0 = I0_4_0; // @[Map2T.scala 15:11]
  assign op_I0_4_1 = I0_4_1; // @[Map2T.scala 15:11]
  assign op_I0_4_2 = I0_4_2; // @[Map2T.scala 15:11]
  assign op_I0_5_0 = I0_5_0; // @[Map2T.scala 15:11]
  assign op_I0_5_1 = I0_5_1; // @[Map2T.scala 15:11]
  assign op_I0_5_2 = I0_5_2; // @[Map2T.scala 15:11]
  assign op_I0_6_0 = I0_6_0; // @[Map2T.scala 15:11]
  assign op_I0_6_1 = I0_6_1; // @[Map2T.scala 15:11]
  assign op_I0_6_2 = I0_6_2; // @[Map2T.scala 15:11]
  assign op_I0_7_0 = I0_7_0; // @[Map2T.scala 15:11]
  assign op_I0_7_1 = I0_7_1; // @[Map2T.scala 15:11]
  assign op_I0_7_2 = I0_7_2; // @[Map2T.scala 15:11]
  assign op_I1_0_0 = I1_0_0; // @[Map2T.scala 16:11]
  assign op_I1_0_1 = I1_0_1; // @[Map2T.scala 16:11]
  assign op_I1_0_2 = I1_0_2; // @[Map2T.scala 16:11]
  assign op_I1_1_0 = I1_1_0; // @[Map2T.scala 16:11]
  assign op_I1_1_1 = I1_1_1; // @[Map2T.scala 16:11]
  assign op_I1_1_2 = I1_1_2; // @[Map2T.scala 16:11]
  assign op_I1_2_0 = I1_2_0; // @[Map2T.scala 16:11]
  assign op_I1_2_1 = I1_2_1; // @[Map2T.scala 16:11]
  assign op_I1_2_2 = I1_2_2; // @[Map2T.scala 16:11]
  assign op_I1_3_0 = I1_3_0; // @[Map2T.scala 16:11]
  assign op_I1_3_1 = I1_3_1; // @[Map2T.scala 16:11]
  assign op_I1_3_2 = I1_3_2; // @[Map2T.scala 16:11]
  assign op_I1_4_0 = I1_4_0; // @[Map2T.scala 16:11]
  assign op_I1_4_1 = I1_4_1; // @[Map2T.scala 16:11]
  assign op_I1_4_2 = I1_4_2; // @[Map2T.scala 16:11]
  assign op_I1_5_0 = I1_5_0; // @[Map2T.scala 16:11]
  assign op_I1_5_1 = I1_5_1; // @[Map2T.scala 16:11]
  assign op_I1_5_2 = I1_5_2; // @[Map2T.scala 16:11]
  assign op_I1_6_0 = I1_6_0; // @[Map2T.scala 16:11]
  assign op_I1_6_1 = I1_6_1; // @[Map2T.scala 16:11]
  assign op_I1_6_2 = I1_6_2; // @[Map2T.scala 16:11]
  assign op_I1_7_0 = I1_7_0; // @[Map2T.scala 16:11]
  assign op_I1_7_1 = I1_7_1; // @[Map2T.scala 16:11]
  assign op_I1_7_2 = I1_7_2; // @[Map2T.scala 16:11]
endmodule
module SSeqTupleAppender_3(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0_0,
  input  [31:0] I0_0_1,
  input  [31:0] I0_0_2,
  input  [31:0] I0_1_0,
  input  [31:0] I0_1_1,
  input  [31:0] I0_1_2,
  input  [31:0] I1_0,
  input  [31:0] I1_1,
  input  [31:0] I1_2,
  output [31:0] O_0_0,
  output [31:0] O_0_1,
  output [31:0] O_0_2,
  output [31:0] O_1_0,
  output [31:0] O_1_1,
  output [31:0] O_1_2,
  output [31:0] O_2_0,
  output [31:0] O_2_1,
  output [31:0] O_2_2
);
  assign valid_down = valid_up; // @[Tuple.scala 28:14]
  assign O_0_0 = I0_0_0; // @[Tuple.scala 24:34]
  assign O_0_1 = I0_0_1; // @[Tuple.scala 24:34]
  assign O_0_2 = I0_0_2; // @[Tuple.scala 24:34]
  assign O_1_0 = I0_1_0; // @[Tuple.scala 24:34]
  assign O_1_1 = I0_1_1; // @[Tuple.scala 24:34]
  assign O_1_2 = I0_1_2; // @[Tuple.scala 24:34]
  assign O_2_0 = I1_0; // @[Tuple.scala 26:32]
  assign O_2_1 = I1_1; // @[Tuple.scala 26:32]
  assign O_2_2 = I1_2; // @[Tuple.scala 26:32]
endmodule
module Map2S_7(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0_0_0,
  input  [31:0] I0_0_0_1,
  input  [31:0] I0_0_0_2,
  input  [31:0] I0_0_1_0,
  input  [31:0] I0_0_1_1,
  input  [31:0] I0_0_1_2,
  input  [31:0] I0_1_0_0,
  input  [31:0] I0_1_0_1,
  input  [31:0] I0_1_0_2,
  input  [31:0] I0_1_1_0,
  input  [31:0] I0_1_1_1,
  input  [31:0] I0_1_1_2,
  input  [31:0] I0_2_0_0,
  input  [31:0] I0_2_0_1,
  input  [31:0] I0_2_0_2,
  input  [31:0] I0_2_1_0,
  input  [31:0] I0_2_1_1,
  input  [31:0] I0_2_1_2,
  input  [31:0] I0_3_0_0,
  input  [31:0] I0_3_0_1,
  input  [31:0] I0_3_0_2,
  input  [31:0] I0_3_1_0,
  input  [31:0] I0_3_1_1,
  input  [31:0] I0_3_1_2,
  input  [31:0] I0_4_0_0,
  input  [31:0] I0_4_0_1,
  input  [31:0] I0_4_0_2,
  input  [31:0] I0_4_1_0,
  input  [31:0] I0_4_1_1,
  input  [31:0] I0_4_1_2,
  input  [31:0] I0_5_0_0,
  input  [31:0] I0_5_0_1,
  input  [31:0] I0_5_0_2,
  input  [31:0] I0_5_1_0,
  input  [31:0] I0_5_1_1,
  input  [31:0] I0_5_1_2,
  input  [31:0] I0_6_0_0,
  input  [31:0] I0_6_0_1,
  input  [31:0] I0_6_0_2,
  input  [31:0] I0_6_1_0,
  input  [31:0] I0_6_1_1,
  input  [31:0] I0_6_1_2,
  input  [31:0] I0_7_0_0,
  input  [31:0] I0_7_0_1,
  input  [31:0] I0_7_0_2,
  input  [31:0] I0_7_1_0,
  input  [31:0] I0_7_1_1,
  input  [31:0] I0_7_1_2,
  input  [31:0] I1_0_0,
  input  [31:0] I1_0_1,
  input  [31:0] I1_0_2,
  input  [31:0] I1_1_0,
  input  [31:0] I1_1_1,
  input  [31:0] I1_1_2,
  input  [31:0] I1_2_0,
  input  [31:0] I1_2_1,
  input  [31:0] I1_2_2,
  input  [31:0] I1_3_0,
  input  [31:0] I1_3_1,
  input  [31:0] I1_3_2,
  input  [31:0] I1_4_0,
  input  [31:0] I1_4_1,
  input  [31:0] I1_4_2,
  input  [31:0] I1_5_0,
  input  [31:0] I1_5_1,
  input  [31:0] I1_5_2,
  input  [31:0] I1_6_0,
  input  [31:0] I1_6_1,
  input  [31:0] I1_6_2,
  input  [31:0] I1_7_0,
  input  [31:0] I1_7_1,
  input  [31:0] I1_7_2,
  output [31:0] O_0_0_0,
  output [31:0] O_0_0_1,
  output [31:0] O_0_0_2,
  output [31:0] O_0_1_0,
  output [31:0] O_0_1_1,
  output [31:0] O_0_1_2,
  output [31:0] O_0_2_0,
  output [31:0] O_0_2_1,
  output [31:0] O_0_2_2,
  output [31:0] O_1_0_0,
  output [31:0] O_1_0_1,
  output [31:0] O_1_0_2,
  output [31:0] O_1_1_0,
  output [31:0] O_1_1_1,
  output [31:0] O_1_1_2,
  output [31:0] O_1_2_0,
  output [31:0] O_1_2_1,
  output [31:0] O_1_2_2,
  output [31:0] O_2_0_0,
  output [31:0] O_2_0_1,
  output [31:0] O_2_0_2,
  output [31:0] O_2_1_0,
  output [31:0] O_2_1_1,
  output [31:0] O_2_1_2,
  output [31:0] O_2_2_0,
  output [31:0] O_2_2_1,
  output [31:0] O_2_2_2,
  output [31:0] O_3_0_0,
  output [31:0] O_3_0_1,
  output [31:0] O_3_0_2,
  output [31:0] O_3_1_0,
  output [31:0] O_3_1_1,
  output [31:0] O_3_1_2,
  output [31:0] O_3_2_0,
  output [31:0] O_3_2_1,
  output [31:0] O_3_2_2,
  output [31:0] O_4_0_0,
  output [31:0] O_4_0_1,
  output [31:0] O_4_0_2,
  output [31:0] O_4_1_0,
  output [31:0] O_4_1_1,
  output [31:0] O_4_1_2,
  output [31:0] O_4_2_0,
  output [31:0] O_4_2_1,
  output [31:0] O_4_2_2,
  output [31:0] O_5_0_0,
  output [31:0] O_5_0_1,
  output [31:0] O_5_0_2,
  output [31:0] O_5_1_0,
  output [31:0] O_5_1_1,
  output [31:0] O_5_1_2,
  output [31:0] O_5_2_0,
  output [31:0] O_5_2_1,
  output [31:0] O_5_2_2,
  output [31:0] O_6_0_0,
  output [31:0] O_6_0_1,
  output [31:0] O_6_0_2,
  output [31:0] O_6_1_0,
  output [31:0] O_6_1_1,
  output [31:0] O_6_1_2,
  output [31:0] O_6_2_0,
  output [31:0] O_6_2_1,
  output [31:0] O_6_2_2,
  output [31:0] O_7_0_0,
  output [31:0] O_7_0_1,
  output [31:0] O_7_0_2,
  output [31:0] O_7_1_0,
  output [31:0] O_7_1_1,
  output [31:0] O_7_1_2,
  output [31:0] O_7_2_0,
  output [31:0] O_7_2_1,
  output [31:0] O_7_2_2
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0_2; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_1_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_1_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_1_2; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_2; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_2; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_1_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_1_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_1_2; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_2_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_2_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_2_2; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_2_2; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  wire  _T_2; // @[Map2S.scala 26:83]
  wire  _T_3; // @[Map2S.scala 26:83]
  wire  _T_4; // @[Map2S.scala 26:83]
  wire  _T_5; // @[Map2S.scala 26:83]
  SSeqTupleAppender_3 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0_0(fst_op_I0_0_0),
    .I0_0_1(fst_op_I0_0_1),
    .I0_0_2(fst_op_I0_0_2),
    .I0_1_0(fst_op_I0_1_0),
    .I0_1_1(fst_op_I0_1_1),
    .I0_1_2(fst_op_I0_1_2),
    .I1_0(fst_op_I1_0),
    .I1_1(fst_op_I1_1),
    .I1_2(fst_op_I1_2),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1),
    .O_0_2(fst_op_O_0_2),
    .O_1_0(fst_op_O_1_0),
    .O_1_1(fst_op_O_1_1),
    .O_1_2(fst_op_O_1_2),
    .O_2_0(fst_op_O_2_0),
    .O_2_1(fst_op_O_2_1),
    .O_2_2(fst_op_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0_0(other_ops_0_I0_0_0),
    .I0_0_1(other_ops_0_I0_0_1),
    .I0_0_2(other_ops_0_I0_0_2),
    .I0_1_0(other_ops_0_I0_1_0),
    .I0_1_1(other_ops_0_I0_1_1),
    .I0_1_2(other_ops_0_I0_1_2),
    .I1_0(other_ops_0_I1_0),
    .I1_1(other_ops_0_I1_1),
    .I1_2(other_ops_0_I1_2),
    .O_0_0(other_ops_0_O_0_0),
    .O_0_1(other_ops_0_O_0_1),
    .O_0_2(other_ops_0_O_0_2),
    .O_1_0(other_ops_0_O_1_0),
    .O_1_1(other_ops_0_O_1_1),
    .O_1_2(other_ops_0_O_1_2),
    .O_2_0(other_ops_0_O_2_0),
    .O_2_1(other_ops_0_O_2_1),
    .O_2_2(other_ops_0_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0_0_0(other_ops_1_I0_0_0),
    .I0_0_1(other_ops_1_I0_0_1),
    .I0_0_2(other_ops_1_I0_0_2),
    .I0_1_0(other_ops_1_I0_1_0),
    .I0_1_1(other_ops_1_I0_1_1),
    .I0_1_2(other_ops_1_I0_1_2),
    .I1_0(other_ops_1_I1_0),
    .I1_1(other_ops_1_I1_1),
    .I1_2(other_ops_1_I1_2),
    .O_0_0(other_ops_1_O_0_0),
    .O_0_1(other_ops_1_O_0_1),
    .O_0_2(other_ops_1_O_0_2),
    .O_1_0(other_ops_1_O_1_0),
    .O_1_1(other_ops_1_O_1_1),
    .O_1_2(other_ops_1_O_1_2),
    .O_2_0(other_ops_1_O_2_0),
    .O_2_1(other_ops_1_O_2_1),
    .O_2_2(other_ops_1_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_2 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0_0_0(other_ops_2_I0_0_0),
    .I0_0_1(other_ops_2_I0_0_1),
    .I0_0_2(other_ops_2_I0_0_2),
    .I0_1_0(other_ops_2_I0_1_0),
    .I0_1_1(other_ops_2_I0_1_1),
    .I0_1_2(other_ops_2_I0_1_2),
    .I1_0(other_ops_2_I1_0),
    .I1_1(other_ops_2_I1_1),
    .I1_2(other_ops_2_I1_2),
    .O_0_0(other_ops_2_O_0_0),
    .O_0_1(other_ops_2_O_0_1),
    .O_0_2(other_ops_2_O_0_2),
    .O_1_0(other_ops_2_O_1_0),
    .O_1_1(other_ops_2_O_1_1),
    .O_1_2(other_ops_2_O_1_2),
    .O_2_0(other_ops_2_O_2_0),
    .O_2_1(other_ops_2_O_2_1),
    .O_2_2(other_ops_2_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_3 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I0_0_0(other_ops_3_I0_0_0),
    .I0_0_1(other_ops_3_I0_0_1),
    .I0_0_2(other_ops_3_I0_0_2),
    .I0_1_0(other_ops_3_I0_1_0),
    .I0_1_1(other_ops_3_I0_1_1),
    .I0_1_2(other_ops_3_I0_1_2),
    .I1_0(other_ops_3_I1_0),
    .I1_1(other_ops_3_I1_1),
    .I1_2(other_ops_3_I1_2),
    .O_0_0(other_ops_3_O_0_0),
    .O_0_1(other_ops_3_O_0_1),
    .O_0_2(other_ops_3_O_0_2),
    .O_1_0(other_ops_3_O_1_0),
    .O_1_1(other_ops_3_O_1_1),
    .O_1_2(other_ops_3_O_1_2),
    .O_2_0(other_ops_3_O_2_0),
    .O_2_1(other_ops_3_O_2_1),
    .O_2_2(other_ops_3_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_4 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I0_0_0(other_ops_4_I0_0_0),
    .I0_0_1(other_ops_4_I0_0_1),
    .I0_0_2(other_ops_4_I0_0_2),
    .I0_1_0(other_ops_4_I0_1_0),
    .I0_1_1(other_ops_4_I0_1_1),
    .I0_1_2(other_ops_4_I0_1_2),
    .I1_0(other_ops_4_I1_0),
    .I1_1(other_ops_4_I1_1),
    .I1_2(other_ops_4_I1_2),
    .O_0_0(other_ops_4_O_0_0),
    .O_0_1(other_ops_4_O_0_1),
    .O_0_2(other_ops_4_O_0_2),
    .O_1_0(other_ops_4_O_1_0),
    .O_1_1(other_ops_4_O_1_1),
    .O_1_2(other_ops_4_O_1_2),
    .O_2_0(other_ops_4_O_2_0),
    .O_2_1(other_ops_4_O_2_1),
    .O_2_2(other_ops_4_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_5 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I0_0_0(other_ops_5_I0_0_0),
    .I0_0_1(other_ops_5_I0_0_1),
    .I0_0_2(other_ops_5_I0_0_2),
    .I0_1_0(other_ops_5_I0_1_0),
    .I0_1_1(other_ops_5_I0_1_1),
    .I0_1_2(other_ops_5_I0_1_2),
    .I1_0(other_ops_5_I1_0),
    .I1_1(other_ops_5_I1_1),
    .I1_2(other_ops_5_I1_2),
    .O_0_0(other_ops_5_O_0_0),
    .O_0_1(other_ops_5_O_0_1),
    .O_0_2(other_ops_5_O_0_2),
    .O_1_0(other_ops_5_O_1_0),
    .O_1_1(other_ops_5_O_1_1),
    .O_1_2(other_ops_5_O_1_2),
    .O_2_0(other_ops_5_O_2_0),
    .O_2_1(other_ops_5_O_2_1),
    .O_2_2(other_ops_5_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_6 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I0_0_0(other_ops_6_I0_0_0),
    .I0_0_1(other_ops_6_I0_0_1),
    .I0_0_2(other_ops_6_I0_0_2),
    .I0_1_0(other_ops_6_I0_1_0),
    .I0_1_1(other_ops_6_I0_1_1),
    .I0_1_2(other_ops_6_I0_1_2),
    .I1_0(other_ops_6_I1_0),
    .I1_1(other_ops_6_I1_1),
    .I1_2(other_ops_6_I1_2),
    .O_0_0(other_ops_6_O_0_0),
    .O_0_1(other_ops_6_O_0_1),
    .O_0_2(other_ops_6_O_0_2),
    .O_1_0(other_ops_6_O_1_0),
    .O_1_1(other_ops_6_O_1_1),
    .O_1_2(other_ops_6_O_1_2),
    .O_2_0(other_ops_6_O_2_0),
    .O_2_1(other_ops_6_O_2_1),
    .O_2_2(other_ops_6_O_2_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[Map2S.scala 26:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[Map2S.scala 26:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_5 & other_ops_6_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[Map2S.scala 19:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[Map2S.scala 19:8]
  assign O_0_0_2 = fst_op_O_0_2; // @[Map2S.scala 19:8]
  assign O_0_1_0 = fst_op_O_1_0; // @[Map2S.scala 19:8]
  assign O_0_1_1 = fst_op_O_1_1; // @[Map2S.scala 19:8]
  assign O_0_1_2 = fst_op_O_1_2; // @[Map2S.scala 19:8]
  assign O_0_2_0 = fst_op_O_2_0; // @[Map2S.scala 19:8]
  assign O_0_2_1 = fst_op_O_2_1; // @[Map2S.scala 19:8]
  assign O_0_2_2 = fst_op_O_2_2; // @[Map2S.scala 19:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[Map2S.scala 24:12]
  assign O_1_0_1 = other_ops_0_O_0_1; // @[Map2S.scala 24:12]
  assign O_1_0_2 = other_ops_0_O_0_2; // @[Map2S.scala 24:12]
  assign O_1_1_0 = other_ops_0_O_1_0; // @[Map2S.scala 24:12]
  assign O_1_1_1 = other_ops_0_O_1_1; // @[Map2S.scala 24:12]
  assign O_1_1_2 = other_ops_0_O_1_2; // @[Map2S.scala 24:12]
  assign O_1_2_0 = other_ops_0_O_2_0; // @[Map2S.scala 24:12]
  assign O_1_2_1 = other_ops_0_O_2_1; // @[Map2S.scala 24:12]
  assign O_1_2_2 = other_ops_0_O_2_2; // @[Map2S.scala 24:12]
  assign O_2_0_0 = other_ops_1_O_0_0; // @[Map2S.scala 24:12]
  assign O_2_0_1 = other_ops_1_O_0_1; // @[Map2S.scala 24:12]
  assign O_2_0_2 = other_ops_1_O_0_2; // @[Map2S.scala 24:12]
  assign O_2_1_0 = other_ops_1_O_1_0; // @[Map2S.scala 24:12]
  assign O_2_1_1 = other_ops_1_O_1_1; // @[Map2S.scala 24:12]
  assign O_2_1_2 = other_ops_1_O_1_2; // @[Map2S.scala 24:12]
  assign O_2_2_0 = other_ops_1_O_2_0; // @[Map2S.scala 24:12]
  assign O_2_2_1 = other_ops_1_O_2_1; // @[Map2S.scala 24:12]
  assign O_2_2_2 = other_ops_1_O_2_2; // @[Map2S.scala 24:12]
  assign O_3_0_0 = other_ops_2_O_0_0; // @[Map2S.scala 24:12]
  assign O_3_0_1 = other_ops_2_O_0_1; // @[Map2S.scala 24:12]
  assign O_3_0_2 = other_ops_2_O_0_2; // @[Map2S.scala 24:12]
  assign O_3_1_0 = other_ops_2_O_1_0; // @[Map2S.scala 24:12]
  assign O_3_1_1 = other_ops_2_O_1_1; // @[Map2S.scala 24:12]
  assign O_3_1_2 = other_ops_2_O_1_2; // @[Map2S.scala 24:12]
  assign O_3_2_0 = other_ops_2_O_2_0; // @[Map2S.scala 24:12]
  assign O_3_2_1 = other_ops_2_O_2_1; // @[Map2S.scala 24:12]
  assign O_3_2_2 = other_ops_2_O_2_2; // @[Map2S.scala 24:12]
  assign O_4_0_0 = other_ops_3_O_0_0; // @[Map2S.scala 24:12]
  assign O_4_0_1 = other_ops_3_O_0_1; // @[Map2S.scala 24:12]
  assign O_4_0_2 = other_ops_3_O_0_2; // @[Map2S.scala 24:12]
  assign O_4_1_0 = other_ops_3_O_1_0; // @[Map2S.scala 24:12]
  assign O_4_1_1 = other_ops_3_O_1_1; // @[Map2S.scala 24:12]
  assign O_4_1_2 = other_ops_3_O_1_2; // @[Map2S.scala 24:12]
  assign O_4_2_0 = other_ops_3_O_2_0; // @[Map2S.scala 24:12]
  assign O_4_2_1 = other_ops_3_O_2_1; // @[Map2S.scala 24:12]
  assign O_4_2_2 = other_ops_3_O_2_2; // @[Map2S.scala 24:12]
  assign O_5_0_0 = other_ops_4_O_0_0; // @[Map2S.scala 24:12]
  assign O_5_0_1 = other_ops_4_O_0_1; // @[Map2S.scala 24:12]
  assign O_5_0_2 = other_ops_4_O_0_2; // @[Map2S.scala 24:12]
  assign O_5_1_0 = other_ops_4_O_1_0; // @[Map2S.scala 24:12]
  assign O_5_1_1 = other_ops_4_O_1_1; // @[Map2S.scala 24:12]
  assign O_5_1_2 = other_ops_4_O_1_2; // @[Map2S.scala 24:12]
  assign O_5_2_0 = other_ops_4_O_2_0; // @[Map2S.scala 24:12]
  assign O_5_2_1 = other_ops_4_O_2_1; // @[Map2S.scala 24:12]
  assign O_5_2_2 = other_ops_4_O_2_2; // @[Map2S.scala 24:12]
  assign O_6_0_0 = other_ops_5_O_0_0; // @[Map2S.scala 24:12]
  assign O_6_0_1 = other_ops_5_O_0_1; // @[Map2S.scala 24:12]
  assign O_6_0_2 = other_ops_5_O_0_2; // @[Map2S.scala 24:12]
  assign O_6_1_0 = other_ops_5_O_1_0; // @[Map2S.scala 24:12]
  assign O_6_1_1 = other_ops_5_O_1_1; // @[Map2S.scala 24:12]
  assign O_6_1_2 = other_ops_5_O_1_2; // @[Map2S.scala 24:12]
  assign O_6_2_0 = other_ops_5_O_2_0; // @[Map2S.scala 24:12]
  assign O_6_2_1 = other_ops_5_O_2_1; // @[Map2S.scala 24:12]
  assign O_6_2_2 = other_ops_5_O_2_2; // @[Map2S.scala 24:12]
  assign O_7_0_0 = other_ops_6_O_0_0; // @[Map2S.scala 24:12]
  assign O_7_0_1 = other_ops_6_O_0_1; // @[Map2S.scala 24:12]
  assign O_7_0_2 = other_ops_6_O_0_2; // @[Map2S.scala 24:12]
  assign O_7_1_0 = other_ops_6_O_1_0; // @[Map2S.scala 24:12]
  assign O_7_1_1 = other_ops_6_O_1_1; // @[Map2S.scala 24:12]
  assign O_7_1_2 = other_ops_6_O_1_2; // @[Map2S.scala 24:12]
  assign O_7_2_0 = other_ops_6_O_2_0; // @[Map2S.scala 24:12]
  assign O_7_2_1 = other_ops_6_O_2_1; // @[Map2S.scala 24:12]
  assign O_7_2_2 = other_ops_6_O_2_2; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0_0 = I0_0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_1 = I0_0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_2 = I0_0_0_2; // @[Map2S.scala 17:13]
  assign fst_op_I0_1_0 = I0_0_1_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1_1 = I0_0_1_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_1_2 = I0_0_1_2; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = I1_0_0; // @[Map2S.scala 18:13]
  assign fst_op_I1_1 = I1_0_1; // @[Map2S.scala 18:13]
  assign fst_op_I1_2 = I1_0_2; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0_0 = I0_1_0_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_0_1 = I0_1_0_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_0_2 = I0_1_0_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1_0 = I0_1_1_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1_1 = I0_1_1_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1_2 = I0_1_1_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I1_0 = I1_1_0; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_1 = I1_1_1; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_2 = I1_1_2; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0_0_0 = I0_2_0_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_0_1 = I0_2_0_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_0_2 = I0_2_0_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1_0 = I0_2_1_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1_1 = I0_2_1_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1_2 = I0_2_1_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1_0 = I1_2_0; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_1 = I1_2_1; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_2 = I1_2_2; // @[Map2S.scala 23:43]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0_0_0 = I0_3_0_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_0_1 = I0_3_0_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_0_2 = I0_3_0_2; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_1_0 = I0_3_1_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_1_1 = I0_3_1_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_1_2 = I0_3_1_2; // @[Map2S.scala 22:43]
  assign other_ops_2_I1_0 = I1_3_0; // @[Map2S.scala 23:43]
  assign other_ops_2_I1_1 = I1_3_1; // @[Map2S.scala 23:43]
  assign other_ops_2_I1_2 = I1_3_2; // @[Map2S.scala 23:43]
  assign other_ops_3_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_3_I0_0_0 = I0_4_0_0; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_0_1 = I0_4_0_1; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_0_2 = I0_4_0_2; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_1_0 = I0_4_1_0; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_1_1 = I0_4_1_1; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_1_2 = I0_4_1_2; // @[Map2S.scala 22:43]
  assign other_ops_3_I1_0 = I1_4_0; // @[Map2S.scala 23:43]
  assign other_ops_3_I1_1 = I1_4_1; // @[Map2S.scala 23:43]
  assign other_ops_3_I1_2 = I1_4_2; // @[Map2S.scala 23:43]
  assign other_ops_4_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_4_I0_0_0 = I0_5_0_0; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_0_1 = I0_5_0_1; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_0_2 = I0_5_0_2; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_1_0 = I0_5_1_0; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_1_1 = I0_5_1_1; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_1_2 = I0_5_1_2; // @[Map2S.scala 22:43]
  assign other_ops_4_I1_0 = I1_5_0; // @[Map2S.scala 23:43]
  assign other_ops_4_I1_1 = I1_5_1; // @[Map2S.scala 23:43]
  assign other_ops_4_I1_2 = I1_5_2; // @[Map2S.scala 23:43]
  assign other_ops_5_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_5_I0_0_0 = I0_6_0_0; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_0_1 = I0_6_0_1; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_0_2 = I0_6_0_2; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_1_0 = I0_6_1_0; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_1_1 = I0_6_1_1; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_1_2 = I0_6_1_2; // @[Map2S.scala 22:43]
  assign other_ops_5_I1_0 = I1_6_0; // @[Map2S.scala 23:43]
  assign other_ops_5_I1_1 = I1_6_1; // @[Map2S.scala 23:43]
  assign other_ops_5_I1_2 = I1_6_2; // @[Map2S.scala 23:43]
  assign other_ops_6_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_6_I0_0_0 = I0_7_0_0; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_0_1 = I0_7_0_1; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_0_2 = I0_7_0_2; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_1_0 = I0_7_1_0; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_1_1 = I0_7_1_1; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_1_2 = I0_7_1_2; // @[Map2S.scala 22:43]
  assign other_ops_6_I1_0 = I1_7_0; // @[Map2S.scala 23:43]
  assign other_ops_6_I1_1 = I1_7_1; // @[Map2S.scala 23:43]
  assign other_ops_6_I1_2 = I1_7_2; // @[Map2S.scala 23:43]
endmodule
module Map2T_7(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0_0_0,
  input  [31:0] I0_0_0_1,
  input  [31:0] I0_0_0_2,
  input  [31:0] I0_0_1_0,
  input  [31:0] I0_0_1_1,
  input  [31:0] I0_0_1_2,
  input  [31:0] I0_1_0_0,
  input  [31:0] I0_1_0_1,
  input  [31:0] I0_1_0_2,
  input  [31:0] I0_1_1_0,
  input  [31:0] I0_1_1_1,
  input  [31:0] I0_1_1_2,
  input  [31:0] I0_2_0_0,
  input  [31:0] I0_2_0_1,
  input  [31:0] I0_2_0_2,
  input  [31:0] I0_2_1_0,
  input  [31:0] I0_2_1_1,
  input  [31:0] I0_2_1_2,
  input  [31:0] I0_3_0_0,
  input  [31:0] I0_3_0_1,
  input  [31:0] I0_3_0_2,
  input  [31:0] I0_3_1_0,
  input  [31:0] I0_3_1_1,
  input  [31:0] I0_3_1_2,
  input  [31:0] I0_4_0_0,
  input  [31:0] I0_4_0_1,
  input  [31:0] I0_4_0_2,
  input  [31:0] I0_4_1_0,
  input  [31:0] I0_4_1_1,
  input  [31:0] I0_4_1_2,
  input  [31:0] I0_5_0_0,
  input  [31:0] I0_5_0_1,
  input  [31:0] I0_5_0_2,
  input  [31:0] I0_5_1_0,
  input  [31:0] I0_5_1_1,
  input  [31:0] I0_5_1_2,
  input  [31:0] I0_6_0_0,
  input  [31:0] I0_6_0_1,
  input  [31:0] I0_6_0_2,
  input  [31:0] I0_6_1_0,
  input  [31:0] I0_6_1_1,
  input  [31:0] I0_6_1_2,
  input  [31:0] I0_7_0_0,
  input  [31:0] I0_7_0_1,
  input  [31:0] I0_7_0_2,
  input  [31:0] I0_7_1_0,
  input  [31:0] I0_7_1_1,
  input  [31:0] I0_7_1_2,
  input  [31:0] I1_0_0,
  input  [31:0] I1_0_1,
  input  [31:0] I1_0_2,
  input  [31:0] I1_1_0,
  input  [31:0] I1_1_1,
  input  [31:0] I1_1_2,
  input  [31:0] I1_2_0,
  input  [31:0] I1_2_1,
  input  [31:0] I1_2_2,
  input  [31:0] I1_3_0,
  input  [31:0] I1_3_1,
  input  [31:0] I1_3_2,
  input  [31:0] I1_4_0,
  input  [31:0] I1_4_1,
  input  [31:0] I1_4_2,
  input  [31:0] I1_5_0,
  input  [31:0] I1_5_1,
  input  [31:0] I1_5_2,
  input  [31:0] I1_6_0,
  input  [31:0] I1_6_1,
  input  [31:0] I1_6_2,
  input  [31:0] I1_7_0,
  input  [31:0] I1_7_1,
  input  [31:0] I1_7_2,
  output [31:0] O_0_0_0,
  output [31:0] O_0_0_1,
  output [31:0] O_0_0_2,
  output [31:0] O_0_1_0,
  output [31:0] O_0_1_1,
  output [31:0] O_0_1_2,
  output [31:0] O_0_2_0,
  output [31:0] O_0_2_1,
  output [31:0] O_0_2_2,
  output [31:0] O_1_0_0,
  output [31:0] O_1_0_1,
  output [31:0] O_1_0_2,
  output [31:0] O_1_1_0,
  output [31:0] O_1_1_1,
  output [31:0] O_1_1_2,
  output [31:0] O_1_2_0,
  output [31:0] O_1_2_1,
  output [31:0] O_1_2_2,
  output [31:0] O_2_0_0,
  output [31:0] O_2_0_1,
  output [31:0] O_2_0_2,
  output [31:0] O_2_1_0,
  output [31:0] O_2_1_1,
  output [31:0] O_2_1_2,
  output [31:0] O_2_2_0,
  output [31:0] O_2_2_1,
  output [31:0] O_2_2_2,
  output [31:0] O_3_0_0,
  output [31:0] O_3_0_1,
  output [31:0] O_3_0_2,
  output [31:0] O_3_1_0,
  output [31:0] O_3_1_1,
  output [31:0] O_3_1_2,
  output [31:0] O_3_2_0,
  output [31:0] O_3_2_1,
  output [31:0] O_3_2_2,
  output [31:0] O_4_0_0,
  output [31:0] O_4_0_1,
  output [31:0] O_4_0_2,
  output [31:0] O_4_1_0,
  output [31:0] O_4_1_1,
  output [31:0] O_4_1_2,
  output [31:0] O_4_2_0,
  output [31:0] O_4_2_1,
  output [31:0] O_4_2_2,
  output [31:0] O_5_0_0,
  output [31:0] O_5_0_1,
  output [31:0] O_5_0_2,
  output [31:0] O_5_1_0,
  output [31:0] O_5_1_1,
  output [31:0] O_5_1_2,
  output [31:0] O_5_2_0,
  output [31:0] O_5_2_1,
  output [31:0] O_5_2_2,
  output [31:0] O_6_0_0,
  output [31:0] O_6_0_1,
  output [31:0] O_6_0_2,
  output [31:0] O_6_1_0,
  output [31:0] O_6_1_1,
  output [31:0] O_6_1_2,
  output [31:0] O_6_2_0,
  output [31:0] O_6_2_1,
  output [31:0] O_6_2_2,
  output [31:0] O_7_0_0,
  output [31:0] O_7_0_1,
  output [31:0] O_7_0_2,
  output [31:0] O_7_1_0,
  output [31:0] O_7_1_1,
  output [31:0] O_7_1_2,
  output [31:0] O_7_2_0,
  output [31:0] O_7_2_1,
  output [31:0] O_7_2_2
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_3_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_3_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_3_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_4_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_4_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_4_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_5_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_5_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_5_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_6_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_6_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_6_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_7_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_7_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_7_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_2_2; // @[Map2T.scala 8:20]
  Map2S_7 op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0_0_0(op_I0_0_0_0),
    .I0_0_0_1(op_I0_0_0_1),
    .I0_0_0_2(op_I0_0_0_2),
    .I0_0_1_0(op_I0_0_1_0),
    .I0_0_1_1(op_I0_0_1_1),
    .I0_0_1_2(op_I0_0_1_2),
    .I0_1_0_0(op_I0_1_0_0),
    .I0_1_0_1(op_I0_1_0_1),
    .I0_1_0_2(op_I0_1_0_2),
    .I0_1_1_0(op_I0_1_1_0),
    .I0_1_1_1(op_I0_1_1_1),
    .I0_1_1_2(op_I0_1_1_2),
    .I0_2_0_0(op_I0_2_0_0),
    .I0_2_0_1(op_I0_2_0_1),
    .I0_2_0_2(op_I0_2_0_2),
    .I0_2_1_0(op_I0_2_1_0),
    .I0_2_1_1(op_I0_2_1_1),
    .I0_2_1_2(op_I0_2_1_2),
    .I0_3_0_0(op_I0_3_0_0),
    .I0_3_0_1(op_I0_3_0_1),
    .I0_3_0_2(op_I0_3_0_2),
    .I0_3_1_0(op_I0_3_1_0),
    .I0_3_1_1(op_I0_3_1_1),
    .I0_3_1_2(op_I0_3_1_2),
    .I0_4_0_0(op_I0_4_0_0),
    .I0_4_0_1(op_I0_4_0_1),
    .I0_4_0_2(op_I0_4_0_2),
    .I0_4_1_0(op_I0_4_1_0),
    .I0_4_1_1(op_I0_4_1_1),
    .I0_4_1_2(op_I0_4_1_2),
    .I0_5_0_0(op_I0_5_0_0),
    .I0_5_0_1(op_I0_5_0_1),
    .I0_5_0_2(op_I0_5_0_2),
    .I0_5_1_0(op_I0_5_1_0),
    .I0_5_1_1(op_I0_5_1_1),
    .I0_5_1_2(op_I0_5_1_2),
    .I0_6_0_0(op_I0_6_0_0),
    .I0_6_0_1(op_I0_6_0_1),
    .I0_6_0_2(op_I0_6_0_2),
    .I0_6_1_0(op_I0_6_1_0),
    .I0_6_1_1(op_I0_6_1_1),
    .I0_6_1_2(op_I0_6_1_2),
    .I0_7_0_0(op_I0_7_0_0),
    .I0_7_0_1(op_I0_7_0_1),
    .I0_7_0_2(op_I0_7_0_2),
    .I0_7_1_0(op_I0_7_1_0),
    .I0_7_1_1(op_I0_7_1_1),
    .I0_7_1_2(op_I0_7_1_2),
    .I1_0_0(op_I1_0_0),
    .I1_0_1(op_I1_0_1),
    .I1_0_2(op_I1_0_2),
    .I1_1_0(op_I1_1_0),
    .I1_1_1(op_I1_1_1),
    .I1_1_2(op_I1_1_2),
    .I1_2_0(op_I1_2_0),
    .I1_2_1(op_I1_2_1),
    .I1_2_2(op_I1_2_2),
    .I1_3_0(op_I1_3_0),
    .I1_3_1(op_I1_3_1),
    .I1_3_2(op_I1_3_2),
    .I1_4_0(op_I1_4_0),
    .I1_4_1(op_I1_4_1),
    .I1_4_2(op_I1_4_2),
    .I1_5_0(op_I1_5_0),
    .I1_5_1(op_I1_5_1),
    .I1_5_2(op_I1_5_2),
    .I1_6_0(op_I1_6_0),
    .I1_6_1(op_I1_6_1),
    .I1_6_2(op_I1_6_2),
    .I1_7_0(op_I1_7_0),
    .I1_7_1(op_I1_7_1),
    .I1_7_2(op_I1_7_2),
    .O_0_0_0(op_O_0_0_0),
    .O_0_0_1(op_O_0_0_1),
    .O_0_0_2(op_O_0_0_2),
    .O_0_1_0(op_O_0_1_0),
    .O_0_1_1(op_O_0_1_1),
    .O_0_1_2(op_O_0_1_2),
    .O_0_2_0(op_O_0_2_0),
    .O_0_2_1(op_O_0_2_1),
    .O_0_2_2(op_O_0_2_2),
    .O_1_0_0(op_O_1_0_0),
    .O_1_0_1(op_O_1_0_1),
    .O_1_0_2(op_O_1_0_2),
    .O_1_1_0(op_O_1_1_0),
    .O_1_1_1(op_O_1_1_1),
    .O_1_1_2(op_O_1_1_2),
    .O_1_2_0(op_O_1_2_0),
    .O_1_2_1(op_O_1_2_1),
    .O_1_2_2(op_O_1_2_2),
    .O_2_0_0(op_O_2_0_0),
    .O_2_0_1(op_O_2_0_1),
    .O_2_0_2(op_O_2_0_2),
    .O_2_1_0(op_O_2_1_0),
    .O_2_1_1(op_O_2_1_1),
    .O_2_1_2(op_O_2_1_2),
    .O_2_2_0(op_O_2_2_0),
    .O_2_2_1(op_O_2_2_1),
    .O_2_2_2(op_O_2_2_2),
    .O_3_0_0(op_O_3_0_0),
    .O_3_0_1(op_O_3_0_1),
    .O_3_0_2(op_O_3_0_2),
    .O_3_1_0(op_O_3_1_0),
    .O_3_1_1(op_O_3_1_1),
    .O_3_1_2(op_O_3_1_2),
    .O_3_2_0(op_O_3_2_0),
    .O_3_2_1(op_O_3_2_1),
    .O_3_2_2(op_O_3_2_2),
    .O_4_0_0(op_O_4_0_0),
    .O_4_0_1(op_O_4_0_1),
    .O_4_0_2(op_O_4_0_2),
    .O_4_1_0(op_O_4_1_0),
    .O_4_1_1(op_O_4_1_1),
    .O_4_1_2(op_O_4_1_2),
    .O_4_2_0(op_O_4_2_0),
    .O_4_2_1(op_O_4_2_1),
    .O_4_2_2(op_O_4_2_2),
    .O_5_0_0(op_O_5_0_0),
    .O_5_0_1(op_O_5_0_1),
    .O_5_0_2(op_O_5_0_2),
    .O_5_1_0(op_O_5_1_0),
    .O_5_1_1(op_O_5_1_1),
    .O_5_1_2(op_O_5_1_2),
    .O_5_2_0(op_O_5_2_0),
    .O_5_2_1(op_O_5_2_1),
    .O_5_2_2(op_O_5_2_2),
    .O_6_0_0(op_O_6_0_0),
    .O_6_0_1(op_O_6_0_1),
    .O_6_0_2(op_O_6_0_2),
    .O_6_1_0(op_O_6_1_0),
    .O_6_1_1(op_O_6_1_1),
    .O_6_1_2(op_O_6_1_2),
    .O_6_2_0(op_O_6_2_0),
    .O_6_2_1(op_O_6_2_1),
    .O_6_2_2(op_O_6_2_2),
    .O_7_0_0(op_O_7_0_0),
    .O_7_0_1(op_O_7_0_1),
    .O_7_0_2(op_O_7_0_2),
    .O_7_1_0(op_O_7_1_0),
    .O_7_1_1(op_O_7_1_1),
    .O_7_1_2(op_O_7_1_2),
    .O_7_2_0(op_O_7_2_0),
    .O_7_2_1(op_O_7_2_1),
    .O_7_2_2(op_O_7_2_2)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_0_0 = op_O_0_0_0; // @[Map2T.scala 17:7]
  assign O_0_0_1 = op_O_0_0_1; // @[Map2T.scala 17:7]
  assign O_0_0_2 = op_O_0_0_2; // @[Map2T.scala 17:7]
  assign O_0_1_0 = op_O_0_1_0; // @[Map2T.scala 17:7]
  assign O_0_1_1 = op_O_0_1_1; // @[Map2T.scala 17:7]
  assign O_0_1_2 = op_O_0_1_2; // @[Map2T.scala 17:7]
  assign O_0_2_0 = op_O_0_2_0; // @[Map2T.scala 17:7]
  assign O_0_2_1 = op_O_0_2_1; // @[Map2T.scala 17:7]
  assign O_0_2_2 = op_O_0_2_2; // @[Map2T.scala 17:7]
  assign O_1_0_0 = op_O_1_0_0; // @[Map2T.scala 17:7]
  assign O_1_0_1 = op_O_1_0_1; // @[Map2T.scala 17:7]
  assign O_1_0_2 = op_O_1_0_2; // @[Map2T.scala 17:7]
  assign O_1_1_0 = op_O_1_1_0; // @[Map2T.scala 17:7]
  assign O_1_1_1 = op_O_1_1_1; // @[Map2T.scala 17:7]
  assign O_1_1_2 = op_O_1_1_2; // @[Map2T.scala 17:7]
  assign O_1_2_0 = op_O_1_2_0; // @[Map2T.scala 17:7]
  assign O_1_2_1 = op_O_1_2_1; // @[Map2T.scala 17:7]
  assign O_1_2_2 = op_O_1_2_2; // @[Map2T.scala 17:7]
  assign O_2_0_0 = op_O_2_0_0; // @[Map2T.scala 17:7]
  assign O_2_0_1 = op_O_2_0_1; // @[Map2T.scala 17:7]
  assign O_2_0_2 = op_O_2_0_2; // @[Map2T.scala 17:7]
  assign O_2_1_0 = op_O_2_1_0; // @[Map2T.scala 17:7]
  assign O_2_1_1 = op_O_2_1_1; // @[Map2T.scala 17:7]
  assign O_2_1_2 = op_O_2_1_2; // @[Map2T.scala 17:7]
  assign O_2_2_0 = op_O_2_2_0; // @[Map2T.scala 17:7]
  assign O_2_2_1 = op_O_2_2_1; // @[Map2T.scala 17:7]
  assign O_2_2_2 = op_O_2_2_2; // @[Map2T.scala 17:7]
  assign O_3_0_0 = op_O_3_0_0; // @[Map2T.scala 17:7]
  assign O_3_0_1 = op_O_3_0_1; // @[Map2T.scala 17:7]
  assign O_3_0_2 = op_O_3_0_2; // @[Map2T.scala 17:7]
  assign O_3_1_0 = op_O_3_1_0; // @[Map2T.scala 17:7]
  assign O_3_1_1 = op_O_3_1_1; // @[Map2T.scala 17:7]
  assign O_3_1_2 = op_O_3_1_2; // @[Map2T.scala 17:7]
  assign O_3_2_0 = op_O_3_2_0; // @[Map2T.scala 17:7]
  assign O_3_2_1 = op_O_3_2_1; // @[Map2T.scala 17:7]
  assign O_3_2_2 = op_O_3_2_2; // @[Map2T.scala 17:7]
  assign O_4_0_0 = op_O_4_0_0; // @[Map2T.scala 17:7]
  assign O_4_0_1 = op_O_4_0_1; // @[Map2T.scala 17:7]
  assign O_4_0_2 = op_O_4_0_2; // @[Map2T.scala 17:7]
  assign O_4_1_0 = op_O_4_1_0; // @[Map2T.scala 17:7]
  assign O_4_1_1 = op_O_4_1_1; // @[Map2T.scala 17:7]
  assign O_4_1_2 = op_O_4_1_2; // @[Map2T.scala 17:7]
  assign O_4_2_0 = op_O_4_2_0; // @[Map2T.scala 17:7]
  assign O_4_2_1 = op_O_4_2_1; // @[Map2T.scala 17:7]
  assign O_4_2_2 = op_O_4_2_2; // @[Map2T.scala 17:7]
  assign O_5_0_0 = op_O_5_0_0; // @[Map2T.scala 17:7]
  assign O_5_0_1 = op_O_5_0_1; // @[Map2T.scala 17:7]
  assign O_5_0_2 = op_O_5_0_2; // @[Map2T.scala 17:7]
  assign O_5_1_0 = op_O_5_1_0; // @[Map2T.scala 17:7]
  assign O_5_1_1 = op_O_5_1_1; // @[Map2T.scala 17:7]
  assign O_5_1_2 = op_O_5_1_2; // @[Map2T.scala 17:7]
  assign O_5_2_0 = op_O_5_2_0; // @[Map2T.scala 17:7]
  assign O_5_2_1 = op_O_5_2_1; // @[Map2T.scala 17:7]
  assign O_5_2_2 = op_O_5_2_2; // @[Map2T.scala 17:7]
  assign O_6_0_0 = op_O_6_0_0; // @[Map2T.scala 17:7]
  assign O_6_0_1 = op_O_6_0_1; // @[Map2T.scala 17:7]
  assign O_6_0_2 = op_O_6_0_2; // @[Map2T.scala 17:7]
  assign O_6_1_0 = op_O_6_1_0; // @[Map2T.scala 17:7]
  assign O_6_1_1 = op_O_6_1_1; // @[Map2T.scala 17:7]
  assign O_6_1_2 = op_O_6_1_2; // @[Map2T.scala 17:7]
  assign O_6_2_0 = op_O_6_2_0; // @[Map2T.scala 17:7]
  assign O_6_2_1 = op_O_6_2_1; // @[Map2T.scala 17:7]
  assign O_6_2_2 = op_O_6_2_2; // @[Map2T.scala 17:7]
  assign O_7_0_0 = op_O_7_0_0; // @[Map2T.scala 17:7]
  assign O_7_0_1 = op_O_7_0_1; // @[Map2T.scala 17:7]
  assign O_7_0_2 = op_O_7_0_2; // @[Map2T.scala 17:7]
  assign O_7_1_0 = op_O_7_1_0; // @[Map2T.scala 17:7]
  assign O_7_1_1 = op_O_7_1_1; // @[Map2T.scala 17:7]
  assign O_7_1_2 = op_O_7_1_2; // @[Map2T.scala 17:7]
  assign O_7_2_0 = op_O_7_2_0; // @[Map2T.scala 17:7]
  assign O_7_2_1 = op_O_7_2_1; // @[Map2T.scala 17:7]
  assign O_7_2_2 = op_O_7_2_2; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0_0_0 = I0_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_0_0_1 = I0_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_0_0_2 = I0_0_0_2; // @[Map2T.scala 15:11]
  assign op_I0_0_1_0 = I0_0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_0_1_1 = I0_0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_0_1_2 = I0_0_1_2; // @[Map2T.scala 15:11]
  assign op_I0_1_0_0 = I0_1_0_0; // @[Map2T.scala 15:11]
  assign op_I0_1_0_1 = I0_1_0_1; // @[Map2T.scala 15:11]
  assign op_I0_1_0_2 = I0_1_0_2; // @[Map2T.scala 15:11]
  assign op_I0_1_1_0 = I0_1_1_0; // @[Map2T.scala 15:11]
  assign op_I0_1_1_1 = I0_1_1_1; // @[Map2T.scala 15:11]
  assign op_I0_1_1_2 = I0_1_1_2; // @[Map2T.scala 15:11]
  assign op_I0_2_0_0 = I0_2_0_0; // @[Map2T.scala 15:11]
  assign op_I0_2_0_1 = I0_2_0_1; // @[Map2T.scala 15:11]
  assign op_I0_2_0_2 = I0_2_0_2; // @[Map2T.scala 15:11]
  assign op_I0_2_1_0 = I0_2_1_0; // @[Map2T.scala 15:11]
  assign op_I0_2_1_1 = I0_2_1_1; // @[Map2T.scala 15:11]
  assign op_I0_2_1_2 = I0_2_1_2; // @[Map2T.scala 15:11]
  assign op_I0_3_0_0 = I0_3_0_0; // @[Map2T.scala 15:11]
  assign op_I0_3_0_1 = I0_3_0_1; // @[Map2T.scala 15:11]
  assign op_I0_3_0_2 = I0_3_0_2; // @[Map2T.scala 15:11]
  assign op_I0_3_1_0 = I0_3_1_0; // @[Map2T.scala 15:11]
  assign op_I0_3_1_1 = I0_3_1_1; // @[Map2T.scala 15:11]
  assign op_I0_3_1_2 = I0_3_1_2; // @[Map2T.scala 15:11]
  assign op_I0_4_0_0 = I0_4_0_0; // @[Map2T.scala 15:11]
  assign op_I0_4_0_1 = I0_4_0_1; // @[Map2T.scala 15:11]
  assign op_I0_4_0_2 = I0_4_0_2; // @[Map2T.scala 15:11]
  assign op_I0_4_1_0 = I0_4_1_0; // @[Map2T.scala 15:11]
  assign op_I0_4_1_1 = I0_4_1_1; // @[Map2T.scala 15:11]
  assign op_I0_4_1_2 = I0_4_1_2; // @[Map2T.scala 15:11]
  assign op_I0_5_0_0 = I0_5_0_0; // @[Map2T.scala 15:11]
  assign op_I0_5_0_1 = I0_5_0_1; // @[Map2T.scala 15:11]
  assign op_I0_5_0_2 = I0_5_0_2; // @[Map2T.scala 15:11]
  assign op_I0_5_1_0 = I0_5_1_0; // @[Map2T.scala 15:11]
  assign op_I0_5_1_1 = I0_5_1_1; // @[Map2T.scala 15:11]
  assign op_I0_5_1_2 = I0_5_1_2; // @[Map2T.scala 15:11]
  assign op_I0_6_0_0 = I0_6_0_0; // @[Map2T.scala 15:11]
  assign op_I0_6_0_1 = I0_6_0_1; // @[Map2T.scala 15:11]
  assign op_I0_6_0_2 = I0_6_0_2; // @[Map2T.scala 15:11]
  assign op_I0_6_1_0 = I0_6_1_0; // @[Map2T.scala 15:11]
  assign op_I0_6_1_1 = I0_6_1_1; // @[Map2T.scala 15:11]
  assign op_I0_6_1_2 = I0_6_1_2; // @[Map2T.scala 15:11]
  assign op_I0_7_0_0 = I0_7_0_0; // @[Map2T.scala 15:11]
  assign op_I0_7_0_1 = I0_7_0_1; // @[Map2T.scala 15:11]
  assign op_I0_7_0_2 = I0_7_0_2; // @[Map2T.scala 15:11]
  assign op_I0_7_1_0 = I0_7_1_0; // @[Map2T.scala 15:11]
  assign op_I0_7_1_1 = I0_7_1_1; // @[Map2T.scala 15:11]
  assign op_I0_7_1_2 = I0_7_1_2; // @[Map2T.scala 15:11]
  assign op_I1_0_0 = I1_0_0; // @[Map2T.scala 16:11]
  assign op_I1_0_1 = I1_0_1; // @[Map2T.scala 16:11]
  assign op_I1_0_2 = I1_0_2; // @[Map2T.scala 16:11]
  assign op_I1_1_0 = I1_1_0; // @[Map2T.scala 16:11]
  assign op_I1_1_1 = I1_1_1; // @[Map2T.scala 16:11]
  assign op_I1_1_2 = I1_1_2; // @[Map2T.scala 16:11]
  assign op_I1_2_0 = I1_2_0; // @[Map2T.scala 16:11]
  assign op_I1_2_1 = I1_2_1; // @[Map2T.scala 16:11]
  assign op_I1_2_2 = I1_2_2; // @[Map2T.scala 16:11]
  assign op_I1_3_0 = I1_3_0; // @[Map2T.scala 16:11]
  assign op_I1_3_1 = I1_3_1; // @[Map2T.scala 16:11]
  assign op_I1_3_2 = I1_3_2; // @[Map2T.scala 16:11]
  assign op_I1_4_0 = I1_4_0; // @[Map2T.scala 16:11]
  assign op_I1_4_1 = I1_4_1; // @[Map2T.scala 16:11]
  assign op_I1_4_2 = I1_4_2; // @[Map2T.scala 16:11]
  assign op_I1_5_0 = I1_5_0; // @[Map2T.scala 16:11]
  assign op_I1_5_1 = I1_5_1; // @[Map2T.scala 16:11]
  assign op_I1_5_2 = I1_5_2; // @[Map2T.scala 16:11]
  assign op_I1_6_0 = I1_6_0; // @[Map2T.scala 16:11]
  assign op_I1_6_1 = I1_6_1; // @[Map2T.scala 16:11]
  assign op_I1_6_2 = I1_6_2; // @[Map2T.scala 16:11]
  assign op_I1_7_0 = I1_7_0; // @[Map2T.scala 16:11]
  assign op_I1_7_1 = I1_7_1; // @[Map2T.scala 16:11]
  assign op_I1_7_2 = I1_7_2; // @[Map2T.scala 16:11]
endmodule
module PartitionS_3(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0_0,
  input  [31:0] I_0_0_1,
  input  [31:0] I_0_0_2,
  input  [31:0] I_0_1_0,
  input  [31:0] I_0_1_1,
  input  [31:0] I_0_1_2,
  input  [31:0] I_0_2_0,
  input  [31:0] I_0_2_1,
  input  [31:0] I_0_2_2,
  input  [31:0] I_1_0_0,
  input  [31:0] I_1_0_1,
  input  [31:0] I_1_0_2,
  input  [31:0] I_1_1_0,
  input  [31:0] I_1_1_1,
  input  [31:0] I_1_1_2,
  input  [31:0] I_1_2_0,
  input  [31:0] I_1_2_1,
  input  [31:0] I_1_2_2,
  input  [31:0] I_2_0_0,
  input  [31:0] I_2_0_1,
  input  [31:0] I_2_0_2,
  input  [31:0] I_2_1_0,
  input  [31:0] I_2_1_1,
  input  [31:0] I_2_1_2,
  input  [31:0] I_2_2_0,
  input  [31:0] I_2_2_1,
  input  [31:0] I_2_2_2,
  input  [31:0] I_3_0_0,
  input  [31:0] I_3_0_1,
  input  [31:0] I_3_0_2,
  input  [31:0] I_3_1_0,
  input  [31:0] I_3_1_1,
  input  [31:0] I_3_1_2,
  input  [31:0] I_3_2_0,
  input  [31:0] I_3_2_1,
  input  [31:0] I_3_2_2,
  input  [31:0] I_4_0_0,
  input  [31:0] I_4_0_1,
  input  [31:0] I_4_0_2,
  input  [31:0] I_4_1_0,
  input  [31:0] I_4_1_1,
  input  [31:0] I_4_1_2,
  input  [31:0] I_4_2_0,
  input  [31:0] I_4_2_1,
  input  [31:0] I_4_2_2,
  input  [31:0] I_5_0_0,
  input  [31:0] I_5_0_1,
  input  [31:0] I_5_0_2,
  input  [31:0] I_5_1_0,
  input  [31:0] I_5_1_1,
  input  [31:0] I_5_1_2,
  input  [31:0] I_5_2_0,
  input  [31:0] I_5_2_1,
  input  [31:0] I_5_2_2,
  input  [31:0] I_6_0_0,
  input  [31:0] I_6_0_1,
  input  [31:0] I_6_0_2,
  input  [31:0] I_6_1_0,
  input  [31:0] I_6_1_1,
  input  [31:0] I_6_1_2,
  input  [31:0] I_6_2_0,
  input  [31:0] I_6_2_1,
  input  [31:0] I_6_2_2,
  input  [31:0] I_7_0_0,
  input  [31:0] I_7_0_1,
  input  [31:0] I_7_0_2,
  input  [31:0] I_7_1_0,
  input  [31:0] I_7_1_1,
  input  [31:0] I_7_1_2,
  input  [31:0] I_7_2_0,
  input  [31:0] I_7_2_1,
  input  [31:0] I_7_2_2,
  output [31:0] O_0_0_0_0,
  output [31:0] O_0_0_0_1,
  output [31:0] O_0_0_0_2,
  output [31:0] O_0_0_1_0,
  output [31:0] O_0_0_1_1,
  output [31:0] O_0_0_1_2,
  output [31:0] O_0_0_2_0,
  output [31:0] O_0_0_2_1,
  output [31:0] O_0_0_2_2,
  output [31:0] O_1_0_0_0,
  output [31:0] O_1_0_0_1,
  output [31:0] O_1_0_0_2,
  output [31:0] O_1_0_1_0,
  output [31:0] O_1_0_1_1,
  output [31:0] O_1_0_1_2,
  output [31:0] O_1_0_2_0,
  output [31:0] O_1_0_2_1,
  output [31:0] O_1_0_2_2,
  output [31:0] O_2_0_0_0,
  output [31:0] O_2_0_0_1,
  output [31:0] O_2_0_0_2,
  output [31:0] O_2_0_1_0,
  output [31:0] O_2_0_1_1,
  output [31:0] O_2_0_1_2,
  output [31:0] O_2_0_2_0,
  output [31:0] O_2_0_2_1,
  output [31:0] O_2_0_2_2,
  output [31:0] O_3_0_0_0,
  output [31:0] O_3_0_0_1,
  output [31:0] O_3_0_0_2,
  output [31:0] O_3_0_1_0,
  output [31:0] O_3_0_1_1,
  output [31:0] O_3_0_1_2,
  output [31:0] O_3_0_2_0,
  output [31:0] O_3_0_2_1,
  output [31:0] O_3_0_2_2,
  output [31:0] O_4_0_0_0,
  output [31:0] O_4_0_0_1,
  output [31:0] O_4_0_0_2,
  output [31:0] O_4_0_1_0,
  output [31:0] O_4_0_1_1,
  output [31:0] O_4_0_1_2,
  output [31:0] O_4_0_2_0,
  output [31:0] O_4_0_2_1,
  output [31:0] O_4_0_2_2,
  output [31:0] O_5_0_0_0,
  output [31:0] O_5_0_0_1,
  output [31:0] O_5_0_0_2,
  output [31:0] O_5_0_1_0,
  output [31:0] O_5_0_1_1,
  output [31:0] O_5_0_1_2,
  output [31:0] O_5_0_2_0,
  output [31:0] O_5_0_2_1,
  output [31:0] O_5_0_2_2,
  output [31:0] O_6_0_0_0,
  output [31:0] O_6_0_0_1,
  output [31:0] O_6_0_0_2,
  output [31:0] O_6_0_1_0,
  output [31:0] O_6_0_1_1,
  output [31:0] O_6_0_1_2,
  output [31:0] O_6_0_2_0,
  output [31:0] O_6_0_2_1,
  output [31:0] O_6_0_2_2,
  output [31:0] O_7_0_0_0,
  output [31:0] O_7_0_0_1,
  output [31:0] O_7_0_0_2,
  output [31:0] O_7_0_1_0,
  output [31:0] O_7_0_1_1,
  output [31:0] O_7_0_1_2,
  output [31:0] O_7_0_2_0,
  output [31:0] O_7_0_2_1,
  output [31:0] O_7_0_2_2
);
  assign valid_down = valid_up; // @[Partition.scala 18:14]
  assign O_0_0_0_0 = I_0_0_0; // @[Partition.scala 15:39]
  assign O_0_0_0_1 = I_0_0_1; // @[Partition.scala 15:39]
  assign O_0_0_0_2 = I_0_0_2; // @[Partition.scala 15:39]
  assign O_0_0_1_0 = I_0_1_0; // @[Partition.scala 15:39]
  assign O_0_0_1_1 = I_0_1_1; // @[Partition.scala 15:39]
  assign O_0_0_1_2 = I_0_1_2; // @[Partition.scala 15:39]
  assign O_0_0_2_0 = I_0_2_0; // @[Partition.scala 15:39]
  assign O_0_0_2_1 = I_0_2_1; // @[Partition.scala 15:39]
  assign O_0_0_2_2 = I_0_2_2; // @[Partition.scala 15:39]
  assign O_1_0_0_0 = I_1_0_0; // @[Partition.scala 15:39]
  assign O_1_0_0_1 = I_1_0_1; // @[Partition.scala 15:39]
  assign O_1_0_0_2 = I_1_0_2; // @[Partition.scala 15:39]
  assign O_1_0_1_0 = I_1_1_0; // @[Partition.scala 15:39]
  assign O_1_0_1_1 = I_1_1_1; // @[Partition.scala 15:39]
  assign O_1_0_1_2 = I_1_1_2; // @[Partition.scala 15:39]
  assign O_1_0_2_0 = I_1_2_0; // @[Partition.scala 15:39]
  assign O_1_0_2_1 = I_1_2_1; // @[Partition.scala 15:39]
  assign O_1_0_2_2 = I_1_2_2; // @[Partition.scala 15:39]
  assign O_2_0_0_0 = I_2_0_0; // @[Partition.scala 15:39]
  assign O_2_0_0_1 = I_2_0_1; // @[Partition.scala 15:39]
  assign O_2_0_0_2 = I_2_0_2; // @[Partition.scala 15:39]
  assign O_2_0_1_0 = I_2_1_0; // @[Partition.scala 15:39]
  assign O_2_0_1_1 = I_2_1_1; // @[Partition.scala 15:39]
  assign O_2_0_1_2 = I_2_1_2; // @[Partition.scala 15:39]
  assign O_2_0_2_0 = I_2_2_0; // @[Partition.scala 15:39]
  assign O_2_0_2_1 = I_2_2_1; // @[Partition.scala 15:39]
  assign O_2_0_2_2 = I_2_2_2; // @[Partition.scala 15:39]
  assign O_3_0_0_0 = I_3_0_0; // @[Partition.scala 15:39]
  assign O_3_0_0_1 = I_3_0_1; // @[Partition.scala 15:39]
  assign O_3_0_0_2 = I_3_0_2; // @[Partition.scala 15:39]
  assign O_3_0_1_0 = I_3_1_0; // @[Partition.scala 15:39]
  assign O_3_0_1_1 = I_3_1_1; // @[Partition.scala 15:39]
  assign O_3_0_1_2 = I_3_1_2; // @[Partition.scala 15:39]
  assign O_3_0_2_0 = I_3_2_0; // @[Partition.scala 15:39]
  assign O_3_0_2_1 = I_3_2_1; // @[Partition.scala 15:39]
  assign O_3_0_2_2 = I_3_2_2; // @[Partition.scala 15:39]
  assign O_4_0_0_0 = I_4_0_0; // @[Partition.scala 15:39]
  assign O_4_0_0_1 = I_4_0_1; // @[Partition.scala 15:39]
  assign O_4_0_0_2 = I_4_0_2; // @[Partition.scala 15:39]
  assign O_4_0_1_0 = I_4_1_0; // @[Partition.scala 15:39]
  assign O_4_0_1_1 = I_4_1_1; // @[Partition.scala 15:39]
  assign O_4_0_1_2 = I_4_1_2; // @[Partition.scala 15:39]
  assign O_4_0_2_0 = I_4_2_0; // @[Partition.scala 15:39]
  assign O_4_0_2_1 = I_4_2_1; // @[Partition.scala 15:39]
  assign O_4_0_2_2 = I_4_2_2; // @[Partition.scala 15:39]
  assign O_5_0_0_0 = I_5_0_0; // @[Partition.scala 15:39]
  assign O_5_0_0_1 = I_5_0_1; // @[Partition.scala 15:39]
  assign O_5_0_0_2 = I_5_0_2; // @[Partition.scala 15:39]
  assign O_5_0_1_0 = I_5_1_0; // @[Partition.scala 15:39]
  assign O_5_0_1_1 = I_5_1_1; // @[Partition.scala 15:39]
  assign O_5_0_1_2 = I_5_1_2; // @[Partition.scala 15:39]
  assign O_5_0_2_0 = I_5_2_0; // @[Partition.scala 15:39]
  assign O_5_0_2_1 = I_5_2_1; // @[Partition.scala 15:39]
  assign O_5_0_2_2 = I_5_2_2; // @[Partition.scala 15:39]
  assign O_6_0_0_0 = I_6_0_0; // @[Partition.scala 15:39]
  assign O_6_0_0_1 = I_6_0_1; // @[Partition.scala 15:39]
  assign O_6_0_0_2 = I_6_0_2; // @[Partition.scala 15:39]
  assign O_6_0_1_0 = I_6_1_0; // @[Partition.scala 15:39]
  assign O_6_0_1_1 = I_6_1_1; // @[Partition.scala 15:39]
  assign O_6_0_1_2 = I_6_1_2; // @[Partition.scala 15:39]
  assign O_6_0_2_0 = I_6_2_0; // @[Partition.scala 15:39]
  assign O_6_0_2_1 = I_6_2_1; // @[Partition.scala 15:39]
  assign O_6_0_2_2 = I_6_2_2; // @[Partition.scala 15:39]
  assign O_7_0_0_0 = I_7_0_0; // @[Partition.scala 15:39]
  assign O_7_0_0_1 = I_7_0_1; // @[Partition.scala 15:39]
  assign O_7_0_0_2 = I_7_0_2; // @[Partition.scala 15:39]
  assign O_7_0_1_0 = I_7_1_0; // @[Partition.scala 15:39]
  assign O_7_0_1_1 = I_7_1_1; // @[Partition.scala 15:39]
  assign O_7_0_1_2 = I_7_1_2; // @[Partition.scala 15:39]
  assign O_7_0_2_0 = I_7_2_0; // @[Partition.scala 15:39]
  assign O_7_0_2_1 = I_7_2_1; // @[Partition.scala 15:39]
  assign O_7_0_2_2 = I_7_2_2; // @[Partition.scala 15:39]
endmodule
module MapT_6(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0_0,
  input  [31:0] I_0_0_1,
  input  [31:0] I_0_0_2,
  input  [31:0] I_0_1_0,
  input  [31:0] I_0_1_1,
  input  [31:0] I_0_1_2,
  input  [31:0] I_0_2_0,
  input  [31:0] I_0_2_1,
  input  [31:0] I_0_2_2,
  input  [31:0] I_1_0_0,
  input  [31:0] I_1_0_1,
  input  [31:0] I_1_0_2,
  input  [31:0] I_1_1_0,
  input  [31:0] I_1_1_1,
  input  [31:0] I_1_1_2,
  input  [31:0] I_1_2_0,
  input  [31:0] I_1_2_1,
  input  [31:0] I_1_2_2,
  input  [31:0] I_2_0_0,
  input  [31:0] I_2_0_1,
  input  [31:0] I_2_0_2,
  input  [31:0] I_2_1_0,
  input  [31:0] I_2_1_1,
  input  [31:0] I_2_1_2,
  input  [31:0] I_2_2_0,
  input  [31:0] I_2_2_1,
  input  [31:0] I_2_2_2,
  input  [31:0] I_3_0_0,
  input  [31:0] I_3_0_1,
  input  [31:0] I_3_0_2,
  input  [31:0] I_3_1_0,
  input  [31:0] I_3_1_1,
  input  [31:0] I_3_1_2,
  input  [31:0] I_3_2_0,
  input  [31:0] I_3_2_1,
  input  [31:0] I_3_2_2,
  input  [31:0] I_4_0_0,
  input  [31:0] I_4_0_1,
  input  [31:0] I_4_0_2,
  input  [31:0] I_4_1_0,
  input  [31:0] I_4_1_1,
  input  [31:0] I_4_1_2,
  input  [31:0] I_4_2_0,
  input  [31:0] I_4_2_1,
  input  [31:0] I_4_2_2,
  input  [31:0] I_5_0_0,
  input  [31:0] I_5_0_1,
  input  [31:0] I_5_0_2,
  input  [31:0] I_5_1_0,
  input  [31:0] I_5_1_1,
  input  [31:0] I_5_1_2,
  input  [31:0] I_5_2_0,
  input  [31:0] I_5_2_1,
  input  [31:0] I_5_2_2,
  input  [31:0] I_6_0_0,
  input  [31:0] I_6_0_1,
  input  [31:0] I_6_0_2,
  input  [31:0] I_6_1_0,
  input  [31:0] I_6_1_1,
  input  [31:0] I_6_1_2,
  input  [31:0] I_6_2_0,
  input  [31:0] I_6_2_1,
  input  [31:0] I_6_2_2,
  input  [31:0] I_7_0_0,
  input  [31:0] I_7_0_1,
  input  [31:0] I_7_0_2,
  input  [31:0] I_7_1_0,
  input  [31:0] I_7_1_1,
  input  [31:0] I_7_1_2,
  input  [31:0] I_7_2_0,
  input  [31:0] I_7_2_1,
  input  [31:0] I_7_2_2,
  output [31:0] O_0_0_0_0,
  output [31:0] O_0_0_0_1,
  output [31:0] O_0_0_0_2,
  output [31:0] O_0_0_1_0,
  output [31:0] O_0_0_1_1,
  output [31:0] O_0_0_1_2,
  output [31:0] O_0_0_2_0,
  output [31:0] O_0_0_2_1,
  output [31:0] O_0_0_2_2,
  output [31:0] O_1_0_0_0,
  output [31:0] O_1_0_0_1,
  output [31:0] O_1_0_0_2,
  output [31:0] O_1_0_1_0,
  output [31:0] O_1_0_1_1,
  output [31:0] O_1_0_1_2,
  output [31:0] O_1_0_2_0,
  output [31:0] O_1_0_2_1,
  output [31:0] O_1_0_2_2,
  output [31:0] O_2_0_0_0,
  output [31:0] O_2_0_0_1,
  output [31:0] O_2_0_0_2,
  output [31:0] O_2_0_1_0,
  output [31:0] O_2_0_1_1,
  output [31:0] O_2_0_1_2,
  output [31:0] O_2_0_2_0,
  output [31:0] O_2_0_2_1,
  output [31:0] O_2_0_2_2,
  output [31:0] O_3_0_0_0,
  output [31:0] O_3_0_0_1,
  output [31:0] O_3_0_0_2,
  output [31:0] O_3_0_1_0,
  output [31:0] O_3_0_1_1,
  output [31:0] O_3_0_1_2,
  output [31:0] O_3_0_2_0,
  output [31:0] O_3_0_2_1,
  output [31:0] O_3_0_2_2,
  output [31:0] O_4_0_0_0,
  output [31:0] O_4_0_0_1,
  output [31:0] O_4_0_0_2,
  output [31:0] O_4_0_1_0,
  output [31:0] O_4_0_1_1,
  output [31:0] O_4_0_1_2,
  output [31:0] O_4_0_2_0,
  output [31:0] O_4_0_2_1,
  output [31:0] O_4_0_2_2,
  output [31:0] O_5_0_0_0,
  output [31:0] O_5_0_0_1,
  output [31:0] O_5_0_0_2,
  output [31:0] O_5_0_1_0,
  output [31:0] O_5_0_1_1,
  output [31:0] O_5_0_1_2,
  output [31:0] O_5_0_2_0,
  output [31:0] O_5_0_2_1,
  output [31:0] O_5_0_2_2,
  output [31:0] O_6_0_0_0,
  output [31:0] O_6_0_0_1,
  output [31:0] O_6_0_0_2,
  output [31:0] O_6_0_1_0,
  output [31:0] O_6_0_1_1,
  output [31:0] O_6_0_1_2,
  output [31:0] O_6_0_2_0,
  output [31:0] O_6_0_2_1,
  output [31:0] O_6_0_2_2,
  output [31:0] O_7_0_0_0,
  output [31:0] O_7_0_0_1,
  output [31:0] O_7_0_0_2,
  output [31:0] O_7_0_1_0,
  output [31:0] O_7_0_1_1,
  output [31:0] O_7_0_1_2,
  output [31:0] O_7_0_2_0,
  output [31:0] O_7_0_2_1,
  output [31:0] O_7_0_2_2
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_0_2_2; // @[MapT.scala 8:20]
  PartitionS_3 op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0(op_I_0_0_0),
    .I_0_0_1(op_I_0_0_1),
    .I_0_0_2(op_I_0_0_2),
    .I_0_1_0(op_I_0_1_0),
    .I_0_1_1(op_I_0_1_1),
    .I_0_1_2(op_I_0_1_2),
    .I_0_2_0(op_I_0_2_0),
    .I_0_2_1(op_I_0_2_1),
    .I_0_2_2(op_I_0_2_2),
    .I_1_0_0(op_I_1_0_0),
    .I_1_0_1(op_I_1_0_1),
    .I_1_0_2(op_I_1_0_2),
    .I_1_1_0(op_I_1_1_0),
    .I_1_1_1(op_I_1_1_1),
    .I_1_1_2(op_I_1_1_2),
    .I_1_2_0(op_I_1_2_0),
    .I_1_2_1(op_I_1_2_1),
    .I_1_2_2(op_I_1_2_2),
    .I_2_0_0(op_I_2_0_0),
    .I_2_0_1(op_I_2_0_1),
    .I_2_0_2(op_I_2_0_2),
    .I_2_1_0(op_I_2_1_0),
    .I_2_1_1(op_I_2_1_1),
    .I_2_1_2(op_I_2_1_2),
    .I_2_2_0(op_I_2_2_0),
    .I_2_2_1(op_I_2_2_1),
    .I_2_2_2(op_I_2_2_2),
    .I_3_0_0(op_I_3_0_0),
    .I_3_0_1(op_I_3_0_1),
    .I_3_0_2(op_I_3_0_2),
    .I_3_1_0(op_I_3_1_0),
    .I_3_1_1(op_I_3_1_1),
    .I_3_1_2(op_I_3_1_2),
    .I_3_2_0(op_I_3_2_0),
    .I_3_2_1(op_I_3_2_1),
    .I_3_2_2(op_I_3_2_2),
    .I_4_0_0(op_I_4_0_0),
    .I_4_0_1(op_I_4_0_1),
    .I_4_0_2(op_I_4_0_2),
    .I_4_1_0(op_I_4_1_0),
    .I_4_1_1(op_I_4_1_1),
    .I_4_1_2(op_I_4_1_2),
    .I_4_2_0(op_I_4_2_0),
    .I_4_2_1(op_I_4_2_1),
    .I_4_2_2(op_I_4_2_2),
    .I_5_0_0(op_I_5_0_0),
    .I_5_0_1(op_I_5_0_1),
    .I_5_0_2(op_I_5_0_2),
    .I_5_1_0(op_I_5_1_0),
    .I_5_1_1(op_I_5_1_1),
    .I_5_1_2(op_I_5_1_2),
    .I_5_2_0(op_I_5_2_0),
    .I_5_2_1(op_I_5_2_1),
    .I_5_2_2(op_I_5_2_2),
    .I_6_0_0(op_I_6_0_0),
    .I_6_0_1(op_I_6_0_1),
    .I_6_0_2(op_I_6_0_2),
    .I_6_1_0(op_I_6_1_0),
    .I_6_1_1(op_I_6_1_1),
    .I_6_1_2(op_I_6_1_2),
    .I_6_2_0(op_I_6_2_0),
    .I_6_2_1(op_I_6_2_1),
    .I_6_2_2(op_I_6_2_2),
    .I_7_0_0(op_I_7_0_0),
    .I_7_0_1(op_I_7_0_1),
    .I_7_0_2(op_I_7_0_2),
    .I_7_1_0(op_I_7_1_0),
    .I_7_1_1(op_I_7_1_1),
    .I_7_1_2(op_I_7_1_2),
    .I_7_2_0(op_I_7_2_0),
    .I_7_2_1(op_I_7_2_1),
    .I_7_2_2(op_I_7_2_2),
    .O_0_0_0_0(op_O_0_0_0_0),
    .O_0_0_0_1(op_O_0_0_0_1),
    .O_0_0_0_2(op_O_0_0_0_2),
    .O_0_0_1_0(op_O_0_0_1_0),
    .O_0_0_1_1(op_O_0_0_1_1),
    .O_0_0_1_2(op_O_0_0_1_2),
    .O_0_0_2_0(op_O_0_0_2_0),
    .O_0_0_2_1(op_O_0_0_2_1),
    .O_0_0_2_2(op_O_0_0_2_2),
    .O_1_0_0_0(op_O_1_0_0_0),
    .O_1_0_0_1(op_O_1_0_0_1),
    .O_1_0_0_2(op_O_1_0_0_2),
    .O_1_0_1_0(op_O_1_0_1_0),
    .O_1_0_1_1(op_O_1_0_1_1),
    .O_1_0_1_2(op_O_1_0_1_2),
    .O_1_0_2_0(op_O_1_0_2_0),
    .O_1_0_2_1(op_O_1_0_2_1),
    .O_1_0_2_2(op_O_1_0_2_2),
    .O_2_0_0_0(op_O_2_0_0_0),
    .O_2_0_0_1(op_O_2_0_0_1),
    .O_2_0_0_2(op_O_2_0_0_2),
    .O_2_0_1_0(op_O_2_0_1_0),
    .O_2_0_1_1(op_O_2_0_1_1),
    .O_2_0_1_2(op_O_2_0_1_2),
    .O_2_0_2_0(op_O_2_0_2_0),
    .O_2_0_2_1(op_O_2_0_2_1),
    .O_2_0_2_2(op_O_2_0_2_2),
    .O_3_0_0_0(op_O_3_0_0_0),
    .O_3_0_0_1(op_O_3_0_0_1),
    .O_3_0_0_2(op_O_3_0_0_2),
    .O_3_0_1_0(op_O_3_0_1_0),
    .O_3_0_1_1(op_O_3_0_1_1),
    .O_3_0_1_2(op_O_3_0_1_2),
    .O_3_0_2_0(op_O_3_0_2_0),
    .O_3_0_2_1(op_O_3_0_2_1),
    .O_3_0_2_2(op_O_3_0_2_2),
    .O_4_0_0_0(op_O_4_0_0_0),
    .O_4_0_0_1(op_O_4_0_0_1),
    .O_4_0_0_2(op_O_4_0_0_2),
    .O_4_0_1_0(op_O_4_0_1_0),
    .O_4_0_1_1(op_O_4_0_1_1),
    .O_4_0_1_2(op_O_4_0_1_2),
    .O_4_0_2_0(op_O_4_0_2_0),
    .O_4_0_2_1(op_O_4_0_2_1),
    .O_4_0_2_2(op_O_4_0_2_2),
    .O_5_0_0_0(op_O_5_0_0_0),
    .O_5_0_0_1(op_O_5_0_0_1),
    .O_5_0_0_2(op_O_5_0_0_2),
    .O_5_0_1_0(op_O_5_0_1_0),
    .O_5_0_1_1(op_O_5_0_1_1),
    .O_5_0_1_2(op_O_5_0_1_2),
    .O_5_0_2_0(op_O_5_0_2_0),
    .O_5_0_2_1(op_O_5_0_2_1),
    .O_5_0_2_2(op_O_5_0_2_2),
    .O_6_0_0_0(op_O_6_0_0_0),
    .O_6_0_0_1(op_O_6_0_0_1),
    .O_6_0_0_2(op_O_6_0_0_2),
    .O_6_0_1_0(op_O_6_0_1_0),
    .O_6_0_1_1(op_O_6_0_1_1),
    .O_6_0_1_2(op_O_6_0_1_2),
    .O_6_0_2_0(op_O_6_0_2_0),
    .O_6_0_2_1(op_O_6_0_2_1),
    .O_6_0_2_2(op_O_6_0_2_2),
    .O_7_0_0_0(op_O_7_0_0_0),
    .O_7_0_0_1(op_O_7_0_0_1),
    .O_7_0_0_2(op_O_7_0_0_2),
    .O_7_0_1_0(op_O_7_0_1_0),
    .O_7_0_1_1(op_O_7_0_1_1),
    .O_7_0_1_2(op_O_7_0_1_2),
    .O_7_0_2_0(op_O_7_0_2_0),
    .O_7_0_2_1(op_O_7_0_2_1),
    .O_7_0_2_2(op_O_7_0_2_2)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0_0 = op_O_0_0_0_0; // @[MapT.scala 15:7]
  assign O_0_0_0_1 = op_O_0_0_0_1; // @[MapT.scala 15:7]
  assign O_0_0_0_2 = op_O_0_0_0_2; // @[MapT.scala 15:7]
  assign O_0_0_1_0 = op_O_0_0_1_0; // @[MapT.scala 15:7]
  assign O_0_0_1_1 = op_O_0_0_1_1; // @[MapT.scala 15:7]
  assign O_0_0_1_2 = op_O_0_0_1_2; // @[MapT.scala 15:7]
  assign O_0_0_2_0 = op_O_0_0_2_0; // @[MapT.scala 15:7]
  assign O_0_0_2_1 = op_O_0_0_2_1; // @[MapT.scala 15:7]
  assign O_0_0_2_2 = op_O_0_0_2_2; // @[MapT.scala 15:7]
  assign O_1_0_0_0 = op_O_1_0_0_0; // @[MapT.scala 15:7]
  assign O_1_0_0_1 = op_O_1_0_0_1; // @[MapT.scala 15:7]
  assign O_1_0_0_2 = op_O_1_0_0_2; // @[MapT.scala 15:7]
  assign O_1_0_1_0 = op_O_1_0_1_0; // @[MapT.scala 15:7]
  assign O_1_0_1_1 = op_O_1_0_1_1; // @[MapT.scala 15:7]
  assign O_1_0_1_2 = op_O_1_0_1_2; // @[MapT.scala 15:7]
  assign O_1_0_2_0 = op_O_1_0_2_0; // @[MapT.scala 15:7]
  assign O_1_0_2_1 = op_O_1_0_2_1; // @[MapT.scala 15:7]
  assign O_1_0_2_2 = op_O_1_0_2_2; // @[MapT.scala 15:7]
  assign O_2_0_0_0 = op_O_2_0_0_0; // @[MapT.scala 15:7]
  assign O_2_0_0_1 = op_O_2_0_0_1; // @[MapT.scala 15:7]
  assign O_2_0_0_2 = op_O_2_0_0_2; // @[MapT.scala 15:7]
  assign O_2_0_1_0 = op_O_2_0_1_0; // @[MapT.scala 15:7]
  assign O_2_0_1_1 = op_O_2_0_1_1; // @[MapT.scala 15:7]
  assign O_2_0_1_2 = op_O_2_0_1_2; // @[MapT.scala 15:7]
  assign O_2_0_2_0 = op_O_2_0_2_0; // @[MapT.scala 15:7]
  assign O_2_0_2_1 = op_O_2_0_2_1; // @[MapT.scala 15:7]
  assign O_2_0_2_2 = op_O_2_0_2_2; // @[MapT.scala 15:7]
  assign O_3_0_0_0 = op_O_3_0_0_0; // @[MapT.scala 15:7]
  assign O_3_0_0_1 = op_O_3_0_0_1; // @[MapT.scala 15:7]
  assign O_3_0_0_2 = op_O_3_0_0_2; // @[MapT.scala 15:7]
  assign O_3_0_1_0 = op_O_3_0_1_0; // @[MapT.scala 15:7]
  assign O_3_0_1_1 = op_O_3_0_1_1; // @[MapT.scala 15:7]
  assign O_3_0_1_2 = op_O_3_0_1_2; // @[MapT.scala 15:7]
  assign O_3_0_2_0 = op_O_3_0_2_0; // @[MapT.scala 15:7]
  assign O_3_0_2_1 = op_O_3_0_2_1; // @[MapT.scala 15:7]
  assign O_3_0_2_2 = op_O_3_0_2_2; // @[MapT.scala 15:7]
  assign O_4_0_0_0 = op_O_4_0_0_0; // @[MapT.scala 15:7]
  assign O_4_0_0_1 = op_O_4_0_0_1; // @[MapT.scala 15:7]
  assign O_4_0_0_2 = op_O_4_0_0_2; // @[MapT.scala 15:7]
  assign O_4_0_1_0 = op_O_4_0_1_0; // @[MapT.scala 15:7]
  assign O_4_0_1_1 = op_O_4_0_1_1; // @[MapT.scala 15:7]
  assign O_4_0_1_2 = op_O_4_0_1_2; // @[MapT.scala 15:7]
  assign O_4_0_2_0 = op_O_4_0_2_0; // @[MapT.scala 15:7]
  assign O_4_0_2_1 = op_O_4_0_2_1; // @[MapT.scala 15:7]
  assign O_4_0_2_2 = op_O_4_0_2_2; // @[MapT.scala 15:7]
  assign O_5_0_0_0 = op_O_5_0_0_0; // @[MapT.scala 15:7]
  assign O_5_0_0_1 = op_O_5_0_0_1; // @[MapT.scala 15:7]
  assign O_5_0_0_2 = op_O_5_0_0_2; // @[MapT.scala 15:7]
  assign O_5_0_1_0 = op_O_5_0_1_0; // @[MapT.scala 15:7]
  assign O_5_0_1_1 = op_O_5_0_1_1; // @[MapT.scala 15:7]
  assign O_5_0_1_2 = op_O_5_0_1_2; // @[MapT.scala 15:7]
  assign O_5_0_2_0 = op_O_5_0_2_0; // @[MapT.scala 15:7]
  assign O_5_0_2_1 = op_O_5_0_2_1; // @[MapT.scala 15:7]
  assign O_5_0_2_2 = op_O_5_0_2_2; // @[MapT.scala 15:7]
  assign O_6_0_0_0 = op_O_6_0_0_0; // @[MapT.scala 15:7]
  assign O_6_0_0_1 = op_O_6_0_0_1; // @[MapT.scala 15:7]
  assign O_6_0_0_2 = op_O_6_0_0_2; // @[MapT.scala 15:7]
  assign O_6_0_1_0 = op_O_6_0_1_0; // @[MapT.scala 15:7]
  assign O_6_0_1_1 = op_O_6_0_1_1; // @[MapT.scala 15:7]
  assign O_6_0_1_2 = op_O_6_0_1_2; // @[MapT.scala 15:7]
  assign O_6_0_2_0 = op_O_6_0_2_0; // @[MapT.scala 15:7]
  assign O_6_0_2_1 = op_O_6_0_2_1; // @[MapT.scala 15:7]
  assign O_6_0_2_2 = op_O_6_0_2_2; // @[MapT.scala 15:7]
  assign O_7_0_0_0 = op_O_7_0_0_0; // @[MapT.scala 15:7]
  assign O_7_0_0_1 = op_O_7_0_0_1; // @[MapT.scala 15:7]
  assign O_7_0_0_2 = op_O_7_0_0_2; // @[MapT.scala 15:7]
  assign O_7_0_1_0 = op_O_7_0_1_0; // @[MapT.scala 15:7]
  assign O_7_0_1_1 = op_O_7_0_1_1; // @[MapT.scala 15:7]
  assign O_7_0_1_2 = op_O_7_0_1_2; // @[MapT.scala 15:7]
  assign O_7_0_2_0 = op_O_7_0_2_0; // @[MapT.scala 15:7]
  assign O_7_0_2_1 = op_O_7_0_2_1; // @[MapT.scala 15:7]
  assign O_7_0_2_2 = op_O_7_0_2_2; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0 = I_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_1 = I_0_0_1; // @[MapT.scala 14:10]
  assign op_I_0_0_2 = I_0_0_2; // @[MapT.scala 14:10]
  assign op_I_0_1_0 = I_0_1_0; // @[MapT.scala 14:10]
  assign op_I_0_1_1 = I_0_1_1; // @[MapT.scala 14:10]
  assign op_I_0_1_2 = I_0_1_2; // @[MapT.scala 14:10]
  assign op_I_0_2_0 = I_0_2_0; // @[MapT.scala 14:10]
  assign op_I_0_2_1 = I_0_2_1; // @[MapT.scala 14:10]
  assign op_I_0_2_2 = I_0_2_2; // @[MapT.scala 14:10]
  assign op_I_1_0_0 = I_1_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_1 = I_1_0_1; // @[MapT.scala 14:10]
  assign op_I_1_0_2 = I_1_0_2; // @[MapT.scala 14:10]
  assign op_I_1_1_0 = I_1_1_0; // @[MapT.scala 14:10]
  assign op_I_1_1_1 = I_1_1_1; // @[MapT.scala 14:10]
  assign op_I_1_1_2 = I_1_1_2; // @[MapT.scala 14:10]
  assign op_I_1_2_0 = I_1_2_0; // @[MapT.scala 14:10]
  assign op_I_1_2_1 = I_1_2_1; // @[MapT.scala 14:10]
  assign op_I_1_2_2 = I_1_2_2; // @[MapT.scala 14:10]
  assign op_I_2_0_0 = I_2_0_0; // @[MapT.scala 14:10]
  assign op_I_2_0_1 = I_2_0_1; // @[MapT.scala 14:10]
  assign op_I_2_0_2 = I_2_0_2; // @[MapT.scala 14:10]
  assign op_I_2_1_0 = I_2_1_0; // @[MapT.scala 14:10]
  assign op_I_2_1_1 = I_2_1_1; // @[MapT.scala 14:10]
  assign op_I_2_1_2 = I_2_1_2; // @[MapT.scala 14:10]
  assign op_I_2_2_0 = I_2_2_0; // @[MapT.scala 14:10]
  assign op_I_2_2_1 = I_2_2_1; // @[MapT.scala 14:10]
  assign op_I_2_2_2 = I_2_2_2; // @[MapT.scala 14:10]
  assign op_I_3_0_0 = I_3_0_0; // @[MapT.scala 14:10]
  assign op_I_3_0_1 = I_3_0_1; // @[MapT.scala 14:10]
  assign op_I_3_0_2 = I_3_0_2; // @[MapT.scala 14:10]
  assign op_I_3_1_0 = I_3_1_0; // @[MapT.scala 14:10]
  assign op_I_3_1_1 = I_3_1_1; // @[MapT.scala 14:10]
  assign op_I_3_1_2 = I_3_1_2; // @[MapT.scala 14:10]
  assign op_I_3_2_0 = I_3_2_0; // @[MapT.scala 14:10]
  assign op_I_3_2_1 = I_3_2_1; // @[MapT.scala 14:10]
  assign op_I_3_2_2 = I_3_2_2; // @[MapT.scala 14:10]
  assign op_I_4_0_0 = I_4_0_0; // @[MapT.scala 14:10]
  assign op_I_4_0_1 = I_4_0_1; // @[MapT.scala 14:10]
  assign op_I_4_0_2 = I_4_0_2; // @[MapT.scala 14:10]
  assign op_I_4_1_0 = I_4_1_0; // @[MapT.scala 14:10]
  assign op_I_4_1_1 = I_4_1_1; // @[MapT.scala 14:10]
  assign op_I_4_1_2 = I_4_1_2; // @[MapT.scala 14:10]
  assign op_I_4_2_0 = I_4_2_0; // @[MapT.scala 14:10]
  assign op_I_4_2_1 = I_4_2_1; // @[MapT.scala 14:10]
  assign op_I_4_2_2 = I_4_2_2; // @[MapT.scala 14:10]
  assign op_I_5_0_0 = I_5_0_0; // @[MapT.scala 14:10]
  assign op_I_5_0_1 = I_5_0_1; // @[MapT.scala 14:10]
  assign op_I_5_0_2 = I_5_0_2; // @[MapT.scala 14:10]
  assign op_I_5_1_0 = I_5_1_0; // @[MapT.scala 14:10]
  assign op_I_5_1_1 = I_5_1_1; // @[MapT.scala 14:10]
  assign op_I_5_1_2 = I_5_1_2; // @[MapT.scala 14:10]
  assign op_I_5_2_0 = I_5_2_0; // @[MapT.scala 14:10]
  assign op_I_5_2_1 = I_5_2_1; // @[MapT.scala 14:10]
  assign op_I_5_2_2 = I_5_2_2; // @[MapT.scala 14:10]
  assign op_I_6_0_0 = I_6_0_0; // @[MapT.scala 14:10]
  assign op_I_6_0_1 = I_6_0_1; // @[MapT.scala 14:10]
  assign op_I_6_0_2 = I_6_0_2; // @[MapT.scala 14:10]
  assign op_I_6_1_0 = I_6_1_0; // @[MapT.scala 14:10]
  assign op_I_6_1_1 = I_6_1_1; // @[MapT.scala 14:10]
  assign op_I_6_1_2 = I_6_1_2; // @[MapT.scala 14:10]
  assign op_I_6_2_0 = I_6_2_0; // @[MapT.scala 14:10]
  assign op_I_6_2_1 = I_6_2_1; // @[MapT.scala 14:10]
  assign op_I_6_2_2 = I_6_2_2; // @[MapT.scala 14:10]
  assign op_I_7_0_0 = I_7_0_0; // @[MapT.scala 14:10]
  assign op_I_7_0_1 = I_7_0_1; // @[MapT.scala 14:10]
  assign op_I_7_0_2 = I_7_0_2; // @[MapT.scala 14:10]
  assign op_I_7_1_0 = I_7_1_0; // @[MapT.scala 14:10]
  assign op_I_7_1_1 = I_7_1_1; // @[MapT.scala 14:10]
  assign op_I_7_1_2 = I_7_1_2; // @[MapT.scala 14:10]
  assign op_I_7_2_0 = I_7_2_0; // @[MapT.scala 14:10]
  assign op_I_7_2_1 = I_7_2_1; // @[MapT.scala 14:10]
  assign op_I_7_2_2 = I_7_2_2; // @[MapT.scala 14:10]
endmodule
module SSeqTupleToSSeq_3(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0,
  input  [31:0] I_0_1,
  input  [31:0] I_0_2,
  input  [31:0] I_1_0,
  input  [31:0] I_1_1,
  input  [31:0] I_1_2,
  input  [31:0] I_2_0,
  input  [31:0] I_2_1,
  input  [31:0] I_2_2,
  output [31:0] O_0_0,
  output [31:0] O_0_1,
  output [31:0] O_0_2,
  output [31:0] O_1_0,
  output [31:0] O_1_1,
  output [31:0] O_1_2,
  output [31:0] O_2_0,
  output [31:0] O_2_1,
  output [31:0] O_2_2
);
  assign valid_down = valid_up; // @[Tuple.scala 42:14]
  assign O_0_0 = I_0_0; // @[Tuple.scala 41:5]
  assign O_0_1 = I_0_1; // @[Tuple.scala 41:5]
  assign O_0_2 = I_0_2; // @[Tuple.scala 41:5]
  assign O_1_0 = I_1_0; // @[Tuple.scala 41:5]
  assign O_1_1 = I_1_1; // @[Tuple.scala 41:5]
  assign O_1_2 = I_1_2; // @[Tuple.scala 41:5]
  assign O_2_0 = I_2_0; // @[Tuple.scala 41:5]
  assign O_2_1 = I_2_1; // @[Tuple.scala 41:5]
  assign O_2_2 = I_2_2; // @[Tuple.scala 41:5]
endmodule
module Remove1S_3(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0_0,
  input  [31:0] I_0_0_1,
  input  [31:0] I_0_0_2,
  input  [31:0] I_0_1_0,
  input  [31:0] I_0_1_1,
  input  [31:0] I_0_1_2,
  input  [31:0] I_0_2_0,
  input  [31:0] I_0_2_1,
  input  [31:0] I_0_2_2,
  output [31:0] O_0_0,
  output [31:0] O_0_1,
  output [31:0] O_0_2,
  output [31:0] O_1_0,
  output [31:0] O_1_1,
  output [31:0] O_1_2,
  output [31:0] O_2_0,
  output [31:0] O_2_1,
  output [31:0] O_2_2
);
  wire  op_inst_valid_up; // @[Remove1S.scala 9:23]
  wire  op_inst_valid_down; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_I_0_0; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_I_0_1; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_I_0_2; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_I_1_0; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_I_1_1; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_I_1_2; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_I_2_0; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_I_2_1; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_I_2_2; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_O_0_0; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_O_0_1; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_O_0_2; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_O_1_0; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_O_1_1; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_O_1_2; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_O_2_0; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_O_2_1; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_O_2_2; // @[Remove1S.scala 9:23]
  SSeqTupleToSSeq_3 op_inst ( // @[Remove1S.scala 9:23]
    .valid_up(op_inst_valid_up),
    .valid_down(op_inst_valid_down),
    .I_0_0(op_inst_I_0_0),
    .I_0_1(op_inst_I_0_1),
    .I_0_2(op_inst_I_0_2),
    .I_1_0(op_inst_I_1_0),
    .I_1_1(op_inst_I_1_1),
    .I_1_2(op_inst_I_1_2),
    .I_2_0(op_inst_I_2_0),
    .I_2_1(op_inst_I_2_1),
    .I_2_2(op_inst_I_2_2),
    .O_0_0(op_inst_O_0_0),
    .O_0_1(op_inst_O_0_1),
    .O_0_2(op_inst_O_0_2),
    .O_1_0(op_inst_O_1_0),
    .O_1_1(op_inst_O_1_1),
    .O_1_2(op_inst_O_1_2),
    .O_2_0(op_inst_O_2_0),
    .O_2_1(op_inst_O_2_1),
    .O_2_2(op_inst_O_2_2)
  );
  assign valid_down = op_inst_valid_down; // @[Remove1S.scala 16:14]
  assign O_0_0 = op_inst_O_0_0; // @[Remove1S.scala 14:5]
  assign O_0_1 = op_inst_O_0_1; // @[Remove1S.scala 14:5]
  assign O_0_2 = op_inst_O_0_2; // @[Remove1S.scala 14:5]
  assign O_1_0 = op_inst_O_1_0; // @[Remove1S.scala 14:5]
  assign O_1_1 = op_inst_O_1_1; // @[Remove1S.scala 14:5]
  assign O_1_2 = op_inst_O_1_2; // @[Remove1S.scala 14:5]
  assign O_2_0 = op_inst_O_2_0; // @[Remove1S.scala 14:5]
  assign O_2_1 = op_inst_O_2_1; // @[Remove1S.scala 14:5]
  assign O_2_2 = op_inst_O_2_2; // @[Remove1S.scala 14:5]
  assign op_inst_valid_up = valid_up; // @[Remove1S.scala 15:20]
  assign op_inst_I_0_0 = I_0_0_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_0_1 = I_0_0_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_0_2 = I_0_0_2; // @[Remove1S.scala 13:13]
  assign op_inst_I_1_0 = I_0_1_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_1_1 = I_0_1_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_1_2 = I_0_1_2; // @[Remove1S.scala 13:13]
  assign op_inst_I_2_0 = I_0_2_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_2_1 = I_0_2_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_2_2 = I_0_2_2; // @[Remove1S.scala 13:13]
endmodule
module MapS_3(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0_0_0,
  input  [31:0] I_0_0_0_1,
  input  [31:0] I_0_0_0_2,
  input  [31:0] I_0_0_1_0,
  input  [31:0] I_0_0_1_1,
  input  [31:0] I_0_0_1_2,
  input  [31:0] I_0_0_2_0,
  input  [31:0] I_0_0_2_1,
  input  [31:0] I_0_0_2_2,
  input  [31:0] I_1_0_0_0,
  input  [31:0] I_1_0_0_1,
  input  [31:0] I_1_0_0_2,
  input  [31:0] I_1_0_1_0,
  input  [31:0] I_1_0_1_1,
  input  [31:0] I_1_0_1_2,
  input  [31:0] I_1_0_2_0,
  input  [31:0] I_1_0_2_1,
  input  [31:0] I_1_0_2_2,
  input  [31:0] I_2_0_0_0,
  input  [31:0] I_2_0_0_1,
  input  [31:0] I_2_0_0_2,
  input  [31:0] I_2_0_1_0,
  input  [31:0] I_2_0_1_1,
  input  [31:0] I_2_0_1_2,
  input  [31:0] I_2_0_2_0,
  input  [31:0] I_2_0_2_1,
  input  [31:0] I_2_0_2_2,
  input  [31:0] I_3_0_0_0,
  input  [31:0] I_3_0_0_1,
  input  [31:0] I_3_0_0_2,
  input  [31:0] I_3_0_1_0,
  input  [31:0] I_3_0_1_1,
  input  [31:0] I_3_0_1_2,
  input  [31:0] I_3_0_2_0,
  input  [31:0] I_3_0_2_1,
  input  [31:0] I_3_0_2_2,
  input  [31:0] I_4_0_0_0,
  input  [31:0] I_4_0_0_1,
  input  [31:0] I_4_0_0_2,
  input  [31:0] I_4_0_1_0,
  input  [31:0] I_4_0_1_1,
  input  [31:0] I_4_0_1_2,
  input  [31:0] I_4_0_2_0,
  input  [31:0] I_4_0_2_1,
  input  [31:0] I_4_0_2_2,
  input  [31:0] I_5_0_0_0,
  input  [31:0] I_5_0_0_1,
  input  [31:0] I_5_0_0_2,
  input  [31:0] I_5_0_1_0,
  input  [31:0] I_5_0_1_1,
  input  [31:0] I_5_0_1_2,
  input  [31:0] I_5_0_2_0,
  input  [31:0] I_5_0_2_1,
  input  [31:0] I_5_0_2_2,
  input  [31:0] I_6_0_0_0,
  input  [31:0] I_6_0_0_1,
  input  [31:0] I_6_0_0_2,
  input  [31:0] I_6_0_1_0,
  input  [31:0] I_6_0_1_1,
  input  [31:0] I_6_0_1_2,
  input  [31:0] I_6_0_2_0,
  input  [31:0] I_6_0_2_1,
  input  [31:0] I_6_0_2_2,
  input  [31:0] I_7_0_0_0,
  input  [31:0] I_7_0_0_1,
  input  [31:0] I_7_0_0_2,
  input  [31:0] I_7_0_1_0,
  input  [31:0] I_7_0_1_1,
  input  [31:0] I_7_0_1_2,
  input  [31:0] I_7_0_2_0,
  input  [31:0] I_7_0_2_1,
  input  [31:0] I_7_0_2_2,
  output [31:0] O_0_0_0,
  output [31:0] O_0_0_1,
  output [31:0] O_0_0_2,
  output [31:0] O_0_1_0,
  output [31:0] O_0_1_1,
  output [31:0] O_0_1_2,
  output [31:0] O_0_2_0,
  output [31:0] O_0_2_1,
  output [31:0] O_0_2_2,
  output [31:0] O_1_0_0,
  output [31:0] O_1_0_1,
  output [31:0] O_1_0_2,
  output [31:0] O_1_1_0,
  output [31:0] O_1_1_1,
  output [31:0] O_1_1_2,
  output [31:0] O_1_2_0,
  output [31:0] O_1_2_1,
  output [31:0] O_1_2_2,
  output [31:0] O_2_0_0,
  output [31:0] O_2_0_1,
  output [31:0] O_2_0_2,
  output [31:0] O_2_1_0,
  output [31:0] O_2_1_1,
  output [31:0] O_2_1_2,
  output [31:0] O_2_2_0,
  output [31:0] O_2_2_1,
  output [31:0] O_2_2_2,
  output [31:0] O_3_0_0,
  output [31:0] O_3_0_1,
  output [31:0] O_3_0_2,
  output [31:0] O_3_1_0,
  output [31:0] O_3_1_1,
  output [31:0] O_3_1_2,
  output [31:0] O_3_2_0,
  output [31:0] O_3_2_1,
  output [31:0] O_3_2_2,
  output [31:0] O_4_0_0,
  output [31:0] O_4_0_1,
  output [31:0] O_4_0_2,
  output [31:0] O_4_1_0,
  output [31:0] O_4_1_1,
  output [31:0] O_4_1_2,
  output [31:0] O_4_2_0,
  output [31:0] O_4_2_1,
  output [31:0] O_4_2_2,
  output [31:0] O_5_0_0,
  output [31:0] O_5_0_1,
  output [31:0] O_5_0_2,
  output [31:0] O_5_1_0,
  output [31:0] O_5_1_1,
  output [31:0] O_5_1_2,
  output [31:0] O_5_2_0,
  output [31:0] O_5_2_1,
  output [31:0] O_5_2_2,
  output [31:0] O_6_0_0,
  output [31:0] O_6_0_1,
  output [31:0] O_6_0_2,
  output [31:0] O_6_1_0,
  output [31:0] O_6_1_1,
  output [31:0] O_6_1_2,
  output [31:0] O_6_2_0,
  output [31:0] O_6_2_1,
  output [31:0] O_6_2_2,
  output [31:0] O_7_0_0,
  output [31:0] O_7_0_1,
  output [31:0] O_7_0_2,
  output [31:0] O_7_1_0,
  output [31:0] O_7_1_1,
  output [31:0] O_7_1_2,
  output [31:0] O_7_2_0,
  output [31:0] O_7_2_1,
  output [31:0] O_7_2_2
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_0_0; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_0_1; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_0_2; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_1_0; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_1_1; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_1_2; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_2_0; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_2_1; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_2_2; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_0_0; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_0_1; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_0_2; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_1_0; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_1_1; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_1_2; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_2_0; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_2_1; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_2_2; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_0_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_0_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_0_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_0_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_0_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_0_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_0_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_0_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_0_2_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_O_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_O_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_O_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_O_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_O_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_O_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_O_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_O_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_0_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_0_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_0_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_0_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_0_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_0_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_0_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_0_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_0_2_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_O_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_O_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_O_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_O_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_O_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_O_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_O_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_O_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_0_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_0_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_0_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_0_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_0_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_0_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_0_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_0_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_0_2_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_O_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_O_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_O_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_O_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_O_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_O_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_O_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_O_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_0_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_0_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_0_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_0_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_0_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_0_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_0_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_0_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_0_2_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_O_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_O_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_O_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_O_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_O_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_O_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_O_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_O_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_0_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_0_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_0_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_0_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_0_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_0_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_0_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_0_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_0_2_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_O_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_O_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_O_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_O_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_O_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_O_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_O_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_O_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_0_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_0_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_0_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_0_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_0_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_0_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_0_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_0_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_0_2_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_O_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_O_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_O_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_O_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_O_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_O_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_O_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_O_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_0_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_0_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_0_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_0_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_0_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_0_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_0_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_0_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_0_2_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_O_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_O_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_O_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_O_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_O_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_O_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_O_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_O_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_O_2_2; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  wire  _T_1; // @[MapS.scala 23:83]
  wire  _T_2; // @[MapS.scala 23:83]
  wire  _T_3; // @[MapS.scala 23:83]
  wire  _T_4; // @[MapS.scala 23:83]
  wire  _T_5; // @[MapS.scala 23:83]
  Remove1S_3 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_0_0(fst_op_I_0_0_0),
    .I_0_0_1(fst_op_I_0_0_1),
    .I_0_0_2(fst_op_I_0_0_2),
    .I_0_1_0(fst_op_I_0_1_0),
    .I_0_1_1(fst_op_I_0_1_1),
    .I_0_1_2(fst_op_I_0_1_2),
    .I_0_2_0(fst_op_I_0_2_0),
    .I_0_2_1(fst_op_I_0_2_1),
    .I_0_2_2(fst_op_I_0_2_2),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1),
    .O_0_2(fst_op_O_0_2),
    .O_1_0(fst_op_O_1_0),
    .O_1_1(fst_op_O_1_1),
    .O_1_2(fst_op_O_1_2),
    .O_2_0(fst_op_O_2_0),
    .O_2_1(fst_op_O_2_1),
    .O_2_2(fst_op_O_2_2)
  );
  Remove1S_3 other_ops_0 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_0_0(other_ops_0_I_0_0_0),
    .I_0_0_1(other_ops_0_I_0_0_1),
    .I_0_0_2(other_ops_0_I_0_0_2),
    .I_0_1_0(other_ops_0_I_0_1_0),
    .I_0_1_1(other_ops_0_I_0_1_1),
    .I_0_1_2(other_ops_0_I_0_1_2),
    .I_0_2_0(other_ops_0_I_0_2_0),
    .I_0_2_1(other_ops_0_I_0_2_1),
    .I_0_2_2(other_ops_0_I_0_2_2),
    .O_0_0(other_ops_0_O_0_0),
    .O_0_1(other_ops_0_O_0_1),
    .O_0_2(other_ops_0_O_0_2),
    .O_1_0(other_ops_0_O_1_0),
    .O_1_1(other_ops_0_O_1_1),
    .O_1_2(other_ops_0_O_1_2),
    .O_2_0(other_ops_0_O_2_0),
    .O_2_1(other_ops_0_O_2_1),
    .O_2_2(other_ops_0_O_2_2)
  );
  Remove1S_3 other_ops_1 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0_0_0(other_ops_1_I_0_0_0),
    .I_0_0_1(other_ops_1_I_0_0_1),
    .I_0_0_2(other_ops_1_I_0_0_2),
    .I_0_1_0(other_ops_1_I_0_1_0),
    .I_0_1_1(other_ops_1_I_0_1_1),
    .I_0_1_2(other_ops_1_I_0_1_2),
    .I_0_2_0(other_ops_1_I_0_2_0),
    .I_0_2_1(other_ops_1_I_0_2_1),
    .I_0_2_2(other_ops_1_I_0_2_2),
    .O_0_0(other_ops_1_O_0_0),
    .O_0_1(other_ops_1_O_0_1),
    .O_0_2(other_ops_1_O_0_2),
    .O_1_0(other_ops_1_O_1_0),
    .O_1_1(other_ops_1_O_1_1),
    .O_1_2(other_ops_1_O_1_2),
    .O_2_0(other_ops_1_O_2_0),
    .O_2_1(other_ops_1_O_2_1),
    .O_2_2(other_ops_1_O_2_2)
  );
  Remove1S_3 other_ops_2 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I_0_0_0(other_ops_2_I_0_0_0),
    .I_0_0_1(other_ops_2_I_0_0_1),
    .I_0_0_2(other_ops_2_I_0_0_2),
    .I_0_1_0(other_ops_2_I_0_1_0),
    .I_0_1_1(other_ops_2_I_0_1_1),
    .I_0_1_2(other_ops_2_I_0_1_2),
    .I_0_2_0(other_ops_2_I_0_2_0),
    .I_0_2_1(other_ops_2_I_0_2_1),
    .I_0_2_2(other_ops_2_I_0_2_2),
    .O_0_0(other_ops_2_O_0_0),
    .O_0_1(other_ops_2_O_0_1),
    .O_0_2(other_ops_2_O_0_2),
    .O_1_0(other_ops_2_O_1_0),
    .O_1_1(other_ops_2_O_1_1),
    .O_1_2(other_ops_2_O_1_2),
    .O_2_0(other_ops_2_O_2_0),
    .O_2_1(other_ops_2_O_2_1),
    .O_2_2(other_ops_2_O_2_2)
  );
  Remove1S_3 other_ops_3 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I_0_0_0(other_ops_3_I_0_0_0),
    .I_0_0_1(other_ops_3_I_0_0_1),
    .I_0_0_2(other_ops_3_I_0_0_2),
    .I_0_1_0(other_ops_3_I_0_1_0),
    .I_0_1_1(other_ops_3_I_0_1_1),
    .I_0_1_2(other_ops_3_I_0_1_2),
    .I_0_2_0(other_ops_3_I_0_2_0),
    .I_0_2_1(other_ops_3_I_0_2_1),
    .I_0_2_2(other_ops_3_I_0_2_2),
    .O_0_0(other_ops_3_O_0_0),
    .O_0_1(other_ops_3_O_0_1),
    .O_0_2(other_ops_3_O_0_2),
    .O_1_0(other_ops_3_O_1_0),
    .O_1_1(other_ops_3_O_1_1),
    .O_1_2(other_ops_3_O_1_2),
    .O_2_0(other_ops_3_O_2_0),
    .O_2_1(other_ops_3_O_2_1),
    .O_2_2(other_ops_3_O_2_2)
  );
  Remove1S_3 other_ops_4 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I_0_0_0(other_ops_4_I_0_0_0),
    .I_0_0_1(other_ops_4_I_0_0_1),
    .I_0_0_2(other_ops_4_I_0_0_2),
    .I_0_1_0(other_ops_4_I_0_1_0),
    .I_0_1_1(other_ops_4_I_0_1_1),
    .I_0_1_2(other_ops_4_I_0_1_2),
    .I_0_2_0(other_ops_4_I_0_2_0),
    .I_0_2_1(other_ops_4_I_0_2_1),
    .I_0_2_2(other_ops_4_I_0_2_2),
    .O_0_0(other_ops_4_O_0_0),
    .O_0_1(other_ops_4_O_0_1),
    .O_0_2(other_ops_4_O_0_2),
    .O_1_0(other_ops_4_O_1_0),
    .O_1_1(other_ops_4_O_1_1),
    .O_1_2(other_ops_4_O_1_2),
    .O_2_0(other_ops_4_O_2_0),
    .O_2_1(other_ops_4_O_2_1),
    .O_2_2(other_ops_4_O_2_2)
  );
  Remove1S_3 other_ops_5 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I_0_0_0(other_ops_5_I_0_0_0),
    .I_0_0_1(other_ops_5_I_0_0_1),
    .I_0_0_2(other_ops_5_I_0_0_2),
    .I_0_1_0(other_ops_5_I_0_1_0),
    .I_0_1_1(other_ops_5_I_0_1_1),
    .I_0_1_2(other_ops_5_I_0_1_2),
    .I_0_2_0(other_ops_5_I_0_2_0),
    .I_0_2_1(other_ops_5_I_0_2_1),
    .I_0_2_2(other_ops_5_I_0_2_2),
    .O_0_0(other_ops_5_O_0_0),
    .O_0_1(other_ops_5_O_0_1),
    .O_0_2(other_ops_5_O_0_2),
    .O_1_0(other_ops_5_O_1_0),
    .O_1_1(other_ops_5_O_1_1),
    .O_1_2(other_ops_5_O_1_2),
    .O_2_0(other_ops_5_O_2_0),
    .O_2_1(other_ops_5_O_2_1),
    .O_2_2(other_ops_5_O_2_2)
  );
  Remove1S_3 other_ops_6 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I_0_0_0(other_ops_6_I_0_0_0),
    .I_0_0_1(other_ops_6_I_0_0_1),
    .I_0_0_2(other_ops_6_I_0_0_2),
    .I_0_1_0(other_ops_6_I_0_1_0),
    .I_0_1_1(other_ops_6_I_0_1_1),
    .I_0_1_2(other_ops_6_I_0_1_2),
    .I_0_2_0(other_ops_6_I_0_2_0),
    .I_0_2_1(other_ops_6_I_0_2_1),
    .I_0_2_2(other_ops_6_I_0_2_2),
    .O_0_0(other_ops_6_O_0_0),
    .O_0_1(other_ops_6_O_0_1),
    .O_0_2(other_ops_6_O_0_2),
    .O_1_0(other_ops_6_O_1_0),
    .O_1_1(other_ops_6_O_1_1),
    .O_1_2(other_ops_6_O_1_2),
    .O_2_0(other_ops_6_O_2_0),
    .O_2_1(other_ops_6_O_2_1),
    .O_2_2(other_ops_6_O_2_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[MapS.scala 23:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[MapS.scala 23:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[MapS.scala 23:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[MapS.scala 23:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T_5 & other_ops_6_valid_down; // @[MapS.scala 23:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[MapS.scala 17:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[MapS.scala 17:8]
  assign O_0_0_2 = fst_op_O_0_2; // @[MapS.scala 17:8]
  assign O_0_1_0 = fst_op_O_1_0; // @[MapS.scala 17:8]
  assign O_0_1_1 = fst_op_O_1_1; // @[MapS.scala 17:8]
  assign O_0_1_2 = fst_op_O_1_2; // @[MapS.scala 17:8]
  assign O_0_2_0 = fst_op_O_2_0; // @[MapS.scala 17:8]
  assign O_0_2_1 = fst_op_O_2_1; // @[MapS.scala 17:8]
  assign O_0_2_2 = fst_op_O_2_2; // @[MapS.scala 17:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[MapS.scala 21:12]
  assign O_1_0_1 = other_ops_0_O_0_1; // @[MapS.scala 21:12]
  assign O_1_0_2 = other_ops_0_O_0_2; // @[MapS.scala 21:12]
  assign O_1_1_0 = other_ops_0_O_1_0; // @[MapS.scala 21:12]
  assign O_1_1_1 = other_ops_0_O_1_1; // @[MapS.scala 21:12]
  assign O_1_1_2 = other_ops_0_O_1_2; // @[MapS.scala 21:12]
  assign O_1_2_0 = other_ops_0_O_2_0; // @[MapS.scala 21:12]
  assign O_1_2_1 = other_ops_0_O_2_1; // @[MapS.scala 21:12]
  assign O_1_2_2 = other_ops_0_O_2_2; // @[MapS.scala 21:12]
  assign O_2_0_0 = other_ops_1_O_0_0; // @[MapS.scala 21:12]
  assign O_2_0_1 = other_ops_1_O_0_1; // @[MapS.scala 21:12]
  assign O_2_0_2 = other_ops_1_O_0_2; // @[MapS.scala 21:12]
  assign O_2_1_0 = other_ops_1_O_1_0; // @[MapS.scala 21:12]
  assign O_2_1_1 = other_ops_1_O_1_1; // @[MapS.scala 21:12]
  assign O_2_1_2 = other_ops_1_O_1_2; // @[MapS.scala 21:12]
  assign O_2_2_0 = other_ops_1_O_2_0; // @[MapS.scala 21:12]
  assign O_2_2_1 = other_ops_1_O_2_1; // @[MapS.scala 21:12]
  assign O_2_2_2 = other_ops_1_O_2_2; // @[MapS.scala 21:12]
  assign O_3_0_0 = other_ops_2_O_0_0; // @[MapS.scala 21:12]
  assign O_3_0_1 = other_ops_2_O_0_1; // @[MapS.scala 21:12]
  assign O_3_0_2 = other_ops_2_O_0_2; // @[MapS.scala 21:12]
  assign O_3_1_0 = other_ops_2_O_1_0; // @[MapS.scala 21:12]
  assign O_3_1_1 = other_ops_2_O_1_1; // @[MapS.scala 21:12]
  assign O_3_1_2 = other_ops_2_O_1_2; // @[MapS.scala 21:12]
  assign O_3_2_0 = other_ops_2_O_2_0; // @[MapS.scala 21:12]
  assign O_3_2_1 = other_ops_2_O_2_1; // @[MapS.scala 21:12]
  assign O_3_2_2 = other_ops_2_O_2_2; // @[MapS.scala 21:12]
  assign O_4_0_0 = other_ops_3_O_0_0; // @[MapS.scala 21:12]
  assign O_4_0_1 = other_ops_3_O_0_1; // @[MapS.scala 21:12]
  assign O_4_0_2 = other_ops_3_O_0_2; // @[MapS.scala 21:12]
  assign O_4_1_0 = other_ops_3_O_1_0; // @[MapS.scala 21:12]
  assign O_4_1_1 = other_ops_3_O_1_1; // @[MapS.scala 21:12]
  assign O_4_1_2 = other_ops_3_O_1_2; // @[MapS.scala 21:12]
  assign O_4_2_0 = other_ops_3_O_2_0; // @[MapS.scala 21:12]
  assign O_4_2_1 = other_ops_3_O_2_1; // @[MapS.scala 21:12]
  assign O_4_2_2 = other_ops_3_O_2_2; // @[MapS.scala 21:12]
  assign O_5_0_0 = other_ops_4_O_0_0; // @[MapS.scala 21:12]
  assign O_5_0_1 = other_ops_4_O_0_1; // @[MapS.scala 21:12]
  assign O_5_0_2 = other_ops_4_O_0_2; // @[MapS.scala 21:12]
  assign O_5_1_0 = other_ops_4_O_1_0; // @[MapS.scala 21:12]
  assign O_5_1_1 = other_ops_4_O_1_1; // @[MapS.scala 21:12]
  assign O_5_1_2 = other_ops_4_O_1_2; // @[MapS.scala 21:12]
  assign O_5_2_0 = other_ops_4_O_2_0; // @[MapS.scala 21:12]
  assign O_5_2_1 = other_ops_4_O_2_1; // @[MapS.scala 21:12]
  assign O_5_2_2 = other_ops_4_O_2_2; // @[MapS.scala 21:12]
  assign O_6_0_0 = other_ops_5_O_0_0; // @[MapS.scala 21:12]
  assign O_6_0_1 = other_ops_5_O_0_1; // @[MapS.scala 21:12]
  assign O_6_0_2 = other_ops_5_O_0_2; // @[MapS.scala 21:12]
  assign O_6_1_0 = other_ops_5_O_1_0; // @[MapS.scala 21:12]
  assign O_6_1_1 = other_ops_5_O_1_1; // @[MapS.scala 21:12]
  assign O_6_1_2 = other_ops_5_O_1_2; // @[MapS.scala 21:12]
  assign O_6_2_0 = other_ops_5_O_2_0; // @[MapS.scala 21:12]
  assign O_6_2_1 = other_ops_5_O_2_1; // @[MapS.scala 21:12]
  assign O_6_2_2 = other_ops_5_O_2_2; // @[MapS.scala 21:12]
  assign O_7_0_0 = other_ops_6_O_0_0; // @[MapS.scala 21:12]
  assign O_7_0_1 = other_ops_6_O_0_1; // @[MapS.scala 21:12]
  assign O_7_0_2 = other_ops_6_O_0_2; // @[MapS.scala 21:12]
  assign O_7_1_0 = other_ops_6_O_1_0; // @[MapS.scala 21:12]
  assign O_7_1_1 = other_ops_6_O_1_1; // @[MapS.scala 21:12]
  assign O_7_1_2 = other_ops_6_O_1_2; // @[MapS.scala 21:12]
  assign O_7_2_0 = other_ops_6_O_2_0; // @[MapS.scala 21:12]
  assign O_7_2_1 = other_ops_6_O_2_1; // @[MapS.scala 21:12]
  assign O_7_2_2 = other_ops_6_O_2_2; // @[MapS.scala 21:12]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_0_0 = I_0_0_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_0_1 = I_0_0_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_0_2 = I_0_0_0_2; // @[MapS.scala 16:12]
  assign fst_op_I_0_1_0 = I_0_0_1_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_1_1 = I_0_0_1_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_1_2 = I_0_0_1_2; // @[MapS.scala 16:12]
  assign fst_op_I_0_2_0 = I_0_0_2_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_2_1 = I_0_0_2_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_2_2 = I_0_0_2_2; // @[MapS.scala 16:12]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_0_0 = I_1_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_0_1 = I_1_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_0_2 = I_1_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1_0 = I_1_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1_1 = I_1_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1_2 = I_1_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2_0 = I_1_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2_1 = I_1_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2_2 = I_1_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0_0_0 = I_2_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_0_1 = I_2_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_0_2 = I_2_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1_0 = I_2_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1_1 = I_2_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1_2 = I_2_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2_0 = I_2_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2_1 = I_2_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2_2 = I_2_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_2_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_2_I_0_0_0 = I_3_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_0_1 = I_3_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_0_2 = I_3_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1_0 = I_3_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1_1 = I_3_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1_2 = I_3_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2_0 = I_3_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2_1 = I_3_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2_2 = I_3_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_3_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_3_I_0_0_0 = I_4_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_0_1 = I_4_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_0_2 = I_4_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_1_0 = I_4_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_1_1 = I_4_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_1_2 = I_4_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_2_0 = I_4_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_2_1 = I_4_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_2_2 = I_4_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_4_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_4_I_0_0_0 = I_5_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_0_1 = I_5_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_0_2 = I_5_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_1_0 = I_5_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_1_1 = I_5_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_1_2 = I_5_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_2_0 = I_5_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_2_1 = I_5_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_2_2 = I_5_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_5_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_5_I_0_0_0 = I_6_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_0_1 = I_6_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_0_2 = I_6_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_1_0 = I_6_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_1_1 = I_6_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_1_2 = I_6_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_2_0 = I_6_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_2_1 = I_6_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_2_2 = I_6_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_6_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_6_I_0_0_0 = I_7_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_0_1 = I_7_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_0_2 = I_7_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_1_0 = I_7_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_1_1 = I_7_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_1_2 = I_7_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_2_0 = I_7_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_2_1 = I_7_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_2_2 = I_7_0_2_2; // @[MapS.scala 20:41]
endmodule
module MapT_7(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0_0_0,
  input  [31:0] I_0_0_0_1,
  input  [31:0] I_0_0_0_2,
  input  [31:0] I_0_0_1_0,
  input  [31:0] I_0_0_1_1,
  input  [31:0] I_0_0_1_2,
  input  [31:0] I_0_0_2_0,
  input  [31:0] I_0_0_2_1,
  input  [31:0] I_0_0_2_2,
  input  [31:0] I_1_0_0_0,
  input  [31:0] I_1_0_0_1,
  input  [31:0] I_1_0_0_2,
  input  [31:0] I_1_0_1_0,
  input  [31:0] I_1_0_1_1,
  input  [31:0] I_1_0_1_2,
  input  [31:0] I_1_0_2_0,
  input  [31:0] I_1_0_2_1,
  input  [31:0] I_1_0_2_2,
  input  [31:0] I_2_0_0_0,
  input  [31:0] I_2_0_0_1,
  input  [31:0] I_2_0_0_2,
  input  [31:0] I_2_0_1_0,
  input  [31:0] I_2_0_1_1,
  input  [31:0] I_2_0_1_2,
  input  [31:0] I_2_0_2_0,
  input  [31:0] I_2_0_2_1,
  input  [31:0] I_2_0_2_2,
  input  [31:0] I_3_0_0_0,
  input  [31:0] I_3_0_0_1,
  input  [31:0] I_3_0_0_2,
  input  [31:0] I_3_0_1_0,
  input  [31:0] I_3_0_1_1,
  input  [31:0] I_3_0_1_2,
  input  [31:0] I_3_0_2_0,
  input  [31:0] I_3_0_2_1,
  input  [31:0] I_3_0_2_2,
  input  [31:0] I_4_0_0_0,
  input  [31:0] I_4_0_0_1,
  input  [31:0] I_4_0_0_2,
  input  [31:0] I_4_0_1_0,
  input  [31:0] I_4_0_1_1,
  input  [31:0] I_4_0_1_2,
  input  [31:0] I_4_0_2_0,
  input  [31:0] I_4_0_2_1,
  input  [31:0] I_4_0_2_2,
  input  [31:0] I_5_0_0_0,
  input  [31:0] I_5_0_0_1,
  input  [31:0] I_5_0_0_2,
  input  [31:0] I_5_0_1_0,
  input  [31:0] I_5_0_1_1,
  input  [31:0] I_5_0_1_2,
  input  [31:0] I_5_0_2_0,
  input  [31:0] I_5_0_2_1,
  input  [31:0] I_5_0_2_2,
  input  [31:0] I_6_0_0_0,
  input  [31:0] I_6_0_0_1,
  input  [31:0] I_6_0_0_2,
  input  [31:0] I_6_0_1_0,
  input  [31:0] I_6_0_1_1,
  input  [31:0] I_6_0_1_2,
  input  [31:0] I_6_0_2_0,
  input  [31:0] I_6_0_2_1,
  input  [31:0] I_6_0_2_2,
  input  [31:0] I_7_0_0_0,
  input  [31:0] I_7_0_0_1,
  input  [31:0] I_7_0_0_2,
  input  [31:0] I_7_0_1_0,
  input  [31:0] I_7_0_1_1,
  input  [31:0] I_7_0_1_2,
  input  [31:0] I_7_0_2_0,
  input  [31:0] I_7_0_2_1,
  input  [31:0] I_7_0_2_2,
  output [31:0] O_0_0_0,
  output [31:0] O_0_0_1,
  output [31:0] O_0_0_2,
  output [31:0] O_0_1_0,
  output [31:0] O_0_1_1,
  output [31:0] O_0_1_2,
  output [31:0] O_0_2_0,
  output [31:0] O_0_2_1,
  output [31:0] O_0_2_2,
  output [31:0] O_1_0_0,
  output [31:0] O_1_0_1,
  output [31:0] O_1_0_2,
  output [31:0] O_1_1_0,
  output [31:0] O_1_1_1,
  output [31:0] O_1_1_2,
  output [31:0] O_1_2_0,
  output [31:0] O_1_2_1,
  output [31:0] O_1_2_2,
  output [31:0] O_2_0_0,
  output [31:0] O_2_0_1,
  output [31:0] O_2_0_2,
  output [31:0] O_2_1_0,
  output [31:0] O_2_1_1,
  output [31:0] O_2_1_2,
  output [31:0] O_2_2_0,
  output [31:0] O_2_2_1,
  output [31:0] O_2_2_2,
  output [31:0] O_3_0_0,
  output [31:0] O_3_0_1,
  output [31:0] O_3_0_2,
  output [31:0] O_3_1_0,
  output [31:0] O_3_1_1,
  output [31:0] O_3_1_2,
  output [31:0] O_3_2_0,
  output [31:0] O_3_2_1,
  output [31:0] O_3_2_2,
  output [31:0] O_4_0_0,
  output [31:0] O_4_0_1,
  output [31:0] O_4_0_2,
  output [31:0] O_4_1_0,
  output [31:0] O_4_1_1,
  output [31:0] O_4_1_2,
  output [31:0] O_4_2_0,
  output [31:0] O_4_2_1,
  output [31:0] O_4_2_2,
  output [31:0] O_5_0_0,
  output [31:0] O_5_0_1,
  output [31:0] O_5_0_2,
  output [31:0] O_5_1_0,
  output [31:0] O_5_1_1,
  output [31:0] O_5_1_2,
  output [31:0] O_5_2_0,
  output [31:0] O_5_2_1,
  output [31:0] O_5_2_2,
  output [31:0] O_6_0_0,
  output [31:0] O_6_0_1,
  output [31:0] O_6_0_2,
  output [31:0] O_6_1_0,
  output [31:0] O_6_1_1,
  output [31:0] O_6_1_2,
  output [31:0] O_6_2_0,
  output [31:0] O_6_2_1,
  output [31:0] O_6_2_2,
  output [31:0] O_7_0_0,
  output [31:0] O_7_0_1,
  output [31:0] O_7_0_2,
  output [31:0] O_7_1_0,
  output [31:0] O_7_1_1,
  output [31:0] O_7_1_2,
  output [31:0] O_7_2_0,
  output [31:0] O_7_2_1,
  output [31:0] O_7_2_2
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_2_2; // @[MapT.scala 8:20]
  MapS_3 op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0_0(op_I_0_0_0_0),
    .I_0_0_0_1(op_I_0_0_0_1),
    .I_0_0_0_2(op_I_0_0_0_2),
    .I_0_0_1_0(op_I_0_0_1_0),
    .I_0_0_1_1(op_I_0_0_1_1),
    .I_0_0_1_2(op_I_0_0_1_2),
    .I_0_0_2_0(op_I_0_0_2_0),
    .I_0_0_2_1(op_I_0_0_2_1),
    .I_0_0_2_2(op_I_0_0_2_2),
    .I_1_0_0_0(op_I_1_0_0_0),
    .I_1_0_0_1(op_I_1_0_0_1),
    .I_1_0_0_2(op_I_1_0_0_2),
    .I_1_0_1_0(op_I_1_0_1_0),
    .I_1_0_1_1(op_I_1_0_1_1),
    .I_1_0_1_2(op_I_1_0_1_2),
    .I_1_0_2_0(op_I_1_0_2_0),
    .I_1_0_2_1(op_I_1_0_2_1),
    .I_1_0_2_2(op_I_1_0_2_2),
    .I_2_0_0_0(op_I_2_0_0_0),
    .I_2_0_0_1(op_I_2_0_0_1),
    .I_2_0_0_2(op_I_2_0_0_2),
    .I_2_0_1_0(op_I_2_0_1_0),
    .I_2_0_1_1(op_I_2_0_1_1),
    .I_2_0_1_2(op_I_2_0_1_2),
    .I_2_0_2_0(op_I_2_0_2_0),
    .I_2_0_2_1(op_I_2_0_2_1),
    .I_2_0_2_2(op_I_2_0_2_2),
    .I_3_0_0_0(op_I_3_0_0_0),
    .I_3_0_0_1(op_I_3_0_0_1),
    .I_3_0_0_2(op_I_3_0_0_2),
    .I_3_0_1_0(op_I_3_0_1_0),
    .I_3_0_1_1(op_I_3_0_1_1),
    .I_3_0_1_2(op_I_3_0_1_2),
    .I_3_0_2_0(op_I_3_0_2_0),
    .I_3_0_2_1(op_I_3_0_2_1),
    .I_3_0_2_2(op_I_3_0_2_2),
    .I_4_0_0_0(op_I_4_0_0_0),
    .I_4_0_0_1(op_I_4_0_0_1),
    .I_4_0_0_2(op_I_4_0_0_2),
    .I_4_0_1_0(op_I_4_0_1_0),
    .I_4_0_1_1(op_I_4_0_1_1),
    .I_4_0_1_2(op_I_4_0_1_2),
    .I_4_0_2_0(op_I_4_0_2_0),
    .I_4_0_2_1(op_I_4_0_2_1),
    .I_4_0_2_2(op_I_4_0_2_2),
    .I_5_0_0_0(op_I_5_0_0_0),
    .I_5_0_0_1(op_I_5_0_0_1),
    .I_5_0_0_2(op_I_5_0_0_2),
    .I_5_0_1_0(op_I_5_0_1_0),
    .I_5_0_1_1(op_I_5_0_1_1),
    .I_5_0_1_2(op_I_5_0_1_2),
    .I_5_0_2_0(op_I_5_0_2_0),
    .I_5_0_2_1(op_I_5_0_2_1),
    .I_5_0_2_2(op_I_5_0_2_2),
    .I_6_0_0_0(op_I_6_0_0_0),
    .I_6_0_0_1(op_I_6_0_0_1),
    .I_6_0_0_2(op_I_6_0_0_2),
    .I_6_0_1_0(op_I_6_0_1_0),
    .I_6_0_1_1(op_I_6_0_1_1),
    .I_6_0_1_2(op_I_6_0_1_2),
    .I_6_0_2_0(op_I_6_0_2_0),
    .I_6_0_2_1(op_I_6_0_2_1),
    .I_6_0_2_2(op_I_6_0_2_2),
    .I_7_0_0_0(op_I_7_0_0_0),
    .I_7_0_0_1(op_I_7_0_0_1),
    .I_7_0_0_2(op_I_7_0_0_2),
    .I_7_0_1_0(op_I_7_0_1_0),
    .I_7_0_1_1(op_I_7_0_1_1),
    .I_7_0_1_2(op_I_7_0_1_2),
    .I_7_0_2_0(op_I_7_0_2_0),
    .I_7_0_2_1(op_I_7_0_2_1),
    .I_7_0_2_2(op_I_7_0_2_2),
    .O_0_0_0(op_O_0_0_0),
    .O_0_0_1(op_O_0_0_1),
    .O_0_0_2(op_O_0_0_2),
    .O_0_1_0(op_O_0_1_0),
    .O_0_1_1(op_O_0_1_1),
    .O_0_1_2(op_O_0_1_2),
    .O_0_2_0(op_O_0_2_0),
    .O_0_2_1(op_O_0_2_1),
    .O_0_2_2(op_O_0_2_2),
    .O_1_0_0(op_O_1_0_0),
    .O_1_0_1(op_O_1_0_1),
    .O_1_0_2(op_O_1_0_2),
    .O_1_1_0(op_O_1_1_0),
    .O_1_1_1(op_O_1_1_1),
    .O_1_1_2(op_O_1_1_2),
    .O_1_2_0(op_O_1_2_0),
    .O_1_2_1(op_O_1_2_1),
    .O_1_2_2(op_O_1_2_2),
    .O_2_0_0(op_O_2_0_0),
    .O_2_0_1(op_O_2_0_1),
    .O_2_0_2(op_O_2_0_2),
    .O_2_1_0(op_O_2_1_0),
    .O_2_1_1(op_O_2_1_1),
    .O_2_1_2(op_O_2_1_2),
    .O_2_2_0(op_O_2_2_0),
    .O_2_2_1(op_O_2_2_1),
    .O_2_2_2(op_O_2_2_2),
    .O_3_0_0(op_O_3_0_0),
    .O_3_0_1(op_O_3_0_1),
    .O_3_0_2(op_O_3_0_2),
    .O_3_1_0(op_O_3_1_0),
    .O_3_1_1(op_O_3_1_1),
    .O_3_1_2(op_O_3_1_2),
    .O_3_2_0(op_O_3_2_0),
    .O_3_2_1(op_O_3_2_1),
    .O_3_2_2(op_O_3_2_2),
    .O_4_0_0(op_O_4_0_0),
    .O_4_0_1(op_O_4_0_1),
    .O_4_0_2(op_O_4_0_2),
    .O_4_1_0(op_O_4_1_0),
    .O_4_1_1(op_O_4_1_1),
    .O_4_1_2(op_O_4_1_2),
    .O_4_2_0(op_O_4_2_0),
    .O_4_2_1(op_O_4_2_1),
    .O_4_2_2(op_O_4_2_2),
    .O_5_0_0(op_O_5_0_0),
    .O_5_0_1(op_O_5_0_1),
    .O_5_0_2(op_O_5_0_2),
    .O_5_1_0(op_O_5_1_0),
    .O_5_1_1(op_O_5_1_1),
    .O_5_1_2(op_O_5_1_2),
    .O_5_2_0(op_O_5_2_0),
    .O_5_2_1(op_O_5_2_1),
    .O_5_2_2(op_O_5_2_2),
    .O_6_0_0(op_O_6_0_0),
    .O_6_0_1(op_O_6_0_1),
    .O_6_0_2(op_O_6_0_2),
    .O_6_1_0(op_O_6_1_0),
    .O_6_1_1(op_O_6_1_1),
    .O_6_1_2(op_O_6_1_2),
    .O_6_2_0(op_O_6_2_0),
    .O_6_2_1(op_O_6_2_1),
    .O_6_2_2(op_O_6_2_2),
    .O_7_0_0(op_O_7_0_0),
    .O_7_0_1(op_O_7_0_1),
    .O_7_0_2(op_O_7_0_2),
    .O_7_1_0(op_O_7_1_0),
    .O_7_1_1(op_O_7_1_1),
    .O_7_1_2(op_O_7_1_2),
    .O_7_2_0(op_O_7_2_0),
    .O_7_2_1(op_O_7_2_1),
    .O_7_2_2(op_O_7_2_2)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0 = op_O_0_0_0; // @[MapT.scala 15:7]
  assign O_0_0_1 = op_O_0_0_1; // @[MapT.scala 15:7]
  assign O_0_0_2 = op_O_0_0_2; // @[MapT.scala 15:7]
  assign O_0_1_0 = op_O_0_1_0; // @[MapT.scala 15:7]
  assign O_0_1_1 = op_O_0_1_1; // @[MapT.scala 15:7]
  assign O_0_1_2 = op_O_0_1_2; // @[MapT.scala 15:7]
  assign O_0_2_0 = op_O_0_2_0; // @[MapT.scala 15:7]
  assign O_0_2_1 = op_O_0_2_1; // @[MapT.scala 15:7]
  assign O_0_2_2 = op_O_0_2_2; // @[MapT.scala 15:7]
  assign O_1_0_0 = op_O_1_0_0; // @[MapT.scala 15:7]
  assign O_1_0_1 = op_O_1_0_1; // @[MapT.scala 15:7]
  assign O_1_0_2 = op_O_1_0_2; // @[MapT.scala 15:7]
  assign O_1_1_0 = op_O_1_1_0; // @[MapT.scala 15:7]
  assign O_1_1_1 = op_O_1_1_1; // @[MapT.scala 15:7]
  assign O_1_1_2 = op_O_1_1_2; // @[MapT.scala 15:7]
  assign O_1_2_0 = op_O_1_2_0; // @[MapT.scala 15:7]
  assign O_1_2_1 = op_O_1_2_1; // @[MapT.scala 15:7]
  assign O_1_2_2 = op_O_1_2_2; // @[MapT.scala 15:7]
  assign O_2_0_0 = op_O_2_0_0; // @[MapT.scala 15:7]
  assign O_2_0_1 = op_O_2_0_1; // @[MapT.scala 15:7]
  assign O_2_0_2 = op_O_2_0_2; // @[MapT.scala 15:7]
  assign O_2_1_0 = op_O_2_1_0; // @[MapT.scala 15:7]
  assign O_2_1_1 = op_O_2_1_1; // @[MapT.scala 15:7]
  assign O_2_1_2 = op_O_2_1_2; // @[MapT.scala 15:7]
  assign O_2_2_0 = op_O_2_2_0; // @[MapT.scala 15:7]
  assign O_2_2_1 = op_O_2_2_1; // @[MapT.scala 15:7]
  assign O_2_2_2 = op_O_2_2_2; // @[MapT.scala 15:7]
  assign O_3_0_0 = op_O_3_0_0; // @[MapT.scala 15:7]
  assign O_3_0_1 = op_O_3_0_1; // @[MapT.scala 15:7]
  assign O_3_0_2 = op_O_3_0_2; // @[MapT.scala 15:7]
  assign O_3_1_0 = op_O_3_1_0; // @[MapT.scala 15:7]
  assign O_3_1_1 = op_O_3_1_1; // @[MapT.scala 15:7]
  assign O_3_1_2 = op_O_3_1_2; // @[MapT.scala 15:7]
  assign O_3_2_0 = op_O_3_2_0; // @[MapT.scala 15:7]
  assign O_3_2_1 = op_O_3_2_1; // @[MapT.scala 15:7]
  assign O_3_2_2 = op_O_3_2_2; // @[MapT.scala 15:7]
  assign O_4_0_0 = op_O_4_0_0; // @[MapT.scala 15:7]
  assign O_4_0_1 = op_O_4_0_1; // @[MapT.scala 15:7]
  assign O_4_0_2 = op_O_4_0_2; // @[MapT.scala 15:7]
  assign O_4_1_0 = op_O_4_1_0; // @[MapT.scala 15:7]
  assign O_4_1_1 = op_O_4_1_1; // @[MapT.scala 15:7]
  assign O_4_1_2 = op_O_4_1_2; // @[MapT.scala 15:7]
  assign O_4_2_0 = op_O_4_2_0; // @[MapT.scala 15:7]
  assign O_4_2_1 = op_O_4_2_1; // @[MapT.scala 15:7]
  assign O_4_2_2 = op_O_4_2_2; // @[MapT.scala 15:7]
  assign O_5_0_0 = op_O_5_0_0; // @[MapT.scala 15:7]
  assign O_5_0_1 = op_O_5_0_1; // @[MapT.scala 15:7]
  assign O_5_0_2 = op_O_5_0_2; // @[MapT.scala 15:7]
  assign O_5_1_0 = op_O_5_1_0; // @[MapT.scala 15:7]
  assign O_5_1_1 = op_O_5_1_1; // @[MapT.scala 15:7]
  assign O_5_1_2 = op_O_5_1_2; // @[MapT.scala 15:7]
  assign O_5_2_0 = op_O_5_2_0; // @[MapT.scala 15:7]
  assign O_5_2_1 = op_O_5_2_1; // @[MapT.scala 15:7]
  assign O_5_2_2 = op_O_5_2_2; // @[MapT.scala 15:7]
  assign O_6_0_0 = op_O_6_0_0; // @[MapT.scala 15:7]
  assign O_6_0_1 = op_O_6_0_1; // @[MapT.scala 15:7]
  assign O_6_0_2 = op_O_6_0_2; // @[MapT.scala 15:7]
  assign O_6_1_0 = op_O_6_1_0; // @[MapT.scala 15:7]
  assign O_6_1_1 = op_O_6_1_1; // @[MapT.scala 15:7]
  assign O_6_1_2 = op_O_6_1_2; // @[MapT.scala 15:7]
  assign O_6_2_0 = op_O_6_2_0; // @[MapT.scala 15:7]
  assign O_6_2_1 = op_O_6_2_1; // @[MapT.scala 15:7]
  assign O_6_2_2 = op_O_6_2_2; // @[MapT.scala 15:7]
  assign O_7_0_0 = op_O_7_0_0; // @[MapT.scala 15:7]
  assign O_7_0_1 = op_O_7_0_1; // @[MapT.scala 15:7]
  assign O_7_0_2 = op_O_7_0_2; // @[MapT.scala 15:7]
  assign O_7_1_0 = op_O_7_1_0; // @[MapT.scala 15:7]
  assign O_7_1_1 = op_O_7_1_1; // @[MapT.scala 15:7]
  assign O_7_1_2 = op_O_7_1_2; // @[MapT.scala 15:7]
  assign O_7_2_0 = op_O_7_2_0; // @[MapT.scala 15:7]
  assign O_7_2_1 = op_O_7_2_1; // @[MapT.scala 15:7]
  assign O_7_2_2 = op_O_7_2_2; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0_0 = I_0_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_0_1 = I_0_0_0_1; // @[MapT.scala 14:10]
  assign op_I_0_0_0_2 = I_0_0_0_2; // @[MapT.scala 14:10]
  assign op_I_0_0_1_0 = I_0_0_1_0; // @[MapT.scala 14:10]
  assign op_I_0_0_1_1 = I_0_0_1_1; // @[MapT.scala 14:10]
  assign op_I_0_0_1_2 = I_0_0_1_2; // @[MapT.scala 14:10]
  assign op_I_0_0_2_0 = I_0_0_2_0; // @[MapT.scala 14:10]
  assign op_I_0_0_2_1 = I_0_0_2_1; // @[MapT.scala 14:10]
  assign op_I_0_0_2_2 = I_0_0_2_2; // @[MapT.scala 14:10]
  assign op_I_1_0_0_0 = I_1_0_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_0_1 = I_1_0_0_1; // @[MapT.scala 14:10]
  assign op_I_1_0_0_2 = I_1_0_0_2; // @[MapT.scala 14:10]
  assign op_I_1_0_1_0 = I_1_0_1_0; // @[MapT.scala 14:10]
  assign op_I_1_0_1_1 = I_1_0_1_1; // @[MapT.scala 14:10]
  assign op_I_1_0_1_2 = I_1_0_1_2; // @[MapT.scala 14:10]
  assign op_I_1_0_2_0 = I_1_0_2_0; // @[MapT.scala 14:10]
  assign op_I_1_0_2_1 = I_1_0_2_1; // @[MapT.scala 14:10]
  assign op_I_1_0_2_2 = I_1_0_2_2; // @[MapT.scala 14:10]
  assign op_I_2_0_0_0 = I_2_0_0_0; // @[MapT.scala 14:10]
  assign op_I_2_0_0_1 = I_2_0_0_1; // @[MapT.scala 14:10]
  assign op_I_2_0_0_2 = I_2_0_0_2; // @[MapT.scala 14:10]
  assign op_I_2_0_1_0 = I_2_0_1_0; // @[MapT.scala 14:10]
  assign op_I_2_0_1_1 = I_2_0_1_1; // @[MapT.scala 14:10]
  assign op_I_2_0_1_2 = I_2_0_1_2; // @[MapT.scala 14:10]
  assign op_I_2_0_2_0 = I_2_0_2_0; // @[MapT.scala 14:10]
  assign op_I_2_0_2_1 = I_2_0_2_1; // @[MapT.scala 14:10]
  assign op_I_2_0_2_2 = I_2_0_2_2; // @[MapT.scala 14:10]
  assign op_I_3_0_0_0 = I_3_0_0_0; // @[MapT.scala 14:10]
  assign op_I_3_0_0_1 = I_3_0_0_1; // @[MapT.scala 14:10]
  assign op_I_3_0_0_2 = I_3_0_0_2; // @[MapT.scala 14:10]
  assign op_I_3_0_1_0 = I_3_0_1_0; // @[MapT.scala 14:10]
  assign op_I_3_0_1_1 = I_3_0_1_1; // @[MapT.scala 14:10]
  assign op_I_3_0_1_2 = I_3_0_1_2; // @[MapT.scala 14:10]
  assign op_I_3_0_2_0 = I_3_0_2_0; // @[MapT.scala 14:10]
  assign op_I_3_0_2_1 = I_3_0_2_1; // @[MapT.scala 14:10]
  assign op_I_3_0_2_2 = I_3_0_2_2; // @[MapT.scala 14:10]
  assign op_I_4_0_0_0 = I_4_0_0_0; // @[MapT.scala 14:10]
  assign op_I_4_0_0_1 = I_4_0_0_1; // @[MapT.scala 14:10]
  assign op_I_4_0_0_2 = I_4_0_0_2; // @[MapT.scala 14:10]
  assign op_I_4_0_1_0 = I_4_0_1_0; // @[MapT.scala 14:10]
  assign op_I_4_0_1_1 = I_4_0_1_1; // @[MapT.scala 14:10]
  assign op_I_4_0_1_2 = I_4_0_1_2; // @[MapT.scala 14:10]
  assign op_I_4_0_2_0 = I_4_0_2_0; // @[MapT.scala 14:10]
  assign op_I_4_0_2_1 = I_4_0_2_1; // @[MapT.scala 14:10]
  assign op_I_4_0_2_2 = I_4_0_2_2; // @[MapT.scala 14:10]
  assign op_I_5_0_0_0 = I_5_0_0_0; // @[MapT.scala 14:10]
  assign op_I_5_0_0_1 = I_5_0_0_1; // @[MapT.scala 14:10]
  assign op_I_5_0_0_2 = I_5_0_0_2; // @[MapT.scala 14:10]
  assign op_I_5_0_1_0 = I_5_0_1_0; // @[MapT.scala 14:10]
  assign op_I_5_0_1_1 = I_5_0_1_1; // @[MapT.scala 14:10]
  assign op_I_5_0_1_2 = I_5_0_1_2; // @[MapT.scala 14:10]
  assign op_I_5_0_2_0 = I_5_0_2_0; // @[MapT.scala 14:10]
  assign op_I_5_0_2_1 = I_5_0_2_1; // @[MapT.scala 14:10]
  assign op_I_5_0_2_2 = I_5_0_2_2; // @[MapT.scala 14:10]
  assign op_I_6_0_0_0 = I_6_0_0_0; // @[MapT.scala 14:10]
  assign op_I_6_0_0_1 = I_6_0_0_1; // @[MapT.scala 14:10]
  assign op_I_6_0_0_2 = I_6_0_0_2; // @[MapT.scala 14:10]
  assign op_I_6_0_1_0 = I_6_0_1_0; // @[MapT.scala 14:10]
  assign op_I_6_0_1_1 = I_6_0_1_1; // @[MapT.scala 14:10]
  assign op_I_6_0_1_2 = I_6_0_1_2; // @[MapT.scala 14:10]
  assign op_I_6_0_2_0 = I_6_0_2_0; // @[MapT.scala 14:10]
  assign op_I_6_0_2_1 = I_6_0_2_1; // @[MapT.scala 14:10]
  assign op_I_6_0_2_2 = I_6_0_2_2; // @[MapT.scala 14:10]
  assign op_I_7_0_0_0 = I_7_0_0_0; // @[MapT.scala 14:10]
  assign op_I_7_0_0_1 = I_7_0_0_1; // @[MapT.scala 14:10]
  assign op_I_7_0_0_2 = I_7_0_0_2; // @[MapT.scala 14:10]
  assign op_I_7_0_1_0 = I_7_0_1_0; // @[MapT.scala 14:10]
  assign op_I_7_0_1_1 = I_7_0_1_1; // @[MapT.scala 14:10]
  assign op_I_7_0_1_2 = I_7_0_1_2; // @[MapT.scala 14:10]
  assign op_I_7_0_2_0 = I_7_0_2_0; // @[MapT.scala 14:10]
  assign op_I_7_0_2_1 = I_7_0_2_1; // @[MapT.scala 14:10]
  assign op_I_7_0_2_2 = I_7_0_2_2; // @[MapT.scala 14:10]
endmodule
module Passthrough(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0_0,
  input  [31:0] I_0_0_1,
  input  [31:0] I_0_0_2,
  input  [31:0] I_0_1_0,
  input  [31:0] I_0_1_1,
  input  [31:0] I_0_1_2,
  input  [31:0] I_0_2_0,
  input  [31:0] I_0_2_1,
  input  [31:0] I_0_2_2,
  input  [31:0] I_1_0_0,
  input  [31:0] I_1_0_1,
  input  [31:0] I_1_0_2,
  input  [31:0] I_1_1_0,
  input  [31:0] I_1_1_1,
  input  [31:0] I_1_1_2,
  input  [31:0] I_1_2_0,
  input  [31:0] I_1_2_1,
  input  [31:0] I_1_2_2,
  input  [31:0] I_2_0_0,
  input  [31:0] I_2_0_1,
  input  [31:0] I_2_0_2,
  input  [31:0] I_2_1_0,
  input  [31:0] I_2_1_1,
  input  [31:0] I_2_1_2,
  input  [31:0] I_2_2_0,
  input  [31:0] I_2_2_1,
  input  [31:0] I_2_2_2,
  input  [31:0] I_3_0_0,
  input  [31:0] I_3_0_1,
  input  [31:0] I_3_0_2,
  input  [31:0] I_3_1_0,
  input  [31:0] I_3_1_1,
  input  [31:0] I_3_1_2,
  input  [31:0] I_3_2_0,
  input  [31:0] I_3_2_1,
  input  [31:0] I_3_2_2,
  input  [31:0] I_4_0_0,
  input  [31:0] I_4_0_1,
  input  [31:0] I_4_0_2,
  input  [31:0] I_4_1_0,
  input  [31:0] I_4_1_1,
  input  [31:0] I_4_1_2,
  input  [31:0] I_4_2_0,
  input  [31:0] I_4_2_1,
  input  [31:0] I_4_2_2,
  input  [31:0] I_5_0_0,
  input  [31:0] I_5_0_1,
  input  [31:0] I_5_0_2,
  input  [31:0] I_5_1_0,
  input  [31:0] I_5_1_1,
  input  [31:0] I_5_1_2,
  input  [31:0] I_5_2_0,
  input  [31:0] I_5_2_1,
  input  [31:0] I_5_2_2,
  input  [31:0] I_6_0_0,
  input  [31:0] I_6_0_1,
  input  [31:0] I_6_0_2,
  input  [31:0] I_6_1_0,
  input  [31:0] I_6_1_1,
  input  [31:0] I_6_1_2,
  input  [31:0] I_6_2_0,
  input  [31:0] I_6_2_1,
  input  [31:0] I_6_2_2,
  input  [31:0] I_7_0_0,
  input  [31:0] I_7_0_1,
  input  [31:0] I_7_0_2,
  input  [31:0] I_7_1_0,
  input  [31:0] I_7_1_1,
  input  [31:0] I_7_1_2,
  input  [31:0] I_7_2_0,
  input  [31:0] I_7_2_1,
  input  [31:0] I_7_2_2,
  output [31:0] O_0_0_0,
  output [31:0] O_0_0_1,
  output [31:0] O_0_0_2,
  output [31:0] O_0_1_0,
  output [31:0] O_0_1_1,
  output [31:0] O_0_1_2,
  output [31:0] O_0_2_0,
  output [31:0] O_0_2_1,
  output [31:0] O_0_2_2,
  output [31:0] O_1_0_0,
  output [31:0] O_1_0_1,
  output [31:0] O_1_0_2,
  output [31:0] O_1_1_0,
  output [31:0] O_1_1_1,
  output [31:0] O_1_1_2,
  output [31:0] O_1_2_0,
  output [31:0] O_1_2_1,
  output [31:0] O_1_2_2,
  output [31:0] O_2_0_0,
  output [31:0] O_2_0_1,
  output [31:0] O_2_0_2,
  output [31:0] O_2_1_0,
  output [31:0] O_2_1_1,
  output [31:0] O_2_1_2,
  output [31:0] O_2_2_0,
  output [31:0] O_2_2_1,
  output [31:0] O_2_2_2,
  output [31:0] O_3_0_0,
  output [31:0] O_3_0_1,
  output [31:0] O_3_0_2,
  output [31:0] O_3_1_0,
  output [31:0] O_3_1_1,
  output [31:0] O_3_1_2,
  output [31:0] O_3_2_0,
  output [31:0] O_3_2_1,
  output [31:0] O_3_2_2,
  output [31:0] O_4_0_0,
  output [31:0] O_4_0_1,
  output [31:0] O_4_0_2,
  output [31:0] O_4_1_0,
  output [31:0] O_4_1_1,
  output [31:0] O_4_1_2,
  output [31:0] O_4_2_0,
  output [31:0] O_4_2_1,
  output [31:0] O_4_2_2,
  output [31:0] O_5_0_0,
  output [31:0] O_5_0_1,
  output [31:0] O_5_0_2,
  output [31:0] O_5_1_0,
  output [31:0] O_5_1_1,
  output [31:0] O_5_1_2,
  output [31:0] O_5_2_0,
  output [31:0] O_5_2_1,
  output [31:0] O_5_2_2,
  output [31:0] O_6_0_0,
  output [31:0] O_6_0_1,
  output [31:0] O_6_0_2,
  output [31:0] O_6_1_0,
  output [31:0] O_6_1_1,
  output [31:0] O_6_1_2,
  output [31:0] O_6_2_0,
  output [31:0] O_6_2_1,
  output [31:0] O_6_2_2,
  output [31:0] O_7_0_0,
  output [31:0] O_7_0_1,
  output [31:0] O_7_0_2,
  output [31:0] O_7_1_0,
  output [31:0] O_7_1_1,
  output [31:0] O_7_1_2,
  output [31:0] O_7_2_0,
  output [31:0] O_7_2_1,
  output [31:0] O_7_2_2
);
  assign valid_down = valid_up; // @[Passthrough.scala 18:14]
  assign O_0_0_0 = I_0_0_0; // @[Passthrough.scala 17:68]
  assign O_0_0_1 = I_0_0_1; // @[Passthrough.scala 17:68]
  assign O_0_0_2 = I_0_0_2; // @[Passthrough.scala 17:68]
  assign O_0_1_0 = I_0_1_0; // @[Passthrough.scala 17:68]
  assign O_0_1_1 = I_0_1_1; // @[Passthrough.scala 17:68]
  assign O_0_1_2 = I_0_1_2; // @[Passthrough.scala 17:68]
  assign O_0_2_0 = I_0_2_0; // @[Passthrough.scala 17:68]
  assign O_0_2_1 = I_0_2_1; // @[Passthrough.scala 17:68]
  assign O_0_2_2 = I_0_2_2; // @[Passthrough.scala 17:68]
  assign O_1_0_0 = I_1_0_0; // @[Passthrough.scala 17:68]
  assign O_1_0_1 = I_1_0_1; // @[Passthrough.scala 17:68]
  assign O_1_0_2 = I_1_0_2; // @[Passthrough.scala 17:68]
  assign O_1_1_0 = I_1_1_0; // @[Passthrough.scala 17:68]
  assign O_1_1_1 = I_1_1_1; // @[Passthrough.scala 17:68]
  assign O_1_1_2 = I_1_1_2; // @[Passthrough.scala 17:68]
  assign O_1_2_0 = I_1_2_0; // @[Passthrough.scala 17:68]
  assign O_1_2_1 = I_1_2_1; // @[Passthrough.scala 17:68]
  assign O_1_2_2 = I_1_2_2; // @[Passthrough.scala 17:68]
  assign O_2_0_0 = I_2_0_0; // @[Passthrough.scala 17:68]
  assign O_2_0_1 = I_2_0_1; // @[Passthrough.scala 17:68]
  assign O_2_0_2 = I_2_0_2; // @[Passthrough.scala 17:68]
  assign O_2_1_0 = I_2_1_0; // @[Passthrough.scala 17:68]
  assign O_2_1_1 = I_2_1_1; // @[Passthrough.scala 17:68]
  assign O_2_1_2 = I_2_1_2; // @[Passthrough.scala 17:68]
  assign O_2_2_0 = I_2_2_0; // @[Passthrough.scala 17:68]
  assign O_2_2_1 = I_2_2_1; // @[Passthrough.scala 17:68]
  assign O_2_2_2 = I_2_2_2; // @[Passthrough.scala 17:68]
  assign O_3_0_0 = I_3_0_0; // @[Passthrough.scala 17:68]
  assign O_3_0_1 = I_3_0_1; // @[Passthrough.scala 17:68]
  assign O_3_0_2 = I_3_0_2; // @[Passthrough.scala 17:68]
  assign O_3_1_0 = I_3_1_0; // @[Passthrough.scala 17:68]
  assign O_3_1_1 = I_3_1_1; // @[Passthrough.scala 17:68]
  assign O_3_1_2 = I_3_1_2; // @[Passthrough.scala 17:68]
  assign O_3_2_0 = I_3_2_0; // @[Passthrough.scala 17:68]
  assign O_3_2_1 = I_3_2_1; // @[Passthrough.scala 17:68]
  assign O_3_2_2 = I_3_2_2; // @[Passthrough.scala 17:68]
  assign O_4_0_0 = I_4_0_0; // @[Passthrough.scala 17:68]
  assign O_4_0_1 = I_4_0_1; // @[Passthrough.scala 17:68]
  assign O_4_0_2 = I_4_0_2; // @[Passthrough.scala 17:68]
  assign O_4_1_0 = I_4_1_0; // @[Passthrough.scala 17:68]
  assign O_4_1_1 = I_4_1_1; // @[Passthrough.scala 17:68]
  assign O_4_1_2 = I_4_1_2; // @[Passthrough.scala 17:68]
  assign O_4_2_0 = I_4_2_0; // @[Passthrough.scala 17:68]
  assign O_4_2_1 = I_4_2_1; // @[Passthrough.scala 17:68]
  assign O_4_2_2 = I_4_2_2; // @[Passthrough.scala 17:68]
  assign O_5_0_0 = I_5_0_0; // @[Passthrough.scala 17:68]
  assign O_5_0_1 = I_5_0_1; // @[Passthrough.scala 17:68]
  assign O_5_0_2 = I_5_0_2; // @[Passthrough.scala 17:68]
  assign O_5_1_0 = I_5_1_0; // @[Passthrough.scala 17:68]
  assign O_5_1_1 = I_5_1_1; // @[Passthrough.scala 17:68]
  assign O_5_1_2 = I_5_1_2; // @[Passthrough.scala 17:68]
  assign O_5_2_0 = I_5_2_0; // @[Passthrough.scala 17:68]
  assign O_5_2_1 = I_5_2_1; // @[Passthrough.scala 17:68]
  assign O_5_2_2 = I_5_2_2; // @[Passthrough.scala 17:68]
  assign O_6_0_0 = I_6_0_0; // @[Passthrough.scala 17:68]
  assign O_6_0_1 = I_6_0_1; // @[Passthrough.scala 17:68]
  assign O_6_0_2 = I_6_0_2; // @[Passthrough.scala 17:68]
  assign O_6_1_0 = I_6_1_0; // @[Passthrough.scala 17:68]
  assign O_6_1_1 = I_6_1_1; // @[Passthrough.scala 17:68]
  assign O_6_1_2 = I_6_1_2; // @[Passthrough.scala 17:68]
  assign O_6_2_0 = I_6_2_0; // @[Passthrough.scala 17:68]
  assign O_6_2_1 = I_6_2_1; // @[Passthrough.scala 17:68]
  assign O_6_2_2 = I_6_2_2; // @[Passthrough.scala 17:68]
  assign O_7_0_0 = I_7_0_0; // @[Passthrough.scala 17:68]
  assign O_7_0_1 = I_7_0_1; // @[Passthrough.scala 17:68]
  assign O_7_0_2 = I_7_0_2; // @[Passthrough.scala 17:68]
  assign O_7_1_0 = I_7_1_0; // @[Passthrough.scala 17:68]
  assign O_7_1_1 = I_7_1_1; // @[Passthrough.scala 17:68]
  assign O_7_1_2 = I_7_1_2; // @[Passthrough.scala 17:68]
  assign O_7_2_0 = I_7_2_0; // @[Passthrough.scala 17:68]
  assign O_7_2_1 = I_7_2_1; // @[Passthrough.scala 17:68]
  assign O_7_2_2 = I_7_2_2; // @[Passthrough.scala 17:68]
endmodule
module Counter_T(
  input         clock,
  input         reset,
  output [31:0] O
);
  reg [31:0] counter_value; // @[Counter.scala 53:30]
  reg [31:0] _RAND_0;
  wire  _T; // @[Counter.scala 61:49]
  wire [31:0] _T_3; // @[Counter.scala 63:70]
  assign _T = counter_value == 32'hef8; // @[Counter.scala 61:49]
  assign _T_3 = counter_value + 32'h8; // @[Counter.scala 63:70]
  assign O = counter_value; // @[Counter.scala 66:5]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  counter_value = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      counter_value <= 32'h0;
    end else if (_T) begin
      counter_value <= 32'h0;
    end else begin
      counter_value <= _T_3;
    end
  end
endmodule
module Counter_TS(
  input         clock,
  input         reset,
  output [31:0] O_0,
  output [31:0] O_1,
  output [31:0] O_2,
  output [31:0] O_3,
  output [31:0] O_4,
  output [31:0] O_5,
  output [31:0] O_6,
  output [31:0] O_7
);
  wire  counter_t_clock; // @[Counter.scala 84:25]
  wire  counter_t_reset; // @[Counter.scala 84:25]
  wire [31:0] counter_t_O; // @[Counter.scala 84:25]
  wire [32:0] _T; // @[Counter.scala 95:49]
  Counter_T counter_t ( // @[Counter.scala 84:25]
    .clock(counter_t_clock),
    .reset(counter_t_reset),
    .O(counter_t_O)
  );
  assign _T = {{1'd0}, counter_t_O}; // @[Counter.scala 95:49]
  assign O_0 = _T[31:0]; // @[Counter.scala 95:12]
  assign O_1 = 32'h1 + counter_t_O; // @[Counter.scala 95:12]
  assign O_2 = 32'h2 + counter_t_O; // @[Counter.scala 95:12]
  assign O_3 = 32'h3 + counter_t_O; // @[Counter.scala 95:12]
  assign O_4 = 32'h4 + counter_t_O; // @[Counter.scala 95:12]
  assign O_5 = 32'h5 + counter_t_O; // @[Counter.scala 95:12]
  assign O_6 = 32'h6 + counter_t_O; // @[Counter.scala 95:12]
  assign O_7 = 32'h7 + counter_t_O; // @[Counter.scala 95:12]
  assign counter_t_clock = clock;
  assign counter_t_reset = reset;
endmodule
module AtomTuple(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0,
  input  [31:0] I1,
  output [31:0] O_t0b,
  output [31:0] O_t1b
);
  assign valid_down = valid_up; // @[Tuple.scala 51:14]
  assign O_t0b = I0; // @[Tuple.scala 49:9]
  assign O_t1b = I1; // @[Tuple.scala 50:9]
endmodule
module Lt(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_t0b,
  input  [31:0] I_t1b,
  output [31:0] O
);
  wire  _T; // @[Arithmetic.scala 462:25]
  assign _T = I_t0b < I_t1b; // @[Arithmetic.scala 462:25]
  assign valid_down = valid_up; // @[Arithmetic.scala 464:14]
  assign O = {{31'd0}, _T}; // @[Arithmetic.scala 462:7]
endmodule
module Not(
  input   valid_up,
  output  valid_down,
  input   I,
  output  O
);
  assign valid_down = valid_up; // @[Arithmetic.scala 45:14]
  assign O = ~I; // @[Arithmetic.scala 44:5]
endmodule
module Module_0(
  output        valid_down,
  input  [31:0] I,
  output        O
);
  wire  n112_valid_up; // @[Top.scala 18:22]
  wire  n112_valid_down; // @[Top.scala 18:22]
  wire [31:0] n112_I0; // @[Top.scala 18:22]
  wire [31:0] n112_I1; // @[Top.scala 18:22]
  wire [31:0] n112_O_t0b; // @[Top.scala 18:22]
  wire [31:0] n112_O_t1b; // @[Top.scala 18:22]
  wire  n113_valid_up; // @[Top.scala 22:22]
  wire  n113_valid_down; // @[Top.scala 22:22]
  wire [31:0] n113_I_t0b; // @[Top.scala 22:22]
  wire [31:0] n113_I_t1b; // @[Top.scala 22:22]
  wire [31:0] n113_O; // @[Top.scala 22:22]
  wire  n114_valid_up; // @[Top.scala 25:22]
  wire  n114_valid_down; // @[Top.scala 25:22]
  wire  n114_I; // @[Top.scala 25:22]
  wire  n114_O; // @[Top.scala 25:22]
  AtomTuple n112 ( // @[Top.scala 18:22]
    .valid_up(n112_valid_up),
    .valid_down(n112_valid_down),
    .I0(n112_I0),
    .I1(n112_I1),
    .O_t0b(n112_O_t0b),
    .O_t1b(n112_O_t1b)
  );
  Lt n113 ( // @[Top.scala 22:22]
    .valid_up(n113_valid_up),
    .valid_down(n113_valid_down),
    .I_t0b(n113_I_t0b),
    .I_t1b(n113_I_t1b),
    .O(n113_O)
  );
  Not n114 ( // @[Top.scala 25:22]
    .valid_up(n114_valid_up),
    .valid_down(n114_valid_down),
    .I(n114_I),
    .O(n114_O)
  );
  assign valid_down = n114_valid_down; // @[Top.scala 29:16]
  assign O = n114_O; // @[Top.scala 28:7]
  assign n112_valid_up = 1'h1; // @[Top.scala 21:19]
  assign n112_I0 = I; // @[Top.scala 19:13]
  assign n112_I1 = 32'h780; // @[Top.scala 20:13]
  assign n113_valid_up = n112_valid_down; // @[Top.scala 24:19]
  assign n113_I_t0b = n112_O_t0b; // @[Top.scala 23:12]
  assign n113_I_t1b = n112_O_t1b; // @[Top.scala 23:12]
  assign n114_valid_up = n113_valid_down; // @[Top.scala 27:19]
  assign n114_I = n113_O[0]; // @[Top.scala 26:12]
endmodule
module MapS_4(
  output        valid_down,
  input  [31:0] I_0,
  input  [31:0] I_1,
  input  [31:0] I_2,
  input  [31:0] I_3,
  input  [31:0] I_4,
  input  [31:0] I_5,
  input  [31:0] I_6,
  input  [31:0] I_7,
  output        O_0,
  output        O_1,
  output        O_2,
  output        O_3,
  output        O_4,
  output        O_5,
  output        O_6,
  output        O_7
);
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I; // @[MapS.scala 9:22]
  wire  fst_op_O; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I; // @[MapS.scala 10:86]
  wire  other_ops_0_O; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I; // @[MapS.scala 10:86]
  wire  other_ops_1_O; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I; // @[MapS.scala 10:86]
  wire  other_ops_2_O; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I; // @[MapS.scala 10:86]
  wire  other_ops_3_O; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I; // @[MapS.scala 10:86]
  wire  other_ops_4_O; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I; // @[MapS.scala 10:86]
  wire  other_ops_5_O; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I; // @[MapS.scala 10:86]
  wire  other_ops_6_O; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  wire  _T_1; // @[MapS.scala 23:83]
  wire  _T_2; // @[MapS.scala 23:83]
  wire  _T_3; // @[MapS.scala 23:83]
  wire  _T_4; // @[MapS.scala 23:83]
  wire  _T_5; // @[MapS.scala 23:83]
  Module_0 fst_op ( // @[MapS.scala 9:22]
    .valid_down(fst_op_valid_down),
    .I(fst_op_I),
    .O(fst_op_O)
  );
  Module_0 other_ops_0 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_0_valid_down),
    .I(other_ops_0_I),
    .O(other_ops_0_O)
  );
  Module_0 other_ops_1 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_1_valid_down),
    .I(other_ops_1_I),
    .O(other_ops_1_O)
  );
  Module_0 other_ops_2 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_2_valid_down),
    .I(other_ops_2_I),
    .O(other_ops_2_O)
  );
  Module_0 other_ops_3 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_3_valid_down),
    .I(other_ops_3_I),
    .O(other_ops_3_O)
  );
  Module_0 other_ops_4 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_4_valid_down),
    .I(other_ops_4_I),
    .O(other_ops_4_O)
  );
  Module_0 other_ops_5 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_5_valid_down),
    .I(other_ops_5_I),
    .O(other_ops_5_O)
  );
  Module_0 other_ops_6 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_6_valid_down),
    .I(other_ops_6_I),
    .O(other_ops_6_O)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[MapS.scala 23:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[MapS.scala 23:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[MapS.scala 23:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[MapS.scala 23:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T_5 & other_ops_6_valid_down; // @[MapS.scala 23:14]
  assign O_0 = fst_op_O; // @[MapS.scala 17:8]
  assign O_1 = other_ops_0_O; // @[MapS.scala 21:12]
  assign O_2 = other_ops_1_O; // @[MapS.scala 21:12]
  assign O_3 = other_ops_2_O; // @[MapS.scala 21:12]
  assign O_4 = other_ops_3_O; // @[MapS.scala 21:12]
  assign O_5 = other_ops_4_O; // @[MapS.scala 21:12]
  assign O_6 = other_ops_5_O; // @[MapS.scala 21:12]
  assign O_7 = other_ops_6_O; // @[MapS.scala 21:12]
  assign fst_op_I = I_0; // @[MapS.scala 16:12]
  assign other_ops_0_I = I_1; // @[MapS.scala 20:41]
  assign other_ops_1_I = I_2; // @[MapS.scala 20:41]
  assign other_ops_2_I = I_3; // @[MapS.scala 20:41]
  assign other_ops_3_I = I_4; // @[MapS.scala 20:41]
  assign other_ops_4_I = I_5; // @[MapS.scala 20:41]
  assign other_ops_5_I = I_6; // @[MapS.scala 20:41]
  assign other_ops_6_I = I_7; // @[MapS.scala 20:41]
endmodule
module MapT_8(
  output        valid_down,
  input  [31:0] I_0,
  input  [31:0] I_1,
  input  [31:0] I_2,
  input  [31:0] I_3,
  input  [31:0] I_4,
  input  [31:0] I_5,
  input  [31:0] I_6,
  input  [31:0] I_7,
  output        O_0,
  output        O_1,
  output        O_2,
  output        O_3,
  output        O_4,
  output        O_5,
  output        O_6,
  output        O_7
);
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [31:0] op_I_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_3; // @[MapT.scala 8:20]
  wire [31:0] op_I_4; // @[MapT.scala 8:20]
  wire [31:0] op_I_5; // @[MapT.scala 8:20]
  wire [31:0] op_I_6; // @[MapT.scala 8:20]
  wire [31:0] op_I_7; // @[MapT.scala 8:20]
  wire  op_O_0; // @[MapT.scala 8:20]
  wire  op_O_1; // @[MapT.scala 8:20]
  wire  op_O_2; // @[MapT.scala 8:20]
  wire  op_O_3; // @[MapT.scala 8:20]
  wire  op_O_4; // @[MapT.scala 8:20]
  wire  op_O_5; // @[MapT.scala 8:20]
  wire  op_O_6; // @[MapT.scala 8:20]
  wire  op_O_7; // @[MapT.scala 8:20]
  MapS_4 op ( // @[MapT.scala 8:20]
    .valid_down(op_valid_down),
    .I_0(op_I_0),
    .I_1(op_I_1),
    .I_2(op_I_2),
    .I_3(op_I_3),
    .I_4(op_I_4),
    .I_5(op_I_5),
    .I_6(op_I_6),
    .I_7(op_I_7),
    .O_0(op_O_0),
    .O_1(op_O_1),
    .O_2(op_O_2),
    .O_3(op_O_3),
    .O_4(op_O_4),
    .O_5(op_O_5),
    .O_6(op_O_6),
    .O_7(op_O_7)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0 = op_O_0; // @[MapT.scala 15:7]
  assign O_1 = op_O_1; // @[MapT.scala 15:7]
  assign O_2 = op_O_2; // @[MapT.scala 15:7]
  assign O_3 = op_O_3; // @[MapT.scala 15:7]
  assign O_4 = op_O_4; // @[MapT.scala 15:7]
  assign O_5 = op_O_5; // @[MapT.scala 15:7]
  assign O_6 = op_O_6; // @[MapT.scala 15:7]
  assign O_7 = op_O_7; // @[MapT.scala 15:7]
  assign op_I_0 = I_0; // @[MapT.scala 14:10]
  assign op_I_1 = I_1; // @[MapT.scala 14:10]
  assign op_I_2 = I_2; // @[MapT.scala 14:10]
  assign op_I_3 = I_3; // @[MapT.scala 14:10]
  assign op_I_4 = I_4; // @[MapT.scala 14:10]
  assign op_I_5 = I_5; // @[MapT.scala 14:10]
  assign op_I_6 = I_6; // @[MapT.scala 14:10]
  assign op_I_7 = I_7; // @[MapT.scala 14:10]
endmodule
module AtomTuple_1(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0,
  input  [7:0]  I1,
  output [31:0] O_t0b,
  output [7:0]  O_t1b
);
  assign valid_down = valid_up; // @[Tuple.scala 51:14]
  assign O_t0b = I0; // @[Tuple.scala 49:9]
  assign O_t1b = I1; // @[Tuple.scala 50:9]
endmodule
module RShift(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_t0b,
  input  [7:0]  I_t1b,
  output [31:0] O
);
  assign valid_down = valid_up; // @[Arithmetic.scala 402:14]
  assign O = I_t0b >> I_t1b; // @[Arithmetic.scala 400:7]
endmodule
module LShift(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_t0b,
  input  [7:0]  I_t1b,
  output [31:0] O
);
  wire [286:0] _GEN_0; // @[Arithmetic.scala 431:25]
  wire [286:0] _T; // @[Arithmetic.scala 431:25]
  assign _GEN_0 = {{255'd0}, I_t0b}; // @[Arithmetic.scala 431:25]
  assign _T = _GEN_0 << I_t1b; // @[Arithmetic.scala 431:25]
  assign valid_down = valid_up; // @[Arithmetic.scala 433:14]
  assign O = _T[31:0]; // @[Arithmetic.scala 431:7]
endmodule
module Eq(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_t0b,
  input  [31:0] I_t1b,
  output [31:0] O
);
  wire  _T; // @[Arithmetic.scala 494:25]
  assign _T = I_t0b == I_t1b; // @[Arithmetic.scala 494:25]
  assign valid_down = valid_up; // @[Arithmetic.scala 496:14]
  assign O = {{31'd0}, _T}; // @[Arithmetic.scala 494:7]
endmodule
module Module_1(
  output        valid_down,
  input  [31:0] I,
  output        O
);
  wire  n120_valid_up; // @[Top.scala 36:22]
  wire  n120_valid_down; // @[Top.scala 36:22]
  wire [31:0] n120_I0; // @[Top.scala 36:22]
  wire [7:0] n120_I1; // @[Top.scala 36:22]
  wire [31:0] n120_O_t0b; // @[Top.scala 36:22]
  wire [7:0] n120_O_t1b; // @[Top.scala 36:22]
  wire  n121_valid_up; // @[Top.scala 40:22]
  wire  n121_valid_down; // @[Top.scala 40:22]
  wire [31:0] n121_I_t0b; // @[Top.scala 40:22]
  wire [7:0] n121_I_t1b; // @[Top.scala 40:22]
  wire [31:0] n121_O; // @[Top.scala 40:22]
  wire  n122_valid_up; // @[Top.scala 43:22]
  wire  n122_valid_down; // @[Top.scala 43:22]
  wire [31:0] n122_I0; // @[Top.scala 43:22]
  wire [7:0] n122_I1; // @[Top.scala 43:22]
  wire [31:0] n122_O_t0b; // @[Top.scala 43:22]
  wire [7:0] n122_O_t1b; // @[Top.scala 43:22]
  wire  n123_valid_up; // @[Top.scala 47:22]
  wire  n123_valid_down; // @[Top.scala 47:22]
  wire [31:0] n123_I_t0b; // @[Top.scala 47:22]
  wire [7:0] n123_I_t1b; // @[Top.scala 47:22]
  wire [31:0] n123_O; // @[Top.scala 47:22]
  wire  n124_valid_up; // @[Top.scala 50:22]
  wire  n124_valid_down; // @[Top.scala 50:22]
  wire [31:0] n124_I0; // @[Top.scala 50:22]
  wire [31:0] n124_I1; // @[Top.scala 50:22]
  wire [31:0] n124_O_t0b; // @[Top.scala 50:22]
  wire [31:0] n124_O_t1b; // @[Top.scala 50:22]
  wire  n125_valid_up; // @[Top.scala 54:22]
  wire  n125_valid_down; // @[Top.scala 54:22]
  wire [31:0] n125_I_t0b; // @[Top.scala 54:22]
  wire [31:0] n125_I_t1b; // @[Top.scala 54:22]
  wire [31:0] n125_O; // @[Top.scala 54:22]
  wire  n126_valid_up; // @[Top.scala 57:22]
  wire  n126_valid_down; // @[Top.scala 57:22]
  wire  n126_I; // @[Top.scala 57:22]
  wire  n126_O; // @[Top.scala 57:22]
  AtomTuple_1 n120 ( // @[Top.scala 36:22]
    .valid_up(n120_valid_up),
    .valid_down(n120_valid_down),
    .I0(n120_I0),
    .I1(n120_I1),
    .O_t0b(n120_O_t0b),
    .O_t1b(n120_O_t1b)
  );
  RShift n121 ( // @[Top.scala 40:22]
    .valid_up(n121_valid_up),
    .valid_down(n121_valid_down),
    .I_t0b(n121_I_t0b),
    .I_t1b(n121_I_t1b),
    .O(n121_O)
  );
  AtomTuple_1 n122 ( // @[Top.scala 43:22]
    .valid_up(n122_valid_up),
    .valid_down(n122_valid_down),
    .I0(n122_I0),
    .I1(n122_I1),
    .O_t0b(n122_O_t0b),
    .O_t1b(n122_O_t1b)
  );
  LShift n123 ( // @[Top.scala 47:22]
    .valid_up(n123_valid_up),
    .valid_down(n123_valid_down),
    .I_t0b(n123_I_t0b),
    .I_t1b(n123_I_t1b),
    .O(n123_O)
  );
  AtomTuple n124 ( // @[Top.scala 50:22]
    .valid_up(n124_valid_up),
    .valid_down(n124_valid_down),
    .I0(n124_I0),
    .I1(n124_I1),
    .O_t0b(n124_O_t0b),
    .O_t1b(n124_O_t1b)
  );
  Eq n125 ( // @[Top.scala 54:22]
    .valid_up(n125_valid_up),
    .valid_down(n125_valid_down),
    .I_t0b(n125_I_t0b),
    .I_t1b(n125_I_t1b),
    .O(n125_O)
  );
  Not n126 ( // @[Top.scala 57:22]
    .valid_up(n126_valid_up),
    .valid_down(n126_valid_down),
    .I(n126_I),
    .O(n126_O)
  );
  assign valid_down = n126_valid_down; // @[Top.scala 61:16]
  assign O = n126_O; // @[Top.scala 60:7]
  assign n120_valid_up = 1'h1; // @[Top.scala 39:19]
  assign n120_I0 = I; // @[Top.scala 37:13]
  assign n120_I1 = 8'h1; // @[Top.scala 38:13]
  assign n121_valid_up = n120_valid_down; // @[Top.scala 42:19]
  assign n121_I_t0b = n120_O_t0b; // @[Top.scala 41:12]
  assign n121_I_t1b = n120_O_t1b; // @[Top.scala 41:12]
  assign n122_valid_up = n121_valid_down; // @[Top.scala 46:19]
  assign n122_I0 = n121_O; // @[Top.scala 44:13]
  assign n122_I1 = 8'h1; // @[Top.scala 45:13]
  assign n123_valid_up = n122_valid_down; // @[Top.scala 49:19]
  assign n123_I_t0b = n122_O_t0b; // @[Top.scala 48:12]
  assign n123_I_t1b = n122_O_t1b; // @[Top.scala 48:12]
  assign n124_valid_up = n123_valid_down; // @[Top.scala 53:19]
  assign n124_I0 = I; // @[Top.scala 51:13]
  assign n124_I1 = n123_O; // @[Top.scala 52:13]
  assign n125_valid_up = n124_valid_down; // @[Top.scala 56:19]
  assign n125_I_t0b = n124_O_t0b; // @[Top.scala 55:12]
  assign n125_I_t1b = n124_O_t1b; // @[Top.scala 55:12]
  assign n126_valid_up = n125_valid_down; // @[Top.scala 59:19]
  assign n126_I = n125_O[0]; // @[Top.scala 58:12]
endmodule
module MapS_5(
  output        valid_down,
  input  [31:0] I_0,
  input  [31:0] I_1,
  input  [31:0] I_2,
  input  [31:0] I_3,
  input  [31:0] I_4,
  input  [31:0] I_5,
  input  [31:0] I_6,
  input  [31:0] I_7,
  output        O_0,
  output        O_1,
  output        O_2,
  output        O_3,
  output        O_4,
  output        O_5,
  output        O_6,
  output        O_7
);
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I; // @[MapS.scala 9:22]
  wire  fst_op_O; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I; // @[MapS.scala 10:86]
  wire  other_ops_0_O; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I; // @[MapS.scala 10:86]
  wire  other_ops_1_O; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I; // @[MapS.scala 10:86]
  wire  other_ops_2_O; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I; // @[MapS.scala 10:86]
  wire  other_ops_3_O; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I; // @[MapS.scala 10:86]
  wire  other_ops_4_O; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I; // @[MapS.scala 10:86]
  wire  other_ops_5_O; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I; // @[MapS.scala 10:86]
  wire  other_ops_6_O; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  wire  _T_1; // @[MapS.scala 23:83]
  wire  _T_2; // @[MapS.scala 23:83]
  wire  _T_3; // @[MapS.scala 23:83]
  wire  _T_4; // @[MapS.scala 23:83]
  wire  _T_5; // @[MapS.scala 23:83]
  Module_1 fst_op ( // @[MapS.scala 9:22]
    .valid_down(fst_op_valid_down),
    .I(fst_op_I),
    .O(fst_op_O)
  );
  Module_1 other_ops_0 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_0_valid_down),
    .I(other_ops_0_I),
    .O(other_ops_0_O)
  );
  Module_1 other_ops_1 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_1_valid_down),
    .I(other_ops_1_I),
    .O(other_ops_1_O)
  );
  Module_1 other_ops_2 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_2_valid_down),
    .I(other_ops_2_I),
    .O(other_ops_2_O)
  );
  Module_1 other_ops_3 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_3_valid_down),
    .I(other_ops_3_I),
    .O(other_ops_3_O)
  );
  Module_1 other_ops_4 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_4_valid_down),
    .I(other_ops_4_I),
    .O(other_ops_4_O)
  );
  Module_1 other_ops_5 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_5_valid_down),
    .I(other_ops_5_I),
    .O(other_ops_5_O)
  );
  Module_1 other_ops_6 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_6_valid_down),
    .I(other_ops_6_I),
    .O(other_ops_6_O)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[MapS.scala 23:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[MapS.scala 23:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[MapS.scala 23:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[MapS.scala 23:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T_5 & other_ops_6_valid_down; // @[MapS.scala 23:14]
  assign O_0 = fst_op_O; // @[MapS.scala 17:8]
  assign O_1 = other_ops_0_O; // @[MapS.scala 21:12]
  assign O_2 = other_ops_1_O; // @[MapS.scala 21:12]
  assign O_3 = other_ops_2_O; // @[MapS.scala 21:12]
  assign O_4 = other_ops_3_O; // @[MapS.scala 21:12]
  assign O_5 = other_ops_4_O; // @[MapS.scala 21:12]
  assign O_6 = other_ops_5_O; // @[MapS.scala 21:12]
  assign O_7 = other_ops_6_O; // @[MapS.scala 21:12]
  assign fst_op_I = I_0; // @[MapS.scala 16:12]
  assign other_ops_0_I = I_1; // @[MapS.scala 20:41]
  assign other_ops_1_I = I_2; // @[MapS.scala 20:41]
  assign other_ops_2_I = I_3; // @[MapS.scala 20:41]
  assign other_ops_3_I = I_4; // @[MapS.scala 20:41]
  assign other_ops_4_I = I_5; // @[MapS.scala 20:41]
  assign other_ops_5_I = I_6; // @[MapS.scala 20:41]
  assign other_ops_6_I = I_7; // @[MapS.scala 20:41]
endmodule
module MapT_9(
  output        valid_down,
  input  [31:0] I_0,
  input  [31:0] I_1,
  input  [31:0] I_2,
  input  [31:0] I_3,
  input  [31:0] I_4,
  input  [31:0] I_5,
  input  [31:0] I_6,
  input  [31:0] I_7,
  output        O_0,
  output        O_1,
  output        O_2,
  output        O_3,
  output        O_4,
  output        O_5,
  output        O_6,
  output        O_7
);
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [31:0] op_I_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_3; // @[MapT.scala 8:20]
  wire [31:0] op_I_4; // @[MapT.scala 8:20]
  wire [31:0] op_I_5; // @[MapT.scala 8:20]
  wire [31:0] op_I_6; // @[MapT.scala 8:20]
  wire [31:0] op_I_7; // @[MapT.scala 8:20]
  wire  op_O_0; // @[MapT.scala 8:20]
  wire  op_O_1; // @[MapT.scala 8:20]
  wire  op_O_2; // @[MapT.scala 8:20]
  wire  op_O_3; // @[MapT.scala 8:20]
  wire  op_O_4; // @[MapT.scala 8:20]
  wire  op_O_5; // @[MapT.scala 8:20]
  wire  op_O_6; // @[MapT.scala 8:20]
  wire  op_O_7; // @[MapT.scala 8:20]
  MapS_5 op ( // @[MapT.scala 8:20]
    .valid_down(op_valid_down),
    .I_0(op_I_0),
    .I_1(op_I_1),
    .I_2(op_I_2),
    .I_3(op_I_3),
    .I_4(op_I_4),
    .I_5(op_I_5),
    .I_6(op_I_6),
    .I_7(op_I_7),
    .O_0(op_O_0),
    .O_1(op_O_1),
    .O_2(op_O_2),
    .O_3(op_O_3),
    .O_4(op_O_4),
    .O_5(op_O_5),
    .O_6(op_O_6),
    .O_7(op_O_7)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0 = op_O_0; // @[MapT.scala 15:7]
  assign O_1 = op_O_1; // @[MapT.scala 15:7]
  assign O_2 = op_O_2; // @[MapT.scala 15:7]
  assign O_3 = op_O_3; // @[MapT.scala 15:7]
  assign O_4 = op_O_4; // @[MapT.scala 15:7]
  assign O_5 = op_O_5; // @[MapT.scala 15:7]
  assign O_6 = op_O_6; // @[MapT.scala 15:7]
  assign O_7 = op_O_7; // @[MapT.scala 15:7]
  assign op_I_0 = I_0; // @[MapT.scala 14:10]
  assign op_I_1 = I_1; // @[MapT.scala 14:10]
  assign op_I_2 = I_2; // @[MapT.scala 14:10]
  assign op_I_3 = I_3; // @[MapT.scala 14:10]
  assign op_I_4 = I_4; // @[MapT.scala 14:10]
  assign op_I_5 = I_5; // @[MapT.scala 14:10]
  assign op_I_6 = I_6; // @[MapT.scala 14:10]
  assign op_I_7 = I_7; // @[MapT.scala 14:10]
endmodule
module AtomTuple_4(
  input   valid_up,
  output  valid_down,
  input   I0,
  input   I1,
  output  O_t0b,
  output  O_t1b
);
  assign valid_down = valid_up; // @[Tuple.scala 51:14]
  assign O_t0b = I0; // @[Tuple.scala 49:9]
  assign O_t1b = I1; // @[Tuple.scala 50:9]
endmodule
module Map2S_8(
  input   valid_up,
  output  valid_down,
  input   I0_0,
  input   I0_1,
  input   I0_2,
  input   I0_3,
  input   I0_4,
  input   I0_5,
  input   I0_6,
  input   I0_7,
  input   I1_0,
  input   I1_1,
  input   I1_2,
  input   I1_3,
  input   I1_4,
  input   I1_5,
  input   I1_6,
  input   I1_7,
  output  O_0_t0b,
  output  O_0_t1b,
  output  O_1_t0b,
  output  O_1_t1b,
  output  O_2_t0b,
  output  O_2_t1b,
  output  O_3_t0b,
  output  O_3_t1b,
  output  O_4_t0b,
  output  O_4_t1b,
  output  O_5_t0b,
  output  O_5_t1b,
  output  O_6_t0b,
  output  O_6_t1b,
  output  O_7_t0b,
  output  O_7_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire  fst_op_I0; // @[Map2S.scala 9:22]
  wire  fst_op_I1; // @[Map2S.scala 9:22]
  wire  fst_op_O_t0b; // @[Map2S.scala 9:22]
  wire  fst_op_O_t1b; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire  other_ops_0_I0; // @[Map2S.scala 10:86]
  wire  other_ops_0_I1; // @[Map2S.scala 10:86]
  wire  other_ops_0_O_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_0_O_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire  other_ops_1_I0; // @[Map2S.scala 10:86]
  wire  other_ops_1_I1; // @[Map2S.scala 10:86]
  wire  other_ops_1_O_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_1_O_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire  other_ops_2_I0; // @[Map2S.scala 10:86]
  wire  other_ops_2_I1; // @[Map2S.scala 10:86]
  wire  other_ops_2_O_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_2_O_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_down; // @[Map2S.scala 10:86]
  wire  other_ops_3_I0; // @[Map2S.scala 10:86]
  wire  other_ops_3_I1; // @[Map2S.scala 10:86]
  wire  other_ops_3_O_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_3_O_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_down; // @[Map2S.scala 10:86]
  wire  other_ops_4_I0; // @[Map2S.scala 10:86]
  wire  other_ops_4_I1; // @[Map2S.scala 10:86]
  wire  other_ops_4_O_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_4_O_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_down; // @[Map2S.scala 10:86]
  wire  other_ops_5_I0; // @[Map2S.scala 10:86]
  wire  other_ops_5_I1; // @[Map2S.scala 10:86]
  wire  other_ops_5_O_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_5_O_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_down; // @[Map2S.scala 10:86]
  wire  other_ops_6_I0; // @[Map2S.scala 10:86]
  wire  other_ops_6_I1; // @[Map2S.scala 10:86]
  wire  other_ops_6_O_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_6_O_t1b; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  wire  _T_2; // @[Map2S.scala 26:83]
  wire  _T_3; // @[Map2S.scala 26:83]
  wire  _T_4; // @[Map2S.scala 26:83]
  wire  _T_5; // @[Map2S.scala 26:83]
  AtomTuple_4 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1(fst_op_I1),
    .O_t0b(fst_op_O_t0b),
    .O_t1b(fst_op_O_t1b)
  );
  AtomTuple_4 other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0(other_ops_0_I0),
    .I1(other_ops_0_I1),
    .O_t0b(other_ops_0_O_t0b),
    .O_t1b(other_ops_0_O_t1b)
  );
  AtomTuple_4 other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0(other_ops_1_I0),
    .I1(other_ops_1_I1),
    .O_t0b(other_ops_1_O_t0b),
    .O_t1b(other_ops_1_O_t1b)
  );
  AtomTuple_4 other_ops_2 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0(other_ops_2_I0),
    .I1(other_ops_2_I1),
    .O_t0b(other_ops_2_O_t0b),
    .O_t1b(other_ops_2_O_t1b)
  );
  AtomTuple_4 other_ops_3 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I0(other_ops_3_I0),
    .I1(other_ops_3_I1),
    .O_t0b(other_ops_3_O_t0b),
    .O_t1b(other_ops_3_O_t1b)
  );
  AtomTuple_4 other_ops_4 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I0(other_ops_4_I0),
    .I1(other_ops_4_I1),
    .O_t0b(other_ops_4_O_t0b),
    .O_t1b(other_ops_4_O_t1b)
  );
  AtomTuple_4 other_ops_5 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I0(other_ops_5_I0),
    .I1(other_ops_5_I1),
    .O_t0b(other_ops_5_O_t0b),
    .O_t1b(other_ops_5_O_t1b)
  );
  AtomTuple_4 other_ops_6 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I0(other_ops_6_I0),
    .I1(other_ops_6_I1),
    .O_t0b(other_ops_6_O_t0b),
    .O_t1b(other_ops_6_O_t1b)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[Map2S.scala 26:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[Map2S.scala 26:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_5 & other_ops_6_valid_down; // @[Map2S.scala 26:14]
  assign O_0_t0b = fst_op_O_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b = fst_op_O_t1b; // @[Map2S.scala 19:8]
  assign O_1_t0b = other_ops_0_O_t0b; // @[Map2S.scala 24:12]
  assign O_1_t1b = other_ops_0_O_t1b; // @[Map2S.scala 24:12]
  assign O_2_t0b = other_ops_1_O_t0b; // @[Map2S.scala 24:12]
  assign O_2_t1b = other_ops_1_O_t1b; // @[Map2S.scala 24:12]
  assign O_3_t0b = other_ops_2_O_t0b; // @[Map2S.scala 24:12]
  assign O_3_t1b = other_ops_2_O_t1b; // @[Map2S.scala 24:12]
  assign O_4_t0b = other_ops_3_O_t0b; // @[Map2S.scala 24:12]
  assign O_4_t1b = other_ops_3_O_t1b; // @[Map2S.scala 24:12]
  assign O_5_t0b = other_ops_4_O_t0b; // @[Map2S.scala 24:12]
  assign O_5_t1b = other_ops_4_O_t1b; // @[Map2S.scala 24:12]
  assign O_6_t0b = other_ops_5_O_t0b; // @[Map2S.scala 24:12]
  assign O_6_t1b = other_ops_5_O_t1b; // @[Map2S.scala 24:12]
  assign O_7_t0b = other_ops_6_O_t0b; // @[Map2S.scala 24:12]
  assign O_7_t1b = other_ops_6_O_t1b; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0 = I0_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I1 = I1_1; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0 = I0_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1 = I1_2; // @[Map2S.scala 23:43]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0 = I0_3; // @[Map2S.scala 22:43]
  assign other_ops_2_I1 = I1_3; // @[Map2S.scala 23:43]
  assign other_ops_3_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_3_I0 = I0_4; // @[Map2S.scala 22:43]
  assign other_ops_3_I1 = I1_4; // @[Map2S.scala 23:43]
  assign other_ops_4_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_4_I0 = I0_5; // @[Map2S.scala 22:43]
  assign other_ops_4_I1 = I1_5; // @[Map2S.scala 23:43]
  assign other_ops_5_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_5_I0 = I0_6; // @[Map2S.scala 22:43]
  assign other_ops_5_I1 = I1_6; // @[Map2S.scala 23:43]
  assign other_ops_6_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_6_I0 = I0_7; // @[Map2S.scala 22:43]
  assign other_ops_6_I1 = I1_7; // @[Map2S.scala 23:43]
endmodule
module Map2T_8(
  input   valid_up,
  output  valid_down,
  input   I0_0,
  input   I0_1,
  input   I0_2,
  input   I0_3,
  input   I0_4,
  input   I0_5,
  input   I0_6,
  input   I0_7,
  input   I1_0,
  input   I1_1,
  input   I1_2,
  input   I1_3,
  input   I1_4,
  input   I1_5,
  input   I1_6,
  input   I1_7,
  output  O_0_t0b,
  output  O_0_t1b,
  output  O_1_t0b,
  output  O_1_t1b,
  output  O_2_t0b,
  output  O_2_t1b,
  output  O_3_t0b,
  output  O_3_t1b,
  output  O_4_t0b,
  output  O_4_t1b,
  output  O_5_t0b,
  output  O_5_t1b,
  output  O_6_t0b,
  output  O_6_t1b,
  output  O_7_t0b,
  output  O_7_t1b
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire  op_I0_0; // @[Map2T.scala 8:20]
  wire  op_I0_1; // @[Map2T.scala 8:20]
  wire  op_I0_2; // @[Map2T.scala 8:20]
  wire  op_I0_3; // @[Map2T.scala 8:20]
  wire  op_I0_4; // @[Map2T.scala 8:20]
  wire  op_I0_5; // @[Map2T.scala 8:20]
  wire  op_I0_6; // @[Map2T.scala 8:20]
  wire  op_I0_7; // @[Map2T.scala 8:20]
  wire  op_I1_0; // @[Map2T.scala 8:20]
  wire  op_I1_1; // @[Map2T.scala 8:20]
  wire  op_I1_2; // @[Map2T.scala 8:20]
  wire  op_I1_3; // @[Map2T.scala 8:20]
  wire  op_I1_4; // @[Map2T.scala 8:20]
  wire  op_I1_5; // @[Map2T.scala 8:20]
  wire  op_I1_6; // @[Map2T.scala 8:20]
  wire  op_I1_7; // @[Map2T.scala 8:20]
  wire  op_O_0_t0b; // @[Map2T.scala 8:20]
  wire  op_O_0_t1b; // @[Map2T.scala 8:20]
  wire  op_O_1_t0b; // @[Map2T.scala 8:20]
  wire  op_O_1_t1b; // @[Map2T.scala 8:20]
  wire  op_O_2_t0b; // @[Map2T.scala 8:20]
  wire  op_O_2_t1b; // @[Map2T.scala 8:20]
  wire  op_O_3_t0b; // @[Map2T.scala 8:20]
  wire  op_O_3_t1b; // @[Map2T.scala 8:20]
  wire  op_O_4_t0b; // @[Map2T.scala 8:20]
  wire  op_O_4_t1b; // @[Map2T.scala 8:20]
  wire  op_O_5_t0b; // @[Map2T.scala 8:20]
  wire  op_O_5_t1b; // @[Map2T.scala 8:20]
  wire  op_O_6_t0b; // @[Map2T.scala 8:20]
  wire  op_O_6_t1b; // @[Map2T.scala 8:20]
  wire  op_O_7_t0b; // @[Map2T.scala 8:20]
  wire  op_O_7_t1b; // @[Map2T.scala 8:20]
  Map2S_8 op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0(op_I0_0),
    .I0_1(op_I0_1),
    .I0_2(op_I0_2),
    .I0_3(op_I0_3),
    .I0_4(op_I0_4),
    .I0_5(op_I0_5),
    .I0_6(op_I0_6),
    .I0_7(op_I0_7),
    .I1_0(op_I1_0),
    .I1_1(op_I1_1),
    .I1_2(op_I1_2),
    .I1_3(op_I1_3),
    .I1_4(op_I1_4),
    .I1_5(op_I1_5),
    .I1_6(op_I1_6),
    .I1_7(op_I1_7),
    .O_0_t0b(op_O_0_t0b),
    .O_0_t1b(op_O_0_t1b),
    .O_1_t0b(op_O_1_t0b),
    .O_1_t1b(op_O_1_t1b),
    .O_2_t0b(op_O_2_t0b),
    .O_2_t1b(op_O_2_t1b),
    .O_3_t0b(op_O_3_t0b),
    .O_3_t1b(op_O_3_t1b),
    .O_4_t0b(op_O_4_t0b),
    .O_4_t1b(op_O_4_t1b),
    .O_5_t0b(op_O_5_t0b),
    .O_5_t1b(op_O_5_t1b),
    .O_6_t0b(op_O_6_t0b),
    .O_6_t1b(op_O_6_t1b),
    .O_7_t0b(op_O_7_t0b),
    .O_7_t1b(op_O_7_t1b)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_t0b = op_O_0_t0b; // @[Map2T.scala 17:7]
  assign O_0_t1b = op_O_0_t1b; // @[Map2T.scala 17:7]
  assign O_1_t0b = op_O_1_t0b; // @[Map2T.scala 17:7]
  assign O_1_t1b = op_O_1_t1b; // @[Map2T.scala 17:7]
  assign O_2_t0b = op_O_2_t0b; // @[Map2T.scala 17:7]
  assign O_2_t1b = op_O_2_t1b; // @[Map2T.scala 17:7]
  assign O_3_t0b = op_O_3_t0b; // @[Map2T.scala 17:7]
  assign O_3_t1b = op_O_3_t1b; // @[Map2T.scala 17:7]
  assign O_4_t0b = op_O_4_t0b; // @[Map2T.scala 17:7]
  assign O_4_t1b = op_O_4_t1b; // @[Map2T.scala 17:7]
  assign O_5_t0b = op_O_5_t0b; // @[Map2T.scala 17:7]
  assign O_5_t1b = op_O_5_t1b; // @[Map2T.scala 17:7]
  assign O_6_t0b = op_O_6_t0b; // @[Map2T.scala 17:7]
  assign O_6_t1b = op_O_6_t1b; // @[Map2T.scala 17:7]
  assign O_7_t0b = op_O_7_t0b; // @[Map2T.scala 17:7]
  assign O_7_t1b = op_O_7_t1b; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0 = I0_0; // @[Map2T.scala 15:11]
  assign op_I0_1 = I0_1; // @[Map2T.scala 15:11]
  assign op_I0_2 = I0_2; // @[Map2T.scala 15:11]
  assign op_I0_3 = I0_3; // @[Map2T.scala 15:11]
  assign op_I0_4 = I0_4; // @[Map2T.scala 15:11]
  assign op_I0_5 = I0_5; // @[Map2T.scala 15:11]
  assign op_I0_6 = I0_6; // @[Map2T.scala 15:11]
  assign op_I0_7 = I0_7; // @[Map2T.scala 15:11]
  assign op_I1_0 = I1_0; // @[Map2T.scala 16:11]
  assign op_I1_1 = I1_1; // @[Map2T.scala 16:11]
  assign op_I1_2 = I1_2; // @[Map2T.scala 16:11]
  assign op_I1_3 = I1_3; // @[Map2T.scala 16:11]
  assign op_I1_4 = I1_4; // @[Map2T.scala 16:11]
  assign op_I1_5 = I1_5; // @[Map2T.scala 16:11]
  assign op_I1_6 = I1_6; // @[Map2T.scala 16:11]
  assign op_I1_7 = I1_7; // @[Map2T.scala 16:11]
endmodule
module PartitionS_4(
  input   valid_up,
  output  valid_down,
  input   I_0_t0b,
  input   I_0_t1b,
  input   I_1_t0b,
  input   I_1_t1b,
  input   I_2_t0b,
  input   I_2_t1b,
  input   I_3_t0b,
  input   I_3_t1b,
  input   I_4_t0b,
  input   I_4_t1b,
  input   I_5_t0b,
  input   I_5_t1b,
  input   I_6_t0b,
  input   I_6_t1b,
  input   I_7_t0b,
  input   I_7_t1b,
  output  O_0_0_t0b,
  output  O_0_0_t1b,
  output  O_1_0_t0b,
  output  O_1_0_t1b,
  output  O_2_0_t0b,
  output  O_2_0_t1b,
  output  O_3_0_t0b,
  output  O_3_0_t1b,
  output  O_4_0_t0b,
  output  O_4_0_t1b,
  output  O_5_0_t0b,
  output  O_5_0_t1b,
  output  O_6_0_t0b,
  output  O_6_0_t1b,
  output  O_7_0_t0b,
  output  O_7_0_t1b
);
  assign valid_down = valid_up; // @[Partition.scala 18:14]
  assign O_0_0_t0b = I_0_t0b; // @[Partition.scala 15:39]
  assign O_0_0_t1b = I_0_t1b; // @[Partition.scala 15:39]
  assign O_1_0_t0b = I_1_t0b; // @[Partition.scala 15:39]
  assign O_1_0_t1b = I_1_t1b; // @[Partition.scala 15:39]
  assign O_2_0_t0b = I_2_t0b; // @[Partition.scala 15:39]
  assign O_2_0_t1b = I_2_t1b; // @[Partition.scala 15:39]
  assign O_3_0_t0b = I_3_t0b; // @[Partition.scala 15:39]
  assign O_3_0_t1b = I_3_t1b; // @[Partition.scala 15:39]
  assign O_4_0_t0b = I_4_t0b; // @[Partition.scala 15:39]
  assign O_4_0_t1b = I_4_t1b; // @[Partition.scala 15:39]
  assign O_5_0_t0b = I_5_t0b; // @[Partition.scala 15:39]
  assign O_5_0_t1b = I_5_t1b; // @[Partition.scala 15:39]
  assign O_6_0_t0b = I_6_t0b; // @[Partition.scala 15:39]
  assign O_6_0_t1b = I_6_t1b; // @[Partition.scala 15:39]
  assign O_7_0_t0b = I_7_t0b; // @[Partition.scala 15:39]
  assign O_7_0_t1b = I_7_t1b; // @[Partition.scala 15:39]
endmodule
module MapT_10(
  input   valid_up,
  output  valid_down,
  input   I_0_t0b,
  input   I_0_t1b,
  input   I_1_t0b,
  input   I_1_t1b,
  input   I_2_t0b,
  input   I_2_t1b,
  input   I_3_t0b,
  input   I_3_t1b,
  input   I_4_t0b,
  input   I_4_t1b,
  input   I_5_t0b,
  input   I_5_t1b,
  input   I_6_t0b,
  input   I_6_t1b,
  input   I_7_t0b,
  input   I_7_t1b,
  output  O_0_0_t0b,
  output  O_0_0_t1b,
  output  O_1_0_t0b,
  output  O_1_0_t1b,
  output  O_2_0_t0b,
  output  O_2_0_t1b,
  output  O_3_0_t0b,
  output  O_3_0_t1b,
  output  O_4_0_t0b,
  output  O_4_0_t1b,
  output  O_5_0_t0b,
  output  O_5_0_t1b,
  output  O_6_0_t0b,
  output  O_6_0_t1b,
  output  O_7_0_t0b,
  output  O_7_0_t1b
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire  op_I_0_t0b; // @[MapT.scala 8:20]
  wire  op_I_0_t1b; // @[MapT.scala 8:20]
  wire  op_I_1_t0b; // @[MapT.scala 8:20]
  wire  op_I_1_t1b; // @[MapT.scala 8:20]
  wire  op_I_2_t0b; // @[MapT.scala 8:20]
  wire  op_I_2_t1b; // @[MapT.scala 8:20]
  wire  op_I_3_t0b; // @[MapT.scala 8:20]
  wire  op_I_3_t1b; // @[MapT.scala 8:20]
  wire  op_I_4_t0b; // @[MapT.scala 8:20]
  wire  op_I_4_t1b; // @[MapT.scala 8:20]
  wire  op_I_5_t0b; // @[MapT.scala 8:20]
  wire  op_I_5_t1b; // @[MapT.scala 8:20]
  wire  op_I_6_t0b; // @[MapT.scala 8:20]
  wire  op_I_6_t1b; // @[MapT.scala 8:20]
  wire  op_I_7_t0b; // @[MapT.scala 8:20]
  wire  op_I_7_t1b; // @[MapT.scala 8:20]
  wire  op_O_0_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_0_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_1_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_1_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_2_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_2_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_3_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_3_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_4_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_4_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_5_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_5_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_6_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_6_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_7_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_7_0_t1b; // @[MapT.scala 8:20]
  PartitionS_4 op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_t0b(op_I_0_t0b),
    .I_0_t1b(op_I_0_t1b),
    .I_1_t0b(op_I_1_t0b),
    .I_1_t1b(op_I_1_t1b),
    .I_2_t0b(op_I_2_t0b),
    .I_2_t1b(op_I_2_t1b),
    .I_3_t0b(op_I_3_t0b),
    .I_3_t1b(op_I_3_t1b),
    .I_4_t0b(op_I_4_t0b),
    .I_4_t1b(op_I_4_t1b),
    .I_5_t0b(op_I_5_t0b),
    .I_5_t1b(op_I_5_t1b),
    .I_6_t0b(op_I_6_t0b),
    .I_6_t1b(op_I_6_t1b),
    .I_7_t0b(op_I_7_t0b),
    .I_7_t1b(op_I_7_t1b),
    .O_0_0_t0b(op_O_0_0_t0b),
    .O_0_0_t1b(op_O_0_0_t1b),
    .O_1_0_t0b(op_O_1_0_t0b),
    .O_1_0_t1b(op_O_1_0_t1b),
    .O_2_0_t0b(op_O_2_0_t0b),
    .O_2_0_t1b(op_O_2_0_t1b),
    .O_3_0_t0b(op_O_3_0_t0b),
    .O_3_0_t1b(op_O_3_0_t1b),
    .O_4_0_t0b(op_O_4_0_t0b),
    .O_4_0_t1b(op_O_4_0_t1b),
    .O_5_0_t0b(op_O_5_0_t0b),
    .O_5_0_t1b(op_O_5_0_t1b),
    .O_6_0_t0b(op_O_6_0_t0b),
    .O_6_0_t1b(op_O_6_0_t1b),
    .O_7_0_t0b(op_O_7_0_t0b),
    .O_7_0_t1b(op_O_7_0_t1b)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_t0b = op_O_0_0_t0b; // @[MapT.scala 15:7]
  assign O_0_0_t1b = op_O_0_0_t1b; // @[MapT.scala 15:7]
  assign O_1_0_t0b = op_O_1_0_t0b; // @[MapT.scala 15:7]
  assign O_1_0_t1b = op_O_1_0_t1b; // @[MapT.scala 15:7]
  assign O_2_0_t0b = op_O_2_0_t0b; // @[MapT.scala 15:7]
  assign O_2_0_t1b = op_O_2_0_t1b; // @[MapT.scala 15:7]
  assign O_3_0_t0b = op_O_3_0_t0b; // @[MapT.scala 15:7]
  assign O_3_0_t1b = op_O_3_0_t1b; // @[MapT.scala 15:7]
  assign O_4_0_t0b = op_O_4_0_t0b; // @[MapT.scala 15:7]
  assign O_4_0_t1b = op_O_4_0_t1b; // @[MapT.scala 15:7]
  assign O_5_0_t0b = op_O_5_0_t0b; // @[MapT.scala 15:7]
  assign O_5_0_t1b = op_O_5_0_t1b; // @[MapT.scala 15:7]
  assign O_6_0_t0b = op_O_6_0_t0b; // @[MapT.scala 15:7]
  assign O_6_0_t1b = op_O_6_0_t1b; // @[MapT.scala 15:7]
  assign O_7_0_t0b = op_O_7_0_t0b; // @[MapT.scala 15:7]
  assign O_7_0_t1b = op_O_7_0_t1b; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_t0b = I_0_t0b; // @[MapT.scala 14:10]
  assign op_I_0_t1b = I_0_t1b; // @[MapT.scala 14:10]
  assign op_I_1_t0b = I_1_t0b; // @[MapT.scala 14:10]
  assign op_I_1_t1b = I_1_t1b; // @[MapT.scala 14:10]
  assign op_I_2_t0b = I_2_t0b; // @[MapT.scala 14:10]
  assign op_I_2_t1b = I_2_t1b; // @[MapT.scala 14:10]
  assign op_I_3_t0b = I_3_t0b; // @[MapT.scala 14:10]
  assign op_I_3_t1b = I_3_t1b; // @[MapT.scala 14:10]
  assign op_I_4_t0b = I_4_t0b; // @[MapT.scala 14:10]
  assign op_I_4_t1b = I_4_t1b; // @[MapT.scala 14:10]
  assign op_I_5_t0b = I_5_t0b; // @[MapT.scala 14:10]
  assign op_I_5_t1b = I_5_t1b; // @[MapT.scala 14:10]
  assign op_I_6_t0b = I_6_t0b; // @[MapT.scala 14:10]
  assign op_I_6_t1b = I_6_t1b; // @[MapT.scala 14:10]
  assign op_I_7_t0b = I_7_t0b; // @[MapT.scala 14:10]
  assign op_I_7_t1b = I_7_t1b; // @[MapT.scala 14:10]
endmodule
module PartitionS_5(
  input   valid_up,
  output  valid_down,
  input   I_0_0_t0b,
  input   I_0_0_t1b,
  input   I_1_0_t0b,
  input   I_1_0_t1b,
  input   I_2_0_t0b,
  input   I_2_0_t1b,
  input   I_3_0_t0b,
  input   I_3_0_t1b,
  input   I_4_0_t0b,
  input   I_4_0_t1b,
  input   I_5_0_t0b,
  input   I_5_0_t1b,
  input   I_6_0_t0b,
  input   I_6_0_t1b,
  input   I_7_0_t0b,
  input   I_7_0_t1b,
  output  O_0_0_0_t0b,
  output  O_0_0_0_t1b,
  output  O_1_0_0_t0b,
  output  O_1_0_0_t1b,
  output  O_2_0_0_t0b,
  output  O_2_0_0_t1b,
  output  O_3_0_0_t0b,
  output  O_3_0_0_t1b,
  output  O_4_0_0_t0b,
  output  O_4_0_0_t1b,
  output  O_5_0_0_t0b,
  output  O_5_0_0_t1b,
  output  O_6_0_0_t0b,
  output  O_6_0_0_t1b,
  output  O_7_0_0_t0b,
  output  O_7_0_0_t1b
);
  assign valid_down = valid_up; // @[Partition.scala 18:14]
  assign O_0_0_0_t0b = I_0_0_t0b; // @[Partition.scala 15:39]
  assign O_0_0_0_t1b = I_0_0_t1b; // @[Partition.scala 15:39]
  assign O_1_0_0_t0b = I_1_0_t0b; // @[Partition.scala 15:39]
  assign O_1_0_0_t1b = I_1_0_t1b; // @[Partition.scala 15:39]
  assign O_2_0_0_t0b = I_2_0_t0b; // @[Partition.scala 15:39]
  assign O_2_0_0_t1b = I_2_0_t1b; // @[Partition.scala 15:39]
  assign O_3_0_0_t0b = I_3_0_t0b; // @[Partition.scala 15:39]
  assign O_3_0_0_t1b = I_3_0_t1b; // @[Partition.scala 15:39]
  assign O_4_0_0_t0b = I_4_0_t0b; // @[Partition.scala 15:39]
  assign O_4_0_0_t1b = I_4_0_t1b; // @[Partition.scala 15:39]
  assign O_5_0_0_t0b = I_5_0_t0b; // @[Partition.scala 15:39]
  assign O_5_0_0_t1b = I_5_0_t1b; // @[Partition.scala 15:39]
  assign O_6_0_0_t0b = I_6_0_t0b; // @[Partition.scala 15:39]
  assign O_6_0_0_t1b = I_6_0_t1b; // @[Partition.scala 15:39]
  assign O_7_0_0_t0b = I_7_0_t0b; // @[Partition.scala 15:39]
  assign O_7_0_0_t1b = I_7_0_t1b; // @[Partition.scala 15:39]
endmodule
module MapT_11(
  input   valid_up,
  output  valid_down,
  input   I_0_0_t0b,
  input   I_0_0_t1b,
  input   I_1_0_t0b,
  input   I_1_0_t1b,
  input   I_2_0_t0b,
  input   I_2_0_t1b,
  input   I_3_0_t0b,
  input   I_3_0_t1b,
  input   I_4_0_t0b,
  input   I_4_0_t1b,
  input   I_5_0_t0b,
  input   I_5_0_t1b,
  input   I_6_0_t0b,
  input   I_6_0_t1b,
  input   I_7_0_t0b,
  input   I_7_0_t1b,
  output  O_0_0_0_t0b,
  output  O_0_0_0_t1b,
  output  O_1_0_0_t0b,
  output  O_1_0_0_t1b,
  output  O_2_0_0_t0b,
  output  O_2_0_0_t1b,
  output  O_3_0_0_t0b,
  output  O_3_0_0_t1b,
  output  O_4_0_0_t0b,
  output  O_4_0_0_t1b,
  output  O_5_0_0_t0b,
  output  O_5_0_0_t1b,
  output  O_6_0_0_t0b,
  output  O_6_0_0_t1b,
  output  O_7_0_0_t0b,
  output  O_7_0_0_t1b
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire  op_I_0_0_t0b; // @[MapT.scala 8:20]
  wire  op_I_0_0_t1b; // @[MapT.scala 8:20]
  wire  op_I_1_0_t0b; // @[MapT.scala 8:20]
  wire  op_I_1_0_t1b; // @[MapT.scala 8:20]
  wire  op_I_2_0_t0b; // @[MapT.scala 8:20]
  wire  op_I_2_0_t1b; // @[MapT.scala 8:20]
  wire  op_I_3_0_t0b; // @[MapT.scala 8:20]
  wire  op_I_3_0_t1b; // @[MapT.scala 8:20]
  wire  op_I_4_0_t0b; // @[MapT.scala 8:20]
  wire  op_I_4_0_t1b; // @[MapT.scala 8:20]
  wire  op_I_5_0_t0b; // @[MapT.scala 8:20]
  wire  op_I_5_0_t1b; // @[MapT.scala 8:20]
  wire  op_I_6_0_t0b; // @[MapT.scala 8:20]
  wire  op_I_6_0_t1b; // @[MapT.scala 8:20]
  wire  op_I_7_0_t0b; // @[MapT.scala 8:20]
  wire  op_I_7_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_0_0_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_0_0_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_1_0_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_1_0_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_2_0_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_2_0_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_3_0_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_3_0_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_4_0_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_4_0_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_5_0_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_5_0_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_6_0_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_6_0_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_7_0_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_7_0_0_t1b; // @[MapT.scala 8:20]
  PartitionS_5 op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_t0b(op_I_0_0_t0b),
    .I_0_0_t1b(op_I_0_0_t1b),
    .I_1_0_t0b(op_I_1_0_t0b),
    .I_1_0_t1b(op_I_1_0_t1b),
    .I_2_0_t0b(op_I_2_0_t0b),
    .I_2_0_t1b(op_I_2_0_t1b),
    .I_3_0_t0b(op_I_3_0_t0b),
    .I_3_0_t1b(op_I_3_0_t1b),
    .I_4_0_t0b(op_I_4_0_t0b),
    .I_4_0_t1b(op_I_4_0_t1b),
    .I_5_0_t0b(op_I_5_0_t0b),
    .I_5_0_t1b(op_I_5_0_t1b),
    .I_6_0_t0b(op_I_6_0_t0b),
    .I_6_0_t1b(op_I_6_0_t1b),
    .I_7_0_t0b(op_I_7_0_t0b),
    .I_7_0_t1b(op_I_7_0_t1b),
    .O_0_0_0_t0b(op_O_0_0_0_t0b),
    .O_0_0_0_t1b(op_O_0_0_0_t1b),
    .O_1_0_0_t0b(op_O_1_0_0_t0b),
    .O_1_0_0_t1b(op_O_1_0_0_t1b),
    .O_2_0_0_t0b(op_O_2_0_0_t0b),
    .O_2_0_0_t1b(op_O_2_0_0_t1b),
    .O_3_0_0_t0b(op_O_3_0_0_t0b),
    .O_3_0_0_t1b(op_O_3_0_0_t1b),
    .O_4_0_0_t0b(op_O_4_0_0_t0b),
    .O_4_0_0_t1b(op_O_4_0_0_t1b),
    .O_5_0_0_t0b(op_O_5_0_0_t0b),
    .O_5_0_0_t1b(op_O_5_0_0_t1b),
    .O_6_0_0_t0b(op_O_6_0_0_t0b),
    .O_6_0_0_t1b(op_O_6_0_0_t1b),
    .O_7_0_0_t0b(op_O_7_0_0_t0b),
    .O_7_0_0_t1b(op_O_7_0_0_t1b)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0_t0b = op_O_0_0_0_t0b; // @[MapT.scala 15:7]
  assign O_0_0_0_t1b = op_O_0_0_0_t1b; // @[MapT.scala 15:7]
  assign O_1_0_0_t0b = op_O_1_0_0_t0b; // @[MapT.scala 15:7]
  assign O_1_0_0_t1b = op_O_1_0_0_t1b; // @[MapT.scala 15:7]
  assign O_2_0_0_t0b = op_O_2_0_0_t0b; // @[MapT.scala 15:7]
  assign O_2_0_0_t1b = op_O_2_0_0_t1b; // @[MapT.scala 15:7]
  assign O_3_0_0_t0b = op_O_3_0_0_t0b; // @[MapT.scala 15:7]
  assign O_3_0_0_t1b = op_O_3_0_0_t1b; // @[MapT.scala 15:7]
  assign O_4_0_0_t0b = op_O_4_0_0_t0b; // @[MapT.scala 15:7]
  assign O_4_0_0_t1b = op_O_4_0_0_t1b; // @[MapT.scala 15:7]
  assign O_5_0_0_t0b = op_O_5_0_0_t0b; // @[MapT.scala 15:7]
  assign O_5_0_0_t1b = op_O_5_0_0_t1b; // @[MapT.scala 15:7]
  assign O_6_0_0_t0b = op_O_6_0_0_t0b; // @[MapT.scala 15:7]
  assign O_6_0_0_t1b = op_O_6_0_0_t1b; // @[MapT.scala 15:7]
  assign O_7_0_0_t0b = op_O_7_0_0_t0b; // @[MapT.scala 15:7]
  assign O_7_0_0_t1b = op_O_7_0_0_t1b; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_t0b = I_0_0_t0b; // @[MapT.scala 14:10]
  assign op_I_0_0_t1b = I_0_0_t1b; // @[MapT.scala 14:10]
  assign op_I_1_0_t0b = I_1_0_t0b; // @[MapT.scala 14:10]
  assign op_I_1_0_t1b = I_1_0_t1b; // @[MapT.scala 14:10]
  assign op_I_2_0_t0b = I_2_0_t0b; // @[MapT.scala 14:10]
  assign op_I_2_0_t1b = I_2_0_t1b; // @[MapT.scala 14:10]
  assign op_I_3_0_t0b = I_3_0_t0b; // @[MapT.scala 14:10]
  assign op_I_3_0_t1b = I_3_0_t1b; // @[MapT.scala 14:10]
  assign op_I_4_0_t0b = I_4_0_t0b; // @[MapT.scala 14:10]
  assign op_I_4_0_t1b = I_4_0_t1b; // @[MapT.scala 14:10]
  assign op_I_5_0_t0b = I_5_0_t0b; // @[MapT.scala 14:10]
  assign op_I_5_0_t1b = I_5_0_t1b; // @[MapT.scala 14:10]
  assign op_I_6_0_t0b = I_6_0_t0b; // @[MapT.scala 14:10]
  assign op_I_6_0_t1b = I_6_0_t1b; // @[MapT.scala 14:10]
  assign op_I_7_0_t0b = I_7_0_t0b; // @[MapT.scala 14:10]
  assign op_I_7_0_t1b = I_7_0_t1b; // @[MapT.scala 14:10]
endmodule
module FIFO_1(
  input   clock,
  input   reset,
  input   valid_up,
  output  valid_down,
  input   I_0_0_0_t0b,
  input   I_0_0_0_t1b,
  input   I_1_0_0_t0b,
  input   I_1_0_0_t1b,
  input   I_2_0_0_t0b,
  input   I_2_0_0_t1b,
  input   I_3_0_0_t0b,
  input   I_3_0_0_t1b,
  input   I_4_0_0_t0b,
  input   I_4_0_0_t1b,
  input   I_5_0_0_t0b,
  input   I_5_0_0_t1b,
  input   I_6_0_0_t0b,
  input   I_6_0_0_t1b,
  input   I_7_0_0_t0b,
  input   I_7_0_0_t1b,
  output  O_0_0_0_t0b,
  output  O_0_0_0_t1b,
  output  O_1_0_0_t0b,
  output  O_1_0_0_t1b,
  output  O_2_0_0_t0b,
  output  O_2_0_0_t1b,
  output  O_3_0_0_t0b,
  output  O_3_0_0_t1b,
  output  O_4_0_0_t0b,
  output  O_4_0_0_t1b,
  output  O_5_0_0_t0b,
  output  O_5_0_0_t1b,
  output  O_6_0_0_t0b,
  output  O_6_0_0_t1b,
  output  O_7_0_0_t0b,
  output  O_7_0_0_t1b
);
  reg  _T__0_0_0_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_0;
  reg  _T__0_0_0_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_1;
  reg  _T__1_0_0_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_2;
  reg  _T__1_0_0_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_3;
  reg  _T__2_0_0_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_4;
  reg  _T__2_0_0_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_5;
  reg  _T__3_0_0_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_6;
  reg  _T__3_0_0_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_7;
  reg  _T__4_0_0_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_8;
  reg  _T__4_0_0_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_9;
  reg  _T__5_0_0_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_10;
  reg  _T__5_0_0_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_11;
  reg  _T__6_0_0_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_12;
  reg  _T__6_0_0_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_13;
  reg  _T__7_0_0_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_14;
  reg  _T__7_0_0_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_15;
  reg  _T_1; // @[FIFO.scala 15:27]
  reg [31:0] _RAND_16;
  assign valid_down = _T_1; // @[FIFO.scala 16:16]
  assign O_0_0_0_t0b = _T__0_0_0_t0b; // @[FIFO.scala 14:7]
  assign O_0_0_0_t1b = _T__0_0_0_t1b; // @[FIFO.scala 14:7]
  assign O_1_0_0_t0b = _T__1_0_0_t0b; // @[FIFO.scala 14:7]
  assign O_1_0_0_t1b = _T__1_0_0_t1b; // @[FIFO.scala 14:7]
  assign O_2_0_0_t0b = _T__2_0_0_t0b; // @[FIFO.scala 14:7]
  assign O_2_0_0_t1b = _T__2_0_0_t1b; // @[FIFO.scala 14:7]
  assign O_3_0_0_t0b = _T__3_0_0_t0b; // @[FIFO.scala 14:7]
  assign O_3_0_0_t1b = _T__3_0_0_t1b; // @[FIFO.scala 14:7]
  assign O_4_0_0_t0b = _T__4_0_0_t0b; // @[FIFO.scala 14:7]
  assign O_4_0_0_t1b = _T__4_0_0_t1b; // @[FIFO.scala 14:7]
  assign O_5_0_0_t0b = _T__5_0_0_t0b; // @[FIFO.scala 14:7]
  assign O_5_0_0_t1b = _T__5_0_0_t1b; // @[FIFO.scala 14:7]
  assign O_6_0_0_t0b = _T__6_0_0_t0b; // @[FIFO.scala 14:7]
  assign O_6_0_0_t1b = _T__6_0_0_t1b; // @[FIFO.scala 14:7]
  assign O_7_0_0_t0b = _T__7_0_0_t0b; // @[FIFO.scala 14:7]
  assign O_7_0_0_t1b = _T__7_0_0_t1b; // @[FIFO.scala 14:7]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T__0_0_0_t0b = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T__0_0_0_t1b = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T__1_0_0_t0b = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T__1_0_0_t1b = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T__2_0_0_t0b = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T__2_0_0_t1b = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T__3_0_0_t0b = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T__3_0_0_t1b = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T__4_0_0_t0b = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T__4_0_0_t1b = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T__5_0_0_t0b = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T__5_0_0_t1b = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T__6_0_0_t0b = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T__6_0_0_t1b = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T__7_0_0_t0b = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T__7_0_0_t1b = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_1 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T__0_0_0_t0b <= I_0_0_0_t0b;
    _T__0_0_0_t1b <= I_0_0_0_t1b;
    _T__1_0_0_t0b <= I_1_0_0_t0b;
    _T__1_0_0_t1b <= I_1_0_0_t1b;
    _T__2_0_0_t0b <= I_2_0_0_t0b;
    _T__2_0_0_t1b <= I_2_0_0_t1b;
    _T__3_0_0_t0b <= I_3_0_0_t0b;
    _T__3_0_0_t1b <= I_3_0_0_t1b;
    _T__4_0_0_t0b <= I_4_0_0_t0b;
    _T__4_0_0_t1b <= I_4_0_0_t1b;
    _T__5_0_0_t0b <= I_5_0_0_t0b;
    _T__5_0_0_t1b <= I_5_0_0_t1b;
    _T__6_0_0_t0b <= I_6_0_0_t0b;
    _T__6_0_0_t1b <= I_6_0_0_t1b;
    _T__7_0_0_t0b <= I_7_0_0_t0b;
    _T__7_0_0_t1b <= I_7_0_0_t1b;
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      _T_1 <= valid_up;
    end
  end
endmodule
module Fst(
  input   valid_up,
  output  valid_down,
  input   I_t0b,
  output  O
);
  assign valid_down = valid_up; // @[Tuple.scala 59:14]
  assign O = I_t0b; // @[Tuple.scala 58:5]
endmodule
module MapS_6(
  input   valid_up,
  output  valid_down,
  input   I_0_t0b,
  output  O_0
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire  fst_op_I_t0b; // @[MapS.scala 9:22]
  wire  fst_op_O; // @[MapS.scala 9:22]
  Fst fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_t0b(fst_op_I_t0b),
    .O(fst_op_O)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0 = fst_op_O; // @[MapS.scala 17:8]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_t0b = I_0_t0b; // @[MapS.scala 16:12]
endmodule
module MapS_7(
  input   valid_up,
  output  valid_down,
  input   I_0_0_t0b,
  output  O_0_0
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire  fst_op_I_0_t0b; // @[MapS.scala 9:22]
  wire  fst_op_O_0; // @[MapS.scala 9:22]
  MapS_6 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_t0b(fst_op_I_0_t0b),
    .O_0(fst_op_O_0)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_t0b = I_0_0_t0b; // @[MapS.scala 16:12]
endmodule
module FIFO_2(
  input   clock,
  input   reset,
  input   valid_up,
  output  valid_down,
  input   I_0_0,
  output  O_0_0
);
  reg  _T_0_0 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_0;
  wire  _T_0_0__T_15_data; // @[FIFO.scala 23:33]
  wire [1:0] _T_0_0__T_15_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_1;
  wire  _T_0_0__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T_0_0__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T_0_0__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T_0_0__T_5_en; // @[FIFO.scala 23:33]
  reg  _T_0_0__T_15_en_pipe_0;
  reg [31:0] _RAND_2;
  reg [1:0] _T_0_0__T_15_addr_pipe_0;
  reg [31:0] _RAND_3;
  reg [1:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_4;
  reg [1:0] value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  reg [1:0] value_2; // @[Counter.scala 29:33]
  reg [31:0] _RAND_6;
  wire  _T_1; // @[FIFO.scala 33:46]
  wire  _T_2; // @[Counter.scala 37:24]
  wire [1:0] _T_4; // @[Counter.scala 38:22]
  wire  _T_6; // @[FIFO.scala 38:39]
  wire [1:0] _T_9; // @[Counter.scala 38:22]
  wire  _T_10; // @[FIFO.scala 42:39]
  wire  _T_16; // @[Counter.scala 37:24]
  wire [1:0] _T_18; // @[Counter.scala 38:22]
  wire  _GEN_8; // @[FIFO.scala 42:57]
  assign _T_0_0__T_15_addr = _T_0_0__T_15_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_0_0__T_15_data = _T_0_0[_T_0_0__T_15_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T_0_0__T_15_data = _T_0_0__T_15_addr >= 2'h3 ? _RAND_1[0:0] : _T_0_0[_T_0_0__T_15_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_0_0__T_5_data = I_0_0;
  assign _T_0_0__T_5_addr = value_2;
  assign _T_0_0__T_5_mask = 1'h1;
  assign _T_0_0__T_5_en = valid_up;
  assign _T_1 = value == 2'h2; // @[FIFO.scala 33:46]
  assign _T_2 = value_2 == 2'h2; // @[Counter.scala 37:24]
  assign _T_4 = value_2 + 2'h1; // @[Counter.scala 38:22]
  assign _T_6 = value < 2'h2; // @[FIFO.scala 38:39]
  assign _T_9 = value + 2'h1; // @[Counter.scala 38:22]
  assign _T_10 = value >= 2'h1; // @[FIFO.scala 42:39]
  assign _T_16 = value_1 == 2'h2; // @[Counter.scala 37:24]
  assign _T_18 = value_1 + 2'h1; // @[Counter.scala 38:22]
  assign _GEN_8 = _T_10 & _T_10; // @[FIFO.scala 42:57]
  assign valid_down = value == 2'h2; // @[FIFO.scala 33:16]
  assign O_0_0 = _T_0_0__T_15_data; // @[FIFO.scala 43:11]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T_0_0[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_0_0__T_15_en_pipe_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_0_0__T_15_addr_pipe_0 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  value = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value_1 = _RAND_5[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  value_2 = _RAND_6[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_0_0__T_5_en & _T_0_0__T_5_mask) begin
      _T_0_0[_T_0_0__T_5_addr] <= _T_0_0__T_5_data; // @[FIFO.scala 23:33]
    end
    _T_0_0__T_15_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T_0_0__T_15_addr_pipe_0 <= value_1;
    end
    if (reset) begin
      value <= 2'h0;
    end else if (valid_up) begin
      if (_T_6) begin
        if (_T_1) begin
          value <= 2'h0;
        end else begin
          value <= _T_9;
        end
      end
    end
    if (reset) begin
      value_1 <= 2'h0;
    end else if (valid_up) begin
      if (_T_10) begin
        if (_T_16) begin
          value_1 <= 2'h0;
        end else begin
          value_1 <= _T_18;
        end
      end
    end
    if (reset) begin
      value_2 <= 2'h0;
    end else if (valid_up) begin
      if (_T_2) begin
        value_2 <= 2'h0;
      end else begin
        value_2 <= _T_4;
      end
    end
  end
endmodule
module Snd(
  input   valid_up,
  output  valid_down,
  input   I_t1b,
  output  O
);
  assign valid_down = valid_up; // @[Tuple.scala 67:14]
  assign O = I_t1b; // @[Tuple.scala 66:5]
endmodule
module MapS_8(
  input   valid_up,
  output  valid_down,
  input   I_0_t1b,
  output  O_0
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire  fst_op_I_t1b; // @[MapS.scala 9:22]
  wire  fst_op_O; // @[MapS.scala 9:22]
  Snd fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_t1b(fst_op_I_t1b),
    .O(fst_op_O)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0 = fst_op_O; // @[MapS.scala 17:8]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_t1b = I_0_t1b; // @[MapS.scala 16:12]
endmodule
module MapS_9(
  input   valid_up,
  output  valid_down,
  input   I_0_0_t1b,
  output  O_0_0
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire  fst_op_I_0_t1b; // @[MapS.scala 9:22]
  wire  fst_op_O_0; // @[MapS.scala 9:22]
  MapS_8 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_t1b(fst_op_I_0_t1b),
    .O_0(fst_op_O_0)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_t1b = I_0_0_t1b; // @[MapS.scala 16:12]
endmodule
module DownS(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_1_0,
  input  [31:0] I_1_1,
  input  [31:0] I_1_2,
  output [31:0] O_0_0,
  output [31:0] O_0_1,
  output [31:0] O_0_2
);
  assign valid_down = valid_up; // @[Downsample.scala 13:14]
  assign O_0_0 = I_1_0; // @[Downsample.scala 12:8]
  assign O_0_1 = I_1_1; // @[Downsample.scala 12:8]
  assign O_0_2 = I_1_2; // @[Downsample.scala 12:8]
endmodule
module DownS_1(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0,
  output [31:0] O_0
);
  assign valid_down = valid_up; // @[Downsample.scala 13:14]
  assign O_0 = I_0; // @[Downsample.scala 12:8]
endmodule
module MapS_10(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0,
  output [31:0] O_0_0
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_0; // @[MapS.scala 9:22]
  DownS_1 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0(fst_op_I_0),
    .O_0(fst_op_O_0)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0 = I_0_0; // @[MapS.scala 16:12]
endmodule
module DownS_2(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_2,
  output [31:0] O_0
);
  assign valid_down = valid_up; // @[Downsample.scala 13:14]
  assign O_0 = I_2; // @[Downsample.scala 12:8]
endmodule
module MapS_11(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_2,
  output [31:0] O_0_0
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_2; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_0; // @[MapS.scala 9:22]
  DownS_2 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_2(fst_op_I_2),
    .O_0(fst_op_O_0)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_2 = I_0_2; // @[MapS.scala 16:12]
endmodule
module Map2S_9(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0,
  input  [31:0] I1_0,
  output [31:0] O_0_t0b,
  output [31:0] O_0_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_t1b; // @[Map2S.scala 9:22]
  AtomTuple fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1(fst_op_I1),
    .O_t0b(fst_op_O_t0b),
    .O_t1b(fst_op_O_t1b)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_t0b = fst_op_O_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b = fst_op_O_t1b; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
endmodule
module Map2S_10(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0_0,
  input  [31:0] I1_0_0,
  output [31:0] O_0_0_t0b,
  output [31:0] O_0_0_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_t1b; // @[Map2S.scala 9:22]
  Map2S_9 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I1_0(fst_op_I1_0),
    .O_0_t0b(fst_op_O_0_t0b),
    .O_0_t1b(fst_op_O_0_t1b)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_t0b = fst_op_O_0_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_t1b = fst_op_O_0_t1b; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = I1_0_0; // @[Map2S.scala 18:13]
endmodule
module Add(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_t0b,
  input  [31:0] I_t1b,
  output [31:0] O
);
  assign valid_down = valid_up; // @[Arithmetic.scala 108:14]
  assign O = I_t0b + I_t1b; // @[Arithmetic.scala 106:7]
endmodule
module MapS_12(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_t0b,
  input  [31:0] I_0_t1b,
  output [31:0] O_0
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_t0b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_t1b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O; // @[MapS.scala 9:22]
  Add fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_t0b(fst_op_I_t0b),
    .I_t1b(fst_op_I_t1b),
    .O(fst_op_O)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0 = fst_op_O; // @[MapS.scala 17:8]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_t0b = I_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_t1b = I_0_t1b; // @[MapS.scala 16:12]
endmodule
module MapS_13(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0_t0b,
  input  [31:0] I_0_0_t1b,
  output [31:0] O_0_0
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_t0b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_t1b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_0; // @[MapS.scala 9:22]
  MapS_12 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_t0b(fst_op_I_0_t0b),
    .I_0_t1b(fst_op_I_0_t1b),
    .O_0(fst_op_O_0)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_t0b = I_0_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_0_t1b = I_0_0_t1b; // @[MapS.scala 16:12]
endmodule
module InitialDelayCounter(
  input   clock,
  input   reset,
  output  valid_down
);
  reg  value; // @[InitialDelayCounter.scala 8:34]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[InitialDelayCounter.scala 17:17]
  wire  _T_4; // @[InitialDelayCounter.scala 17:53]
  assign _T_1 = value < 1'h1; // @[InitialDelayCounter.scala 17:17]
  assign _T_4 = value + 1'h1; // @[InitialDelayCounter.scala 17:53]
  assign valid_down = value; // @[InitialDelayCounter.scala 16:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 1'h0;
    end else if (_T_1) begin
      value <= _T_4;
    end
  end
endmodule
module Module_2(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I,
  output [31:0] O_t0b,
  output [7:0]  O_t1b
);
  wire  InitialDelayCounter_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_valid_down; // @[Const.scala 11:33]
  wire  n182_valid_up; // @[Top.scala 68:22]
  wire  n182_valid_down; // @[Top.scala 68:22]
  wire [31:0] n182_I0; // @[Top.scala 68:22]
  wire [7:0] n182_I1; // @[Top.scala 68:22]
  wire [31:0] n182_O_t0b; // @[Top.scala 68:22]
  wire [7:0] n182_O_t1b; // @[Top.scala 68:22]
  InitialDelayCounter InitialDelayCounter ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_clock),
    .reset(InitialDelayCounter_reset),
    .valid_down(InitialDelayCounter_valid_down)
  );
  AtomTuple_1 n182 ( // @[Top.scala 68:22]
    .valid_up(n182_valid_up),
    .valid_down(n182_valid_down),
    .I0(n182_I0),
    .I1(n182_I1),
    .O_t0b(n182_O_t0b),
    .O_t1b(n182_O_t1b)
  );
  assign valid_down = n182_valid_down; // @[Top.scala 73:16]
  assign O_t0b = n182_O_t0b; // @[Top.scala 72:7]
  assign O_t1b = n182_O_t1b; // @[Top.scala 72:7]
  assign InitialDelayCounter_clock = clock;
  assign InitialDelayCounter_reset = reset;
  assign n182_valid_up = valid_up & InitialDelayCounter_valid_down; // @[Top.scala 71:19]
  assign n182_I0 = I; // @[Top.scala 69:13]
  assign n182_I1 = 8'h1; // @[Top.scala 70:13]
endmodule
module MapS_14(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0,
  output [31:0] O_0_t0b,
  output [7:0]  O_0_t1b
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_t1b; // @[MapS.scala 9:22]
  Module_2 fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I(fst_op_I),
    .O_t0b(fst_op_O_t0b),
    .O_t1b(fst_op_O_t1b)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0_t0b = fst_op_O_t0b; // @[MapS.scala 17:8]
  assign O_0_t1b = fst_op_O_t1b; // @[MapS.scala 17:8]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I = I_0; // @[MapS.scala 16:12]
endmodule
module MapS_15(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0,
  output [31:0] O_0_0_t0b,
  output [7:0]  O_0_0_t1b
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_0_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0_t1b; // @[MapS.scala 9:22]
  MapS_14 fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0(fst_op_I_0),
    .O_0_t0b(fst_op_O_0_t0b),
    .O_0_t1b(fst_op_O_0_t1b)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0_0_t0b = fst_op_O_0_t0b; // @[MapS.scala 17:8]
  assign O_0_0_t1b = fst_op_O_0_t1b; // @[MapS.scala 17:8]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0 = I_0_0; // @[MapS.scala 16:12]
endmodule
module MapS_16(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_t0b,
  input  [7:0]  I_0_t1b,
  output [31:0] O_0
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_t1b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O; // @[MapS.scala 9:22]
  RShift fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_t0b(fst_op_I_t0b),
    .I_t1b(fst_op_I_t1b),
    .O(fst_op_O)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0 = fst_op_O; // @[MapS.scala 17:8]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_t0b = I_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_t1b = I_0_t1b; // @[MapS.scala 16:12]
endmodule
module MapS_17(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0_t0b,
  input  [7:0]  I_0_0_t1b,
  output [31:0] O_0_0
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_t1b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_0; // @[MapS.scala 9:22]
  MapS_16 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_t0b(fst_op_I_0_t0b),
    .I_0_t1b(fst_op_I_0_t1b),
    .O_0(fst_op_O_0)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_t0b = I_0_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_0_t1b = I_0_0_t1b; // @[MapS.scala 16:12]
endmodule
module DownS_3(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_1,
  output [31:0] O_0
);
  assign valid_down = valid_up; // @[Downsample.scala 13:14]
  assign O_0 = I_1; // @[Downsample.scala 12:8]
endmodule
module MapS_18(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_1,
  output [31:0] O_0_0
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_1; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_0; // @[MapS.scala 9:22]
  DownS_3 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_1(fst_op_I_1),
    .O_0(fst_op_O_0)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_1 = I_0_1; // @[MapS.scala 16:12]
endmodule
module DownS_4(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0,
  input  [31:0] I_0_1,
  input  [31:0] I_0_2,
  output [31:0] O_0_0,
  output [31:0] O_0_1,
  output [31:0] O_0_2
);
  assign valid_down = valid_up; // @[Downsample.scala 13:14]
  assign O_0_0 = I_0_0; // @[Downsample.scala 12:8]
  assign O_0_1 = I_0_1; // @[Downsample.scala 12:8]
  assign O_0_2 = I_0_2; // @[Downsample.scala 12:8]
endmodule
module DownS_6(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_2_0,
  input  [31:0] I_2_1,
  input  [31:0] I_2_2,
  output [31:0] O_0_0,
  output [31:0] O_0_1,
  output [31:0] O_0_2
);
  assign valid_down = valid_up; // @[Downsample.scala 13:14]
  assign O_0_0 = I_2_0; // @[Downsample.scala 12:8]
  assign O_0_1 = I_2_1; // @[Downsample.scala 12:8]
  assign O_0_2 = I_2_2; // @[Downsample.scala 12:8]
endmodule
module AtomTuple_10(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0,
  input  [31:0] I1_t0b,
  input  [31:0] I1_t1b,
  output [31:0] O_t0b,
  output [31:0] O_t1b_t0b,
  output [31:0] O_t1b_t1b
);
  assign valid_down = valid_up; // @[Tuple.scala 51:14]
  assign O_t0b = I0; // @[Tuple.scala 49:9]
  assign O_t1b_t0b = I1_t0b; // @[Tuple.scala 50:9]
  assign O_t1b_t1b = I1_t1b; // @[Tuple.scala 50:9]
endmodule
module Map2S_15(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0,
  input  [31:0] I1_0_t0b,
  input  [31:0] I1_0_t1b,
  output [31:0] O_0_t0b,
  output [31:0] O_0_t1b_t0b,
  output [31:0] O_0_t1b_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_t1b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_t1b_t1b; // @[Map2S.scala 9:22]
  AtomTuple_10 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1_t0b(fst_op_I1_t0b),
    .I1_t1b(fst_op_I1_t1b),
    .O_t0b(fst_op_O_t0b),
    .O_t1b_t0b(fst_op_O_t1b_t0b),
    .O_t1b_t1b(fst_op_O_t1b_t1b)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_t0b = fst_op_O_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b_t0b = fst_op_O_t1b_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b_t1b = fst_op_O_t1b_t1b; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1_t0b = I1_0_t0b; // @[Map2S.scala 18:13]
  assign fst_op_I1_t1b = I1_0_t1b; // @[Map2S.scala 18:13]
endmodule
module Map2S_16(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0_0,
  input  [31:0] I1_0_0_t0b,
  input  [31:0] I1_0_0_t1b,
  output [31:0] O_0_0_t0b,
  output [31:0] O_0_0_t1b_t0b,
  output [31:0] O_0_0_t1b_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_0_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_0_t1b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_t1b_t1b; // @[Map2S.scala 9:22]
  Map2S_15 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I1_0_t0b(fst_op_I1_0_t0b),
    .I1_0_t1b(fst_op_I1_0_t1b),
    .O_0_t0b(fst_op_O_0_t0b),
    .O_0_t1b_t0b(fst_op_O_0_t1b_t0b),
    .O_0_t1b_t1b(fst_op_O_0_t1b_t1b)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_t0b = fst_op_O_0_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_t1b_t0b = fst_op_O_0_t1b_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_t1b_t1b = fst_op_O_0_t1b_t1b; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1_0_t0b = I1_0_0_t0b; // @[Map2S.scala 18:13]
  assign fst_op_I1_0_t1b = I1_0_0_t1b; // @[Map2S.scala 18:13]
endmodule
module FIFO_4(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0_t0b,
  input  [31:0] I_0_0_t1b_t0b,
  input  [31:0] I_0_0_t1b_t1b,
  output [31:0] O_0_0_t0b,
  output [31:0] O_0_0_t1b_t0b,
  output [31:0] O_0_0_t1b_t1b
);
  reg [31:0] _T_0_0_t0b [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_0;
  wire [31:0] _T_0_0_t0b__T_15_data; // @[FIFO.scala 23:33]
  wire [1:0] _T_0_0_t0b__T_15_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_1;
  wire [31:0] _T_0_0_t0b__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T_0_0_t0b__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T_0_0_t0b__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T_0_0_t0b__T_5_en; // @[FIFO.scala 23:33]
  reg  _T_0_0_t0b__T_15_en_pipe_0;
  reg [31:0] _RAND_2;
  reg [1:0] _T_0_0_t0b__T_15_addr_pipe_0;
  reg [31:0] _RAND_3;
  reg [31:0] _T_0_0_t1b_t0b [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_4;
  wire [31:0] _T_0_0_t1b_t0b__T_15_data; // @[FIFO.scala 23:33]
  wire [1:0] _T_0_0_t1b_t0b__T_15_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_5;
  wire [31:0] _T_0_0_t1b_t0b__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T_0_0_t1b_t0b__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T_0_0_t1b_t0b__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T_0_0_t1b_t0b__T_5_en; // @[FIFO.scala 23:33]
  reg  _T_0_0_t1b_t0b__T_15_en_pipe_0;
  reg [31:0] _RAND_6;
  reg [1:0] _T_0_0_t1b_t0b__T_15_addr_pipe_0;
  reg [31:0] _RAND_7;
  reg [31:0] _T_0_0_t1b_t1b [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_8;
  wire [31:0] _T_0_0_t1b_t1b__T_15_data; // @[FIFO.scala 23:33]
  wire [1:0] _T_0_0_t1b_t1b__T_15_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_9;
  wire [31:0] _T_0_0_t1b_t1b__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T_0_0_t1b_t1b__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T_0_0_t1b_t1b__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T_0_0_t1b_t1b__T_5_en; // @[FIFO.scala 23:33]
  reg  _T_0_0_t1b_t1b__T_15_en_pipe_0;
  reg [31:0] _RAND_10;
  reg [1:0] _T_0_0_t1b_t1b__T_15_addr_pipe_0;
  reg [31:0] _RAND_11;
  reg [1:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_12;
  reg [1:0] value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_13;
  reg [1:0] value_2; // @[Counter.scala 29:33]
  reg [31:0] _RAND_14;
  wire  _T_1; // @[FIFO.scala 33:46]
  wire  _T_2; // @[Counter.scala 37:24]
  wire [1:0] _T_4; // @[Counter.scala 38:22]
  wire  _T_6; // @[FIFO.scala 38:39]
  wire [1:0] _T_9; // @[Counter.scala 38:22]
  wire  _T_10; // @[FIFO.scala 42:39]
  wire  _T_16; // @[Counter.scala 37:24]
  wire [1:0] _T_18; // @[Counter.scala 38:22]
  wire  _GEN_8; // @[FIFO.scala 42:57]
  assign _T_0_0_t0b__T_15_addr = _T_0_0_t0b__T_15_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_0_0_t0b__T_15_data = _T_0_0_t0b[_T_0_0_t0b__T_15_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T_0_0_t0b__T_15_data = _T_0_0_t0b__T_15_addr >= 2'h3 ? _RAND_1[31:0] : _T_0_0_t0b[_T_0_0_t0b__T_15_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_0_0_t0b__T_5_data = I_0_0_t0b;
  assign _T_0_0_t0b__T_5_addr = value_2;
  assign _T_0_0_t0b__T_5_mask = 1'h1;
  assign _T_0_0_t0b__T_5_en = valid_up;
  assign _T_0_0_t1b_t0b__T_15_addr = _T_0_0_t1b_t0b__T_15_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_0_0_t1b_t0b__T_15_data = _T_0_0_t1b_t0b[_T_0_0_t1b_t0b__T_15_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T_0_0_t1b_t0b__T_15_data = _T_0_0_t1b_t0b__T_15_addr >= 2'h3 ? _RAND_5[31:0] : _T_0_0_t1b_t0b[_T_0_0_t1b_t0b__T_15_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_0_0_t1b_t0b__T_5_data = I_0_0_t1b_t0b;
  assign _T_0_0_t1b_t0b__T_5_addr = value_2;
  assign _T_0_0_t1b_t0b__T_5_mask = 1'h1;
  assign _T_0_0_t1b_t0b__T_5_en = valid_up;
  assign _T_0_0_t1b_t1b__T_15_addr = _T_0_0_t1b_t1b__T_15_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_0_0_t1b_t1b__T_15_data = _T_0_0_t1b_t1b[_T_0_0_t1b_t1b__T_15_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T_0_0_t1b_t1b__T_15_data = _T_0_0_t1b_t1b__T_15_addr >= 2'h3 ? _RAND_9[31:0] : _T_0_0_t1b_t1b[_T_0_0_t1b_t1b__T_15_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_0_0_t1b_t1b__T_5_data = I_0_0_t1b_t1b;
  assign _T_0_0_t1b_t1b__T_5_addr = value_2;
  assign _T_0_0_t1b_t1b__T_5_mask = 1'h1;
  assign _T_0_0_t1b_t1b__T_5_en = valid_up;
  assign _T_1 = value == 2'h2; // @[FIFO.scala 33:46]
  assign _T_2 = value_2 == 2'h2; // @[Counter.scala 37:24]
  assign _T_4 = value_2 + 2'h1; // @[Counter.scala 38:22]
  assign _T_6 = value < 2'h2; // @[FIFO.scala 38:39]
  assign _T_9 = value + 2'h1; // @[Counter.scala 38:22]
  assign _T_10 = value >= 2'h1; // @[FIFO.scala 42:39]
  assign _T_16 = value_1 == 2'h2; // @[Counter.scala 37:24]
  assign _T_18 = value_1 + 2'h1; // @[Counter.scala 38:22]
  assign _GEN_8 = _T_10 & _T_10; // @[FIFO.scala 42:57]
  assign valid_down = value == 2'h2; // @[FIFO.scala 33:16]
  assign O_0_0_t0b = _T_0_0_t0b__T_15_data; // @[FIFO.scala 43:11]
  assign O_0_0_t1b_t0b = _T_0_0_t1b_t0b__T_15_data; // @[FIFO.scala 43:11]
  assign O_0_0_t1b_t1b = _T_0_0_t1b_t1b__T_15_data; // @[FIFO.scala 43:11]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T_0_0_t0b[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_0_0_t0b__T_15_en_pipe_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_0_0_t0b__T_15_addr_pipe_0 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T_0_0_t1b_t0b[initvar] = _RAND_4[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_0_0_t1b_t0b__T_15_en_pipe_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_0_0_t1b_t0b__T_15_addr_pipe_0 = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T_0_0_t1b_t1b[initvar] = _RAND_8[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_9 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_0_0_t1b_t1b__T_15_en_pipe_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_0_0_t1b_t1b__T_15_addr_pipe_0 = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  value = _RAND_12[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  value_1 = _RAND_13[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  value_2 = _RAND_14[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_0_0_t0b__T_5_en & _T_0_0_t0b__T_5_mask) begin
      _T_0_0_t0b[_T_0_0_t0b__T_5_addr] <= _T_0_0_t0b__T_5_data; // @[FIFO.scala 23:33]
    end
    _T_0_0_t0b__T_15_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T_0_0_t0b__T_15_addr_pipe_0 <= value_1;
    end
    if(_T_0_0_t1b_t0b__T_5_en & _T_0_0_t1b_t0b__T_5_mask) begin
      _T_0_0_t1b_t0b[_T_0_0_t1b_t0b__T_5_addr] <= _T_0_0_t1b_t0b__T_5_data; // @[FIFO.scala 23:33]
    end
    _T_0_0_t1b_t0b__T_15_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T_0_0_t1b_t0b__T_15_addr_pipe_0 <= value_1;
    end
    if(_T_0_0_t1b_t1b__T_5_en & _T_0_0_t1b_t1b__T_5_mask) begin
      _T_0_0_t1b_t1b[_T_0_0_t1b_t1b__T_5_addr] <= _T_0_0_t1b_t1b__T_5_data; // @[FIFO.scala 23:33]
    end
    _T_0_0_t1b_t1b__T_15_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T_0_0_t1b_t1b__T_15_addr_pipe_0 <= value_1;
    end
    if (reset) begin
      value <= 2'h0;
    end else if (valid_up) begin
      if (_T_6) begin
        if (_T_1) begin
          value <= 2'h0;
        end else begin
          value <= _T_9;
        end
      end
    end
    if (reset) begin
      value_1 <= 2'h0;
    end else if (valid_up) begin
      if (_T_10) begin
        if (_T_16) begin
          value_1 <= 2'h0;
        end else begin
          value_1 <= _T_18;
        end
      end
    end
    if (reset) begin
      value_2 <= 2'h0;
    end else if (valid_up) begin
      if (_T_2) begin
        value_2 <= 2'h0;
      end else begin
        value_2 <= _T_4;
      end
    end
  end
endmodule
module FIFO_5(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0,
  output [31:0] O_0_0
);
  reg [31:0] _T_0_0 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_0;
  wire [31:0] _T_0_0__T_15_data; // @[FIFO.scala 23:33]
  wire [1:0] _T_0_0__T_15_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_1;
  wire [31:0] _T_0_0__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T_0_0__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T_0_0__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T_0_0__T_5_en; // @[FIFO.scala 23:33]
  reg  _T_0_0__T_15_en_pipe_0;
  reg [31:0] _RAND_2;
  reg [1:0] _T_0_0__T_15_addr_pipe_0;
  reg [31:0] _RAND_3;
  reg [1:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_4;
  reg [1:0] value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  reg [1:0] value_2; // @[Counter.scala 29:33]
  reg [31:0] _RAND_6;
  wire  _T_1; // @[FIFO.scala 33:46]
  wire  _T_2; // @[Counter.scala 37:24]
  wire [1:0] _T_4; // @[Counter.scala 38:22]
  wire  _T_6; // @[FIFO.scala 38:39]
  wire [1:0] _T_9; // @[Counter.scala 38:22]
  wire  _T_10; // @[FIFO.scala 42:39]
  wire  _T_16; // @[Counter.scala 37:24]
  wire [1:0] _T_18; // @[Counter.scala 38:22]
  wire  _GEN_8; // @[FIFO.scala 42:57]
  assign _T_0_0__T_15_addr = _T_0_0__T_15_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_0_0__T_15_data = _T_0_0[_T_0_0__T_15_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T_0_0__T_15_data = _T_0_0__T_15_addr >= 2'h3 ? _RAND_1[31:0] : _T_0_0[_T_0_0__T_15_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_0_0__T_5_data = I_0_0;
  assign _T_0_0__T_5_addr = value_2;
  assign _T_0_0__T_5_mask = 1'h1;
  assign _T_0_0__T_5_en = valid_up;
  assign _T_1 = value == 2'h2; // @[FIFO.scala 33:46]
  assign _T_2 = value_2 == 2'h2; // @[Counter.scala 37:24]
  assign _T_4 = value_2 + 2'h1; // @[Counter.scala 38:22]
  assign _T_6 = value < 2'h2; // @[FIFO.scala 38:39]
  assign _T_9 = value + 2'h1; // @[Counter.scala 38:22]
  assign _T_10 = value >= 2'h1; // @[FIFO.scala 42:39]
  assign _T_16 = value_1 == 2'h2; // @[Counter.scala 37:24]
  assign _T_18 = value_1 + 2'h1; // @[Counter.scala 38:22]
  assign _GEN_8 = _T_10 & _T_10; // @[FIFO.scala 42:57]
  assign valid_down = value == 2'h2; // @[FIFO.scala 33:16]
  assign O_0_0 = _T_0_0__T_15_data; // @[FIFO.scala 43:11]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T_0_0[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_0_0__T_15_en_pipe_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_0_0__T_15_addr_pipe_0 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  value = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value_1 = _RAND_5[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  value_2 = _RAND_6[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_0_0__T_5_en & _T_0_0__T_5_mask) begin
      _T_0_0[_T_0_0__T_5_addr] <= _T_0_0__T_5_data; // @[FIFO.scala 23:33]
    end
    _T_0_0__T_15_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T_0_0__T_15_addr_pipe_0 <= value_1;
    end
    if (reset) begin
      value <= 2'h0;
    end else if (valid_up) begin
      if (_T_6) begin
        if (_T_1) begin
          value <= 2'h0;
        end else begin
          value <= _T_9;
        end
      end
    end
    if (reset) begin
      value_1 <= 2'h0;
    end else if (valid_up) begin
      if (_T_10) begin
        if (_T_16) begin
          value_1 <= 2'h0;
        end else begin
          value_1 <= _T_18;
        end
      end
    end
    if (reset) begin
      value_2 <= 2'h0;
    end else if (valid_up) begin
      if (_T_2) begin
        value_2 <= 2'h0;
      end else begin
        value_2 <= _T_4;
      end
    end
  end
endmodule
module Map2S_17(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0,
  input  [31:0] I1_0,
  output [31:0] O_0_0,
  output [31:0] O_0_1
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_1; // @[Map2S.scala 9:22]
  SSeqTupleCreator fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1(fst_op_I1),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0 = fst_op_O_0; // @[Map2S.scala 19:8]
  assign O_0_1 = fst_op_O_1; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
endmodule
module Map2S_18(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0_0,
  input  [31:0] I1_0_0,
  output [31:0] O_0_0_0,
  output [31:0] O_0_0_1
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_1; // @[Map2S.scala 9:22]
  Map2S_17 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I1_0(fst_op_I1_0),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[Map2S.scala 19:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = I1_0_0; // @[Map2S.scala 18:13]
endmodule
module Map2S_19(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0_0,
  input  [31:0] I0_0_1,
  input  [31:0] I1_0,
  output [31:0] O_0_0,
  output [31:0] O_0_1,
  output [31:0] O_0_2
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_2; // @[Map2S.scala 9:22]
  SSeqTupleAppender fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I0_1(fst_op_I0_1),
    .I1(fst_op_I1),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1),
    .O_2(fst_op_O_2)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0 = fst_op_O_0; // @[Map2S.scala 19:8]
  assign O_0_1 = fst_op_O_1; // @[Map2S.scala 19:8]
  assign O_0_2 = fst_op_O_2; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1 = I0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
endmodule
module Map2S_20(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0_0_0,
  input  [31:0] I0_0_0_1,
  input  [31:0] I1_0_0,
  output [31:0] O_0_0_0,
  output [31:0] O_0_0_1,
  output [31:0] O_0_0_2
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_2; // @[Map2S.scala 9:22]
  Map2S_19 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0_0(fst_op_I0_0_0),
    .I0_0_1(fst_op_I0_0_1),
    .I1_0(fst_op_I1_0),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1),
    .O_0_2(fst_op_O_0_2)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[Map2S.scala 19:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[Map2S.scala 19:8]
  assign O_0_0_2 = fst_op_O_0_2; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0_0 = I0_0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_1 = I0_0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = I1_0_0; // @[Map2S.scala 18:13]
endmodule
module SSeqTupleAppender_5(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0,
  input  [31:0] I0_1,
  input  [31:0] I0_2,
  input  [31:0] I1,
  output [31:0] O_0,
  output [31:0] O_1,
  output [31:0] O_2,
  output [31:0] O_3
);
  assign valid_down = valid_up; // @[Tuple.scala 28:14]
  assign O_0 = I0_0; // @[Tuple.scala 24:34]
  assign O_1 = I0_1; // @[Tuple.scala 24:34]
  assign O_2 = I0_2; // @[Tuple.scala 24:34]
  assign O_3 = I1; // @[Tuple.scala 26:32]
endmodule
module Map2S_21(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0_0,
  input  [31:0] I0_0_1,
  input  [31:0] I0_0_2,
  input  [31:0] I1_0,
  output [31:0] O_0_0,
  output [31:0] O_0_1,
  output [31:0] O_0_2,
  output [31:0] O_0_3
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_2; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_2; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_3; // @[Map2S.scala 9:22]
  SSeqTupleAppender_5 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I0_1(fst_op_I0_1),
    .I0_2(fst_op_I0_2),
    .I1(fst_op_I1),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1),
    .O_2(fst_op_O_2),
    .O_3(fst_op_O_3)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0 = fst_op_O_0; // @[Map2S.scala 19:8]
  assign O_0_1 = fst_op_O_1; // @[Map2S.scala 19:8]
  assign O_0_2 = fst_op_O_2; // @[Map2S.scala 19:8]
  assign O_0_3 = fst_op_O_3; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1 = I0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_2 = I0_0_2; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
endmodule
module Map2S_22(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0_0_0,
  input  [31:0] I0_0_0_1,
  input  [31:0] I0_0_0_2,
  input  [31:0] I1_0_0,
  output [31:0] O_0_0_0,
  output [31:0] O_0_0_1,
  output [31:0] O_0_0_2,
  output [31:0] O_0_0_3
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0_2; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_2; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_3; // @[Map2S.scala 9:22]
  Map2S_21 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0_0(fst_op_I0_0_0),
    .I0_0_1(fst_op_I0_0_1),
    .I0_0_2(fst_op_I0_0_2),
    .I1_0(fst_op_I1_0),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1),
    .O_0_2(fst_op_O_0_2),
    .O_0_3(fst_op_O_0_3)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[Map2S.scala 19:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[Map2S.scala 19:8]
  assign O_0_0_2 = fst_op_O_0_2; // @[Map2S.scala 19:8]
  assign O_0_0_3 = fst_op_O_0_3; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0_0 = I0_0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_1 = I0_0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_2 = I0_0_0_2; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = I1_0_0; // @[Map2S.scala 18:13]
endmodule
module SSeqTupleToSSeq_4(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0,
  input  [31:0] I_1,
  input  [31:0] I_2,
  input  [31:0] I_3,
  output [31:0] O_0,
  output [31:0] O_1,
  output [31:0] O_2,
  output [31:0] O_3
);
  assign valid_down = valid_up; // @[Tuple.scala 42:14]
  assign O_0 = I_0; // @[Tuple.scala 41:5]
  assign O_1 = I_1; // @[Tuple.scala 41:5]
  assign O_2 = I_2; // @[Tuple.scala 41:5]
  assign O_3 = I_3; // @[Tuple.scala 41:5]
endmodule
module Remove1S_4(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0,
  input  [31:0] I_0_1,
  input  [31:0] I_0_2,
  input  [31:0] I_0_3,
  output [31:0] O_0,
  output [31:0] O_1,
  output [31:0] O_2,
  output [31:0] O_3
);
  wire  op_inst_valid_up; // @[Remove1S.scala 9:23]
  wire  op_inst_valid_down; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_I_0; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_I_1; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_I_2; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_I_3; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_O_0; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_O_1; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_O_2; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_O_3; // @[Remove1S.scala 9:23]
  SSeqTupleToSSeq_4 op_inst ( // @[Remove1S.scala 9:23]
    .valid_up(op_inst_valid_up),
    .valid_down(op_inst_valid_down),
    .I_0(op_inst_I_0),
    .I_1(op_inst_I_1),
    .I_2(op_inst_I_2),
    .I_3(op_inst_I_3),
    .O_0(op_inst_O_0),
    .O_1(op_inst_O_1),
    .O_2(op_inst_O_2),
    .O_3(op_inst_O_3)
  );
  assign valid_down = op_inst_valid_down; // @[Remove1S.scala 16:14]
  assign O_0 = op_inst_O_0; // @[Remove1S.scala 14:5]
  assign O_1 = op_inst_O_1; // @[Remove1S.scala 14:5]
  assign O_2 = op_inst_O_2; // @[Remove1S.scala 14:5]
  assign O_3 = op_inst_O_3; // @[Remove1S.scala 14:5]
  assign op_inst_valid_up = valid_up; // @[Remove1S.scala 15:20]
  assign op_inst_I_0 = I_0_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_1 = I_0_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_2 = I_0_2; // @[Remove1S.scala 13:13]
  assign op_inst_I_3 = I_0_3; // @[Remove1S.scala 13:13]
endmodule
module MapS_27(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0_0,
  input  [31:0] I_0_0_1,
  input  [31:0] I_0_0_2,
  input  [31:0] I_0_0_3,
  output [31:0] O_0_0,
  output [31:0] O_0_1,
  output [31:0] O_0_2,
  output [31:0] O_0_3
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_0; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_1; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_2; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_3; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_0; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_1; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_2; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_3; // @[MapS.scala 9:22]
  Remove1S_4 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_0(fst_op_I_0_0),
    .I_0_1(fst_op_I_0_1),
    .I_0_2(fst_op_I_0_2),
    .I_0_3(fst_op_I_0_3),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1),
    .O_2(fst_op_O_2),
    .O_3(fst_op_O_3)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign O_0_1 = fst_op_O_1; // @[MapS.scala 17:8]
  assign O_0_2 = fst_op_O_2; // @[MapS.scala 17:8]
  assign O_0_3 = fst_op_O_3; // @[MapS.scala 17:8]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_0 = I_0_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_1 = I_0_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_2 = I_0_0_2; // @[MapS.scala 16:12]
  assign fst_op_I_0_3 = I_0_0_3; // @[MapS.scala 16:12]
endmodule
module AddNoValid(
  input  [31:0] I_t0b,
  input  [31:0] I_t1b,
  output [31:0] O
);
  assign O = I_t0b + I_t1b; // @[Arithmetic.scala 122:7]
endmodule
module ReduceS(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0,
  input  [31:0] I_1,
  input  [31:0] I_2,
  input  [31:0] I_3,
  output [31:0] O_0
);
  wire [31:0] AddNoValid_I_t0b; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_I_t1b; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_O; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_1_I_t0b; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_1_I_t1b; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_1_O; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_2_I_t0b; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_2_I_t1b; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_2_O; // @[ReduceS.scala 20:43]
  reg [31:0] _T; // @[ReduceS.scala 27:24]
  reg [31:0] _RAND_0;
  reg [31:0] _T_1; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_1;
  reg [31:0] _T_2; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_2;
  reg [31:0] _T_3; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_3;
  reg [31:0] _T_4; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_4;
  reg  _T_5; // @[ReduceS.scala 47:32]
  reg [31:0] _RAND_5;
  reg  _T_6; // @[ReduceS.scala 47:24]
  reg [31:0] _RAND_6;
  AddNoValid AddNoValid ( // @[ReduceS.scala 20:43]
    .I_t0b(AddNoValid_I_t0b),
    .I_t1b(AddNoValid_I_t1b),
    .O(AddNoValid_O)
  );
  AddNoValid AddNoValid_1 ( // @[ReduceS.scala 20:43]
    .I_t0b(AddNoValid_1_I_t0b),
    .I_t1b(AddNoValid_1_I_t1b),
    .O(AddNoValid_1_O)
  );
  AddNoValid AddNoValid_2 ( // @[ReduceS.scala 20:43]
    .I_t0b(AddNoValid_2_I_t0b),
    .I_t1b(AddNoValid_2_I_t1b),
    .O(AddNoValid_2_O)
  );
  assign valid_down = _T_6; // @[ReduceS.scala 47:14]
  assign O_0 = _T; // @[ReduceS.scala 27:14]
  assign AddNoValid_I_t0b = _T_4; // @[ReduceS.scala 43:18]
  assign AddNoValid_I_t1b = AddNoValid_1_O; // @[ReduceS.scala 36:18]
  assign AddNoValid_1_I_t0b = AddNoValid_2_O; // @[ReduceS.scala 31:18]
  assign AddNoValid_1_I_t1b = _T_2; // @[ReduceS.scala 43:18]
  assign AddNoValid_2_I_t0b = _T_3; // @[ReduceS.scala 43:18]
  assign AddNoValid_2_I_t1b = _T_1; // @[ReduceS.scala 43:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_2 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_3 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_4 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_6 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T <= AddNoValid_O;
    _T_1 <= I_0;
    _T_2 <= I_1;
    _T_3 <= I_2;
    _T_4 <= I_3;
    if (reset) begin
      _T_5 <= 1'h0;
    end else begin
      _T_5 <= valid_up;
    end
    _T_6 <= _T_5;
  end
endmodule
module MapS_28(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0,
  input  [31:0] I_0_1,
  input  [31:0] I_0_2,
  input  [31:0] I_0_3,
  output [31:0] O_0_0
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_1; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_2; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_3; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_0; // @[MapS.scala 9:22]
  ReduceS fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0(fst_op_I_0),
    .I_1(fst_op_I_1),
    .I_2(fst_op_I_2),
    .I_3(fst_op_I_3),
    .O_0(fst_op_O_0)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0 = I_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_1 = I_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_2 = I_0_2; // @[MapS.scala 16:12]
  assign fst_op_I_3 = I_0_3; // @[MapS.scala 16:12]
endmodule
module InitialDelayCounter_2(
  input   clock,
  input   reset,
  output  valid_down
);
  reg [1:0] value; // @[InitialDelayCounter.scala 8:34]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[InitialDelayCounter.scala 17:17]
  wire [1:0] _T_4; // @[InitialDelayCounter.scala 17:53]
  assign _T_1 = value < 2'h3; // @[InitialDelayCounter.scala 17:17]
  assign _T_4 = value + 2'h1; // @[InitialDelayCounter.scala 17:53]
  assign valid_down = value == 2'h3; // @[InitialDelayCounter.scala 16:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 2'h0;
    end else if (_T_1) begin
      value <= _T_4;
    end
  end
endmodule
module Module_4(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I,
  output [31:0] O_t0b,
  output [7:0]  O_t1b
);
  wire  InitialDelayCounter_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_valid_down; // @[Const.scala 11:33]
  wire  n274_valid_up; // @[Top.scala 92:22]
  wire  n274_valid_down; // @[Top.scala 92:22]
  wire [31:0] n274_I0; // @[Top.scala 92:22]
  wire [7:0] n274_I1; // @[Top.scala 92:22]
  wire [31:0] n274_O_t0b; // @[Top.scala 92:22]
  wire [7:0] n274_O_t1b; // @[Top.scala 92:22]
  InitialDelayCounter_2 InitialDelayCounter ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_clock),
    .reset(InitialDelayCounter_reset),
    .valid_down(InitialDelayCounter_valid_down)
  );
  AtomTuple_1 n274 ( // @[Top.scala 92:22]
    .valid_up(n274_valid_up),
    .valid_down(n274_valid_down),
    .I0(n274_I0),
    .I1(n274_I1),
    .O_t0b(n274_O_t0b),
    .O_t1b(n274_O_t1b)
  );
  assign valid_down = n274_valid_down; // @[Top.scala 97:16]
  assign O_t0b = n274_O_t0b; // @[Top.scala 96:7]
  assign O_t1b = n274_O_t1b; // @[Top.scala 96:7]
  assign InitialDelayCounter_clock = clock;
  assign InitialDelayCounter_reset = reset;
  assign n274_valid_up = valid_up & InitialDelayCounter_valid_down; // @[Top.scala 95:19]
  assign n274_I0 = I; // @[Top.scala 93:13]
  assign n274_I1 = 8'h2; // @[Top.scala 94:13]
endmodule
module MapS_29(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0,
  output [31:0] O_0_t0b,
  output [7:0]  O_0_t1b
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_t1b; // @[MapS.scala 9:22]
  Module_4 fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I(fst_op_I),
    .O_t0b(fst_op_O_t0b),
    .O_t1b(fst_op_O_t1b)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0_t0b = fst_op_O_t0b; // @[MapS.scala 17:8]
  assign O_0_t1b = fst_op_O_t1b; // @[MapS.scala 17:8]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I = I_0; // @[MapS.scala 16:12]
endmodule
module MapS_30(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0,
  output [31:0] O_0_0_t0b,
  output [7:0]  O_0_0_t1b
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_0_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0_t1b; // @[MapS.scala 9:22]
  MapS_29 fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0(fst_op_I_0),
    .O_0_t0b(fst_op_O_0_t0b),
    .O_0_t1b(fst_op_O_0_t1b)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0_0_t0b = fst_op_O_0_t0b; // @[MapS.scala 17:8]
  assign O_0_0_t1b = fst_op_O_0_t1b; // @[MapS.scala 17:8]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0 = I_0_0; // @[MapS.scala 16:12]
endmodule
module ReduceS_1(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0,
  input  [31:0] I_1,
  input  [31:0] I_2,
  input  [31:0] I_3,
  output [31:0] O_0
);
  wire [31:0] AddNoValid_I_t0b; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_I_t1b; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_O; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_1_I_t0b; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_1_I_t1b; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_1_O; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_2_I_t0b; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_2_I_t1b; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_2_O; // @[ReduceS.scala 20:43]
  reg [31:0] _T; // @[ReduceS.scala 27:24]
  reg [31:0] _RAND_0;
  reg [31:0] _T_1; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_1;
  reg [31:0] _T_2; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_2;
  reg [31:0] _T_3; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_3;
  reg [31:0] _T_4; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_4;
  reg  _T_5; // @[ReduceS.scala 47:32]
  reg [31:0] _RAND_5;
  reg  _T_6; // @[ReduceS.scala 47:24]
  reg [31:0] _RAND_6;
  AddNoValid AddNoValid ( // @[ReduceS.scala 20:43]
    .I_t0b(AddNoValid_I_t0b),
    .I_t1b(AddNoValid_I_t1b),
    .O(AddNoValid_O)
  );
  AddNoValid AddNoValid_1 ( // @[ReduceS.scala 20:43]
    .I_t0b(AddNoValid_1_I_t0b),
    .I_t1b(AddNoValid_1_I_t1b),
    .O(AddNoValid_1_O)
  );
  AddNoValid AddNoValid_2 ( // @[ReduceS.scala 20:43]
    .I_t0b(AddNoValid_2_I_t0b),
    .I_t1b(AddNoValid_2_I_t1b),
    .O(AddNoValid_2_O)
  );
  assign valid_down = _T_6; // @[ReduceS.scala 47:14]
  assign O_0 = _T; // @[ReduceS.scala 27:14]
  assign AddNoValid_I_t0b = _T_3; // @[ReduceS.scala 43:18]
  assign AddNoValid_I_t1b = AddNoValid_1_O; // @[ReduceS.scala 36:18]
  assign AddNoValid_1_I_t0b = AddNoValid_2_O; // @[ReduceS.scala 31:18]
  assign AddNoValid_1_I_t1b = _T_2; // @[ReduceS.scala 43:18]
  assign AddNoValid_2_I_t0b = _T_1; // @[ReduceS.scala 43:18]
  assign AddNoValid_2_I_t1b = _T_4; // @[ReduceS.scala 43:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_2 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_3 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_4 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_6 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T <= AddNoValid_O;
    _T_1 <= I_0;
    _T_2 <= I_1;
    _T_3 <= I_2;
    _T_4 <= I_3;
    if (reset) begin
      _T_5 <= 1'h0;
    end else begin
      _T_5 <= valid_up;
    end
    _T_6 <= _T_5;
  end
endmodule
module MapS_38(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0,
  input  [31:0] I_0_1,
  input  [31:0] I_0_2,
  input  [31:0] I_0_3,
  output [31:0] O_0_0
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_1; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_2; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_3; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_0; // @[MapS.scala 9:22]
  ReduceS_1 fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0(fst_op_I_0),
    .I_1(fst_op_I_1),
    .I_2(fst_op_I_2),
    .I_3(fst_op_I_3),
    .O_0(fst_op_O_0)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0 = I_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_1 = I_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_2 = I_0_2; // @[MapS.scala 16:12]
  assign fst_op_I_3 = I_0_3; // @[MapS.scala 16:12]
endmodule
module AtomTuple_15(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_t0b,
  input  [31:0] I0_t1b_t0b,
  input  [31:0] I0_t1b_t1b,
  input  [31:0] I1_t0b,
  input  [31:0] I1_t1b_t0b,
  input  [31:0] I1_t1b_t1b,
  output [31:0] O_t0b_t0b,
  output [31:0] O_t0b_t1b_t0b,
  output [31:0] O_t0b_t1b_t1b,
  output [31:0] O_t1b_t0b,
  output [31:0] O_t1b_t1b_t0b,
  output [31:0] O_t1b_t1b_t1b
);
  assign valid_down = valid_up; // @[Tuple.scala 51:14]
  assign O_t0b_t0b = I0_t0b; // @[Tuple.scala 49:9]
  assign O_t0b_t1b_t0b = I0_t1b_t0b; // @[Tuple.scala 49:9]
  assign O_t0b_t1b_t1b = I0_t1b_t1b; // @[Tuple.scala 49:9]
  assign O_t1b_t0b = I1_t0b; // @[Tuple.scala 50:9]
  assign O_t1b_t1b_t0b = I1_t1b_t0b; // @[Tuple.scala 50:9]
  assign O_t1b_t1b_t1b = I1_t1b_t1b; // @[Tuple.scala 50:9]
endmodule
module Map2S_33(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0_t0b,
  input  [31:0] I0_0_t1b_t0b,
  input  [31:0] I0_0_t1b_t1b,
  input  [31:0] I1_0_t0b,
  input  [31:0] I1_0_t1b_t0b,
  input  [31:0] I1_0_t1b_t1b,
  output [31:0] O_0_t0b_t0b,
  output [31:0] O_0_t0b_t1b_t0b,
  output [31:0] O_0_t0b_t1b_t1b,
  output [31:0] O_0_t1b_t0b,
  output [31:0] O_0_t1b_t1b_t0b,
  output [31:0] O_0_t1b_t1b_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_t1b_t1b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_t1b_t1b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_t0b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_t0b_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_t0b_t1b_t1b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_t1b_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_t1b_t1b_t1b; // @[Map2S.scala 9:22]
  AtomTuple_15 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_t0b(fst_op_I0_t0b),
    .I0_t1b_t0b(fst_op_I0_t1b_t0b),
    .I0_t1b_t1b(fst_op_I0_t1b_t1b),
    .I1_t0b(fst_op_I1_t0b),
    .I1_t1b_t0b(fst_op_I1_t1b_t0b),
    .I1_t1b_t1b(fst_op_I1_t1b_t1b),
    .O_t0b_t0b(fst_op_O_t0b_t0b),
    .O_t0b_t1b_t0b(fst_op_O_t0b_t1b_t0b),
    .O_t0b_t1b_t1b(fst_op_O_t0b_t1b_t1b),
    .O_t1b_t0b(fst_op_O_t1b_t0b),
    .O_t1b_t1b_t0b(fst_op_O_t1b_t1b_t0b),
    .O_t1b_t1b_t1b(fst_op_O_t1b_t1b_t1b)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_t0b_t0b = fst_op_O_t0b_t0b; // @[Map2S.scala 19:8]
  assign O_0_t0b_t1b_t0b = fst_op_O_t0b_t1b_t0b; // @[Map2S.scala 19:8]
  assign O_0_t0b_t1b_t1b = fst_op_O_t0b_t1b_t1b; // @[Map2S.scala 19:8]
  assign O_0_t1b_t0b = fst_op_O_t1b_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b_t1b_t0b = fst_op_O_t1b_t1b_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b_t1b_t1b = fst_op_O_t1b_t1b_t1b; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_t0b = I0_0_t0b; // @[Map2S.scala 17:13]
  assign fst_op_I0_t1b_t0b = I0_0_t1b_t0b; // @[Map2S.scala 17:13]
  assign fst_op_I0_t1b_t1b = I0_0_t1b_t1b; // @[Map2S.scala 17:13]
  assign fst_op_I1_t0b = I1_0_t0b; // @[Map2S.scala 18:13]
  assign fst_op_I1_t1b_t0b = I1_0_t1b_t0b; // @[Map2S.scala 18:13]
  assign fst_op_I1_t1b_t1b = I1_0_t1b_t1b; // @[Map2S.scala 18:13]
endmodule
module Map2S_34(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0_0_t0b,
  input  [31:0] I0_0_0_t1b_t0b,
  input  [31:0] I0_0_0_t1b_t1b,
  input  [31:0] I1_0_0_t0b,
  input  [31:0] I1_0_0_t1b_t0b,
  input  [31:0] I1_0_0_t1b_t1b,
  output [31:0] O_0_0_t0b_t0b,
  output [31:0] O_0_0_t0b_t1b_t0b,
  output [31:0] O_0_0_t0b_t1b_t1b,
  output [31:0] O_0_0_t1b_t0b,
  output [31:0] O_0_0_t1b_t1b_t0b,
  output [31:0] O_0_0_t1b_t1b_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0_t1b_t1b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_0_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_0_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_0_t1b_t1b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_t0b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_t0b_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_t0b_t1b_t1b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_t1b_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_t1b_t1b_t1b; // @[Map2S.scala 9:22]
  Map2S_33 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0_t0b(fst_op_I0_0_t0b),
    .I0_0_t1b_t0b(fst_op_I0_0_t1b_t0b),
    .I0_0_t1b_t1b(fst_op_I0_0_t1b_t1b),
    .I1_0_t0b(fst_op_I1_0_t0b),
    .I1_0_t1b_t0b(fst_op_I1_0_t1b_t0b),
    .I1_0_t1b_t1b(fst_op_I1_0_t1b_t1b),
    .O_0_t0b_t0b(fst_op_O_0_t0b_t0b),
    .O_0_t0b_t1b_t0b(fst_op_O_0_t0b_t1b_t0b),
    .O_0_t0b_t1b_t1b(fst_op_O_0_t0b_t1b_t1b),
    .O_0_t1b_t0b(fst_op_O_0_t1b_t0b),
    .O_0_t1b_t1b_t0b(fst_op_O_0_t1b_t1b_t0b),
    .O_0_t1b_t1b_t1b(fst_op_O_0_t1b_t1b_t1b)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_t0b_t0b = fst_op_O_0_t0b_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_t0b_t1b_t0b = fst_op_O_0_t0b_t1b_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_t0b_t1b_t1b = fst_op_O_0_t0b_t1b_t1b; // @[Map2S.scala 19:8]
  assign O_0_0_t1b_t0b = fst_op_O_0_t1b_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_t1b_t1b_t0b = fst_op_O_0_t1b_t1b_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_t1b_t1b_t1b = fst_op_O_0_t1b_t1b_t1b; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0_t0b = I0_0_0_t0b; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_t1b_t0b = I0_0_0_t1b_t0b; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_t1b_t1b = I0_0_0_t1b_t1b; // @[Map2S.scala 17:13]
  assign fst_op_I1_0_t0b = I1_0_0_t0b; // @[Map2S.scala 18:13]
  assign fst_op_I1_0_t1b_t0b = I1_0_0_t1b_t0b; // @[Map2S.scala 18:13]
  assign fst_op_I1_0_t1b_t1b = I1_0_0_t1b_t1b; // @[Map2S.scala 18:13]
endmodule
module AtomTuple_16(
  input         valid_up,
  output        valid_down,
  input         I0,
  input  [31:0] I1_t0b_t0b,
  input  [31:0] I1_t0b_t1b_t0b,
  input  [31:0] I1_t0b_t1b_t1b,
  input  [31:0] I1_t1b_t0b,
  input  [31:0] I1_t1b_t1b_t0b,
  input  [31:0] I1_t1b_t1b_t1b,
  output        O_t0b,
  output [31:0] O_t1b_t0b_t0b,
  output [31:0] O_t1b_t0b_t1b_t0b,
  output [31:0] O_t1b_t0b_t1b_t1b,
  output [31:0] O_t1b_t1b_t0b,
  output [31:0] O_t1b_t1b_t1b_t0b,
  output [31:0] O_t1b_t1b_t1b_t1b
);
  assign valid_down = valid_up; // @[Tuple.scala 51:14]
  assign O_t0b = I0; // @[Tuple.scala 49:9]
  assign O_t1b_t0b_t0b = I1_t0b_t0b; // @[Tuple.scala 50:9]
  assign O_t1b_t0b_t1b_t0b = I1_t0b_t1b_t0b; // @[Tuple.scala 50:9]
  assign O_t1b_t0b_t1b_t1b = I1_t0b_t1b_t1b; // @[Tuple.scala 50:9]
  assign O_t1b_t1b_t0b = I1_t1b_t0b; // @[Tuple.scala 50:9]
  assign O_t1b_t1b_t1b_t0b = I1_t1b_t1b_t0b; // @[Tuple.scala 50:9]
  assign O_t1b_t1b_t1b_t1b = I1_t1b_t1b_t1b; // @[Tuple.scala 50:9]
endmodule
module Map2S_35(
  input         valid_up,
  output        valid_down,
  input         I0_0,
  input  [31:0] I1_0_t0b_t0b,
  input  [31:0] I1_0_t0b_t1b_t0b,
  input  [31:0] I1_0_t0b_t1b_t1b,
  input  [31:0] I1_0_t1b_t0b,
  input  [31:0] I1_0_t1b_t1b_t0b,
  input  [31:0] I1_0_t1b_t1b_t1b,
  output        O_0_t0b,
  output [31:0] O_0_t1b_t0b_t0b,
  output [31:0] O_0_t1b_t0b_t1b_t0b,
  output [31:0] O_0_t1b_t0b_t1b_t1b,
  output [31:0] O_0_t1b_t1b_t0b,
  output [31:0] O_0_t1b_t1b_t1b_t0b,
  output [31:0] O_0_t1b_t1b_t1b_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire  fst_op_I0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_t0b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_t0b_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_t0b_t1b_t1b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_t1b_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_t1b_t1b_t1b; // @[Map2S.scala 9:22]
  wire  fst_op_O_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_t1b_t0b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_t1b_t0b_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_t1b_t0b_t1b_t1b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_t1b_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_t1b_t1b_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_t1b_t1b_t1b_t1b; // @[Map2S.scala 9:22]
  AtomTuple_16 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1_t0b_t0b(fst_op_I1_t0b_t0b),
    .I1_t0b_t1b_t0b(fst_op_I1_t0b_t1b_t0b),
    .I1_t0b_t1b_t1b(fst_op_I1_t0b_t1b_t1b),
    .I1_t1b_t0b(fst_op_I1_t1b_t0b),
    .I1_t1b_t1b_t0b(fst_op_I1_t1b_t1b_t0b),
    .I1_t1b_t1b_t1b(fst_op_I1_t1b_t1b_t1b),
    .O_t0b(fst_op_O_t0b),
    .O_t1b_t0b_t0b(fst_op_O_t1b_t0b_t0b),
    .O_t1b_t0b_t1b_t0b(fst_op_O_t1b_t0b_t1b_t0b),
    .O_t1b_t0b_t1b_t1b(fst_op_O_t1b_t0b_t1b_t1b),
    .O_t1b_t1b_t0b(fst_op_O_t1b_t1b_t0b),
    .O_t1b_t1b_t1b_t0b(fst_op_O_t1b_t1b_t1b_t0b),
    .O_t1b_t1b_t1b_t1b(fst_op_O_t1b_t1b_t1b_t1b)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_t0b = fst_op_O_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b_t0b_t0b = fst_op_O_t1b_t0b_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b_t0b_t1b_t0b = fst_op_O_t1b_t0b_t1b_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b_t0b_t1b_t1b = fst_op_O_t1b_t0b_t1b_t1b; // @[Map2S.scala 19:8]
  assign O_0_t1b_t1b_t0b = fst_op_O_t1b_t1b_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b_t1b_t1b_t0b = fst_op_O_t1b_t1b_t1b_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b_t1b_t1b_t1b = fst_op_O_t1b_t1b_t1b_t1b; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1_t0b_t0b = I1_0_t0b_t0b; // @[Map2S.scala 18:13]
  assign fst_op_I1_t0b_t1b_t0b = I1_0_t0b_t1b_t0b; // @[Map2S.scala 18:13]
  assign fst_op_I1_t0b_t1b_t1b = I1_0_t0b_t1b_t1b; // @[Map2S.scala 18:13]
  assign fst_op_I1_t1b_t0b = I1_0_t1b_t0b; // @[Map2S.scala 18:13]
  assign fst_op_I1_t1b_t1b_t0b = I1_0_t1b_t1b_t0b; // @[Map2S.scala 18:13]
  assign fst_op_I1_t1b_t1b_t1b = I1_0_t1b_t1b_t1b; // @[Map2S.scala 18:13]
endmodule
module Map2S_36(
  input         valid_up,
  output        valid_down,
  input         I0_0_0,
  input  [31:0] I1_0_0_t0b_t0b,
  input  [31:0] I1_0_0_t0b_t1b_t0b,
  input  [31:0] I1_0_0_t0b_t1b_t1b,
  input  [31:0] I1_0_0_t1b_t0b,
  input  [31:0] I1_0_0_t1b_t1b_t0b,
  input  [31:0] I1_0_0_t1b_t1b_t1b,
  output        O_0_0_t0b,
  output [31:0] O_0_0_t1b_t0b_t0b,
  output [31:0] O_0_0_t1b_t0b_t1b_t0b,
  output [31:0] O_0_0_t1b_t0b_t1b_t1b,
  output [31:0] O_0_0_t1b_t1b_t0b,
  output [31:0] O_0_0_t1b_t1b_t1b_t0b,
  output [31:0] O_0_0_t1b_t1b_t1b_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire  fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_0_t0b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_0_t0b_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_0_t0b_t1b_t1b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_0_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_0_t1b_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_0_t1b_t1b_t1b; // @[Map2S.scala 9:22]
  wire  fst_op_O_0_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_t1b_t0b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_t1b_t0b_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_t1b_t0b_t1b_t1b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_t1b_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_t1b_t1b_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_t1b_t1b_t1b_t1b; // @[Map2S.scala 9:22]
  Map2S_35 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I1_0_t0b_t0b(fst_op_I1_0_t0b_t0b),
    .I1_0_t0b_t1b_t0b(fst_op_I1_0_t0b_t1b_t0b),
    .I1_0_t0b_t1b_t1b(fst_op_I1_0_t0b_t1b_t1b),
    .I1_0_t1b_t0b(fst_op_I1_0_t1b_t0b),
    .I1_0_t1b_t1b_t0b(fst_op_I1_0_t1b_t1b_t0b),
    .I1_0_t1b_t1b_t1b(fst_op_I1_0_t1b_t1b_t1b),
    .O_0_t0b(fst_op_O_0_t0b),
    .O_0_t1b_t0b_t0b(fst_op_O_0_t1b_t0b_t0b),
    .O_0_t1b_t0b_t1b_t0b(fst_op_O_0_t1b_t0b_t1b_t0b),
    .O_0_t1b_t0b_t1b_t1b(fst_op_O_0_t1b_t0b_t1b_t1b),
    .O_0_t1b_t1b_t0b(fst_op_O_0_t1b_t1b_t0b),
    .O_0_t1b_t1b_t1b_t0b(fst_op_O_0_t1b_t1b_t1b_t0b),
    .O_0_t1b_t1b_t1b_t1b(fst_op_O_0_t1b_t1b_t1b_t1b)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_t0b = fst_op_O_0_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_t1b_t0b_t0b = fst_op_O_0_t1b_t0b_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_t1b_t0b_t1b_t0b = fst_op_O_0_t1b_t0b_t1b_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_t1b_t0b_t1b_t1b = fst_op_O_0_t1b_t0b_t1b_t1b; // @[Map2S.scala 19:8]
  assign O_0_0_t1b_t1b_t0b = fst_op_O_0_t1b_t1b_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_t1b_t1b_t1b_t0b = fst_op_O_0_t1b_t1b_t1b_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_t1b_t1b_t1b_t1b = fst_op_O_0_t1b_t1b_t1b_t1b; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1_0_t0b_t0b = I1_0_0_t0b_t0b; // @[Map2S.scala 18:13]
  assign fst_op_I1_0_t0b_t1b_t0b = I1_0_0_t0b_t1b_t0b; // @[Map2S.scala 18:13]
  assign fst_op_I1_0_t0b_t1b_t1b = I1_0_0_t0b_t1b_t1b; // @[Map2S.scala 18:13]
  assign fst_op_I1_0_t1b_t0b = I1_0_0_t1b_t0b; // @[Map2S.scala 18:13]
  assign fst_op_I1_0_t1b_t1b_t0b = I1_0_0_t1b_t1b_t0b; // @[Map2S.scala 18:13]
  assign fst_op_I1_0_t1b_t1b_t1b = I1_0_0_t1b_t1b_t1b; // @[Map2S.scala 18:13]
endmodule
module If(
  input         valid_up,
  output        valid_down,
  input         I_t0b,
  input  [31:0] I_t1b_t0b_t0b,
  input  [31:0] I_t1b_t0b_t1b_t0b,
  input  [31:0] I_t1b_t0b_t1b_t1b,
  input  [31:0] I_t1b_t1b_t0b,
  input  [31:0] I_t1b_t1b_t1b_t0b,
  input  [31:0] I_t1b_t1b_t1b_t1b,
  output [31:0] O_t0b,
  output [31:0] O_t1b_t0b,
  output [31:0] O_t1b_t1b
);
  assign valid_down = valid_up; // @[Arithmetic.scala 525:14]
  assign O_t0b = I_t0b ? I_t1b_t0b_t0b : I_t1b_t1b_t0b; // @[Arithmetic.scala 523:9 Arithmetic.scala 524:20]
  assign O_t1b_t0b = I_t0b ? I_t1b_t0b_t1b_t0b : I_t1b_t1b_t1b_t0b; // @[Arithmetic.scala 523:9 Arithmetic.scala 524:20]
  assign O_t1b_t1b = I_t0b ? I_t1b_t0b_t1b_t1b : I_t1b_t1b_t1b_t1b; // @[Arithmetic.scala 523:9 Arithmetic.scala 524:20]
endmodule
module MapS_43(
  input         valid_up,
  output        valid_down,
  input         I_0_t0b,
  input  [31:0] I_0_t1b_t0b_t0b,
  input  [31:0] I_0_t1b_t0b_t1b_t0b,
  input  [31:0] I_0_t1b_t0b_t1b_t1b,
  input  [31:0] I_0_t1b_t1b_t0b,
  input  [31:0] I_0_t1b_t1b_t1b_t0b,
  input  [31:0] I_0_t1b_t1b_t1b_t1b,
  output [31:0] O_0_t0b,
  output [31:0] O_0_t1b_t0b,
  output [31:0] O_0_t1b_t1b
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire  fst_op_I_t0b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_t1b_t0b_t0b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_t1b_t0b_t1b_t0b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_t1b_t0b_t1b_t1b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_t1b_t1b_t0b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_t1b_t1b_t1b_t0b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_t1b_t1b_t1b_t1b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_t0b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_t1b_t0b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_t1b_t1b; // @[MapS.scala 9:22]
  If fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_t0b(fst_op_I_t0b),
    .I_t1b_t0b_t0b(fst_op_I_t1b_t0b_t0b),
    .I_t1b_t0b_t1b_t0b(fst_op_I_t1b_t0b_t1b_t0b),
    .I_t1b_t0b_t1b_t1b(fst_op_I_t1b_t0b_t1b_t1b),
    .I_t1b_t1b_t0b(fst_op_I_t1b_t1b_t0b),
    .I_t1b_t1b_t1b_t0b(fst_op_I_t1b_t1b_t1b_t0b),
    .I_t1b_t1b_t1b_t1b(fst_op_I_t1b_t1b_t1b_t1b),
    .O_t0b(fst_op_O_t0b),
    .O_t1b_t0b(fst_op_O_t1b_t0b),
    .O_t1b_t1b(fst_op_O_t1b_t1b)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0_t0b = fst_op_O_t0b; // @[MapS.scala 17:8]
  assign O_0_t1b_t0b = fst_op_O_t1b_t0b; // @[MapS.scala 17:8]
  assign O_0_t1b_t1b = fst_op_O_t1b_t1b; // @[MapS.scala 17:8]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_t0b = I_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_t1b_t0b_t0b = I_0_t1b_t0b_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_t1b_t0b_t1b_t0b = I_0_t1b_t0b_t1b_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_t1b_t0b_t1b_t1b = I_0_t1b_t0b_t1b_t1b; // @[MapS.scala 16:12]
  assign fst_op_I_t1b_t1b_t0b = I_0_t1b_t1b_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_t1b_t1b_t1b_t0b = I_0_t1b_t1b_t1b_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_t1b_t1b_t1b_t1b = I_0_t1b_t1b_t1b_t1b; // @[MapS.scala 16:12]
endmodule
module MapS_44(
  input         valid_up,
  output        valid_down,
  input         I_0_0_t0b,
  input  [31:0] I_0_0_t1b_t0b_t0b,
  input  [31:0] I_0_0_t1b_t0b_t1b_t0b,
  input  [31:0] I_0_0_t1b_t0b_t1b_t1b,
  input  [31:0] I_0_0_t1b_t1b_t0b,
  input  [31:0] I_0_0_t1b_t1b_t1b_t0b,
  input  [31:0] I_0_0_t1b_t1b_t1b_t1b,
  output [31:0] O_0_0_t0b,
  output [31:0] O_0_0_t1b_t0b,
  output [31:0] O_0_0_t1b_t1b
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire  fst_op_I_0_t0b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_t1b_t0b_t0b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_t1b_t0b_t1b_t0b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_t1b_t0b_t1b_t1b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_t1b_t1b_t0b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_t1b_t1b_t1b_t0b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_t1b_t1b_t1b_t1b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_0_t0b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_0_t1b_t0b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_0_t1b_t1b; // @[MapS.scala 9:22]
  MapS_43 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_t0b(fst_op_I_0_t0b),
    .I_0_t1b_t0b_t0b(fst_op_I_0_t1b_t0b_t0b),
    .I_0_t1b_t0b_t1b_t0b(fst_op_I_0_t1b_t0b_t1b_t0b),
    .I_0_t1b_t0b_t1b_t1b(fst_op_I_0_t1b_t0b_t1b_t1b),
    .I_0_t1b_t1b_t0b(fst_op_I_0_t1b_t1b_t0b),
    .I_0_t1b_t1b_t1b_t0b(fst_op_I_0_t1b_t1b_t1b_t0b),
    .I_0_t1b_t1b_t1b_t1b(fst_op_I_0_t1b_t1b_t1b_t1b),
    .O_0_t0b(fst_op_O_0_t0b),
    .O_0_t1b_t0b(fst_op_O_0_t1b_t0b),
    .O_0_t1b_t1b(fst_op_O_0_t1b_t1b)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0_0_t0b = fst_op_O_0_t0b; // @[MapS.scala 17:8]
  assign O_0_0_t1b_t0b = fst_op_O_0_t1b_t0b; // @[MapS.scala 17:8]
  assign O_0_0_t1b_t1b = fst_op_O_0_t1b_t1b; // @[MapS.scala 17:8]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_t0b = I_0_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_0_t1b_t0b_t0b = I_0_0_t1b_t0b_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_0_t1b_t0b_t1b_t0b = I_0_0_t1b_t0b_t1b_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_0_t1b_t0b_t1b_t1b = I_0_0_t1b_t0b_t1b_t1b; // @[MapS.scala 16:12]
  assign fst_op_I_0_t1b_t1b_t0b = I_0_0_t1b_t1b_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_0_t1b_t1b_t1b_t0b = I_0_0_t1b_t1b_t1b_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_0_t1b_t1b_t1b_t1b = I_0_0_t1b_t1b_t1b_t1b; // @[MapS.scala 16:12]
endmodule
module Module_6(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0_0,
  input  [31:0] I0_0_1,
  input  [31:0] I0_0_2,
  input  [31:0] I0_1_0,
  input  [31:0] I0_1_1,
  input  [31:0] I0_1_2,
  input  [31:0] I0_2_0,
  input  [31:0] I0_2_1,
  input  [31:0] I0_2_2,
  input         I1_0_0_t0b,
  input         I1_0_0_t1b,
  output [31:0] O_0_0_t0b,
  output [31:0] O_0_0_t1b_t0b,
  output [31:0] O_0_0_t1b_t1b
);
  wire  n152_valid_up; // @[Top.scala 116:22]
  wire  n152_valid_down; // @[Top.scala 116:22]
  wire  n152_I_0_0_t0b; // @[Top.scala 116:22]
  wire  n152_O_0_0; // @[Top.scala 116:22]
  wire  n430_clock; // @[Top.scala 119:22]
  wire  n430_reset; // @[Top.scala 119:22]
  wire  n430_valid_up; // @[Top.scala 119:22]
  wire  n430_valid_down; // @[Top.scala 119:22]
  wire  n430_I_0_0; // @[Top.scala 119:22]
  wire  n430_O_0_0; // @[Top.scala 119:22]
  wire  n157_valid_up; // @[Top.scala 122:22]
  wire  n157_valid_down; // @[Top.scala 122:22]
  wire  n157_I_0_0_t1b; // @[Top.scala 122:22]
  wire  n157_O_0_0; // @[Top.scala 122:22]
  wire  n360_clock; // @[Top.scala 125:22]
  wire  n360_reset; // @[Top.scala 125:22]
  wire  n360_valid_up; // @[Top.scala 125:22]
  wire  n360_valid_down; // @[Top.scala 125:22]
  wire  n360_I_0_0; // @[Top.scala 125:22]
  wire  n360_O_0_0; // @[Top.scala 125:22]
  wire  n159_valid_up; // @[Top.scala 128:22]
  wire  n159_valid_down; // @[Top.scala 128:22]
  wire [31:0] n159_I_1_0; // @[Top.scala 128:22]
  wire [31:0] n159_I_1_1; // @[Top.scala 128:22]
  wire [31:0] n159_I_1_2; // @[Top.scala 128:22]
  wire [31:0] n159_O_0_0; // @[Top.scala 128:22]
  wire [31:0] n159_O_0_1; // @[Top.scala 128:22]
  wire [31:0] n159_O_0_2; // @[Top.scala 128:22]
  wire  n162_valid_up; // @[Top.scala 131:22]
  wire  n162_valid_down; // @[Top.scala 131:22]
  wire [31:0] n162_I_0_0; // @[Top.scala 131:22]
  wire [31:0] n162_O_0_0; // @[Top.scala 131:22]
  wire  n165_valid_up; // @[Top.scala 134:22]
  wire  n165_valid_down; // @[Top.scala 134:22]
  wire [31:0] n165_I_0_2; // @[Top.scala 134:22]
  wire [31:0] n165_O_0_0; // @[Top.scala 134:22]
  wire  n166_valid_up; // @[Top.scala 137:22]
  wire  n166_valid_down; // @[Top.scala 137:22]
  wire [31:0] n166_I0_0_0; // @[Top.scala 137:22]
  wire [31:0] n166_I1_0_0; // @[Top.scala 137:22]
  wire [31:0] n166_O_0_0_t0b; // @[Top.scala 137:22]
  wire [31:0] n166_O_0_0_t1b; // @[Top.scala 137:22]
  wire  n177_valid_up; // @[Top.scala 141:22]
  wire  n177_valid_down; // @[Top.scala 141:22]
  wire [31:0] n177_I_0_0_t0b; // @[Top.scala 141:22]
  wire [31:0] n177_I_0_0_t1b; // @[Top.scala 141:22]
  wire [31:0] n177_O_0_0; // @[Top.scala 141:22]
  wire  n184_clock; // @[Top.scala 144:22]
  wire  n184_reset; // @[Top.scala 144:22]
  wire  n184_valid_up; // @[Top.scala 144:22]
  wire  n184_valid_down; // @[Top.scala 144:22]
  wire [31:0] n184_I_0_0; // @[Top.scala 144:22]
  wire [31:0] n184_O_0_0_t0b; // @[Top.scala 144:22]
  wire [7:0] n184_O_0_0_t1b; // @[Top.scala 144:22]
  wire  n189_valid_up; // @[Top.scala 147:22]
  wire  n189_valid_down; // @[Top.scala 147:22]
  wire [31:0] n189_I_0_0_t0b; // @[Top.scala 147:22]
  wire [7:0] n189_I_0_0_t1b; // @[Top.scala 147:22]
  wire [31:0] n189_O_0_0; // @[Top.scala 147:22]
  wire  n192_valid_up; // @[Top.scala 150:22]
  wire  n192_valid_down; // @[Top.scala 150:22]
  wire [31:0] n192_I_0_1; // @[Top.scala 150:22]
  wire [31:0] n192_O_0_0; // @[Top.scala 150:22]
  wire  n193_valid_up; // @[Top.scala 153:22]
  wire  n193_valid_down; // @[Top.scala 153:22]
  wire [31:0] n193_I_0_0; // @[Top.scala 153:22]
  wire [31:0] n193_I_0_1; // @[Top.scala 153:22]
  wire [31:0] n193_I_0_2; // @[Top.scala 153:22]
  wire [31:0] n193_O_0_0; // @[Top.scala 153:22]
  wire [31:0] n193_O_0_1; // @[Top.scala 153:22]
  wire [31:0] n193_O_0_2; // @[Top.scala 153:22]
  wire  n196_valid_up; // @[Top.scala 156:22]
  wire  n196_valid_down; // @[Top.scala 156:22]
  wire [31:0] n196_I_0_1; // @[Top.scala 156:22]
  wire [31:0] n196_O_0_0; // @[Top.scala 156:22]
  wire  n197_valid_up; // @[Top.scala 159:22]
  wire  n197_valid_down; // @[Top.scala 159:22]
  wire [31:0] n197_I_2_0; // @[Top.scala 159:22]
  wire [31:0] n197_I_2_1; // @[Top.scala 159:22]
  wire [31:0] n197_I_2_2; // @[Top.scala 159:22]
  wire [31:0] n197_O_0_0; // @[Top.scala 159:22]
  wire [31:0] n197_O_0_1; // @[Top.scala 159:22]
  wire [31:0] n197_O_0_2; // @[Top.scala 159:22]
  wire  n200_valid_up; // @[Top.scala 162:22]
  wire  n200_valid_down; // @[Top.scala 162:22]
  wire [31:0] n200_I_0_1; // @[Top.scala 162:22]
  wire [31:0] n200_O_0_0; // @[Top.scala 162:22]
  wire  n201_valid_up; // @[Top.scala 165:22]
  wire  n201_valid_down; // @[Top.scala 165:22]
  wire [31:0] n201_I0_0_0; // @[Top.scala 165:22]
  wire [31:0] n201_I1_0_0; // @[Top.scala 165:22]
  wire [31:0] n201_O_0_0_t0b; // @[Top.scala 165:22]
  wire [31:0] n201_O_0_0_t1b; // @[Top.scala 165:22]
  wire  n212_valid_up; // @[Top.scala 169:22]
  wire  n212_valid_down; // @[Top.scala 169:22]
  wire [31:0] n212_I_0_0_t0b; // @[Top.scala 169:22]
  wire [31:0] n212_I_0_0_t1b; // @[Top.scala 169:22]
  wire [31:0] n212_O_0_0; // @[Top.scala 169:22]
  wire  n219_clock; // @[Top.scala 172:22]
  wire  n219_reset; // @[Top.scala 172:22]
  wire  n219_valid_up; // @[Top.scala 172:22]
  wire  n219_valid_down; // @[Top.scala 172:22]
  wire [31:0] n219_I_0_0; // @[Top.scala 172:22]
  wire [31:0] n219_O_0_0_t0b; // @[Top.scala 172:22]
  wire [7:0] n219_O_0_0_t1b; // @[Top.scala 172:22]
  wire  n224_valid_up; // @[Top.scala 175:22]
  wire  n224_valid_down; // @[Top.scala 175:22]
  wire [31:0] n224_I_0_0_t0b; // @[Top.scala 175:22]
  wire [7:0] n224_I_0_0_t1b; // @[Top.scala 175:22]
  wire [31:0] n224_O_0_0; // @[Top.scala 175:22]
  wire  n225_valid_up; // @[Top.scala 178:22]
  wire  n225_valid_down; // @[Top.scala 178:22]
  wire [31:0] n225_I0_0_0; // @[Top.scala 178:22]
  wire [31:0] n225_I1_0_0; // @[Top.scala 178:22]
  wire [31:0] n225_O_0_0_t0b; // @[Top.scala 178:22]
  wire [31:0] n225_O_0_0_t1b; // @[Top.scala 178:22]
  wire  n232_valid_up; // @[Top.scala 182:22]
  wire  n232_valid_down; // @[Top.scala 182:22]
  wire [31:0] n232_I0_0_0; // @[Top.scala 182:22]
  wire [31:0] n232_I1_0_0_t0b; // @[Top.scala 182:22]
  wire [31:0] n232_I1_0_0_t1b; // @[Top.scala 182:22]
  wire [31:0] n232_O_0_0_t0b; // @[Top.scala 182:22]
  wire [31:0] n232_O_0_0_t1b_t0b; // @[Top.scala 182:22]
  wire [31:0] n232_O_0_0_t1b_t1b; // @[Top.scala 182:22]
  wire  n352_clock; // @[Top.scala 186:22]
  wire  n352_reset; // @[Top.scala 186:22]
  wire  n352_valid_up; // @[Top.scala 186:22]
  wire  n352_valid_down; // @[Top.scala 186:22]
  wire [31:0] n352_I_0_0_t0b; // @[Top.scala 186:22]
  wire [31:0] n352_I_0_0_t1b_t0b; // @[Top.scala 186:22]
  wire [31:0] n352_I_0_0_t1b_t1b; // @[Top.scala 186:22]
  wire [31:0] n352_O_0_0_t0b; // @[Top.scala 186:22]
  wire [31:0] n352_O_0_0_t1b_t0b; // @[Top.scala 186:22]
  wire [31:0] n352_O_0_0_t1b_t1b; // @[Top.scala 186:22]
  wire  n344_clock; // @[Top.scala 189:22]
  wire  n344_reset; // @[Top.scala 189:22]
  wire  n344_valid_up; // @[Top.scala 189:22]
  wire  n344_valid_down; // @[Top.scala 189:22]
  wire [31:0] n344_I_0_0; // @[Top.scala 189:22]
  wire [31:0] n344_O_0_0; // @[Top.scala 189:22]
  wire  n239_valid_up; // @[Top.scala 192:22]
  wire  n239_valid_down; // @[Top.scala 192:22]
  wire [31:0] n239_I0_0_0; // @[Top.scala 192:22]
  wire [31:0] n239_I1_0_0; // @[Top.scala 192:22]
  wire [31:0] n239_O_0_0_0; // @[Top.scala 192:22]
  wire [31:0] n239_O_0_0_1; // @[Top.scala 192:22]
  wire  n246_valid_up; // @[Top.scala 196:22]
  wire  n246_valid_down; // @[Top.scala 196:22]
  wire [31:0] n246_I0_0_0_0; // @[Top.scala 196:22]
  wire [31:0] n246_I0_0_0_1; // @[Top.scala 196:22]
  wire [31:0] n246_I1_0_0; // @[Top.scala 196:22]
  wire [31:0] n246_O_0_0_0; // @[Top.scala 196:22]
  wire [31:0] n246_O_0_0_1; // @[Top.scala 196:22]
  wire [31:0] n246_O_0_0_2; // @[Top.scala 196:22]
  wire  n253_valid_up; // @[Top.scala 200:22]
  wire  n253_valid_down; // @[Top.scala 200:22]
  wire [31:0] n253_I0_0_0_0; // @[Top.scala 200:22]
  wire [31:0] n253_I0_0_0_1; // @[Top.scala 200:22]
  wire [31:0] n253_I0_0_0_2; // @[Top.scala 200:22]
  wire [31:0] n253_I1_0_0; // @[Top.scala 200:22]
  wire [31:0] n253_O_0_0_0; // @[Top.scala 200:22]
  wire [31:0] n253_O_0_0_1; // @[Top.scala 200:22]
  wire [31:0] n253_O_0_0_2; // @[Top.scala 200:22]
  wire [31:0] n253_O_0_0_3; // @[Top.scala 200:22]
  wire  n264_valid_up; // @[Top.scala 204:22]
  wire  n264_valid_down; // @[Top.scala 204:22]
  wire [31:0] n264_I_0_0_0; // @[Top.scala 204:22]
  wire [31:0] n264_I_0_0_1; // @[Top.scala 204:22]
  wire [31:0] n264_I_0_0_2; // @[Top.scala 204:22]
  wire [31:0] n264_I_0_0_3; // @[Top.scala 204:22]
  wire [31:0] n264_O_0_0; // @[Top.scala 204:22]
  wire [31:0] n264_O_0_1; // @[Top.scala 204:22]
  wire [31:0] n264_O_0_2; // @[Top.scala 204:22]
  wire [31:0] n264_O_0_3; // @[Top.scala 204:22]
  wire  n269_clock; // @[Top.scala 207:22]
  wire  n269_reset; // @[Top.scala 207:22]
  wire  n269_valid_up; // @[Top.scala 207:22]
  wire  n269_valid_down; // @[Top.scala 207:22]
  wire [31:0] n269_I_0_0; // @[Top.scala 207:22]
  wire [31:0] n269_I_0_1; // @[Top.scala 207:22]
  wire [31:0] n269_I_0_2; // @[Top.scala 207:22]
  wire [31:0] n269_I_0_3; // @[Top.scala 207:22]
  wire [31:0] n269_O_0_0; // @[Top.scala 207:22]
  wire  n276_clock; // @[Top.scala 210:22]
  wire  n276_reset; // @[Top.scala 210:22]
  wire  n276_valid_up; // @[Top.scala 210:22]
  wire  n276_valid_down; // @[Top.scala 210:22]
  wire [31:0] n276_I_0_0; // @[Top.scala 210:22]
  wire [31:0] n276_O_0_0_t0b; // @[Top.scala 210:22]
  wire [7:0] n276_O_0_0_t1b; // @[Top.scala 210:22]
  wire  n281_valid_up; // @[Top.scala 213:22]
  wire  n281_valid_down; // @[Top.scala 213:22]
  wire [31:0] n281_I_0_0_t0b; // @[Top.scala 213:22]
  wire [7:0] n281_I_0_0_t1b; // @[Top.scala 213:22]
  wire [31:0] n281_O_0_0; // @[Top.scala 213:22]
  wire  n284_valid_up; // @[Top.scala 216:22]
  wire  n284_valid_down; // @[Top.scala 216:22]
  wire [31:0] n284_I_0_0; // @[Top.scala 216:22]
  wire [31:0] n284_O_0_0; // @[Top.scala 216:22]
  wire  n287_valid_up; // @[Top.scala 219:22]
  wire  n287_valid_down; // @[Top.scala 219:22]
  wire [31:0] n287_I_0_2; // @[Top.scala 219:22]
  wire [31:0] n287_O_0_0; // @[Top.scala 219:22]
  wire  n288_valid_up; // @[Top.scala 222:22]
  wire  n288_valid_down; // @[Top.scala 222:22]
  wire [31:0] n288_I0_0_0; // @[Top.scala 222:22]
  wire [31:0] n288_I1_0_0; // @[Top.scala 222:22]
  wire [31:0] n288_O_0_0_0; // @[Top.scala 222:22]
  wire [31:0] n288_O_0_0_1; // @[Top.scala 222:22]
  wire  n297_valid_up; // @[Top.scala 226:22]
  wire  n297_valid_down; // @[Top.scala 226:22]
  wire [31:0] n297_I_0_0; // @[Top.scala 226:22]
  wire [31:0] n297_O_0_0; // @[Top.scala 226:22]
  wire  n298_valid_up; // @[Top.scala 229:22]
  wire  n298_valid_down; // @[Top.scala 229:22]
  wire [31:0] n298_I0_0_0_0; // @[Top.scala 229:22]
  wire [31:0] n298_I0_0_0_1; // @[Top.scala 229:22]
  wire [31:0] n298_I1_0_0; // @[Top.scala 229:22]
  wire [31:0] n298_O_0_0_0; // @[Top.scala 229:22]
  wire [31:0] n298_O_0_0_1; // @[Top.scala 229:22]
  wire [31:0] n298_O_0_0_2; // @[Top.scala 229:22]
  wire  n307_valid_up; // @[Top.scala 233:22]
  wire  n307_valid_down; // @[Top.scala 233:22]
  wire [31:0] n307_I_0_2; // @[Top.scala 233:22]
  wire [31:0] n307_O_0_0; // @[Top.scala 233:22]
  wire  n308_valid_up; // @[Top.scala 236:22]
  wire  n308_valid_down; // @[Top.scala 236:22]
  wire [31:0] n308_I0_0_0_0; // @[Top.scala 236:22]
  wire [31:0] n308_I0_0_0_1; // @[Top.scala 236:22]
  wire [31:0] n308_I0_0_0_2; // @[Top.scala 236:22]
  wire [31:0] n308_I1_0_0; // @[Top.scala 236:22]
  wire [31:0] n308_O_0_0_0; // @[Top.scala 236:22]
  wire [31:0] n308_O_0_0_1; // @[Top.scala 236:22]
  wire [31:0] n308_O_0_0_2; // @[Top.scala 236:22]
  wire [31:0] n308_O_0_0_3; // @[Top.scala 236:22]
  wire  n319_valid_up; // @[Top.scala 240:22]
  wire  n319_valid_down; // @[Top.scala 240:22]
  wire [31:0] n319_I_0_0_0; // @[Top.scala 240:22]
  wire [31:0] n319_I_0_0_1; // @[Top.scala 240:22]
  wire [31:0] n319_I_0_0_2; // @[Top.scala 240:22]
  wire [31:0] n319_I_0_0_3; // @[Top.scala 240:22]
  wire [31:0] n319_O_0_0; // @[Top.scala 240:22]
  wire [31:0] n319_O_0_1; // @[Top.scala 240:22]
  wire [31:0] n319_O_0_2; // @[Top.scala 240:22]
  wire [31:0] n319_O_0_3; // @[Top.scala 240:22]
  wire  n324_clock; // @[Top.scala 243:22]
  wire  n324_reset; // @[Top.scala 243:22]
  wire  n324_valid_up; // @[Top.scala 243:22]
  wire  n324_valid_down; // @[Top.scala 243:22]
  wire [31:0] n324_I_0_0; // @[Top.scala 243:22]
  wire [31:0] n324_I_0_1; // @[Top.scala 243:22]
  wire [31:0] n324_I_0_2; // @[Top.scala 243:22]
  wire [31:0] n324_I_0_3; // @[Top.scala 243:22]
  wire [31:0] n324_O_0_0; // @[Top.scala 243:22]
  wire  n331_clock; // @[Top.scala 246:22]
  wire  n331_reset; // @[Top.scala 246:22]
  wire  n331_valid_up; // @[Top.scala 246:22]
  wire  n331_valid_down; // @[Top.scala 246:22]
  wire [31:0] n331_I_0_0; // @[Top.scala 246:22]
  wire [31:0] n331_O_0_0_t0b; // @[Top.scala 246:22]
  wire [7:0] n331_O_0_0_t1b; // @[Top.scala 246:22]
  wire  n336_valid_up; // @[Top.scala 249:22]
  wire  n336_valid_down; // @[Top.scala 249:22]
  wire [31:0] n336_I_0_0_t0b; // @[Top.scala 249:22]
  wire [7:0] n336_I_0_0_t1b; // @[Top.scala 249:22]
  wire [31:0] n336_O_0_0; // @[Top.scala 249:22]
  wire  n337_valid_up; // @[Top.scala 252:22]
  wire  n337_valid_down; // @[Top.scala 252:22]
  wire [31:0] n337_I0_0_0; // @[Top.scala 252:22]
  wire [31:0] n337_I1_0_0; // @[Top.scala 252:22]
  wire [31:0] n337_O_0_0_t0b; // @[Top.scala 252:22]
  wire [31:0] n337_O_0_0_t1b; // @[Top.scala 252:22]
  wire  n345_valid_up; // @[Top.scala 256:22]
  wire  n345_valid_down; // @[Top.scala 256:22]
  wire [31:0] n345_I0_0_0; // @[Top.scala 256:22]
  wire [31:0] n345_I1_0_0_t0b; // @[Top.scala 256:22]
  wire [31:0] n345_I1_0_0_t1b; // @[Top.scala 256:22]
  wire [31:0] n345_O_0_0_t0b; // @[Top.scala 256:22]
  wire [31:0] n345_O_0_0_t1b_t0b; // @[Top.scala 256:22]
  wire [31:0] n345_O_0_0_t1b_t1b; // @[Top.scala 256:22]
  wire  n353_valid_up; // @[Top.scala 260:22]
  wire  n353_valid_down; // @[Top.scala 260:22]
  wire [31:0] n353_I0_0_0_t0b; // @[Top.scala 260:22]
  wire [31:0] n353_I0_0_0_t1b_t0b; // @[Top.scala 260:22]
  wire [31:0] n353_I0_0_0_t1b_t1b; // @[Top.scala 260:22]
  wire [31:0] n353_I1_0_0_t0b; // @[Top.scala 260:22]
  wire [31:0] n353_I1_0_0_t1b_t0b; // @[Top.scala 260:22]
  wire [31:0] n353_I1_0_0_t1b_t1b; // @[Top.scala 260:22]
  wire [31:0] n353_O_0_0_t0b_t0b; // @[Top.scala 260:22]
  wire [31:0] n353_O_0_0_t0b_t1b_t0b; // @[Top.scala 260:22]
  wire [31:0] n353_O_0_0_t0b_t1b_t1b; // @[Top.scala 260:22]
  wire [31:0] n353_O_0_0_t1b_t0b; // @[Top.scala 260:22]
  wire [31:0] n353_O_0_0_t1b_t1b_t0b; // @[Top.scala 260:22]
  wire [31:0] n353_O_0_0_t1b_t1b_t1b; // @[Top.scala 260:22]
  wire  n361_valid_up; // @[Top.scala 264:22]
  wire  n361_valid_down; // @[Top.scala 264:22]
  wire  n361_I0_0_0; // @[Top.scala 264:22]
  wire [31:0] n361_I1_0_0_t0b_t0b; // @[Top.scala 264:22]
  wire [31:0] n361_I1_0_0_t0b_t1b_t0b; // @[Top.scala 264:22]
  wire [31:0] n361_I1_0_0_t0b_t1b_t1b; // @[Top.scala 264:22]
  wire [31:0] n361_I1_0_0_t1b_t0b; // @[Top.scala 264:22]
  wire [31:0] n361_I1_0_0_t1b_t1b_t0b; // @[Top.scala 264:22]
  wire [31:0] n361_I1_0_0_t1b_t1b_t1b; // @[Top.scala 264:22]
  wire  n361_O_0_0_t0b; // @[Top.scala 264:22]
  wire [31:0] n361_O_0_0_t1b_t0b_t0b; // @[Top.scala 264:22]
  wire [31:0] n361_O_0_0_t1b_t0b_t1b_t0b; // @[Top.scala 264:22]
  wire [31:0] n361_O_0_0_t1b_t0b_t1b_t1b; // @[Top.scala 264:22]
  wire [31:0] n361_O_0_0_t1b_t1b_t0b; // @[Top.scala 264:22]
  wire [31:0] n361_O_0_0_t1b_t1b_t1b_t0b; // @[Top.scala 264:22]
  wire [31:0] n361_O_0_0_t1b_t1b_t1b_t1b; // @[Top.scala 264:22]
  wire  n372_valid_up; // @[Top.scala 268:22]
  wire  n372_valid_down; // @[Top.scala 268:22]
  wire  n372_I_0_0_t0b; // @[Top.scala 268:22]
  wire [31:0] n372_I_0_0_t1b_t0b_t0b; // @[Top.scala 268:22]
  wire [31:0] n372_I_0_0_t1b_t0b_t1b_t0b; // @[Top.scala 268:22]
  wire [31:0] n372_I_0_0_t1b_t0b_t1b_t1b; // @[Top.scala 268:22]
  wire [31:0] n372_I_0_0_t1b_t1b_t0b; // @[Top.scala 268:22]
  wire [31:0] n372_I_0_0_t1b_t1b_t1b_t0b; // @[Top.scala 268:22]
  wire [31:0] n372_I_0_0_t1b_t1b_t1b_t1b; // @[Top.scala 268:22]
  wire [31:0] n372_O_0_0_t0b; // @[Top.scala 268:22]
  wire [31:0] n372_O_0_0_t1b_t0b; // @[Top.scala 268:22]
  wire [31:0] n372_O_0_0_t1b_t1b; // @[Top.scala 268:22]
  wire  n410_clock; // @[Top.scala 271:22]
  wire  n410_reset; // @[Top.scala 271:22]
  wire  n410_valid_up; // @[Top.scala 271:22]
  wire  n410_valid_down; // @[Top.scala 271:22]
  wire  n410_I_0_0; // @[Top.scala 271:22]
  wire  n410_O_0_0; // @[Top.scala 271:22]
  wire  n373_clock; // @[Top.scala 274:22]
  wire  n373_reset; // @[Top.scala 274:22]
  wire  n373_valid_up; // @[Top.scala 274:22]
  wire  n373_valid_down; // @[Top.scala 274:22]
  wire [31:0] n373_I_0_0; // @[Top.scala 274:22]
  wire [31:0] n373_O_0_0; // @[Top.scala 274:22]
  wire  n374_valid_up; // @[Top.scala 277:22]
  wire  n374_valid_down; // @[Top.scala 277:22]
  wire [31:0] n374_I0_0_0; // @[Top.scala 277:22]
  wire [31:0] n374_I1_0_0; // @[Top.scala 277:22]
  wire [31:0] n374_O_0_0_t0b; // @[Top.scala 277:22]
  wire [31:0] n374_O_0_0_t1b; // @[Top.scala 277:22]
  wire  n381_valid_up; // @[Top.scala 281:22]
  wire  n381_valid_down; // @[Top.scala 281:22]
  wire [31:0] n381_I0_0_0; // @[Top.scala 281:22]
  wire [31:0] n381_I1_0_0_t0b; // @[Top.scala 281:22]
  wire [31:0] n381_I1_0_0_t1b; // @[Top.scala 281:22]
  wire [31:0] n381_O_0_0_t0b; // @[Top.scala 281:22]
  wire [31:0] n381_O_0_0_t1b_t0b; // @[Top.scala 281:22]
  wire [31:0] n381_O_0_0_t1b_t1b; // @[Top.scala 281:22]
  wire  n388_valid_up; // @[Top.scala 285:22]
  wire  n388_valid_down; // @[Top.scala 285:22]
  wire [31:0] n388_I0_0_0; // @[Top.scala 285:22]
  wire [31:0] n388_I1_0_0; // @[Top.scala 285:22]
  wire [31:0] n388_O_0_0_t0b; // @[Top.scala 285:22]
  wire [31:0] n388_O_0_0_t1b; // @[Top.scala 285:22]
  wire  n395_valid_up; // @[Top.scala 289:22]
  wire  n395_valid_down; // @[Top.scala 289:22]
  wire [31:0] n395_I0_0_0; // @[Top.scala 289:22]
  wire [31:0] n395_I1_0_0_t0b; // @[Top.scala 289:22]
  wire [31:0] n395_I1_0_0_t1b; // @[Top.scala 289:22]
  wire [31:0] n395_O_0_0_t0b; // @[Top.scala 289:22]
  wire [31:0] n395_O_0_0_t1b_t0b; // @[Top.scala 289:22]
  wire [31:0] n395_O_0_0_t1b_t1b; // @[Top.scala 289:22]
  wire  n402_clock; // @[Top.scala 293:22]
  wire  n402_reset; // @[Top.scala 293:22]
  wire  n402_valid_up; // @[Top.scala 293:22]
  wire  n402_valid_down; // @[Top.scala 293:22]
  wire [31:0] n402_I_0_0_t0b; // @[Top.scala 293:22]
  wire [31:0] n402_I_0_0_t1b_t0b; // @[Top.scala 293:22]
  wire [31:0] n402_I_0_0_t1b_t1b; // @[Top.scala 293:22]
  wire [31:0] n402_O_0_0_t0b; // @[Top.scala 293:22]
  wire [31:0] n402_O_0_0_t1b_t0b; // @[Top.scala 293:22]
  wire [31:0] n402_O_0_0_t1b_t1b; // @[Top.scala 293:22]
  wire  n403_valid_up; // @[Top.scala 296:22]
  wire  n403_valid_down; // @[Top.scala 296:22]
  wire [31:0] n403_I0_0_0_t0b; // @[Top.scala 296:22]
  wire [31:0] n403_I0_0_0_t1b_t0b; // @[Top.scala 296:22]
  wire [31:0] n403_I0_0_0_t1b_t1b; // @[Top.scala 296:22]
  wire [31:0] n403_I1_0_0_t0b; // @[Top.scala 296:22]
  wire [31:0] n403_I1_0_0_t1b_t0b; // @[Top.scala 296:22]
  wire [31:0] n403_I1_0_0_t1b_t1b; // @[Top.scala 296:22]
  wire [31:0] n403_O_0_0_t0b_t0b; // @[Top.scala 296:22]
  wire [31:0] n403_O_0_0_t0b_t1b_t0b; // @[Top.scala 296:22]
  wire [31:0] n403_O_0_0_t0b_t1b_t1b; // @[Top.scala 296:22]
  wire [31:0] n403_O_0_0_t1b_t0b; // @[Top.scala 296:22]
  wire [31:0] n403_O_0_0_t1b_t1b_t0b; // @[Top.scala 296:22]
  wire [31:0] n403_O_0_0_t1b_t1b_t1b; // @[Top.scala 296:22]
  wire  n411_valid_up; // @[Top.scala 300:22]
  wire  n411_valid_down; // @[Top.scala 300:22]
  wire  n411_I0_0_0; // @[Top.scala 300:22]
  wire [31:0] n411_I1_0_0_t0b_t0b; // @[Top.scala 300:22]
  wire [31:0] n411_I1_0_0_t0b_t1b_t0b; // @[Top.scala 300:22]
  wire [31:0] n411_I1_0_0_t0b_t1b_t1b; // @[Top.scala 300:22]
  wire [31:0] n411_I1_0_0_t1b_t0b; // @[Top.scala 300:22]
  wire [31:0] n411_I1_0_0_t1b_t1b_t0b; // @[Top.scala 300:22]
  wire [31:0] n411_I1_0_0_t1b_t1b_t1b; // @[Top.scala 300:22]
  wire  n411_O_0_0_t0b; // @[Top.scala 300:22]
  wire [31:0] n411_O_0_0_t1b_t0b_t0b; // @[Top.scala 300:22]
  wire [31:0] n411_O_0_0_t1b_t0b_t1b_t0b; // @[Top.scala 300:22]
  wire [31:0] n411_O_0_0_t1b_t0b_t1b_t1b; // @[Top.scala 300:22]
  wire [31:0] n411_O_0_0_t1b_t1b_t0b; // @[Top.scala 300:22]
  wire [31:0] n411_O_0_0_t1b_t1b_t1b_t0b; // @[Top.scala 300:22]
  wire [31:0] n411_O_0_0_t1b_t1b_t1b_t1b; // @[Top.scala 300:22]
  wire  n422_valid_up; // @[Top.scala 304:22]
  wire  n422_valid_down; // @[Top.scala 304:22]
  wire  n422_I_0_0_t0b; // @[Top.scala 304:22]
  wire [31:0] n422_I_0_0_t1b_t0b_t0b; // @[Top.scala 304:22]
  wire [31:0] n422_I_0_0_t1b_t0b_t1b_t0b; // @[Top.scala 304:22]
  wire [31:0] n422_I_0_0_t1b_t0b_t1b_t1b; // @[Top.scala 304:22]
  wire [31:0] n422_I_0_0_t1b_t1b_t0b; // @[Top.scala 304:22]
  wire [31:0] n422_I_0_0_t1b_t1b_t1b_t0b; // @[Top.scala 304:22]
  wire [31:0] n422_I_0_0_t1b_t1b_t1b_t1b; // @[Top.scala 304:22]
  wire [31:0] n422_O_0_0_t0b; // @[Top.scala 304:22]
  wire [31:0] n422_O_0_0_t1b_t0b; // @[Top.scala 304:22]
  wire [31:0] n422_O_0_0_t1b_t1b; // @[Top.scala 304:22]
  wire  n423_valid_up; // @[Top.scala 307:22]
  wire  n423_valid_down; // @[Top.scala 307:22]
  wire [31:0] n423_I0_0_0_t0b; // @[Top.scala 307:22]
  wire [31:0] n423_I0_0_0_t1b_t0b; // @[Top.scala 307:22]
  wire [31:0] n423_I0_0_0_t1b_t1b; // @[Top.scala 307:22]
  wire [31:0] n423_I1_0_0_t0b; // @[Top.scala 307:22]
  wire [31:0] n423_I1_0_0_t1b_t0b; // @[Top.scala 307:22]
  wire [31:0] n423_I1_0_0_t1b_t1b; // @[Top.scala 307:22]
  wire [31:0] n423_O_0_0_t0b_t0b; // @[Top.scala 307:22]
  wire [31:0] n423_O_0_0_t0b_t1b_t0b; // @[Top.scala 307:22]
  wire [31:0] n423_O_0_0_t0b_t1b_t1b; // @[Top.scala 307:22]
  wire [31:0] n423_O_0_0_t1b_t0b; // @[Top.scala 307:22]
  wire [31:0] n423_O_0_0_t1b_t1b_t0b; // @[Top.scala 307:22]
  wire [31:0] n423_O_0_0_t1b_t1b_t1b; // @[Top.scala 307:22]
  wire  n431_valid_up; // @[Top.scala 311:22]
  wire  n431_valid_down; // @[Top.scala 311:22]
  wire  n431_I0_0_0; // @[Top.scala 311:22]
  wire [31:0] n431_I1_0_0_t0b_t0b; // @[Top.scala 311:22]
  wire [31:0] n431_I1_0_0_t0b_t1b_t0b; // @[Top.scala 311:22]
  wire [31:0] n431_I1_0_0_t0b_t1b_t1b; // @[Top.scala 311:22]
  wire [31:0] n431_I1_0_0_t1b_t0b; // @[Top.scala 311:22]
  wire [31:0] n431_I1_0_0_t1b_t1b_t0b; // @[Top.scala 311:22]
  wire [31:0] n431_I1_0_0_t1b_t1b_t1b; // @[Top.scala 311:22]
  wire  n431_O_0_0_t0b; // @[Top.scala 311:22]
  wire [31:0] n431_O_0_0_t1b_t0b_t0b; // @[Top.scala 311:22]
  wire [31:0] n431_O_0_0_t1b_t0b_t1b_t0b; // @[Top.scala 311:22]
  wire [31:0] n431_O_0_0_t1b_t0b_t1b_t1b; // @[Top.scala 311:22]
  wire [31:0] n431_O_0_0_t1b_t1b_t0b; // @[Top.scala 311:22]
  wire [31:0] n431_O_0_0_t1b_t1b_t1b_t0b; // @[Top.scala 311:22]
  wire [31:0] n431_O_0_0_t1b_t1b_t1b_t1b; // @[Top.scala 311:22]
  wire  n442_valid_up; // @[Top.scala 315:22]
  wire  n442_valid_down; // @[Top.scala 315:22]
  wire  n442_I_0_0_t0b; // @[Top.scala 315:22]
  wire [31:0] n442_I_0_0_t1b_t0b_t0b; // @[Top.scala 315:22]
  wire [31:0] n442_I_0_0_t1b_t0b_t1b_t0b; // @[Top.scala 315:22]
  wire [31:0] n442_I_0_0_t1b_t0b_t1b_t1b; // @[Top.scala 315:22]
  wire [31:0] n442_I_0_0_t1b_t1b_t0b; // @[Top.scala 315:22]
  wire [31:0] n442_I_0_0_t1b_t1b_t1b_t0b; // @[Top.scala 315:22]
  wire [31:0] n442_I_0_0_t1b_t1b_t1b_t1b; // @[Top.scala 315:22]
  wire [31:0] n442_O_0_0_t0b; // @[Top.scala 315:22]
  wire [31:0] n442_O_0_0_t1b_t0b; // @[Top.scala 315:22]
  wire [31:0] n442_O_0_0_t1b_t1b; // @[Top.scala 315:22]
  MapS_7 n152 ( // @[Top.scala 116:22]
    .valid_up(n152_valid_up),
    .valid_down(n152_valid_down),
    .I_0_0_t0b(n152_I_0_0_t0b),
    .O_0_0(n152_O_0_0)
  );
  FIFO_2 n430 ( // @[Top.scala 119:22]
    .clock(n430_clock),
    .reset(n430_reset),
    .valid_up(n430_valid_up),
    .valid_down(n430_valid_down),
    .I_0_0(n430_I_0_0),
    .O_0_0(n430_O_0_0)
  );
  MapS_9 n157 ( // @[Top.scala 122:22]
    .valid_up(n157_valid_up),
    .valid_down(n157_valid_down),
    .I_0_0_t1b(n157_I_0_0_t1b),
    .O_0_0(n157_O_0_0)
  );
  FIFO_2 n360 ( // @[Top.scala 125:22]
    .clock(n360_clock),
    .reset(n360_reset),
    .valid_up(n360_valid_up),
    .valid_down(n360_valid_down),
    .I_0_0(n360_I_0_0),
    .O_0_0(n360_O_0_0)
  );
  DownS n159 ( // @[Top.scala 128:22]
    .valid_up(n159_valid_up),
    .valid_down(n159_valid_down),
    .I_1_0(n159_I_1_0),
    .I_1_1(n159_I_1_1),
    .I_1_2(n159_I_1_2),
    .O_0_0(n159_O_0_0),
    .O_0_1(n159_O_0_1),
    .O_0_2(n159_O_0_2)
  );
  MapS_10 n162 ( // @[Top.scala 131:22]
    .valid_up(n162_valid_up),
    .valid_down(n162_valid_down),
    .I_0_0(n162_I_0_0),
    .O_0_0(n162_O_0_0)
  );
  MapS_11 n165 ( // @[Top.scala 134:22]
    .valid_up(n165_valid_up),
    .valid_down(n165_valid_down),
    .I_0_2(n165_I_0_2),
    .O_0_0(n165_O_0_0)
  );
  Map2S_10 n166 ( // @[Top.scala 137:22]
    .valid_up(n166_valid_up),
    .valid_down(n166_valid_down),
    .I0_0_0(n166_I0_0_0),
    .I1_0_0(n166_I1_0_0),
    .O_0_0_t0b(n166_O_0_0_t0b),
    .O_0_0_t1b(n166_O_0_0_t1b)
  );
  MapS_13 n177 ( // @[Top.scala 141:22]
    .valid_up(n177_valid_up),
    .valid_down(n177_valid_down),
    .I_0_0_t0b(n177_I_0_0_t0b),
    .I_0_0_t1b(n177_I_0_0_t1b),
    .O_0_0(n177_O_0_0)
  );
  MapS_15 n184 ( // @[Top.scala 144:22]
    .clock(n184_clock),
    .reset(n184_reset),
    .valid_up(n184_valid_up),
    .valid_down(n184_valid_down),
    .I_0_0(n184_I_0_0),
    .O_0_0_t0b(n184_O_0_0_t0b),
    .O_0_0_t1b(n184_O_0_0_t1b)
  );
  MapS_17 n189 ( // @[Top.scala 147:22]
    .valid_up(n189_valid_up),
    .valid_down(n189_valid_down),
    .I_0_0_t0b(n189_I_0_0_t0b),
    .I_0_0_t1b(n189_I_0_0_t1b),
    .O_0_0(n189_O_0_0)
  );
  MapS_18 n192 ( // @[Top.scala 150:22]
    .valid_up(n192_valid_up),
    .valid_down(n192_valid_down),
    .I_0_1(n192_I_0_1),
    .O_0_0(n192_O_0_0)
  );
  DownS_4 n193 ( // @[Top.scala 153:22]
    .valid_up(n193_valid_up),
    .valid_down(n193_valid_down),
    .I_0_0(n193_I_0_0),
    .I_0_1(n193_I_0_1),
    .I_0_2(n193_I_0_2),
    .O_0_0(n193_O_0_0),
    .O_0_1(n193_O_0_1),
    .O_0_2(n193_O_0_2)
  );
  MapS_18 n196 ( // @[Top.scala 156:22]
    .valid_up(n196_valid_up),
    .valid_down(n196_valid_down),
    .I_0_1(n196_I_0_1),
    .O_0_0(n196_O_0_0)
  );
  DownS_6 n197 ( // @[Top.scala 159:22]
    .valid_up(n197_valid_up),
    .valid_down(n197_valid_down),
    .I_2_0(n197_I_2_0),
    .I_2_1(n197_I_2_1),
    .I_2_2(n197_I_2_2),
    .O_0_0(n197_O_0_0),
    .O_0_1(n197_O_0_1),
    .O_0_2(n197_O_0_2)
  );
  MapS_18 n200 ( // @[Top.scala 162:22]
    .valid_up(n200_valid_up),
    .valid_down(n200_valid_down),
    .I_0_1(n200_I_0_1),
    .O_0_0(n200_O_0_0)
  );
  Map2S_10 n201 ( // @[Top.scala 165:22]
    .valid_up(n201_valid_up),
    .valid_down(n201_valid_down),
    .I0_0_0(n201_I0_0_0),
    .I1_0_0(n201_I1_0_0),
    .O_0_0_t0b(n201_O_0_0_t0b),
    .O_0_0_t1b(n201_O_0_0_t1b)
  );
  MapS_13 n212 ( // @[Top.scala 169:22]
    .valid_up(n212_valid_up),
    .valid_down(n212_valid_down),
    .I_0_0_t0b(n212_I_0_0_t0b),
    .I_0_0_t1b(n212_I_0_0_t1b),
    .O_0_0(n212_O_0_0)
  );
  MapS_15 n219 ( // @[Top.scala 172:22]
    .clock(n219_clock),
    .reset(n219_reset),
    .valid_up(n219_valid_up),
    .valid_down(n219_valid_down),
    .I_0_0(n219_I_0_0),
    .O_0_0_t0b(n219_O_0_0_t0b),
    .O_0_0_t1b(n219_O_0_0_t1b)
  );
  MapS_17 n224 ( // @[Top.scala 175:22]
    .valid_up(n224_valid_up),
    .valid_down(n224_valid_down),
    .I_0_0_t0b(n224_I_0_0_t0b),
    .I_0_0_t1b(n224_I_0_0_t1b),
    .O_0_0(n224_O_0_0)
  );
  Map2S_10 n225 ( // @[Top.scala 178:22]
    .valid_up(n225_valid_up),
    .valid_down(n225_valid_down),
    .I0_0_0(n225_I0_0_0),
    .I1_0_0(n225_I1_0_0),
    .O_0_0_t0b(n225_O_0_0_t0b),
    .O_0_0_t1b(n225_O_0_0_t1b)
  );
  Map2S_16 n232 ( // @[Top.scala 182:22]
    .valid_up(n232_valid_up),
    .valid_down(n232_valid_down),
    .I0_0_0(n232_I0_0_0),
    .I1_0_0_t0b(n232_I1_0_0_t0b),
    .I1_0_0_t1b(n232_I1_0_0_t1b),
    .O_0_0_t0b(n232_O_0_0_t0b),
    .O_0_0_t1b_t0b(n232_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(n232_O_0_0_t1b_t1b)
  );
  FIFO_4 n352 ( // @[Top.scala 186:22]
    .clock(n352_clock),
    .reset(n352_reset),
    .valid_up(n352_valid_up),
    .valid_down(n352_valid_down),
    .I_0_0_t0b(n352_I_0_0_t0b),
    .I_0_0_t1b_t0b(n352_I_0_0_t1b_t0b),
    .I_0_0_t1b_t1b(n352_I_0_0_t1b_t1b),
    .O_0_0_t0b(n352_O_0_0_t0b),
    .O_0_0_t1b_t0b(n352_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(n352_O_0_0_t1b_t1b)
  );
  FIFO_5 n344 ( // @[Top.scala 189:22]
    .clock(n344_clock),
    .reset(n344_reset),
    .valid_up(n344_valid_up),
    .valid_down(n344_valid_down),
    .I_0_0(n344_I_0_0),
    .O_0_0(n344_O_0_0)
  );
  Map2S_18 n239 ( // @[Top.scala 192:22]
    .valid_up(n239_valid_up),
    .valid_down(n239_valid_down),
    .I0_0_0(n239_I0_0_0),
    .I1_0_0(n239_I1_0_0),
    .O_0_0_0(n239_O_0_0_0),
    .O_0_0_1(n239_O_0_0_1)
  );
  Map2S_20 n246 ( // @[Top.scala 196:22]
    .valid_up(n246_valid_up),
    .valid_down(n246_valid_down),
    .I0_0_0_0(n246_I0_0_0_0),
    .I0_0_0_1(n246_I0_0_0_1),
    .I1_0_0(n246_I1_0_0),
    .O_0_0_0(n246_O_0_0_0),
    .O_0_0_1(n246_O_0_0_1),
    .O_0_0_2(n246_O_0_0_2)
  );
  Map2S_22 n253 ( // @[Top.scala 200:22]
    .valid_up(n253_valid_up),
    .valid_down(n253_valid_down),
    .I0_0_0_0(n253_I0_0_0_0),
    .I0_0_0_1(n253_I0_0_0_1),
    .I0_0_0_2(n253_I0_0_0_2),
    .I1_0_0(n253_I1_0_0),
    .O_0_0_0(n253_O_0_0_0),
    .O_0_0_1(n253_O_0_0_1),
    .O_0_0_2(n253_O_0_0_2),
    .O_0_0_3(n253_O_0_0_3)
  );
  MapS_27 n264 ( // @[Top.scala 204:22]
    .valid_up(n264_valid_up),
    .valid_down(n264_valid_down),
    .I_0_0_0(n264_I_0_0_0),
    .I_0_0_1(n264_I_0_0_1),
    .I_0_0_2(n264_I_0_0_2),
    .I_0_0_3(n264_I_0_0_3),
    .O_0_0(n264_O_0_0),
    .O_0_1(n264_O_0_1),
    .O_0_2(n264_O_0_2),
    .O_0_3(n264_O_0_3)
  );
  MapS_28 n269 ( // @[Top.scala 207:22]
    .clock(n269_clock),
    .reset(n269_reset),
    .valid_up(n269_valid_up),
    .valid_down(n269_valid_down),
    .I_0_0(n269_I_0_0),
    .I_0_1(n269_I_0_1),
    .I_0_2(n269_I_0_2),
    .I_0_3(n269_I_0_3),
    .O_0_0(n269_O_0_0)
  );
  MapS_30 n276 ( // @[Top.scala 210:22]
    .clock(n276_clock),
    .reset(n276_reset),
    .valid_up(n276_valid_up),
    .valid_down(n276_valid_down),
    .I_0_0(n276_I_0_0),
    .O_0_0_t0b(n276_O_0_0_t0b),
    .O_0_0_t1b(n276_O_0_0_t1b)
  );
  MapS_17 n281 ( // @[Top.scala 213:22]
    .valid_up(n281_valid_up),
    .valid_down(n281_valid_down),
    .I_0_0_t0b(n281_I_0_0_t0b),
    .I_0_0_t1b(n281_I_0_0_t1b),
    .O_0_0(n281_O_0_0)
  );
  MapS_10 n284 ( // @[Top.scala 216:22]
    .valid_up(n284_valid_up),
    .valid_down(n284_valid_down),
    .I_0_0(n284_I_0_0),
    .O_0_0(n284_O_0_0)
  );
  MapS_11 n287 ( // @[Top.scala 219:22]
    .valid_up(n287_valid_up),
    .valid_down(n287_valid_down),
    .I_0_2(n287_I_0_2),
    .O_0_0(n287_O_0_0)
  );
  Map2S_18 n288 ( // @[Top.scala 222:22]
    .valid_up(n288_valid_up),
    .valid_down(n288_valid_down),
    .I0_0_0(n288_I0_0_0),
    .I1_0_0(n288_I1_0_0),
    .O_0_0_0(n288_O_0_0_0),
    .O_0_0_1(n288_O_0_0_1)
  );
  MapS_10 n297 ( // @[Top.scala 226:22]
    .valid_up(n297_valid_up),
    .valid_down(n297_valid_down),
    .I_0_0(n297_I_0_0),
    .O_0_0(n297_O_0_0)
  );
  Map2S_20 n298 ( // @[Top.scala 229:22]
    .valid_up(n298_valid_up),
    .valid_down(n298_valid_down),
    .I0_0_0_0(n298_I0_0_0_0),
    .I0_0_0_1(n298_I0_0_0_1),
    .I1_0_0(n298_I1_0_0),
    .O_0_0_0(n298_O_0_0_0),
    .O_0_0_1(n298_O_0_0_1),
    .O_0_0_2(n298_O_0_0_2)
  );
  MapS_11 n307 ( // @[Top.scala 233:22]
    .valid_up(n307_valid_up),
    .valid_down(n307_valid_down),
    .I_0_2(n307_I_0_2),
    .O_0_0(n307_O_0_0)
  );
  Map2S_22 n308 ( // @[Top.scala 236:22]
    .valid_up(n308_valid_up),
    .valid_down(n308_valid_down),
    .I0_0_0_0(n308_I0_0_0_0),
    .I0_0_0_1(n308_I0_0_0_1),
    .I0_0_0_2(n308_I0_0_0_2),
    .I1_0_0(n308_I1_0_0),
    .O_0_0_0(n308_O_0_0_0),
    .O_0_0_1(n308_O_0_0_1),
    .O_0_0_2(n308_O_0_0_2),
    .O_0_0_3(n308_O_0_0_3)
  );
  MapS_27 n319 ( // @[Top.scala 240:22]
    .valid_up(n319_valid_up),
    .valid_down(n319_valid_down),
    .I_0_0_0(n319_I_0_0_0),
    .I_0_0_1(n319_I_0_0_1),
    .I_0_0_2(n319_I_0_0_2),
    .I_0_0_3(n319_I_0_0_3),
    .O_0_0(n319_O_0_0),
    .O_0_1(n319_O_0_1),
    .O_0_2(n319_O_0_2),
    .O_0_3(n319_O_0_3)
  );
  MapS_38 n324 ( // @[Top.scala 243:22]
    .clock(n324_clock),
    .reset(n324_reset),
    .valid_up(n324_valid_up),
    .valid_down(n324_valid_down),
    .I_0_0(n324_I_0_0),
    .I_0_1(n324_I_0_1),
    .I_0_2(n324_I_0_2),
    .I_0_3(n324_I_0_3),
    .O_0_0(n324_O_0_0)
  );
  MapS_30 n331 ( // @[Top.scala 246:22]
    .clock(n331_clock),
    .reset(n331_reset),
    .valid_up(n331_valid_up),
    .valid_down(n331_valid_down),
    .I_0_0(n331_I_0_0),
    .O_0_0_t0b(n331_O_0_0_t0b),
    .O_0_0_t1b(n331_O_0_0_t1b)
  );
  MapS_17 n336 ( // @[Top.scala 249:22]
    .valid_up(n336_valid_up),
    .valid_down(n336_valid_down),
    .I_0_0_t0b(n336_I_0_0_t0b),
    .I_0_0_t1b(n336_I_0_0_t1b),
    .O_0_0(n336_O_0_0)
  );
  Map2S_10 n337 ( // @[Top.scala 252:22]
    .valid_up(n337_valid_up),
    .valid_down(n337_valid_down),
    .I0_0_0(n337_I0_0_0),
    .I1_0_0(n337_I1_0_0),
    .O_0_0_t0b(n337_O_0_0_t0b),
    .O_0_0_t1b(n337_O_0_0_t1b)
  );
  Map2S_16 n345 ( // @[Top.scala 256:22]
    .valid_up(n345_valid_up),
    .valid_down(n345_valid_down),
    .I0_0_0(n345_I0_0_0),
    .I1_0_0_t0b(n345_I1_0_0_t0b),
    .I1_0_0_t1b(n345_I1_0_0_t1b),
    .O_0_0_t0b(n345_O_0_0_t0b),
    .O_0_0_t1b_t0b(n345_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(n345_O_0_0_t1b_t1b)
  );
  Map2S_34 n353 ( // @[Top.scala 260:22]
    .valid_up(n353_valid_up),
    .valid_down(n353_valid_down),
    .I0_0_0_t0b(n353_I0_0_0_t0b),
    .I0_0_0_t1b_t0b(n353_I0_0_0_t1b_t0b),
    .I0_0_0_t1b_t1b(n353_I0_0_0_t1b_t1b),
    .I1_0_0_t0b(n353_I1_0_0_t0b),
    .I1_0_0_t1b_t0b(n353_I1_0_0_t1b_t0b),
    .I1_0_0_t1b_t1b(n353_I1_0_0_t1b_t1b),
    .O_0_0_t0b_t0b(n353_O_0_0_t0b_t0b),
    .O_0_0_t0b_t1b_t0b(n353_O_0_0_t0b_t1b_t0b),
    .O_0_0_t0b_t1b_t1b(n353_O_0_0_t0b_t1b_t1b),
    .O_0_0_t1b_t0b(n353_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b_t0b(n353_O_0_0_t1b_t1b_t0b),
    .O_0_0_t1b_t1b_t1b(n353_O_0_0_t1b_t1b_t1b)
  );
  Map2S_36 n361 ( // @[Top.scala 264:22]
    .valid_up(n361_valid_up),
    .valid_down(n361_valid_down),
    .I0_0_0(n361_I0_0_0),
    .I1_0_0_t0b_t0b(n361_I1_0_0_t0b_t0b),
    .I1_0_0_t0b_t1b_t0b(n361_I1_0_0_t0b_t1b_t0b),
    .I1_0_0_t0b_t1b_t1b(n361_I1_0_0_t0b_t1b_t1b),
    .I1_0_0_t1b_t0b(n361_I1_0_0_t1b_t0b),
    .I1_0_0_t1b_t1b_t0b(n361_I1_0_0_t1b_t1b_t0b),
    .I1_0_0_t1b_t1b_t1b(n361_I1_0_0_t1b_t1b_t1b),
    .O_0_0_t0b(n361_O_0_0_t0b),
    .O_0_0_t1b_t0b_t0b(n361_O_0_0_t1b_t0b_t0b),
    .O_0_0_t1b_t0b_t1b_t0b(n361_O_0_0_t1b_t0b_t1b_t0b),
    .O_0_0_t1b_t0b_t1b_t1b(n361_O_0_0_t1b_t0b_t1b_t1b),
    .O_0_0_t1b_t1b_t0b(n361_O_0_0_t1b_t1b_t0b),
    .O_0_0_t1b_t1b_t1b_t0b(n361_O_0_0_t1b_t1b_t1b_t0b),
    .O_0_0_t1b_t1b_t1b_t1b(n361_O_0_0_t1b_t1b_t1b_t1b)
  );
  MapS_44 n372 ( // @[Top.scala 268:22]
    .valid_up(n372_valid_up),
    .valid_down(n372_valid_down),
    .I_0_0_t0b(n372_I_0_0_t0b),
    .I_0_0_t1b_t0b_t0b(n372_I_0_0_t1b_t0b_t0b),
    .I_0_0_t1b_t0b_t1b_t0b(n372_I_0_0_t1b_t0b_t1b_t0b),
    .I_0_0_t1b_t0b_t1b_t1b(n372_I_0_0_t1b_t0b_t1b_t1b),
    .I_0_0_t1b_t1b_t0b(n372_I_0_0_t1b_t1b_t0b),
    .I_0_0_t1b_t1b_t1b_t0b(n372_I_0_0_t1b_t1b_t1b_t0b),
    .I_0_0_t1b_t1b_t1b_t1b(n372_I_0_0_t1b_t1b_t1b_t1b),
    .O_0_0_t0b(n372_O_0_0_t0b),
    .O_0_0_t1b_t0b(n372_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(n372_O_0_0_t1b_t1b)
  );
  FIFO_2 n410 ( // @[Top.scala 271:22]
    .clock(n410_clock),
    .reset(n410_reset),
    .valid_up(n410_valid_up),
    .valid_down(n410_valid_down),
    .I_0_0(n410_I_0_0),
    .O_0_0(n410_O_0_0)
  );
  FIFO_5 n373 ( // @[Top.scala 274:22]
    .clock(n373_clock),
    .reset(n373_reset),
    .valid_up(n373_valid_up),
    .valid_down(n373_valid_down),
    .I_0_0(n373_I_0_0),
    .O_0_0(n373_O_0_0)
  );
  Map2S_10 n374 ( // @[Top.scala 277:22]
    .valid_up(n374_valid_up),
    .valid_down(n374_valid_down),
    .I0_0_0(n374_I0_0_0),
    .I1_0_0(n374_I1_0_0),
    .O_0_0_t0b(n374_O_0_0_t0b),
    .O_0_0_t1b(n374_O_0_0_t1b)
  );
  Map2S_16 n381 ( // @[Top.scala 281:22]
    .valid_up(n381_valid_up),
    .valid_down(n381_valid_down),
    .I0_0_0(n381_I0_0_0),
    .I1_0_0_t0b(n381_I1_0_0_t0b),
    .I1_0_0_t1b(n381_I1_0_0_t1b),
    .O_0_0_t0b(n381_O_0_0_t0b),
    .O_0_0_t1b_t0b(n381_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(n381_O_0_0_t1b_t1b)
  );
  Map2S_10 n388 ( // @[Top.scala 285:22]
    .valid_up(n388_valid_up),
    .valid_down(n388_valid_down),
    .I0_0_0(n388_I0_0_0),
    .I1_0_0(n388_I1_0_0),
    .O_0_0_t0b(n388_O_0_0_t0b),
    .O_0_0_t1b(n388_O_0_0_t1b)
  );
  Map2S_16 n395 ( // @[Top.scala 289:22]
    .valid_up(n395_valid_up),
    .valid_down(n395_valid_down),
    .I0_0_0(n395_I0_0_0),
    .I1_0_0_t0b(n395_I1_0_0_t0b),
    .I1_0_0_t1b(n395_I1_0_0_t1b),
    .O_0_0_t0b(n395_O_0_0_t0b),
    .O_0_0_t1b_t0b(n395_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(n395_O_0_0_t1b_t1b)
  );
  FIFO_4 n402 ( // @[Top.scala 293:22]
    .clock(n402_clock),
    .reset(n402_reset),
    .valid_up(n402_valid_up),
    .valid_down(n402_valid_down),
    .I_0_0_t0b(n402_I_0_0_t0b),
    .I_0_0_t1b_t0b(n402_I_0_0_t1b_t0b),
    .I_0_0_t1b_t1b(n402_I_0_0_t1b_t1b),
    .O_0_0_t0b(n402_O_0_0_t0b),
    .O_0_0_t1b_t0b(n402_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(n402_O_0_0_t1b_t1b)
  );
  Map2S_34 n403 ( // @[Top.scala 296:22]
    .valid_up(n403_valid_up),
    .valid_down(n403_valid_down),
    .I0_0_0_t0b(n403_I0_0_0_t0b),
    .I0_0_0_t1b_t0b(n403_I0_0_0_t1b_t0b),
    .I0_0_0_t1b_t1b(n403_I0_0_0_t1b_t1b),
    .I1_0_0_t0b(n403_I1_0_0_t0b),
    .I1_0_0_t1b_t0b(n403_I1_0_0_t1b_t0b),
    .I1_0_0_t1b_t1b(n403_I1_0_0_t1b_t1b),
    .O_0_0_t0b_t0b(n403_O_0_0_t0b_t0b),
    .O_0_0_t0b_t1b_t0b(n403_O_0_0_t0b_t1b_t0b),
    .O_0_0_t0b_t1b_t1b(n403_O_0_0_t0b_t1b_t1b),
    .O_0_0_t1b_t0b(n403_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b_t0b(n403_O_0_0_t1b_t1b_t0b),
    .O_0_0_t1b_t1b_t1b(n403_O_0_0_t1b_t1b_t1b)
  );
  Map2S_36 n411 ( // @[Top.scala 300:22]
    .valid_up(n411_valid_up),
    .valid_down(n411_valid_down),
    .I0_0_0(n411_I0_0_0),
    .I1_0_0_t0b_t0b(n411_I1_0_0_t0b_t0b),
    .I1_0_0_t0b_t1b_t0b(n411_I1_0_0_t0b_t1b_t0b),
    .I1_0_0_t0b_t1b_t1b(n411_I1_0_0_t0b_t1b_t1b),
    .I1_0_0_t1b_t0b(n411_I1_0_0_t1b_t0b),
    .I1_0_0_t1b_t1b_t0b(n411_I1_0_0_t1b_t1b_t0b),
    .I1_0_0_t1b_t1b_t1b(n411_I1_0_0_t1b_t1b_t1b),
    .O_0_0_t0b(n411_O_0_0_t0b),
    .O_0_0_t1b_t0b_t0b(n411_O_0_0_t1b_t0b_t0b),
    .O_0_0_t1b_t0b_t1b_t0b(n411_O_0_0_t1b_t0b_t1b_t0b),
    .O_0_0_t1b_t0b_t1b_t1b(n411_O_0_0_t1b_t0b_t1b_t1b),
    .O_0_0_t1b_t1b_t0b(n411_O_0_0_t1b_t1b_t0b),
    .O_0_0_t1b_t1b_t1b_t0b(n411_O_0_0_t1b_t1b_t1b_t0b),
    .O_0_0_t1b_t1b_t1b_t1b(n411_O_0_0_t1b_t1b_t1b_t1b)
  );
  MapS_44 n422 ( // @[Top.scala 304:22]
    .valid_up(n422_valid_up),
    .valid_down(n422_valid_down),
    .I_0_0_t0b(n422_I_0_0_t0b),
    .I_0_0_t1b_t0b_t0b(n422_I_0_0_t1b_t0b_t0b),
    .I_0_0_t1b_t0b_t1b_t0b(n422_I_0_0_t1b_t0b_t1b_t0b),
    .I_0_0_t1b_t0b_t1b_t1b(n422_I_0_0_t1b_t0b_t1b_t1b),
    .I_0_0_t1b_t1b_t0b(n422_I_0_0_t1b_t1b_t0b),
    .I_0_0_t1b_t1b_t1b_t0b(n422_I_0_0_t1b_t1b_t1b_t0b),
    .I_0_0_t1b_t1b_t1b_t1b(n422_I_0_0_t1b_t1b_t1b_t1b),
    .O_0_0_t0b(n422_O_0_0_t0b),
    .O_0_0_t1b_t0b(n422_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(n422_O_0_0_t1b_t1b)
  );
  Map2S_34 n423 ( // @[Top.scala 307:22]
    .valid_up(n423_valid_up),
    .valid_down(n423_valid_down),
    .I0_0_0_t0b(n423_I0_0_0_t0b),
    .I0_0_0_t1b_t0b(n423_I0_0_0_t1b_t0b),
    .I0_0_0_t1b_t1b(n423_I0_0_0_t1b_t1b),
    .I1_0_0_t0b(n423_I1_0_0_t0b),
    .I1_0_0_t1b_t0b(n423_I1_0_0_t1b_t0b),
    .I1_0_0_t1b_t1b(n423_I1_0_0_t1b_t1b),
    .O_0_0_t0b_t0b(n423_O_0_0_t0b_t0b),
    .O_0_0_t0b_t1b_t0b(n423_O_0_0_t0b_t1b_t0b),
    .O_0_0_t0b_t1b_t1b(n423_O_0_0_t0b_t1b_t1b),
    .O_0_0_t1b_t0b(n423_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b_t0b(n423_O_0_0_t1b_t1b_t0b),
    .O_0_0_t1b_t1b_t1b(n423_O_0_0_t1b_t1b_t1b)
  );
  Map2S_36 n431 ( // @[Top.scala 311:22]
    .valid_up(n431_valid_up),
    .valid_down(n431_valid_down),
    .I0_0_0(n431_I0_0_0),
    .I1_0_0_t0b_t0b(n431_I1_0_0_t0b_t0b),
    .I1_0_0_t0b_t1b_t0b(n431_I1_0_0_t0b_t1b_t0b),
    .I1_0_0_t0b_t1b_t1b(n431_I1_0_0_t0b_t1b_t1b),
    .I1_0_0_t1b_t0b(n431_I1_0_0_t1b_t0b),
    .I1_0_0_t1b_t1b_t0b(n431_I1_0_0_t1b_t1b_t0b),
    .I1_0_0_t1b_t1b_t1b(n431_I1_0_0_t1b_t1b_t1b),
    .O_0_0_t0b(n431_O_0_0_t0b),
    .O_0_0_t1b_t0b_t0b(n431_O_0_0_t1b_t0b_t0b),
    .O_0_0_t1b_t0b_t1b_t0b(n431_O_0_0_t1b_t0b_t1b_t0b),
    .O_0_0_t1b_t0b_t1b_t1b(n431_O_0_0_t1b_t0b_t1b_t1b),
    .O_0_0_t1b_t1b_t0b(n431_O_0_0_t1b_t1b_t0b),
    .O_0_0_t1b_t1b_t1b_t0b(n431_O_0_0_t1b_t1b_t1b_t0b),
    .O_0_0_t1b_t1b_t1b_t1b(n431_O_0_0_t1b_t1b_t1b_t1b)
  );
  MapS_44 n442 ( // @[Top.scala 315:22]
    .valid_up(n442_valid_up),
    .valid_down(n442_valid_down),
    .I_0_0_t0b(n442_I_0_0_t0b),
    .I_0_0_t1b_t0b_t0b(n442_I_0_0_t1b_t0b_t0b),
    .I_0_0_t1b_t0b_t1b_t0b(n442_I_0_0_t1b_t0b_t1b_t0b),
    .I_0_0_t1b_t0b_t1b_t1b(n442_I_0_0_t1b_t0b_t1b_t1b),
    .I_0_0_t1b_t1b_t0b(n442_I_0_0_t1b_t1b_t0b),
    .I_0_0_t1b_t1b_t1b_t0b(n442_I_0_0_t1b_t1b_t1b_t0b),
    .I_0_0_t1b_t1b_t1b_t1b(n442_I_0_0_t1b_t1b_t1b_t1b),
    .O_0_0_t0b(n442_O_0_0_t0b),
    .O_0_0_t1b_t0b(n442_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(n442_O_0_0_t1b_t1b)
  );
  assign valid_down = n442_valid_down; // @[Top.scala 319:16]
  assign O_0_0_t0b = n442_O_0_0_t0b; // @[Top.scala 318:7]
  assign O_0_0_t1b_t0b = n442_O_0_0_t1b_t0b; // @[Top.scala 318:7]
  assign O_0_0_t1b_t1b = n442_O_0_0_t1b_t1b; // @[Top.scala 318:7]
  assign n152_valid_up = valid_up; // @[Top.scala 118:19]
  assign n152_I_0_0_t0b = I1_0_0_t0b; // @[Top.scala 117:12]
  assign n430_clock = clock;
  assign n430_reset = reset;
  assign n430_valid_up = n152_valid_down; // @[Top.scala 121:19]
  assign n430_I_0_0 = n152_O_0_0; // @[Top.scala 120:12]
  assign n157_valid_up = valid_up; // @[Top.scala 124:19]
  assign n157_I_0_0_t1b = I1_0_0_t1b; // @[Top.scala 123:12]
  assign n360_clock = clock;
  assign n360_reset = reset;
  assign n360_valid_up = n157_valid_down; // @[Top.scala 127:19]
  assign n360_I_0_0 = n157_O_0_0; // @[Top.scala 126:12]
  assign n159_valid_up = valid_up; // @[Top.scala 130:19]
  assign n159_I_1_0 = I0_1_0; // @[Top.scala 129:12]
  assign n159_I_1_1 = I0_1_1; // @[Top.scala 129:12]
  assign n159_I_1_2 = I0_1_2; // @[Top.scala 129:12]
  assign n162_valid_up = n159_valid_down; // @[Top.scala 133:19]
  assign n162_I_0_0 = n159_O_0_0; // @[Top.scala 132:12]
  assign n165_valid_up = n159_valid_down; // @[Top.scala 136:19]
  assign n165_I_0_2 = n159_O_0_2; // @[Top.scala 135:12]
  assign n166_valid_up = n162_valid_down & n165_valid_down; // @[Top.scala 140:19]
  assign n166_I0_0_0 = n162_O_0_0; // @[Top.scala 138:13]
  assign n166_I1_0_0 = n165_O_0_0; // @[Top.scala 139:13]
  assign n177_valid_up = n166_valid_down; // @[Top.scala 143:19]
  assign n177_I_0_0_t0b = n166_O_0_0_t0b; // @[Top.scala 142:12]
  assign n177_I_0_0_t1b = n166_O_0_0_t1b; // @[Top.scala 142:12]
  assign n184_clock = clock;
  assign n184_reset = reset;
  assign n184_valid_up = n177_valid_down; // @[Top.scala 146:19]
  assign n184_I_0_0 = n177_O_0_0; // @[Top.scala 145:12]
  assign n189_valid_up = n184_valid_down; // @[Top.scala 149:19]
  assign n189_I_0_0_t0b = n184_O_0_0_t0b; // @[Top.scala 148:12]
  assign n189_I_0_0_t1b = n184_O_0_0_t1b; // @[Top.scala 148:12]
  assign n192_valid_up = n159_valid_down; // @[Top.scala 152:19]
  assign n192_I_0_1 = n159_O_0_1; // @[Top.scala 151:12]
  assign n193_valid_up = valid_up; // @[Top.scala 155:19]
  assign n193_I_0_0 = I0_0_0; // @[Top.scala 154:12]
  assign n193_I_0_1 = I0_0_1; // @[Top.scala 154:12]
  assign n193_I_0_2 = I0_0_2; // @[Top.scala 154:12]
  assign n196_valid_up = n193_valid_down; // @[Top.scala 158:19]
  assign n196_I_0_1 = n193_O_0_1; // @[Top.scala 157:12]
  assign n197_valid_up = valid_up; // @[Top.scala 161:19]
  assign n197_I_2_0 = I0_2_0; // @[Top.scala 160:12]
  assign n197_I_2_1 = I0_2_1; // @[Top.scala 160:12]
  assign n197_I_2_2 = I0_2_2; // @[Top.scala 160:12]
  assign n200_valid_up = n197_valid_down; // @[Top.scala 164:19]
  assign n200_I_0_1 = n197_O_0_1; // @[Top.scala 163:12]
  assign n201_valid_up = n196_valid_down & n200_valid_down; // @[Top.scala 168:19]
  assign n201_I0_0_0 = n196_O_0_0; // @[Top.scala 166:13]
  assign n201_I1_0_0 = n200_O_0_0; // @[Top.scala 167:13]
  assign n212_valid_up = n201_valid_down; // @[Top.scala 171:19]
  assign n212_I_0_0_t0b = n201_O_0_0_t0b; // @[Top.scala 170:12]
  assign n212_I_0_0_t1b = n201_O_0_0_t1b; // @[Top.scala 170:12]
  assign n219_clock = clock;
  assign n219_reset = reset;
  assign n219_valid_up = n212_valid_down; // @[Top.scala 174:19]
  assign n219_I_0_0 = n212_O_0_0; // @[Top.scala 173:12]
  assign n224_valid_up = n219_valid_down; // @[Top.scala 177:19]
  assign n224_I_0_0_t0b = n219_O_0_0_t0b; // @[Top.scala 176:12]
  assign n224_I_0_0_t1b = n219_O_0_0_t1b; // @[Top.scala 176:12]
  assign n225_valid_up = n192_valid_down & n224_valid_down; // @[Top.scala 181:19]
  assign n225_I0_0_0 = n192_O_0_0; // @[Top.scala 179:13]
  assign n225_I1_0_0 = n224_O_0_0; // @[Top.scala 180:13]
  assign n232_valid_up = n189_valid_down & n225_valid_down; // @[Top.scala 185:19]
  assign n232_I0_0_0 = n189_O_0_0; // @[Top.scala 183:13]
  assign n232_I1_0_0_t0b = n225_O_0_0_t0b; // @[Top.scala 184:13]
  assign n232_I1_0_0_t1b = n225_O_0_0_t1b; // @[Top.scala 184:13]
  assign n352_clock = clock;
  assign n352_reset = reset;
  assign n352_valid_up = n232_valid_down; // @[Top.scala 188:19]
  assign n352_I_0_0_t0b = n232_O_0_0_t0b; // @[Top.scala 187:12]
  assign n352_I_0_0_t1b_t0b = n232_O_0_0_t1b_t0b; // @[Top.scala 187:12]
  assign n352_I_0_0_t1b_t1b = n232_O_0_0_t1b_t1b; // @[Top.scala 187:12]
  assign n344_clock = clock;
  assign n344_reset = reset;
  assign n344_valid_up = n192_valid_down; // @[Top.scala 191:19]
  assign n344_I_0_0 = n192_O_0_0; // @[Top.scala 190:12]
  assign n239_valid_up = n162_valid_down & n196_valid_down; // @[Top.scala 195:19]
  assign n239_I0_0_0 = n162_O_0_0; // @[Top.scala 193:13]
  assign n239_I1_0_0 = n196_O_0_0; // @[Top.scala 194:13]
  assign n246_valid_up = n239_valid_down & n165_valid_down; // @[Top.scala 199:19]
  assign n246_I0_0_0_0 = n239_O_0_0_0; // @[Top.scala 197:13]
  assign n246_I0_0_0_1 = n239_O_0_0_1; // @[Top.scala 197:13]
  assign n246_I1_0_0 = n165_O_0_0; // @[Top.scala 198:13]
  assign n253_valid_up = n246_valid_down & n200_valid_down; // @[Top.scala 203:19]
  assign n253_I0_0_0_0 = n246_O_0_0_0; // @[Top.scala 201:13]
  assign n253_I0_0_0_1 = n246_O_0_0_1; // @[Top.scala 201:13]
  assign n253_I0_0_0_2 = n246_O_0_0_2; // @[Top.scala 201:13]
  assign n253_I1_0_0 = n200_O_0_0; // @[Top.scala 202:13]
  assign n264_valid_up = n253_valid_down; // @[Top.scala 206:19]
  assign n264_I_0_0_0 = n253_O_0_0_0; // @[Top.scala 205:12]
  assign n264_I_0_0_1 = n253_O_0_0_1; // @[Top.scala 205:12]
  assign n264_I_0_0_2 = n253_O_0_0_2; // @[Top.scala 205:12]
  assign n264_I_0_0_3 = n253_O_0_0_3; // @[Top.scala 205:12]
  assign n269_clock = clock;
  assign n269_reset = reset;
  assign n269_valid_up = n264_valid_down; // @[Top.scala 209:19]
  assign n269_I_0_0 = n264_O_0_0; // @[Top.scala 208:12]
  assign n269_I_0_1 = n264_O_0_1; // @[Top.scala 208:12]
  assign n269_I_0_2 = n264_O_0_2; // @[Top.scala 208:12]
  assign n269_I_0_3 = n264_O_0_3; // @[Top.scala 208:12]
  assign n276_clock = clock;
  assign n276_reset = reset;
  assign n276_valid_up = n269_valid_down; // @[Top.scala 212:19]
  assign n276_I_0_0 = n269_O_0_0; // @[Top.scala 211:12]
  assign n281_valid_up = n276_valid_down; // @[Top.scala 215:19]
  assign n281_I_0_0_t0b = n276_O_0_0_t0b; // @[Top.scala 214:12]
  assign n281_I_0_0_t1b = n276_O_0_0_t1b; // @[Top.scala 214:12]
  assign n284_valid_up = n193_valid_down; // @[Top.scala 218:19]
  assign n284_I_0_0 = n193_O_0_0; // @[Top.scala 217:12]
  assign n287_valid_up = n193_valid_down; // @[Top.scala 221:19]
  assign n287_I_0_2 = n193_O_0_2; // @[Top.scala 220:12]
  assign n288_valid_up = n284_valid_down & n287_valid_down; // @[Top.scala 225:19]
  assign n288_I0_0_0 = n284_O_0_0; // @[Top.scala 223:13]
  assign n288_I1_0_0 = n287_O_0_0; // @[Top.scala 224:13]
  assign n297_valid_up = n197_valid_down; // @[Top.scala 228:19]
  assign n297_I_0_0 = n197_O_0_0; // @[Top.scala 227:12]
  assign n298_valid_up = n288_valid_down & n297_valid_down; // @[Top.scala 232:19]
  assign n298_I0_0_0_0 = n288_O_0_0_0; // @[Top.scala 230:13]
  assign n298_I0_0_0_1 = n288_O_0_0_1; // @[Top.scala 230:13]
  assign n298_I1_0_0 = n297_O_0_0; // @[Top.scala 231:13]
  assign n307_valid_up = n197_valid_down; // @[Top.scala 235:19]
  assign n307_I_0_2 = n197_O_0_2; // @[Top.scala 234:12]
  assign n308_valid_up = n298_valid_down & n307_valid_down; // @[Top.scala 239:19]
  assign n308_I0_0_0_0 = n298_O_0_0_0; // @[Top.scala 237:13]
  assign n308_I0_0_0_1 = n298_O_0_0_1; // @[Top.scala 237:13]
  assign n308_I0_0_0_2 = n298_O_0_0_2; // @[Top.scala 237:13]
  assign n308_I1_0_0 = n307_O_0_0; // @[Top.scala 238:13]
  assign n319_valid_up = n308_valid_down; // @[Top.scala 242:19]
  assign n319_I_0_0_0 = n308_O_0_0_0; // @[Top.scala 241:12]
  assign n319_I_0_0_1 = n308_O_0_0_1; // @[Top.scala 241:12]
  assign n319_I_0_0_2 = n308_O_0_0_2; // @[Top.scala 241:12]
  assign n319_I_0_0_3 = n308_O_0_0_3; // @[Top.scala 241:12]
  assign n324_clock = clock;
  assign n324_reset = reset;
  assign n324_valid_up = n319_valid_down; // @[Top.scala 245:19]
  assign n324_I_0_0 = n319_O_0_0; // @[Top.scala 244:12]
  assign n324_I_0_1 = n319_O_0_1; // @[Top.scala 244:12]
  assign n324_I_0_2 = n319_O_0_2; // @[Top.scala 244:12]
  assign n324_I_0_3 = n319_O_0_3; // @[Top.scala 244:12]
  assign n331_clock = clock;
  assign n331_reset = reset;
  assign n331_valid_up = n324_valid_down; // @[Top.scala 248:19]
  assign n331_I_0_0 = n324_O_0_0; // @[Top.scala 247:12]
  assign n336_valid_up = n331_valid_down; // @[Top.scala 251:19]
  assign n336_I_0_0_t0b = n331_O_0_0_t0b; // @[Top.scala 250:12]
  assign n336_I_0_0_t1b = n331_O_0_0_t1b; // @[Top.scala 250:12]
  assign n337_valid_up = n281_valid_down & n336_valid_down; // @[Top.scala 255:19]
  assign n337_I0_0_0 = n281_O_0_0; // @[Top.scala 253:13]
  assign n337_I1_0_0 = n336_O_0_0; // @[Top.scala 254:13]
  assign n345_valid_up = n344_valid_down & n337_valid_down; // @[Top.scala 259:19]
  assign n345_I0_0_0 = n344_O_0_0; // @[Top.scala 257:13]
  assign n345_I1_0_0_t0b = n337_O_0_0_t0b; // @[Top.scala 258:13]
  assign n345_I1_0_0_t1b = n337_O_0_0_t1b; // @[Top.scala 258:13]
  assign n353_valid_up = n352_valid_down & n345_valid_down; // @[Top.scala 263:19]
  assign n353_I0_0_0_t0b = n352_O_0_0_t0b; // @[Top.scala 261:13]
  assign n353_I0_0_0_t1b_t0b = n352_O_0_0_t1b_t0b; // @[Top.scala 261:13]
  assign n353_I0_0_0_t1b_t1b = n352_O_0_0_t1b_t1b; // @[Top.scala 261:13]
  assign n353_I1_0_0_t0b = n345_O_0_0_t0b; // @[Top.scala 262:13]
  assign n353_I1_0_0_t1b_t0b = n345_O_0_0_t1b_t0b; // @[Top.scala 262:13]
  assign n353_I1_0_0_t1b_t1b = n345_O_0_0_t1b_t1b; // @[Top.scala 262:13]
  assign n361_valid_up = n360_valid_down & n353_valid_down; // @[Top.scala 267:19]
  assign n361_I0_0_0 = n360_O_0_0; // @[Top.scala 265:13]
  assign n361_I1_0_0_t0b_t0b = n353_O_0_0_t0b_t0b; // @[Top.scala 266:13]
  assign n361_I1_0_0_t0b_t1b_t0b = n353_O_0_0_t0b_t1b_t0b; // @[Top.scala 266:13]
  assign n361_I1_0_0_t0b_t1b_t1b = n353_O_0_0_t0b_t1b_t1b; // @[Top.scala 266:13]
  assign n361_I1_0_0_t1b_t0b = n353_O_0_0_t1b_t0b; // @[Top.scala 266:13]
  assign n361_I1_0_0_t1b_t1b_t0b = n353_O_0_0_t1b_t1b_t0b; // @[Top.scala 266:13]
  assign n361_I1_0_0_t1b_t1b_t1b = n353_O_0_0_t1b_t1b_t1b; // @[Top.scala 266:13]
  assign n372_valid_up = n361_valid_down; // @[Top.scala 270:19]
  assign n372_I_0_0_t0b = n361_O_0_0_t0b; // @[Top.scala 269:12]
  assign n372_I_0_0_t1b_t0b_t0b = n361_O_0_0_t1b_t0b_t0b; // @[Top.scala 269:12]
  assign n372_I_0_0_t1b_t0b_t1b_t0b = n361_O_0_0_t1b_t0b_t1b_t0b; // @[Top.scala 269:12]
  assign n372_I_0_0_t1b_t0b_t1b_t1b = n361_O_0_0_t1b_t0b_t1b_t1b; // @[Top.scala 269:12]
  assign n372_I_0_0_t1b_t1b_t0b = n361_O_0_0_t1b_t1b_t0b; // @[Top.scala 269:12]
  assign n372_I_0_0_t1b_t1b_t1b_t0b = n361_O_0_0_t1b_t1b_t1b_t0b; // @[Top.scala 269:12]
  assign n372_I_0_0_t1b_t1b_t1b_t1b = n361_O_0_0_t1b_t1b_t1b_t1b; // @[Top.scala 269:12]
  assign n410_clock = clock;
  assign n410_reset = reset;
  assign n410_valid_up = n157_valid_down; // @[Top.scala 273:19]
  assign n410_I_0_0 = n157_O_0_0; // @[Top.scala 272:12]
  assign n373_clock = clock;
  assign n373_reset = reset;
  assign n373_valid_up = n192_valid_down; // @[Top.scala 276:19]
  assign n373_I_0_0 = n192_O_0_0; // @[Top.scala 275:12]
  assign n374_valid_up = n281_valid_down & n373_valid_down; // @[Top.scala 280:19]
  assign n374_I0_0_0 = n281_O_0_0; // @[Top.scala 278:13]
  assign n374_I1_0_0 = n373_O_0_0; // @[Top.scala 279:13]
  assign n381_valid_up = n336_valid_down & n374_valid_down; // @[Top.scala 284:19]
  assign n381_I0_0_0 = n336_O_0_0; // @[Top.scala 282:13]
  assign n381_I1_0_0_t0b = n374_O_0_0_t0b; // @[Top.scala 283:13]
  assign n381_I1_0_0_t1b = n374_O_0_0_t1b; // @[Top.scala 283:13]
  assign n388_valid_up = n192_valid_down & n189_valid_down; // @[Top.scala 288:19]
  assign n388_I0_0_0 = n192_O_0_0; // @[Top.scala 286:13]
  assign n388_I1_0_0 = n189_O_0_0; // @[Top.scala 287:13]
  assign n395_valid_up = n224_valid_down & n388_valid_down; // @[Top.scala 292:19]
  assign n395_I0_0_0 = n224_O_0_0; // @[Top.scala 290:13]
  assign n395_I1_0_0_t0b = n388_O_0_0_t0b; // @[Top.scala 291:13]
  assign n395_I1_0_0_t1b = n388_O_0_0_t1b; // @[Top.scala 291:13]
  assign n402_clock = clock;
  assign n402_reset = reset;
  assign n402_valid_up = n395_valid_down; // @[Top.scala 295:19]
  assign n402_I_0_0_t0b = n395_O_0_0_t0b; // @[Top.scala 294:12]
  assign n402_I_0_0_t1b_t0b = n395_O_0_0_t1b_t0b; // @[Top.scala 294:12]
  assign n402_I_0_0_t1b_t1b = n395_O_0_0_t1b_t1b; // @[Top.scala 294:12]
  assign n403_valid_up = n381_valid_down & n402_valid_down; // @[Top.scala 299:19]
  assign n403_I0_0_0_t0b = n381_O_0_0_t0b; // @[Top.scala 297:13]
  assign n403_I0_0_0_t1b_t0b = n381_O_0_0_t1b_t0b; // @[Top.scala 297:13]
  assign n403_I0_0_0_t1b_t1b = n381_O_0_0_t1b_t1b; // @[Top.scala 297:13]
  assign n403_I1_0_0_t0b = n402_O_0_0_t0b; // @[Top.scala 298:13]
  assign n403_I1_0_0_t1b_t0b = n402_O_0_0_t1b_t0b; // @[Top.scala 298:13]
  assign n403_I1_0_0_t1b_t1b = n402_O_0_0_t1b_t1b; // @[Top.scala 298:13]
  assign n411_valid_up = n410_valid_down & n403_valid_down; // @[Top.scala 303:19]
  assign n411_I0_0_0 = n410_O_0_0; // @[Top.scala 301:13]
  assign n411_I1_0_0_t0b_t0b = n403_O_0_0_t0b_t0b; // @[Top.scala 302:13]
  assign n411_I1_0_0_t0b_t1b_t0b = n403_O_0_0_t0b_t1b_t0b; // @[Top.scala 302:13]
  assign n411_I1_0_0_t0b_t1b_t1b = n403_O_0_0_t0b_t1b_t1b; // @[Top.scala 302:13]
  assign n411_I1_0_0_t1b_t0b = n403_O_0_0_t1b_t0b; // @[Top.scala 302:13]
  assign n411_I1_0_0_t1b_t1b_t0b = n403_O_0_0_t1b_t1b_t0b; // @[Top.scala 302:13]
  assign n411_I1_0_0_t1b_t1b_t1b = n403_O_0_0_t1b_t1b_t1b; // @[Top.scala 302:13]
  assign n422_valid_up = n411_valid_down; // @[Top.scala 306:19]
  assign n422_I_0_0_t0b = n411_O_0_0_t0b; // @[Top.scala 305:12]
  assign n422_I_0_0_t1b_t0b_t0b = n411_O_0_0_t1b_t0b_t0b; // @[Top.scala 305:12]
  assign n422_I_0_0_t1b_t0b_t1b_t0b = n411_O_0_0_t1b_t0b_t1b_t0b; // @[Top.scala 305:12]
  assign n422_I_0_0_t1b_t0b_t1b_t1b = n411_O_0_0_t1b_t0b_t1b_t1b; // @[Top.scala 305:12]
  assign n422_I_0_0_t1b_t1b_t0b = n411_O_0_0_t1b_t1b_t0b; // @[Top.scala 305:12]
  assign n422_I_0_0_t1b_t1b_t1b_t0b = n411_O_0_0_t1b_t1b_t1b_t0b; // @[Top.scala 305:12]
  assign n422_I_0_0_t1b_t1b_t1b_t1b = n411_O_0_0_t1b_t1b_t1b_t1b; // @[Top.scala 305:12]
  assign n423_valid_up = n372_valid_down & n422_valid_down; // @[Top.scala 310:19]
  assign n423_I0_0_0_t0b = n372_O_0_0_t0b; // @[Top.scala 308:13]
  assign n423_I0_0_0_t1b_t0b = n372_O_0_0_t1b_t0b; // @[Top.scala 308:13]
  assign n423_I0_0_0_t1b_t1b = n372_O_0_0_t1b_t1b; // @[Top.scala 308:13]
  assign n423_I1_0_0_t0b = n422_O_0_0_t0b; // @[Top.scala 309:13]
  assign n423_I1_0_0_t1b_t0b = n422_O_0_0_t1b_t0b; // @[Top.scala 309:13]
  assign n423_I1_0_0_t1b_t1b = n422_O_0_0_t1b_t1b; // @[Top.scala 309:13]
  assign n431_valid_up = n430_valid_down & n423_valid_down; // @[Top.scala 314:19]
  assign n431_I0_0_0 = n430_O_0_0; // @[Top.scala 312:13]
  assign n431_I1_0_0_t0b_t0b = n423_O_0_0_t0b_t0b; // @[Top.scala 313:13]
  assign n431_I1_0_0_t0b_t1b_t0b = n423_O_0_0_t0b_t1b_t0b; // @[Top.scala 313:13]
  assign n431_I1_0_0_t0b_t1b_t1b = n423_O_0_0_t0b_t1b_t1b; // @[Top.scala 313:13]
  assign n431_I1_0_0_t1b_t0b = n423_O_0_0_t1b_t0b; // @[Top.scala 313:13]
  assign n431_I1_0_0_t1b_t1b_t0b = n423_O_0_0_t1b_t1b_t0b; // @[Top.scala 313:13]
  assign n431_I1_0_0_t1b_t1b_t1b = n423_O_0_0_t1b_t1b_t1b; // @[Top.scala 313:13]
  assign n442_valid_up = n431_valid_down; // @[Top.scala 317:19]
  assign n442_I_0_0_t0b = n431_O_0_0_t0b; // @[Top.scala 316:12]
  assign n442_I_0_0_t1b_t0b_t0b = n431_O_0_0_t1b_t0b_t0b; // @[Top.scala 316:12]
  assign n442_I_0_0_t1b_t0b_t1b_t0b = n431_O_0_0_t1b_t0b_t1b_t0b; // @[Top.scala 316:12]
  assign n442_I_0_0_t1b_t0b_t1b_t1b = n431_O_0_0_t1b_t0b_t1b_t1b; // @[Top.scala 316:12]
  assign n442_I_0_0_t1b_t1b_t0b = n431_O_0_0_t1b_t1b_t0b; // @[Top.scala 316:12]
  assign n442_I_0_0_t1b_t1b_t1b_t0b = n431_O_0_0_t1b_t1b_t1b_t0b; // @[Top.scala 316:12]
  assign n442_I_0_0_t1b_t1b_t1b_t1b = n431_O_0_0_t1b_t1b_t1b_t1b; // @[Top.scala 316:12]
endmodule
module Map2S_53(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0_0_0,
  input  [31:0] I0_0_0_1,
  input  [31:0] I0_0_0_2,
  input  [31:0] I0_0_1_0,
  input  [31:0] I0_0_1_1,
  input  [31:0] I0_0_1_2,
  input  [31:0] I0_0_2_0,
  input  [31:0] I0_0_2_1,
  input  [31:0] I0_0_2_2,
  input  [31:0] I0_1_0_0,
  input  [31:0] I0_1_0_1,
  input  [31:0] I0_1_0_2,
  input  [31:0] I0_1_1_0,
  input  [31:0] I0_1_1_1,
  input  [31:0] I0_1_1_2,
  input  [31:0] I0_1_2_0,
  input  [31:0] I0_1_2_1,
  input  [31:0] I0_1_2_2,
  input  [31:0] I0_2_0_0,
  input  [31:0] I0_2_0_1,
  input  [31:0] I0_2_0_2,
  input  [31:0] I0_2_1_0,
  input  [31:0] I0_2_1_1,
  input  [31:0] I0_2_1_2,
  input  [31:0] I0_2_2_0,
  input  [31:0] I0_2_2_1,
  input  [31:0] I0_2_2_2,
  input  [31:0] I0_3_0_0,
  input  [31:0] I0_3_0_1,
  input  [31:0] I0_3_0_2,
  input  [31:0] I0_3_1_0,
  input  [31:0] I0_3_1_1,
  input  [31:0] I0_3_1_2,
  input  [31:0] I0_3_2_0,
  input  [31:0] I0_3_2_1,
  input  [31:0] I0_3_2_2,
  input  [31:0] I0_4_0_0,
  input  [31:0] I0_4_0_1,
  input  [31:0] I0_4_0_2,
  input  [31:0] I0_4_1_0,
  input  [31:0] I0_4_1_1,
  input  [31:0] I0_4_1_2,
  input  [31:0] I0_4_2_0,
  input  [31:0] I0_4_2_1,
  input  [31:0] I0_4_2_2,
  input  [31:0] I0_5_0_0,
  input  [31:0] I0_5_0_1,
  input  [31:0] I0_5_0_2,
  input  [31:0] I0_5_1_0,
  input  [31:0] I0_5_1_1,
  input  [31:0] I0_5_1_2,
  input  [31:0] I0_5_2_0,
  input  [31:0] I0_5_2_1,
  input  [31:0] I0_5_2_2,
  input  [31:0] I0_6_0_0,
  input  [31:0] I0_6_0_1,
  input  [31:0] I0_6_0_2,
  input  [31:0] I0_6_1_0,
  input  [31:0] I0_6_1_1,
  input  [31:0] I0_6_1_2,
  input  [31:0] I0_6_2_0,
  input  [31:0] I0_6_2_1,
  input  [31:0] I0_6_2_2,
  input  [31:0] I0_7_0_0,
  input  [31:0] I0_7_0_1,
  input  [31:0] I0_7_0_2,
  input  [31:0] I0_7_1_0,
  input  [31:0] I0_7_1_1,
  input  [31:0] I0_7_1_2,
  input  [31:0] I0_7_2_0,
  input  [31:0] I0_7_2_1,
  input  [31:0] I0_7_2_2,
  input         I1_0_0_0_t0b,
  input         I1_0_0_0_t1b,
  input         I1_1_0_0_t0b,
  input         I1_1_0_0_t1b,
  input         I1_2_0_0_t0b,
  input         I1_2_0_0_t1b,
  input         I1_3_0_0_t0b,
  input         I1_3_0_0_t1b,
  input         I1_4_0_0_t0b,
  input         I1_4_0_0_t1b,
  input         I1_5_0_0_t0b,
  input         I1_5_0_0_t1b,
  input         I1_6_0_0_t0b,
  input         I1_6_0_0_t1b,
  input         I1_7_0_0_t0b,
  input         I1_7_0_0_t1b,
  output [31:0] O_0_0_0_t0b,
  output [31:0] O_0_0_0_t1b_t0b,
  output [31:0] O_0_0_0_t1b_t1b,
  output [31:0] O_1_0_0_t0b,
  output [31:0] O_1_0_0_t1b_t0b,
  output [31:0] O_1_0_0_t1b_t1b,
  output [31:0] O_2_0_0_t0b,
  output [31:0] O_2_0_0_t1b_t0b,
  output [31:0] O_2_0_0_t1b_t1b,
  output [31:0] O_3_0_0_t0b,
  output [31:0] O_3_0_0_t1b_t0b,
  output [31:0] O_3_0_0_t1b_t1b,
  output [31:0] O_4_0_0_t0b,
  output [31:0] O_4_0_0_t1b_t0b,
  output [31:0] O_4_0_0_t1b_t1b,
  output [31:0] O_5_0_0_t0b,
  output [31:0] O_5_0_0_t1b_t0b,
  output [31:0] O_5_0_0_t1b_t1b,
  output [31:0] O_6_0_0_t0b,
  output [31:0] O_6_0_0_t1b_t0b,
  output [31:0] O_6_0_0_t1b_t1b,
  output [31:0] O_7_0_0_t0b,
  output [31:0] O_7_0_0_t1b_t0b,
  output [31:0] O_7_0_0_t1b_t1b
);
  wire  fst_op_clock; // @[Map2S.scala 9:22]
  wire  fst_op_reset; // @[Map2S.scala 9:22]
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0_2; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_1_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_1_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_1_2; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_2_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_2_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_2_2; // @[Map2S.scala 9:22]
  wire  fst_op_I1_0_0_t0b; // @[Map2S.scala 9:22]
  wire  fst_op_I1_0_0_t1b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_0_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_0_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_0_t1b_t1b; // @[Map2S.scala 9:22]
  wire  other_ops_0_clock; // @[Map2S.scala 10:86]
  wire  other_ops_0_reset; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_0_I1_0_0_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_0_I1_0_0_t1b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_0_0_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_0_0_t1b_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_0_0_t1b_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_1_clock; // @[Map2S.scala 10:86]
  wire  other_ops_1_reset; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_1_I1_0_0_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_1_I1_0_0_t1b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_0_0_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_0_0_t1b_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_0_0_t1b_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_2_clock; // @[Map2S.scala 10:86]
  wire  other_ops_2_reset; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_2_I1_0_0_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_2_I1_0_0_t1b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_0_0_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_0_0_t1b_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_0_0_t1b_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_3_clock; // @[Map2S.scala 10:86]
  wire  other_ops_3_reset; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_3_I1_0_0_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_3_I1_0_0_t1b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_0_0_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_0_0_t1b_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_0_0_t1b_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_4_clock; // @[Map2S.scala 10:86]
  wire  other_ops_4_reset; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_4_I1_0_0_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_4_I1_0_0_t1b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_0_0_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_0_0_t1b_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_0_0_t1b_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_5_clock; // @[Map2S.scala 10:86]
  wire  other_ops_5_reset; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_5_I1_0_0_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_5_I1_0_0_t1b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_0_0_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_0_0_t1b_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_0_0_t1b_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_6_clock; // @[Map2S.scala 10:86]
  wire  other_ops_6_reset; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_6_I1_0_0_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_6_I1_0_0_t1b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_0_0_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_0_0_t1b_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_0_0_t1b_t1b; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  wire  _T_2; // @[Map2S.scala 26:83]
  wire  _T_3; // @[Map2S.scala 26:83]
  wire  _T_4; // @[Map2S.scala 26:83]
  wire  _T_5; // @[Map2S.scala 26:83]
  Module_6 fst_op ( // @[Map2S.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0_0(fst_op_I0_0_0),
    .I0_0_1(fst_op_I0_0_1),
    .I0_0_2(fst_op_I0_0_2),
    .I0_1_0(fst_op_I0_1_0),
    .I0_1_1(fst_op_I0_1_1),
    .I0_1_2(fst_op_I0_1_2),
    .I0_2_0(fst_op_I0_2_0),
    .I0_2_1(fst_op_I0_2_1),
    .I0_2_2(fst_op_I0_2_2),
    .I1_0_0_t0b(fst_op_I1_0_0_t0b),
    .I1_0_0_t1b(fst_op_I1_0_0_t1b),
    .O_0_0_t0b(fst_op_O_0_0_t0b),
    .O_0_0_t1b_t0b(fst_op_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(fst_op_O_0_0_t1b_t1b)
  );
  Module_6 other_ops_0 ( // @[Map2S.scala 10:86]
    .clock(other_ops_0_clock),
    .reset(other_ops_0_reset),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0_0(other_ops_0_I0_0_0),
    .I0_0_1(other_ops_0_I0_0_1),
    .I0_0_2(other_ops_0_I0_0_2),
    .I0_1_0(other_ops_0_I0_1_0),
    .I0_1_1(other_ops_0_I0_1_1),
    .I0_1_2(other_ops_0_I0_1_2),
    .I0_2_0(other_ops_0_I0_2_0),
    .I0_2_1(other_ops_0_I0_2_1),
    .I0_2_2(other_ops_0_I0_2_2),
    .I1_0_0_t0b(other_ops_0_I1_0_0_t0b),
    .I1_0_0_t1b(other_ops_0_I1_0_0_t1b),
    .O_0_0_t0b(other_ops_0_O_0_0_t0b),
    .O_0_0_t1b_t0b(other_ops_0_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(other_ops_0_O_0_0_t1b_t1b)
  );
  Module_6 other_ops_1 ( // @[Map2S.scala 10:86]
    .clock(other_ops_1_clock),
    .reset(other_ops_1_reset),
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0_0_0(other_ops_1_I0_0_0),
    .I0_0_1(other_ops_1_I0_0_1),
    .I0_0_2(other_ops_1_I0_0_2),
    .I0_1_0(other_ops_1_I0_1_0),
    .I0_1_1(other_ops_1_I0_1_1),
    .I0_1_2(other_ops_1_I0_1_2),
    .I0_2_0(other_ops_1_I0_2_0),
    .I0_2_1(other_ops_1_I0_2_1),
    .I0_2_2(other_ops_1_I0_2_2),
    .I1_0_0_t0b(other_ops_1_I1_0_0_t0b),
    .I1_0_0_t1b(other_ops_1_I1_0_0_t1b),
    .O_0_0_t0b(other_ops_1_O_0_0_t0b),
    .O_0_0_t1b_t0b(other_ops_1_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(other_ops_1_O_0_0_t1b_t1b)
  );
  Module_6 other_ops_2 ( // @[Map2S.scala 10:86]
    .clock(other_ops_2_clock),
    .reset(other_ops_2_reset),
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0_0_0(other_ops_2_I0_0_0),
    .I0_0_1(other_ops_2_I0_0_1),
    .I0_0_2(other_ops_2_I0_0_2),
    .I0_1_0(other_ops_2_I0_1_0),
    .I0_1_1(other_ops_2_I0_1_1),
    .I0_1_2(other_ops_2_I0_1_2),
    .I0_2_0(other_ops_2_I0_2_0),
    .I0_2_1(other_ops_2_I0_2_1),
    .I0_2_2(other_ops_2_I0_2_2),
    .I1_0_0_t0b(other_ops_2_I1_0_0_t0b),
    .I1_0_0_t1b(other_ops_2_I1_0_0_t1b),
    .O_0_0_t0b(other_ops_2_O_0_0_t0b),
    .O_0_0_t1b_t0b(other_ops_2_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(other_ops_2_O_0_0_t1b_t1b)
  );
  Module_6 other_ops_3 ( // @[Map2S.scala 10:86]
    .clock(other_ops_3_clock),
    .reset(other_ops_3_reset),
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I0_0_0(other_ops_3_I0_0_0),
    .I0_0_1(other_ops_3_I0_0_1),
    .I0_0_2(other_ops_3_I0_0_2),
    .I0_1_0(other_ops_3_I0_1_0),
    .I0_1_1(other_ops_3_I0_1_1),
    .I0_1_2(other_ops_3_I0_1_2),
    .I0_2_0(other_ops_3_I0_2_0),
    .I0_2_1(other_ops_3_I0_2_1),
    .I0_2_2(other_ops_3_I0_2_2),
    .I1_0_0_t0b(other_ops_3_I1_0_0_t0b),
    .I1_0_0_t1b(other_ops_3_I1_0_0_t1b),
    .O_0_0_t0b(other_ops_3_O_0_0_t0b),
    .O_0_0_t1b_t0b(other_ops_3_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(other_ops_3_O_0_0_t1b_t1b)
  );
  Module_6 other_ops_4 ( // @[Map2S.scala 10:86]
    .clock(other_ops_4_clock),
    .reset(other_ops_4_reset),
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I0_0_0(other_ops_4_I0_0_0),
    .I0_0_1(other_ops_4_I0_0_1),
    .I0_0_2(other_ops_4_I0_0_2),
    .I0_1_0(other_ops_4_I0_1_0),
    .I0_1_1(other_ops_4_I0_1_1),
    .I0_1_2(other_ops_4_I0_1_2),
    .I0_2_0(other_ops_4_I0_2_0),
    .I0_2_1(other_ops_4_I0_2_1),
    .I0_2_2(other_ops_4_I0_2_2),
    .I1_0_0_t0b(other_ops_4_I1_0_0_t0b),
    .I1_0_0_t1b(other_ops_4_I1_0_0_t1b),
    .O_0_0_t0b(other_ops_4_O_0_0_t0b),
    .O_0_0_t1b_t0b(other_ops_4_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(other_ops_4_O_0_0_t1b_t1b)
  );
  Module_6 other_ops_5 ( // @[Map2S.scala 10:86]
    .clock(other_ops_5_clock),
    .reset(other_ops_5_reset),
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I0_0_0(other_ops_5_I0_0_0),
    .I0_0_1(other_ops_5_I0_0_1),
    .I0_0_2(other_ops_5_I0_0_2),
    .I0_1_0(other_ops_5_I0_1_0),
    .I0_1_1(other_ops_5_I0_1_1),
    .I0_1_2(other_ops_5_I0_1_2),
    .I0_2_0(other_ops_5_I0_2_0),
    .I0_2_1(other_ops_5_I0_2_1),
    .I0_2_2(other_ops_5_I0_2_2),
    .I1_0_0_t0b(other_ops_5_I1_0_0_t0b),
    .I1_0_0_t1b(other_ops_5_I1_0_0_t1b),
    .O_0_0_t0b(other_ops_5_O_0_0_t0b),
    .O_0_0_t1b_t0b(other_ops_5_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(other_ops_5_O_0_0_t1b_t1b)
  );
  Module_6 other_ops_6 ( // @[Map2S.scala 10:86]
    .clock(other_ops_6_clock),
    .reset(other_ops_6_reset),
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I0_0_0(other_ops_6_I0_0_0),
    .I0_0_1(other_ops_6_I0_0_1),
    .I0_0_2(other_ops_6_I0_0_2),
    .I0_1_0(other_ops_6_I0_1_0),
    .I0_1_1(other_ops_6_I0_1_1),
    .I0_1_2(other_ops_6_I0_1_2),
    .I0_2_0(other_ops_6_I0_2_0),
    .I0_2_1(other_ops_6_I0_2_1),
    .I0_2_2(other_ops_6_I0_2_2),
    .I1_0_0_t0b(other_ops_6_I1_0_0_t0b),
    .I1_0_0_t1b(other_ops_6_I1_0_0_t1b),
    .O_0_0_t0b(other_ops_6_O_0_0_t0b),
    .O_0_0_t1b_t0b(other_ops_6_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(other_ops_6_O_0_0_t1b_t1b)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[Map2S.scala 26:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[Map2S.scala 26:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_5 & other_ops_6_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_0_t0b = fst_op_O_0_0_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_0_t1b_t0b = fst_op_O_0_0_t1b_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_0_t1b_t1b = fst_op_O_0_0_t1b_t1b; // @[Map2S.scala 19:8]
  assign O_1_0_0_t0b = other_ops_0_O_0_0_t0b; // @[Map2S.scala 24:12]
  assign O_1_0_0_t1b_t0b = other_ops_0_O_0_0_t1b_t0b; // @[Map2S.scala 24:12]
  assign O_1_0_0_t1b_t1b = other_ops_0_O_0_0_t1b_t1b; // @[Map2S.scala 24:12]
  assign O_2_0_0_t0b = other_ops_1_O_0_0_t0b; // @[Map2S.scala 24:12]
  assign O_2_0_0_t1b_t0b = other_ops_1_O_0_0_t1b_t0b; // @[Map2S.scala 24:12]
  assign O_2_0_0_t1b_t1b = other_ops_1_O_0_0_t1b_t1b; // @[Map2S.scala 24:12]
  assign O_3_0_0_t0b = other_ops_2_O_0_0_t0b; // @[Map2S.scala 24:12]
  assign O_3_0_0_t1b_t0b = other_ops_2_O_0_0_t1b_t0b; // @[Map2S.scala 24:12]
  assign O_3_0_0_t1b_t1b = other_ops_2_O_0_0_t1b_t1b; // @[Map2S.scala 24:12]
  assign O_4_0_0_t0b = other_ops_3_O_0_0_t0b; // @[Map2S.scala 24:12]
  assign O_4_0_0_t1b_t0b = other_ops_3_O_0_0_t1b_t0b; // @[Map2S.scala 24:12]
  assign O_4_0_0_t1b_t1b = other_ops_3_O_0_0_t1b_t1b; // @[Map2S.scala 24:12]
  assign O_5_0_0_t0b = other_ops_4_O_0_0_t0b; // @[Map2S.scala 24:12]
  assign O_5_0_0_t1b_t0b = other_ops_4_O_0_0_t1b_t0b; // @[Map2S.scala 24:12]
  assign O_5_0_0_t1b_t1b = other_ops_4_O_0_0_t1b_t1b; // @[Map2S.scala 24:12]
  assign O_6_0_0_t0b = other_ops_5_O_0_0_t0b; // @[Map2S.scala 24:12]
  assign O_6_0_0_t1b_t0b = other_ops_5_O_0_0_t1b_t0b; // @[Map2S.scala 24:12]
  assign O_6_0_0_t1b_t1b = other_ops_5_O_0_0_t1b_t1b; // @[Map2S.scala 24:12]
  assign O_7_0_0_t0b = other_ops_6_O_0_0_t0b; // @[Map2S.scala 24:12]
  assign O_7_0_0_t1b_t0b = other_ops_6_O_0_0_t1b_t0b; // @[Map2S.scala 24:12]
  assign O_7_0_0_t1b_t1b = other_ops_6_O_0_0_t1b_t1b; // @[Map2S.scala 24:12]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0_0 = I0_0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_1 = I0_0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_2 = I0_0_0_2; // @[Map2S.scala 17:13]
  assign fst_op_I0_1_0 = I0_0_1_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1_1 = I0_0_1_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_1_2 = I0_0_1_2; // @[Map2S.scala 17:13]
  assign fst_op_I0_2_0 = I0_0_2_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_2_1 = I0_0_2_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_2_2 = I0_0_2_2; // @[Map2S.scala 17:13]
  assign fst_op_I1_0_0_t0b = I1_0_0_0_t0b; // @[Map2S.scala 18:13]
  assign fst_op_I1_0_0_t1b = I1_0_0_0_t1b; // @[Map2S.scala 18:13]
  assign other_ops_0_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_0_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0_0 = I0_1_0_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_0_1 = I0_1_0_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_0_2 = I0_1_0_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1_0 = I0_1_1_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1_1 = I0_1_1_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1_2 = I0_1_1_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_2_0 = I0_1_2_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_2_1 = I0_1_2_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_2_2 = I0_1_2_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I1_0_0_t0b = I1_1_0_0_t0b; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_0_0_t1b = I1_1_0_0_t1b; // @[Map2S.scala 23:43]
  assign other_ops_1_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_1_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0_0_0 = I0_2_0_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_0_1 = I0_2_0_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_0_2 = I0_2_0_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1_0 = I0_2_1_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1_1 = I0_2_1_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1_2 = I0_2_1_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_2_0 = I0_2_2_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_2_1 = I0_2_2_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_2_2 = I0_2_2_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1_0_0_t0b = I1_2_0_0_t0b; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_0_0_t1b = I1_2_0_0_t1b; // @[Map2S.scala 23:43]
  assign other_ops_2_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_2_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0_0_0 = I0_3_0_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_0_1 = I0_3_0_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_0_2 = I0_3_0_2; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_1_0 = I0_3_1_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_1_1 = I0_3_1_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_1_2 = I0_3_1_2; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_2_0 = I0_3_2_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_2_1 = I0_3_2_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_2_2 = I0_3_2_2; // @[Map2S.scala 22:43]
  assign other_ops_2_I1_0_0_t0b = I1_3_0_0_t0b; // @[Map2S.scala 23:43]
  assign other_ops_2_I1_0_0_t1b = I1_3_0_0_t1b; // @[Map2S.scala 23:43]
  assign other_ops_3_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_3_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_3_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_3_I0_0_0 = I0_4_0_0; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_0_1 = I0_4_0_1; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_0_2 = I0_4_0_2; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_1_0 = I0_4_1_0; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_1_1 = I0_4_1_1; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_1_2 = I0_4_1_2; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_2_0 = I0_4_2_0; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_2_1 = I0_4_2_1; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_2_2 = I0_4_2_2; // @[Map2S.scala 22:43]
  assign other_ops_3_I1_0_0_t0b = I1_4_0_0_t0b; // @[Map2S.scala 23:43]
  assign other_ops_3_I1_0_0_t1b = I1_4_0_0_t1b; // @[Map2S.scala 23:43]
  assign other_ops_4_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_4_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_4_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_4_I0_0_0 = I0_5_0_0; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_0_1 = I0_5_0_1; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_0_2 = I0_5_0_2; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_1_0 = I0_5_1_0; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_1_1 = I0_5_1_1; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_1_2 = I0_5_1_2; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_2_0 = I0_5_2_0; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_2_1 = I0_5_2_1; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_2_2 = I0_5_2_2; // @[Map2S.scala 22:43]
  assign other_ops_4_I1_0_0_t0b = I1_5_0_0_t0b; // @[Map2S.scala 23:43]
  assign other_ops_4_I1_0_0_t1b = I1_5_0_0_t1b; // @[Map2S.scala 23:43]
  assign other_ops_5_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_5_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_5_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_5_I0_0_0 = I0_6_0_0; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_0_1 = I0_6_0_1; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_0_2 = I0_6_0_2; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_1_0 = I0_6_1_0; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_1_1 = I0_6_1_1; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_1_2 = I0_6_1_2; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_2_0 = I0_6_2_0; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_2_1 = I0_6_2_1; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_2_2 = I0_6_2_2; // @[Map2S.scala 22:43]
  assign other_ops_5_I1_0_0_t0b = I1_6_0_0_t0b; // @[Map2S.scala 23:43]
  assign other_ops_5_I1_0_0_t1b = I1_6_0_0_t1b; // @[Map2S.scala 23:43]
  assign other_ops_6_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_6_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_6_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_6_I0_0_0 = I0_7_0_0; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_0_1 = I0_7_0_1; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_0_2 = I0_7_0_2; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_1_0 = I0_7_1_0; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_1_1 = I0_7_1_1; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_1_2 = I0_7_1_2; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_2_0 = I0_7_2_0; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_2_1 = I0_7_2_1; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_2_2 = I0_7_2_2; // @[Map2S.scala 22:43]
  assign other_ops_6_I1_0_0_t0b = I1_7_0_0_t0b; // @[Map2S.scala 23:43]
  assign other_ops_6_I1_0_0_t1b = I1_7_0_0_t1b; // @[Map2S.scala 23:43]
endmodule
module Map2T_9(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0_0_0,
  input  [31:0] I0_0_0_1,
  input  [31:0] I0_0_0_2,
  input  [31:0] I0_0_1_0,
  input  [31:0] I0_0_1_1,
  input  [31:0] I0_0_1_2,
  input  [31:0] I0_0_2_0,
  input  [31:0] I0_0_2_1,
  input  [31:0] I0_0_2_2,
  input  [31:0] I0_1_0_0,
  input  [31:0] I0_1_0_1,
  input  [31:0] I0_1_0_2,
  input  [31:0] I0_1_1_0,
  input  [31:0] I0_1_1_1,
  input  [31:0] I0_1_1_2,
  input  [31:0] I0_1_2_0,
  input  [31:0] I0_1_2_1,
  input  [31:0] I0_1_2_2,
  input  [31:0] I0_2_0_0,
  input  [31:0] I0_2_0_1,
  input  [31:0] I0_2_0_2,
  input  [31:0] I0_2_1_0,
  input  [31:0] I0_2_1_1,
  input  [31:0] I0_2_1_2,
  input  [31:0] I0_2_2_0,
  input  [31:0] I0_2_2_1,
  input  [31:0] I0_2_2_2,
  input  [31:0] I0_3_0_0,
  input  [31:0] I0_3_0_1,
  input  [31:0] I0_3_0_2,
  input  [31:0] I0_3_1_0,
  input  [31:0] I0_3_1_1,
  input  [31:0] I0_3_1_2,
  input  [31:0] I0_3_2_0,
  input  [31:0] I0_3_2_1,
  input  [31:0] I0_3_2_2,
  input  [31:0] I0_4_0_0,
  input  [31:0] I0_4_0_1,
  input  [31:0] I0_4_0_2,
  input  [31:0] I0_4_1_0,
  input  [31:0] I0_4_1_1,
  input  [31:0] I0_4_1_2,
  input  [31:0] I0_4_2_0,
  input  [31:0] I0_4_2_1,
  input  [31:0] I0_4_2_2,
  input  [31:0] I0_5_0_0,
  input  [31:0] I0_5_0_1,
  input  [31:0] I0_5_0_2,
  input  [31:0] I0_5_1_0,
  input  [31:0] I0_5_1_1,
  input  [31:0] I0_5_1_2,
  input  [31:0] I0_5_2_0,
  input  [31:0] I0_5_2_1,
  input  [31:0] I0_5_2_2,
  input  [31:0] I0_6_0_0,
  input  [31:0] I0_6_0_1,
  input  [31:0] I0_6_0_2,
  input  [31:0] I0_6_1_0,
  input  [31:0] I0_6_1_1,
  input  [31:0] I0_6_1_2,
  input  [31:0] I0_6_2_0,
  input  [31:0] I0_6_2_1,
  input  [31:0] I0_6_2_2,
  input  [31:0] I0_7_0_0,
  input  [31:0] I0_7_0_1,
  input  [31:0] I0_7_0_2,
  input  [31:0] I0_7_1_0,
  input  [31:0] I0_7_1_1,
  input  [31:0] I0_7_1_2,
  input  [31:0] I0_7_2_0,
  input  [31:0] I0_7_2_1,
  input  [31:0] I0_7_2_2,
  input         I1_0_0_0_t0b,
  input         I1_0_0_0_t1b,
  input         I1_1_0_0_t0b,
  input         I1_1_0_0_t1b,
  input         I1_2_0_0_t0b,
  input         I1_2_0_0_t1b,
  input         I1_3_0_0_t0b,
  input         I1_3_0_0_t1b,
  input         I1_4_0_0_t0b,
  input         I1_4_0_0_t1b,
  input         I1_5_0_0_t0b,
  input         I1_5_0_0_t1b,
  input         I1_6_0_0_t0b,
  input         I1_6_0_0_t1b,
  input         I1_7_0_0_t0b,
  input         I1_7_0_0_t1b,
  output [31:0] O_0_0_0_t0b,
  output [31:0] O_0_0_0_t1b_t0b,
  output [31:0] O_0_0_0_t1b_t1b,
  output [31:0] O_1_0_0_t0b,
  output [31:0] O_1_0_0_t1b_t0b,
  output [31:0] O_1_0_0_t1b_t1b,
  output [31:0] O_2_0_0_t0b,
  output [31:0] O_2_0_0_t1b_t0b,
  output [31:0] O_2_0_0_t1b_t1b,
  output [31:0] O_3_0_0_t0b,
  output [31:0] O_3_0_0_t1b_t0b,
  output [31:0] O_3_0_0_t1b_t1b,
  output [31:0] O_4_0_0_t0b,
  output [31:0] O_4_0_0_t1b_t0b,
  output [31:0] O_4_0_0_t1b_t1b,
  output [31:0] O_5_0_0_t0b,
  output [31:0] O_5_0_0_t1b_t0b,
  output [31:0] O_5_0_0_t1b_t1b,
  output [31:0] O_6_0_0_t0b,
  output [31:0] O_6_0_0_t1b_t0b,
  output [31:0] O_6_0_0_t1b_t1b,
  output [31:0] O_7_0_0_t0b,
  output [31:0] O_7_0_0_t1b_t0b,
  output [31:0] O_7_0_0_t1b_t1b
);
  wire  op_clock; // @[Map2T.scala 8:20]
  wire  op_reset; // @[Map2T.scala 8:20]
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7_2_2; // @[Map2T.scala 8:20]
  wire  op_I1_0_0_0_t0b; // @[Map2T.scala 8:20]
  wire  op_I1_0_0_0_t1b; // @[Map2T.scala 8:20]
  wire  op_I1_1_0_0_t0b; // @[Map2T.scala 8:20]
  wire  op_I1_1_0_0_t1b; // @[Map2T.scala 8:20]
  wire  op_I1_2_0_0_t0b; // @[Map2T.scala 8:20]
  wire  op_I1_2_0_0_t1b; // @[Map2T.scala 8:20]
  wire  op_I1_3_0_0_t0b; // @[Map2T.scala 8:20]
  wire  op_I1_3_0_0_t1b; // @[Map2T.scala 8:20]
  wire  op_I1_4_0_0_t0b; // @[Map2T.scala 8:20]
  wire  op_I1_4_0_0_t1b; // @[Map2T.scala 8:20]
  wire  op_I1_5_0_0_t0b; // @[Map2T.scala 8:20]
  wire  op_I1_5_0_0_t1b; // @[Map2T.scala 8:20]
  wire  op_I1_6_0_0_t0b; // @[Map2T.scala 8:20]
  wire  op_I1_6_0_0_t1b; // @[Map2T.scala 8:20]
  wire  op_I1_7_0_0_t0b; // @[Map2T.scala 8:20]
  wire  op_I1_7_0_0_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_0_0_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_0_0_t1b_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_0_0_t1b_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_0_0_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_0_0_t1b_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_0_0_t1b_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_0_0_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_0_0_t1b_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_0_0_t1b_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_0_0_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_0_0_t1b_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_0_0_t1b_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_0_0_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_0_0_t1b_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_0_0_t1b_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_0_0_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_0_0_t1b_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_0_0_t1b_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_0_0_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_0_0_t1b_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_0_0_t1b_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_0_0_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_0_0_t1b_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_0_0_t1b_t1b; // @[Map2T.scala 8:20]
  Map2S_53 op ( // @[Map2T.scala 8:20]
    .clock(op_clock),
    .reset(op_reset),
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0_0_0(op_I0_0_0_0),
    .I0_0_0_1(op_I0_0_0_1),
    .I0_0_0_2(op_I0_0_0_2),
    .I0_0_1_0(op_I0_0_1_0),
    .I0_0_1_1(op_I0_0_1_1),
    .I0_0_1_2(op_I0_0_1_2),
    .I0_0_2_0(op_I0_0_2_0),
    .I0_0_2_1(op_I0_0_2_1),
    .I0_0_2_2(op_I0_0_2_2),
    .I0_1_0_0(op_I0_1_0_0),
    .I0_1_0_1(op_I0_1_0_1),
    .I0_1_0_2(op_I0_1_0_2),
    .I0_1_1_0(op_I0_1_1_0),
    .I0_1_1_1(op_I0_1_1_1),
    .I0_1_1_2(op_I0_1_1_2),
    .I0_1_2_0(op_I0_1_2_0),
    .I0_1_2_1(op_I0_1_2_1),
    .I0_1_2_2(op_I0_1_2_2),
    .I0_2_0_0(op_I0_2_0_0),
    .I0_2_0_1(op_I0_2_0_1),
    .I0_2_0_2(op_I0_2_0_2),
    .I0_2_1_0(op_I0_2_1_0),
    .I0_2_1_1(op_I0_2_1_1),
    .I0_2_1_2(op_I0_2_1_2),
    .I0_2_2_0(op_I0_2_2_0),
    .I0_2_2_1(op_I0_2_2_1),
    .I0_2_2_2(op_I0_2_2_2),
    .I0_3_0_0(op_I0_3_0_0),
    .I0_3_0_1(op_I0_3_0_1),
    .I0_3_0_2(op_I0_3_0_2),
    .I0_3_1_0(op_I0_3_1_0),
    .I0_3_1_1(op_I0_3_1_1),
    .I0_3_1_2(op_I0_3_1_2),
    .I0_3_2_0(op_I0_3_2_0),
    .I0_3_2_1(op_I0_3_2_1),
    .I0_3_2_2(op_I0_3_2_2),
    .I0_4_0_0(op_I0_4_0_0),
    .I0_4_0_1(op_I0_4_0_1),
    .I0_4_0_2(op_I0_4_0_2),
    .I0_4_1_0(op_I0_4_1_0),
    .I0_4_1_1(op_I0_4_1_1),
    .I0_4_1_2(op_I0_4_1_2),
    .I0_4_2_0(op_I0_4_2_0),
    .I0_4_2_1(op_I0_4_2_1),
    .I0_4_2_2(op_I0_4_2_2),
    .I0_5_0_0(op_I0_5_0_0),
    .I0_5_0_1(op_I0_5_0_1),
    .I0_5_0_2(op_I0_5_0_2),
    .I0_5_1_0(op_I0_5_1_0),
    .I0_5_1_1(op_I0_5_1_1),
    .I0_5_1_2(op_I0_5_1_2),
    .I0_5_2_0(op_I0_5_2_0),
    .I0_5_2_1(op_I0_5_2_1),
    .I0_5_2_2(op_I0_5_2_2),
    .I0_6_0_0(op_I0_6_0_0),
    .I0_6_0_1(op_I0_6_0_1),
    .I0_6_0_2(op_I0_6_0_2),
    .I0_6_1_0(op_I0_6_1_0),
    .I0_6_1_1(op_I0_6_1_1),
    .I0_6_1_2(op_I0_6_1_2),
    .I0_6_2_0(op_I0_6_2_0),
    .I0_6_2_1(op_I0_6_2_1),
    .I0_6_2_2(op_I0_6_2_2),
    .I0_7_0_0(op_I0_7_0_0),
    .I0_7_0_1(op_I0_7_0_1),
    .I0_7_0_2(op_I0_7_0_2),
    .I0_7_1_0(op_I0_7_1_0),
    .I0_7_1_1(op_I0_7_1_1),
    .I0_7_1_2(op_I0_7_1_2),
    .I0_7_2_0(op_I0_7_2_0),
    .I0_7_2_1(op_I0_7_2_1),
    .I0_7_2_2(op_I0_7_2_2),
    .I1_0_0_0_t0b(op_I1_0_0_0_t0b),
    .I1_0_0_0_t1b(op_I1_0_0_0_t1b),
    .I1_1_0_0_t0b(op_I1_1_0_0_t0b),
    .I1_1_0_0_t1b(op_I1_1_0_0_t1b),
    .I1_2_0_0_t0b(op_I1_2_0_0_t0b),
    .I1_2_0_0_t1b(op_I1_2_0_0_t1b),
    .I1_3_0_0_t0b(op_I1_3_0_0_t0b),
    .I1_3_0_0_t1b(op_I1_3_0_0_t1b),
    .I1_4_0_0_t0b(op_I1_4_0_0_t0b),
    .I1_4_0_0_t1b(op_I1_4_0_0_t1b),
    .I1_5_0_0_t0b(op_I1_5_0_0_t0b),
    .I1_5_0_0_t1b(op_I1_5_0_0_t1b),
    .I1_6_0_0_t0b(op_I1_6_0_0_t0b),
    .I1_6_0_0_t1b(op_I1_6_0_0_t1b),
    .I1_7_0_0_t0b(op_I1_7_0_0_t0b),
    .I1_7_0_0_t1b(op_I1_7_0_0_t1b),
    .O_0_0_0_t0b(op_O_0_0_0_t0b),
    .O_0_0_0_t1b_t0b(op_O_0_0_0_t1b_t0b),
    .O_0_0_0_t1b_t1b(op_O_0_0_0_t1b_t1b),
    .O_1_0_0_t0b(op_O_1_0_0_t0b),
    .O_1_0_0_t1b_t0b(op_O_1_0_0_t1b_t0b),
    .O_1_0_0_t1b_t1b(op_O_1_0_0_t1b_t1b),
    .O_2_0_0_t0b(op_O_2_0_0_t0b),
    .O_2_0_0_t1b_t0b(op_O_2_0_0_t1b_t0b),
    .O_2_0_0_t1b_t1b(op_O_2_0_0_t1b_t1b),
    .O_3_0_0_t0b(op_O_3_0_0_t0b),
    .O_3_0_0_t1b_t0b(op_O_3_0_0_t1b_t0b),
    .O_3_0_0_t1b_t1b(op_O_3_0_0_t1b_t1b),
    .O_4_0_0_t0b(op_O_4_0_0_t0b),
    .O_4_0_0_t1b_t0b(op_O_4_0_0_t1b_t0b),
    .O_4_0_0_t1b_t1b(op_O_4_0_0_t1b_t1b),
    .O_5_0_0_t0b(op_O_5_0_0_t0b),
    .O_5_0_0_t1b_t0b(op_O_5_0_0_t1b_t0b),
    .O_5_0_0_t1b_t1b(op_O_5_0_0_t1b_t1b),
    .O_6_0_0_t0b(op_O_6_0_0_t0b),
    .O_6_0_0_t1b_t0b(op_O_6_0_0_t1b_t0b),
    .O_6_0_0_t1b_t1b(op_O_6_0_0_t1b_t1b),
    .O_7_0_0_t0b(op_O_7_0_0_t0b),
    .O_7_0_0_t1b_t0b(op_O_7_0_0_t1b_t0b),
    .O_7_0_0_t1b_t1b(op_O_7_0_0_t1b_t1b)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_0_0_t0b = op_O_0_0_0_t0b; // @[Map2T.scala 17:7]
  assign O_0_0_0_t1b_t0b = op_O_0_0_0_t1b_t0b; // @[Map2T.scala 17:7]
  assign O_0_0_0_t1b_t1b = op_O_0_0_0_t1b_t1b; // @[Map2T.scala 17:7]
  assign O_1_0_0_t0b = op_O_1_0_0_t0b; // @[Map2T.scala 17:7]
  assign O_1_0_0_t1b_t0b = op_O_1_0_0_t1b_t0b; // @[Map2T.scala 17:7]
  assign O_1_0_0_t1b_t1b = op_O_1_0_0_t1b_t1b; // @[Map2T.scala 17:7]
  assign O_2_0_0_t0b = op_O_2_0_0_t0b; // @[Map2T.scala 17:7]
  assign O_2_0_0_t1b_t0b = op_O_2_0_0_t1b_t0b; // @[Map2T.scala 17:7]
  assign O_2_0_0_t1b_t1b = op_O_2_0_0_t1b_t1b; // @[Map2T.scala 17:7]
  assign O_3_0_0_t0b = op_O_3_0_0_t0b; // @[Map2T.scala 17:7]
  assign O_3_0_0_t1b_t0b = op_O_3_0_0_t1b_t0b; // @[Map2T.scala 17:7]
  assign O_3_0_0_t1b_t1b = op_O_3_0_0_t1b_t1b; // @[Map2T.scala 17:7]
  assign O_4_0_0_t0b = op_O_4_0_0_t0b; // @[Map2T.scala 17:7]
  assign O_4_0_0_t1b_t0b = op_O_4_0_0_t1b_t0b; // @[Map2T.scala 17:7]
  assign O_4_0_0_t1b_t1b = op_O_4_0_0_t1b_t1b; // @[Map2T.scala 17:7]
  assign O_5_0_0_t0b = op_O_5_0_0_t0b; // @[Map2T.scala 17:7]
  assign O_5_0_0_t1b_t0b = op_O_5_0_0_t1b_t0b; // @[Map2T.scala 17:7]
  assign O_5_0_0_t1b_t1b = op_O_5_0_0_t1b_t1b; // @[Map2T.scala 17:7]
  assign O_6_0_0_t0b = op_O_6_0_0_t0b; // @[Map2T.scala 17:7]
  assign O_6_0_0_t1b_t0b = op_O_6_0_0_t1b_t0b; // @[Map2T.scala 17:7]
  assign O_6_0_0_t1b_t1b = op_O_6_0_0_t1b_t1b; // @[Map2T.scala 17:7]
  assign O_7_0_0_t0b = op_O_7_0_0_t0b; // @[Map2T.scala 17:7]
  assign O_7_0_0_t1b_t0b = op_O_7_0_0_t1b_t0b; // @[Map2T.scala 17:7]
  assign O_7_0_0_t1b_t1b = op_O_7_0_0_t1b_t1b; // @[Map2T.scala 17:7]
  assign op_clock = clock;
  assign op_reset = reset;
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0_0_0 = I0_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_0_0_1 = I0_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_0_0_2 = I0_0_0_2; // @[Map2T.scala 15:11]
  assign op_I0_0_1_0 = I0_0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_0_1_1 = I0_0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_0_1_2 = I0_0_1_2; // @[Map2T.scala 15:11]
  assign op_I0_0_2_0 = I0_0_2_0; // @[Map2T.scala 15:11]
  assign op_I0_0_2_1 = I0_0_2_1; // @[Map2T.scala 15:11]
  assign op_I0_0_2_2 = I0_0_2_2; // @[Map2T.scala 15:11]
  assign op_I0_1_0_0 = I0_1_0_0; // @[Map2T.scala 15:11]
  assign op_I0_1_0_1 = I0_1_0_1; // @[Map2T.scala 15:11]
  assign op_I0_1_0_2 = I0_1_0_2; // @[Map2T.scala 15:11]
  assign op_I0_1_1_0 = I0_1_1_0; // @[Map2T.scala 15:11]
  assign op_I0_1_1_1 = I0_1_1_1; // @[Map2T.scala 15:11]
  assign op_I0_1_1_2 = I0_1_1_2; // @[Map2T.scala 15:11]
  assign op_I0_1_2_0 = I0_1_2_0; // @[Map2T.scala 15:11]
  assign op_I0_1_2_1 = I0_1_2_1; // @[Map2T.scala 15:11]
  assign op_I0_1_2_2 = I0_1_2_2; // @[Map2T.scala 15:11]
  assign op_I0_2_0_0 = I0_2_0_0; // @[Map2T.scala 15:11]
  assign op_I0_2_0_1 = I0_2_0_1; // @[Map2T.scala 15:11]
  assign op_I0_2_0_2 = I0_2_0_2; // @[Map2T.scala 15:11]
  assign op_I0_2_1_0 = I0_2_1_0; // @[Map2T.scala 15:11]
  assign op_I0_2_1_1 = I0_2_1_1; // @[Map2T.scala 15:11]
  assign op_I0_2_1_2 = I0_2_1_2; // @[Map2T.scala 15:11]
  assign op_I0_2_2_0 = I0_2_2_0; // @[Map2T.scala 15:11]
  assign op_I0_2_2_1 = I0_2_2_1; // @[Map2T.scala 15:11]
  assign op_I0_2_2_2 = I0_2_2_2; // @[Map2T.scala 15:11]
  assign op_I0_3_0_0 = I0_3_0_0; // @[Map2T.scala 15:11]
  assign op_I0_3_0_1 = I0_3_0_1; // @[Map2T.scala 15:11]
  assign op_I0_3_0_2 = I0_3_0_2; // @[Map2T.scala 15:11]
  assign op_I0_3_1_0 = I0_3_1_0; // @[Map2T.scala 15:11]
  assign op_I0_3_1_1 = I0_3_1_1; // @[Map2T.scala 15:11]
  assign op_I0_3_1_2 = I0_3_1_2; // @[Map2T.scala 15:11]
  assign op_I0_3_2_0 = I0_3_2_0; // @[Map2T.scala 15:11]
  assign op_I0_3_2_1 = I0_3_2_1; // @[Map2T.scala 15:11]
  assign op_I0_3_2_2 = I0_3_2_2; // @[Map2T.scala 15:11]
  assign op_I0_4_0_0 = I0_4_0_0; // @[Map2T.scala 15:11]
  assign op_I0_4_0_1 = I0_4_0_1; // @[Map2T.scala 15:11]
  assign op_I0_4_0_2 = I0_4_0_2; // @[Map2T.scala 15:11]
  assign op_I0_4_1_0 = I0_4_1_0; // @[Map2T.scala 15:11]
  assign op_I0_4_1_1 = I0_4_1_1; // @[Map2T.scala 15:11]
  assign op_I0_4_1_2 = I0_4_1_2; // @[Map2T.scala 15:11]
  assign op_I0_4_2_0 = I0_4_2_0; // @[Map2T.scala 15:11]
  assign op_I0_4_2_1 = I0_4_2_1; // @[Map2T.scala 15:11]
  assign op_I0_4_2_2 = I0_4_2_2; // @[Map2T.scala 15:11]
  assign op_I0_5_0_0 = I0_5_0_0; // @[Map2T.scala 15:11]
  assign op_I0_5_0_1 = I0_5_0_1; // @[Map2T.scala 15:11]
  assign op_I0_5_0_2 = I0_5_0_2; // @[Map2T.scala 15:11]
  assign op_I0_5_1_0 = I0_5_1_0; // @[Map2T.scala 15:11]
  assign op_I0_5_1_1 = I0_5_1_1; // @[Map2T.scala 15:11]
  assign op_I0_5_1_2 = I0_5_1_2; // @[Map2T.scala 15:11]
  assign op_I0_5_2_0 = I0_5_2_0; // @[Map2T.scala 15:11]
  assign op_I0_5_2_1 = I0_5_2_1; // @[Map2T.scala 15:11]
  assign op_I0_5_2_2 = I0_5_2_2; // @[Map2T.scala 15:11]
  assign op_I0_6_0_0 = I0_6_0_0; // @[Map2T.scala 15:11]
  assign op_I0_6_0_1 = I0_6_0_1; // @[Map2T.scala 15:11]
  assign op_I0_6_0_2 = I0_6_0_2; // @[Map2T.scala 15:11]
  assign op_I0_6_1_0 = I0_6_1_0; // @[Map2T.scala 15:11]
  assign op_I0_6_1_1 = I0_6_1_1; // @[Map2T.scala 15:11]
  assign op_I0_6_1_2 = I0_6_1_2; // @[Map2T.scala 15:11]
  assign op_I0_6_2_0 = I0_6_2_0; // @[Map2T.scala 15:11]
  assign op_I0_6_2_1 = I0_6_2_1; // @[Map2T.scala 15:11]
  assign op_I0_6_2_2 = I0_6_2_2; // @[Map2T.scala 15:11]
  assign op_I0_7_0_0 = I0_7_0_0; // @[Map2T.scala 15:11]
  assign op_I0_7_0_1 = I0_7_0_1; // @[Map2T.scala 15:11]
  assign op_I0_7_0_2 = I0_7_0_2; // @[Map2T.scala 15:11]
  assign op_I0_7_1_0 = I0_7_1_0; // @[Map2T.scala 15:11]
  assign op_I0_7_1_1 = I0_7_1_1; // @[Map2T.scala 15:11]
  assign op_I0_7_1_2 = I0_7_1_2; // @[Map2T.scala 15:11]
  assign op_I0_7_2_0 = I0_7_2_0; // @[Map2T.scala 15:11]
  assign op_I0_7_2_1 = I0_7_2_1; // @[Map2T.scala 15:11]
  assign op_I0_7_2_2 = I0_7_2_2; // @[Map2T.scala 15:11]
  assign op_I1_0_0_0_t0b = I1_0_0_0_t0b; // @[Map2T.scala 16:11]
  assign op_I1_0_0_0_t1b = I1_0_0_0_t1b; // @[Map2T.scala 16:11]
  assign op_I1_1_0_0_t0b = I1_1_0_0_t0b; // @[Map2T.scala 16:11]
  assign op_I1_1_0_0_t1b = I1_1_0_0_t1b; // @[Map2T.scala 16:11]
  assign op_I1_2_0_0_t0b = I1_2_0_0_t0b; // @[Map2T.scala 16:11]
  assign op_I1_2_0_0_t1b = I1_2_0_0_t1b; // @[Map2T.scala 16:11]
  assign op_I1_3_0_0_t0b = I1_3_0_0_t0b; // @[Map2T.scala 16:11]
  assign op_I1_3_0_0_t1b = I1_3_0_0_t1b; // @[Map2T.scala 16:11]
  assign op_I1_4_0_0_t0b = I1_4_0_0_t0b; // @[Map2T.scala 16:11]
  assign op_I1_4_0_0_t1b = I1_4_0_0_t1b; // @[Map2T.scala 16:11]
  assign op_I1_5_0_0_t0b = I1_5_0_0_t0b; // @[Map2T.scala 16:11]
  assign op_I1_5_0_0_t1b = I1_5_0_0_t1b; // @[Map2T.scala 16:11]
  assign op_I1_6_0_0_t0b = I1_6_0_0_t0b; // @[Map2T.scala 16:11]
  assign op_I1_6_0_0_t1b = I1_6_0_0_t1b; // @[Map2T.scala 16:11]
  assign op_I1_7_0_0_t0b = I1_7_0_0_t0b; // @[Map2T.scala 16:11]
  assign op_I1_7_0_0_t1b = I1_7_0_0_t1b; // @[Map2T.scala 16:11]
endmodule
module Module_7(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0_0,
  input  [31:0] I_0_0_1,
  input  [31:0] I_0_0_2,
  input  [31:0] I_0_1_0,
  input  [31:0] I_0_1_1,
  input  [31:0] I_0_1_2,
  input  [31:0] I_0_2_0,
  input  [31:0] I_0_2_1,
  input  [31:0] I_0_2_2,
  input  [31:0] I_1_0_0,
  input  [31:0] I_1_0_1,
  input  [31:0] I_1_0_2,
  input  [31:0] I_1_1_0,
  input  [31:0] I_1_1_1,
  input  [31:0] I_1_1_2,
  input  [31:0] I_1_2_0,
  input  [31:0] I_1_2_1,
  input  [31:0] I_1_2_2,
  input  [31:0] I_2_0_0,
  input  [31:0] I_2_0_1,
  input  [31:0] I_2_0_2,
  input  [31:0] I_2_1_0,
  input  [31:0] I_2_1_1,
  input  [31:0] I_2_1_2,
  input  [31:0] I_2_2_0,
  input  [31:0] I_2_2_1,
  input  [31:0] I_2_2_2,
  input  [31:0] I_3_0_0,
  input  [31:0] I_3_0_1,
  input  [31:0] I_3_0_2,
  input  [31:0] I_3_1_0,
  input  [31:0] I_3_1_1,
  input  [31:0] I_3_1_2,
  input  [31:0] I_3_2_0,
  input  [31:0] I_3_2_1,
  input  [31:0] I_3_2_2,
  input  [31:0] I_4_0_0,
  input  [31:0] I_4_0_1,
  input  [31:0] I_4_0_2,
  input  [31:0] I_4_1_0,
  input  [31:0] I_4_1_1,
  input  [31:0] I_4_1_2,
  input  [31:0] I_4_2_0,
  input  [31:0] I_4_2_1,
  input  [31:0] I_4_2_2,
  input  [31:0] I_5_0_0,
  input  [31:0] I_5_0_1,
  input  [31:0] I_5_0_2,
  input  [31:0] I_5_1_0,
  input  [31:0] I_5_1_1,
  input  [31:0] I_5_1_2,
  input  [31:0] I_5_2_0,
  input  [31:0] I_5_2_1,
  input  [31:0] I_5_2_2,
  input  [31:0] I_6_0_0,
  input  [31:0] I_6_0_1,
  input  [31:0] I_6_0_2,
  input  [31:0] I_6_1_0,
  input  [31:0] I_6_1_1,
  input  [31:0] I_6_1_2,
  input  [31:0] I_6_2_0,
  input  [31:0] I_6_2_1,
  input  [31:0] I_6_2_2,
  input  [31:0] I_7_0_0,
  input  [31:0] I_7_0_1,
  input  [31:0] I_7_0_2,
  input  [31:0] I_7_1_0,
  input  [31:0] I_7_1_1,
  input  [31:0] I_7_1_2,
  input  [31:0] I_7_2_0,
  input  [31:0] I_7_2_1,
  input  [31:0] I_7_2_2,
  output [31:0] O_0_0_0_t0b,
  output [31:0] O_0_0_0_t1b_t0b,
  output [31:0] O_0_0_0_t1b_t1b,
  output [31:0] O_1_0_0_t0b,
  output [31:0] O_1_0_0_t1b_t0b,
  output [31:0] O_1_0_0_t1b_t1b,
  output [31:0] O_2_0_0_t0b,
  output [31:0] O_2_0_0_t1b_t0b,
  output [31:0] O_2_0_0_t1b_t1b,
  output [31:0] O_3_0_0_t0b,
  output [31:0] O_3_0_0_t1b_t0b,
  output [31:0] O_3_0_0_t1b_t1b,
  output [31:0] O_4_0_0_t0b,
  output [31:0] O_4_0_0_t1b_t0b,
  output [31:0] O_4_0_0_t1b_t1b,
  output [31:0] O_5_0_0_t0b,
  output [31:0] O_5_0_0_t1b_t0b,
  output [31:0] O_5_0_0_t1b_t1b,
  output [31:0] O_6_0_0_t0b,
  output [31:0] O_6_0_0_t1b_t0b,
  output [31:0] O_6_0_0_t1b_t1b,
  output [31:0] O_7_0_0_t0b,
  output [31:0] O_7_0_0_t1b_t0b,
  output [31:0] O_7_0_0_t1b_t1b
);
  wire  counter108_clock; // @[Top.scala 325:28]
  wire  counter108_reset; // @[Top.scala 325:28]
  wire [31:0] counter108_O_0; // @[Top.scala 325:28]
  wire [31:0] counter108_O_1; // @[Top.scala 325:28]
  wire [31:0] counter108_O_2; // @[Top.scala 325:28]
  wire [31:0] counter108_O_3; // @[Top.scala 325:28]
  wire [31:0] counter108_O_4; // @[Top.scala 325:28]
  wire [31:0] counter108_O_5; // @[Top.scala 325:28]
  wire [31:0] counter108_O_6; // @[Top.scala 325:28]
  wire [31:0] counter108_O_7; // @[Top.scala 325:28]
  wire  n116_valid_down; // @[Top.scala 327:22]
  wire [31:0] n116_I_0; // @[Top.scala 327:22]
  wire [31:0] n116_I_1; // @[Top.scala 327:22]
  wire [31:0] n116_I_2; // @[Top.scala 327:22]
  wire [31:0] n116_I_3; // @[Top.scala 327:22]
  wire [31:0] n116_I_4; // @[Top.scala 327:22]
  wire [31:0] n116_I_5; // @[Top.scala 327:22]
  wire [31:0] n116_I_6; // @[Top.scala 327:22]
  wire [31:0] n116_I_7; // @[Top.scala 327:22]
  wire  n116_O_0; // @[Top.scala 327:22]
  wire  n116_O_1; // @[Top.scala 327:22]
  wire  n116_O_2; // @[Top.scala 327:22]
  wire  n116_O_3; // @[Top.scala 327:22]
  wire  n116_O_4; // @[Top.scala 327:22]
  wire  n116_O_5; // @[Top.scala 327:22]
  wire  n116_O_6; // @[Top.scala 327:22]
  wire  n116_O_7; // @[Top.scala 327:22]
  wire  n128_valid_down; // @[Top.scala 330:22]
  wire [31:0] n128_I_0; // @[Top.scala 330:22]
  wire [31:0] n128_I_1; // @[Top.scala 330:22]
  wire [31:0] n128_I_2; // @[Top.scala 330:22]
  wire [31:0] n128_I_3; // @[Top.scala 330:22]
  wire [31:0] n128_I_4; // @[Top.scala 330:22]
  wire [31:0] n128_I_5; // @[Top.scala 330:22]
  wire [31:0] n128_I_6; // @[Top.scala 330:22]
  wire [31:0] n128_I_7; // @[Top.scala 330:22]
  wire  n128_O_0; // @[Top.scala 330:22]
  wire  n128_O_1; // @[Top.scala 330:22]
  wire  n128_O_2; // @[Top.scala 330:22]
  wire  n128_O_3; // @[Top.scala 330:22]
  wire  n128_O_4; // @[Top.scala 330:22]
  wire  n128_O_5; // @[Top.scala 330:22]
  wire  n128_O_6; // @[Top.scala 330:22]
  wire  n128_O_7; // @[Top.scala 330:22]
  wire  n129_valid_up; // @[Top.scala 333:22]
  wire  n129_valid_down; // @[Top.scala 333:22]
  wire  n129_I0_0; // @[Top.scala 333:22]
  wire  n129_I0_1; // @[Top.scala 333:22]
  wire  n129_I0_2; // @[Top.scala 333:22]
  wire  n129_I0_3; // @[Top.scala 333:22]
  wire  n129_I0_4; // @[Top.scala 333:22]
  wire  n129_I0_5; // @[Top.scala 333:22]
  wire  n129_I0_6; // @[Top.scala 333:22]
  wire  n129_I0_7; // @[Top.scala 333:22]
  wire  n129_I1_0; // @[Top.scala 333:22]
  wire  n129_I1_1; // @[Top.scala 333:22]
  wire  n129_I1_2; // @[Top.scala 333:22]
  wire  n129_I1_3; // @[Top.scala 333:22]
  wire  n129_I1_4; // @[Top.scala 333:22]
  wire  n129_I1_5; // @[Top.scala 333:22]
  wire  n129_I1_6; // @[Top.scala 333:22]
  wire  n129_I1_7; // @[Top.scala 333:22]
  wire  n129_O_0_t0b; // @[Top.scala 333:22]
  wire  n129_O_0_t1b; // @[Top.scala 333:22]
  wire  n129_O_1_t0b; // @[Top.scala 333:22]
  wire  n129_O_1_t1b; // @[Top.scala 333:22]
  wire  n129_O_2_t0b; // @[Top.scala 333:22]
  wire  n129_O_2_t1b; // @[Top.scala 333:22]
  wire  n129_O_3_t0b; // @[Top.scala 333:22]
  wire  n129_O_3_t1b; // @[Top.scala 333:22]
  wire  n129_O_4_t0b; // @[Top.scala 333:22]
  wire  n129_O_4_t1b; // @[Top.scala 333:22]
  wire  n129_O_5_t0b; // @[Top.scala 333:22]
  wire  n129_O_5_t1b; // @[Top.scala 333:22]
  wire  n129_O_6_t0b; // @[Top.scala 333:22]
  wire  n129_O_6_t1b; // @[Top.scala 333:22]
  wire  n129_O_7_t0b; // @[Top.scala 333:22]
  wire  n129_O_7_t1b; // @[Top.scala 333:22]
  wire  n138_valid_up; // @[Top.scala 337:22]
  wire  n138_valid_down; // @[Top.scala 337:22]
  wire  n138_I_0_t0b; // @[Top.scala 337:22]
  wire  n138_I_0_t1b; // @[Top.scala 337:22]
  wire  n138_I_1_t0b; // @[Top.scala 337:22]
  wire  n138_I_1_t1b; // @[Top.scala 337:22]
  wire  n138_I_2_t0b; // @[Top.scala 337:22]
  wire  n138_I_2_t1b; // @[Top.scala 337:22]
  wire  n138_I_3_t0b; // @[Top.scala 337:22]
  wire  n138_I_3_t1b; // @[Top.scala 337:22]
  wire  n138_I_4_t0b; // @[Top.scala 337:22]
  wire  n138_I_4_t1b; // @[Top.scala 337:22]
  wire  n138_I_5_t0b; // @[Top.scala 337:22]
  wire  n138_I_5_t1b; // @[Top.scala 337:22]
  wire  n138_I_6_t0b; // @[Top.scala 337:22]
  wire  n138_I_6_t1b; // @[Top.scala 337:22]
  wire  n138_I_7_t0b; // @[Top.scala 337:22]
  wire  n138_I_7_t1b; // @[Top.scala 337:22]
  wire  n138_O_0_0_t0b; // @[Top.scala 337:22]
  wire  n138_O_0_0_t1b; // @[Top.scala 337:22]
  wire  n138_O_1_0_t0b; // @[Top.scala 337:22]
  wire  n138_O_1_0_t1b; // @[Top.scala 337:22]
  wire  n138_O_2_0_t0b; // @[Top.scala 337:22]
  wire  n138_O_2_0_t1b; // @[Top.scala 337:22]
  wire  n138_O_3_0_t0b; // @[Top.scala 337:22]
  wire  n138_O_3_0_t1b; // @[Top.scala 337:22]
  wire  n138_O_4_0_t0b; // @[Top.scala 337:22]
  wire  n138_O_4_0_t1b; // @[Top.scala 337:22]
  wire  n138_O_5_0_t0b; // @[Top.scala 337:22]
  wire  n138_O_5_0_t1b; // @[Top.scala 337:22]
  wire  n138_O_6_0_t0b; // @[Top.scala 337:22]
  wire  n138_O_6_0_t1b; // @[Top.scala 337:22]
  wire  n138_O_7_0_t0b; // @[Top.scala 337:22]
  wire  n138_O_7_0_t1b; // @[Top.scala 337:22]
  wire  n141_valid_up; // @[Top.scala 340:22]
  wire  n141_valid_down; // @[Top.scala 340:22]
  wire  n141_I_0_0_t0b; // @[Top.scala 340:22]
  wire  n141_I_0_0_t1b; // @[Top.scala 340:22]
  wire  n141_I_1_0_t0b; // @[Top.scala 340:22]
  wire  n141_I_1_0_t1b; // @[Top.scala 340:22]
  wire  n141_I_2_0_t0b; // @[Top.scala 340:22]
  wire  n141_I_2_0_t1b; // @[Top.scala 340:22]
  wire  n141_I_3_0_t0b; // @[Top.scala 340:22]
  wire  n141_I_3_0_t1b; // @[Top.scala 340:22]
  wire  n141_I_4_0_t0b; // @[Top.scala 340:22]
  wire  n141_I_4_0_t1b; // @[Top.scala 340:22]
  wire  n141_I_5_0_t0b; // @[Top.scala 340:22]
  wire  n141_I_5_0_t1b; // @[Top.scala 340:22]
  wire  n141_I_6_0_t0b; // @[Top.scala 340:22]
  wire  n141_I_6_0_t1b; // @[Top.scala 340:22]
  wire  n141_I_7_0_t0b; // @[Top.scala 340:22]
  wire  n141_I_7_0_t1b; // @[Top.scala 340:22]
  wire  n141_O_0_0_0_t0b; // @[Top.scala 340:22]
  wire  n141_O_0_0_0_t1b; // @[Top.scala 340:22]
  wire  n141_O_1_0_0_t0b; // @[Top.scala 340:22]
  wire  n141_O_1_0_0_t1b; // @[Top.scala 340:22]
  wire  n141_O_2_0_0_t0b; // @[Top.scala 340:22]
  wire  n141_O_2_0_0_t1b; // @[Top.scala 340:22]
  wire  n141_O_3_0_0_t0b; // @[Top.scala 340:22]
  wire  n141_O_3_0_0_t1b; // @[Top.scala 340:22]
  wire  n141_O_4_0_0_t0b; // @[Top.scala 340:22]
  wire  n141_O_4_0_0_t1b; // @[Top.scala 340:22]
  wire  n141_O_5_0_0_t0b; // @[Top.scala 340:22]
  wire  n141_O_5_0_0_t1b; // @[Top.scala 340:22]
  wire  n141_O_6_0_0_t0b; // @[Top.scala 340:22]
  wire  n141_O_6_0_0_t1b; // @[Top.scala 340:22]
  wire  n141_O_7_0_0_t0b; // @[Top.scala 340:22]
  wire  n141_O_7_0_0_t1b; // @[Top.scala 340:22]
  wire  n142_clock; // @[Top.scala 343:22]
  wire  n142_reset; // @[Top.scala 343:22]
  wire  n142_valid_up; // @[Top.scala 343:22]
  wire  n142_valid_down; // @[Top.scala 343:22]
  wire  n142_I_0_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_I_0_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_I_1_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_I_1_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_I_2_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_I_2_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_I_3_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_I_3_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_I_4_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_I_4_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_I_5_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_I_5_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_I_6_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_I_6_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_I_7_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_I_7_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_O_0_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_O_0_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_O_1_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_O_1_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_O_2_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_O_2_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_O_3_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_O_3_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_O_4_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_O_4_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_O_5_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_O_5_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_O_6_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_O_6_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_O_7_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_O_7_0_0_t1b; // @[Top.scala 343:22]
  wire  n143_clock; // @[Top.scala 346:22]
  wire  n143_reset; // @[Top.scala 346:22]
  wire  n143_valid_up; // @[Top.scala 346:22]
  wire  n143_valid_down; // @[Top.scala 346:22]
  wire [31:0] n143_I0_0_0_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_0_0_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_0_0_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_0_1_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_0_1_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_0_1_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_0_2_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_0_2_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_0_2_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_1_0_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_1_0_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_1_0_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_1_1_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_1_1_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_1_1_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_1_2_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_1_2_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_1_2_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_2_0_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_2_0_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_2_0_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_2_1_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_2_1_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_2_1_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_2_2_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_2_2_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_2_2_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_3_0_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_3_0_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_3_0_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_3_1_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_3_1_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_3_1_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_3_2_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_3_2_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_3_2_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_4_0_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_4_0_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_4_0_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_4_1_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_4_1_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_4_1_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_4_2_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_4_2_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_4_2_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_5_0_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_5_0_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_5_0_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_5_1_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_5_1_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_5_1_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_5_2_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_5_2_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_5_2_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_6_0_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_6_0_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_6_0_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_6_1_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_6_1_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_6_1_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_6_2_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_6_2_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_6_2_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_7_0_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_7_0_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_7_0_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_7_1_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_7_1_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_7_1_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_7_2_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_7_2_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_7_2_2; // @[Top.scala 346:22]
  wire  n143_I1_0_0_0_t0b; // @[Top.scala 346:22]
  wire  n143_I1_0_0_0_t1b; // @[Top.scala 346:22]
  wire  n143_I1_1_0_0_t0b; // @[Top.scala 346:22]
  wire  n143_I1_1_0_0_t1b; // @[Top.scala 346:22]
  wire  n143_I1_2_0_0_t0b; // @[Top.scala 346:22]
  wire  n143_I1_2_0_0_t1b; // @[Top.scala 346:22]
  wire  n143_I1_3_0_0_t0b; // @[Top.scala 346:22]
  wire  n143_I1_3_0_0_t1b; // @[Top.scala 346:22]
  wire  n143_I1_4_0_0_t0b; // @[Top.scala 346:22]
  wire  n143_I1_4_0_0_t1b; // @[Top.scala 346:22]
  wire  n143_I1_5_0_0_t0b; // @[Top.scala 346:22]
  wire  n143_I1_5_0_0_t1b; // @[Top.scala 346:22]
  wire  n143_I1_6_0_0_t0b; // @[Top.scala 346:22]
  wire  n143_I1_6_0_0_t1b; // @[Top.scala 346:22]
  wire  n143_I1_7_0_0_t0b; // @[Top.scala 346:22]
  wire  n143_I1_7_0_0_t1b; // @[Top.scala 346:22]
  wire [31:0] n143_O_0_0_0_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_0_0_0_t1b_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_0_0_0_t1b_t1b; // @[Top.scala 346:22]
  wire [31:0] n143_O_1_0_0_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_1_0_0_t1b_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_1_0_0_t1b_t1b; // @[Top.scala 346:22]
  wire [31:0] n143_O_2_0_0_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_2_0_0_t1b_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_2_0_0_t1b_t1b; // @[Top.scala 346:22]
  wire [31:0] n143_O_3_0_0_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_3_0_0_t1b_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_3_0_0_t1b_t1b; // @[Top.scala 346:22]
  wire [31:0] n143_O_4_0_0_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_4_0_0_t1b_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_4_0_0_t1b_t1b; // @[Top.scala 346:22]
  wire [31:0] n143_O_5_0_0_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_5_0_0_t1b_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_5_0_0_t1b_t1b; // @[Top.scala 346:22]
  wire [31:0] n143_O_6_0_0_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_6_0_0_t1b_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_6_0_0_t1b_t1b; // @[Top.scala 346:22]
  wire [31:0] n143_O_7_0_0_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_7_0_0_t1b_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_7_0_0_t1b_t1b; // @[Top.scala 346:22]
  Counter_TS counter108 ( // @[Top.scala 325:28]
    .clock(counter108_clock),
    .reset(counter108_reset),
    .O_0(counter108_O_0),
    .O_1(counter108_O_1),
    .O_2(counter108_O_2),
    .O_3(counter108_O_3),
    .O_4(counter108_O_4),
    .O_5(counter108_O_5),
    .O_6(counter108_O_6),
    .O_7(counter108_O_7)
  );
  MapT_8 n116 ( // @[Top.scala 327:22]
    .valid_down(n116_valid_down),
    .I_0(n116_I_0),
    .I_1(n116_I_1),
    .I_2(n116_I_2),
    .I_3(n116_I_3),
    .I_4(n116_I_4),
    .I_5(n116_I_5),
    .I_6(n116_I_6),
    .I_7(n116_I_7),
    .O_0(n116_O_0),
    .O_1(n116_O_1),
    .O_2(n116_O_2),
    .O_3(n116_O_3),
    .O_4(n116_O_4),
    .O_5(n116_O_5),
    .O_6(n116_O_6),
    .O_7(n116_O_7)
  );
  MapT_9 n128 ( // @[Top.scala 330:22]
    .valid_down(n128_valid_down),
    .I_0(n128_I_0),
    .I_1(n128_I_1),
    .I_2(n128_I_2),
    .I_3(n128_I_3),
    .I_4(n128_I_4),
    .I_5(n128_I_5),
    .I_6(n128_I_6),
    .I_7(n128_I_7),
    .O_0(n128_O_0),
    .O_1(n128_O_1),
    .O_2(n128_O_2),
    .O_3(n128_O_3),
    .O_4(n128_O_4),
    .O_5(n128_O_5),
    .O_6(n128_O_6),
    .O_7(n128_O_7)
  );
  Map2T_8 n129 ( // @[Top.scala 333:22]
    .valid_up(n129_valid_up),
    .valid_down(n129_valid_down),
    .I0_0(n129_I0_0),
    .I0_1(n129_I0_1),
    .I0_2(n129_I0_2),
    .I0_3(n129_I0_3),
    .I0_4(n129_I0_4),
    .I0_5(n129_I0_5),
    .I0_6(n129_I0_6),
    .I0_7(n129_I0_7),
    .I1_0(n129_I1_0),
    .I1_1(n129_I1_1),
    .I1_2(n129_I1_2),
    .I1_3(n129_I1_3),
    .I1_4(n129_I1_4),
    .I1_5(n129_I1_5),
    .I1_6(n129_I1_6),
    .I1_7(n129_I1_7),
    .O_0_t0b(n129_O_0_t0b),
    .O_0_t1b(n129_O_0_t1b),
    .O_1_t0b(n129_O_1_t0b),
    .O_1_t1b(n129_O_1_t1b),
    .O_2_t0b(n129_O_2_t0b),
    .O_2_t1b(n129_O_2_t1b),
    .O_3_t0b(n129_O_3_t0b),
    .O_3_t1b(n129_O_3_t1b),
    .O_4_t0b(n129_O_4_t0b),
    .O_4_t1b(n129_O_4_t1b),
    .O_5_t0b(n129_O_5_t0b),
    .O_5_t1b(n129_O_5_t1b),
    .O_6_t0b(n129_O_6_t0b),
    .O_6_t1b(n129_O_6_t1b),
    .O_7_t0b(n129_O_7_t0b),
    .O_7_t1b(n129_O_7_t1b)
  );
  MapT_10 n138 ( // @[Top.scala 337:22]
    .valid_up(n138_valid_up),
    .valid_down(n138_valid_down),
    .I_0_t0b(n138_I_0_t0b),
    .I_0_t1b(n138_I_0_t1b),
    .I_1_t0b(n138_I_1_t0b),
    .I_1_t1b(n138_I_1_t1b),
    .I_2_t0b(n138_I_2_t0b),
    .I_2_t1b(n138_I_2_t1b),
    .I_3_t0b(n138_I_3_t0b),
    .I_3_t1b(n138_I_3_t1b),
    .I_4_t0b(n138_I_4_t0b),
    .I_4_t1b(n138_I_4_t1b),
    .I_5_t0b(n138_I_5_t0b),
    .I_5_t1b(n138_I_5_t1b),
    .I_6_t0b(n138_I_6_t0b),
    .I_6_t1b(n138_I_6_t1b),
    .I_7_t0b(n138_I_7_t0b),
    .I_7_t1b(n138_I_7_t1b),
    .O_0_0_t0b(n138_O_0_0_t0b),
    .O_0_0_t1b(n138_O_0_0_t1b),
    .O_1_0_t0b(n138_O_1_0_t0b),
    .O_1_0_t1b(n138_O_1_0_t1b),
    .O_2_0_t0b(n138_O_2_0_t0b),
    .O_2_0_t1b(n138_O_2_0_t1b),
    .O_3_0_t0b(n138_O_3_0_t0b),
    .O_3_0_t1b(n138_O_3_0_t1b),
    .O_4_0_t0b(n138_O_4_0_t0b),
    .O_4_0_t1b(n138_O_4_0_t1b),
    .O_5_0_t0b(n138_O_5_0_t0b),
    .O_5_0_t1b(n138_O_5_0_t1b),
    .O_6_0_t0b(n138_O_6_0_t0b),
    .O_6_0_t1b(n138_O_6_0_t1b),
    .O_7_0_t0b(n138_O_7_0_t0b),
    .O_7_0_t1b(n138_O_7_0_t1b)
  );
  MapT_11 n141 ( // @[Top.scala 340:22]
    .valid_up(n141_valid_up),
    .valid_down(n141_valid_down),
    .I_0_0_t0b(n141_I_0_0_t0b),
    .I_0_0_t1b(n141_I_0_0_t1b),
    .I_1_0_t0b(n141_I_1_0_t0b),
    .I_1_0_t1b(n141_I_1_0_t1b),
    .I_2_0_t0b(n141_I_2_0_t0b),
    .I_2_0_t1b(n141_I_2_0_t1b),
    .I_3_0_t0b(n141_I_3_0_t0b),
    .I_3_0_t1b(n141_I_3_0_t1b),
    .I_4_0_t0b(n141_I_4_0_t0b),
    .I_4_0_t1b(n141_I_4_0_t1b),
    .I_5_0_t0b(n141_I_5_0_t0b),
    .I_5_0_t1b(n141_I_5_0_t1b),
    .I_6_0_t0b(n141_I_6_0_t0b),
    .I_6_0_t1b(n141_I_6_0_t1b),
    .I_7_0_t0b(n141_I_7_0_t0b),
    .I_7_0_t1b(n141_I_7_0_t1b),
    .O_0_0_0_t0b(n141_O_0_0_0_t0b),
    .O_0_0_0_t1b(n141_O_0_0_0_t1b),
    .O_1_0_0_t0b(n141_O_1_0_0_t0b),
    .O_1_0_0_t1b(n141_O_1_0_0_t1b),
    .O_2_0_0_t0b(n141_O_2_0_0_t0b),
    .O_2_0_0_t1b(n141_O_2_0_0_t1b),
    .O_3_0_0_t0b(n141_O_3_0_0_t0b),
    .O_3_0_0_t1b(n141_O_3_0_0_t1b),
    .O_4_0_0_t0b(n141_O_4_0_0_t0b),
    .O_4_0_0_t1b(n141_O_4_0_0_t1b),
    .O_5_0_0_t0b(n141_O_5_0_0_t0b),
    .O_5_0_0_t1b(n141_O_5_0_0_t1b),
    .O_6_0_0_t0b(n141_O_6_0_0_t0b),
    .O_6_0_0_t1b(n141_O_6_0_0_t1b),
    .O_7_0_0_t0b(n141_O_7_0_0_t0b),
    .O_7_0_0_t1b(n141_O_7_0_0_t1b)
  );
  FIFO_1 n142 ( // @[Top.scala 343:22]
    .clock(n142_clock),
    .reset(n142_reset),
    .valid_up(n142_valid_up),
    .valid_down(n142_valid_down),
    .I_0_0_0_t0b(n142_I_0_0_0_t0b),
    .I_0_0_0_t1b(n142_I_0_0_0_t1b),
    .I_1_0_0_t0b(n142_I_1_0_0_t0b),
    .I_1_0_0_t1b(n142_I_1_0_0_t1b),
    .I_2_0_0_t0b(n142_I_2_0_0_t0b),
    .I_2_0_0_t1b(n142_I_2_0_0_t1b),
    .I_3_0_0_t0b(n142_I_3_0_0_t0b),
    .I_3_0_0_t1b(n142_I_3_0_0_t1b),
    .I_4_0_0_t0b(n142_I_4_0_0_t0b),
    .I_4_0_0_t1b(n142_I_4_0_0_t1b),
    .I_5_0_0_t0b(n142_I_5_0_0_t0b),
    .I_5_0_0_t1b(n142_I_5_0_0_t1b),
    .I_6_0_0_t0b(n142_I_6_0_0_t0b),
    .I_6_0_0_t1b(n142_I_6_0_0_t1b),
    .I_7_0_0_t0b(n142_I_7_0_0_t0b),
    .I_7_0_0_t1b(n142_I_7_0_0_t1b),
    .O_0_0_0_t0b(n142_O_0_0_0_t0b),
    .O_0_0_0_t1b(n142_O_0_0_0_t1b),
    .O_1_0_0_t0b(n142_O_1_0_0_t0b),
    .O_1_0_0_t1b(n142_O_1_0_0_t1b),
    .O_2_0_0_t0b(n142_O_2_0_0_t0b),
    .O_2_0_0_t1b(n142_O_2_0_0_t1b),
    .O_3_0_0_t0b(n142_O_3_0_0_t0b),
    .O_3_0_0_t1b(n142_O_3_0_0_t1b),
    .O_4_0_0_t0b(n142_O_4_0_0_t0b),
    .O_4_0_0_t1b(n142_O_4_0_0_t1b),
    .O_5_0_0_t0b(n142_O_5_0_0_t0b),
    .O_5_0_0_t1b(n142_O_5_0_0_t1b),
    .O_6_0_0_t0b(n142_O_6_0_0_t0b),
    .O_6_0_0_t1b(n142_O_6_0_0_t1b),
    .O_7_0_0_t0b(n142_O_7_0_0_t0b),
    .O_7_0_0_t1b(n142_O_7_0_0_t1b)
  );
  Map2T_9 n143 ( // @[Top.scala 346:22]
    .clock(n143_clock),
    .reset(n143_reset),
    .valid_up(n143_valid_up),
    .valid_down(n143_valid_down),
    .I0_0_0_0(n143_I0_0_0_0),
    .I0_0_0_1(n143_I0_0_0_1),
    .I0_0_0_2(n143_I0_0_0_2),
    .I0_0_1_0(n143_I0_0_1_0),
    .I0_0_1_1(n143_I0_0_1_1),
    .I0_0_1_2(n143_I0_0_1_2),
    .I0_0_2_0(n143_I0_0_2_0),
    .I0_0_2_1(n143_I0_0_2_1),
    .I0_0_2_2(n143_I0_0_2_2),
    .I0_1_0_0(n143_I0_1_0_0),
    .I0_1_0_1(n143_I0_1_0_1),
    .I0_1_0_2(n143_I0_1_0_2),
    .I0_1_1_0(n143_I0_1_1_0),
    .I0_1_1_1(n143_I0_1_1_1),
    .I0_1_1_2(n143_I0_1_1_2),
    .I0_1_2_0(n143_I0_1_2_0),
    .I0_1_2_1(n143_I0_1_2_1),
    .I0_1_2_2(n143_I0_1_2_2),
    .I0_2_0_0(n143_I0_2_0_0),
    .I0_2_0_1(n143_I0_2_0_1),
    .I0_2_0_2(n143_I0_2_0_2),
    .I0_2_1_0(n143_I0_2_1_0),
    .I0_2_1_1(n143_I0_2_1_1),
    .I0_2_1_2(n143_I0_2_1_2),
    .I0_2_2_0(n143_I0_2_2_0),
    .I0_2_2_1(n143_I0_2_2_1),
    .I0_2_2_2(n143_I0_2_2_2),
    .I0_3_0_0(n143_I0_3_0_0),
    .I0_3_0_1(n143_I0_3_0_1),
    .I0_3_0_2(n143_I0_3_0_2),
    .I0_3_1_0(n143_I0_3_1_0),
    .I0_3_1_1(n143_I0_3_1_1),
    .I0_3_1_2(n143_I0_3_1_2),
    .I0_3_2_0(n143_I0_3_2_0),
    .I0_3_2_1(n143_I0_3_2_1),
    .I0_3_2_2(n143_I0_3_2_2),
    .I0_4_0_0(n143_I0_4_0_0),
    .I0_4_0_1(n143_I0_4_0_1),
    .I0_4_0_2(n143_I0_4_0_2),
    .I0_4_1_0(n143_I0_4_1_0),
    .I0_4_1_1(n143_I0_4_1_1),
    .I0_4_1_2(n143_I0_4_1_2),
    .I0_4_2_0(n143_I0_4_2_0),
    .I0_4_2_1(n143_I0_4_2_1),
    .I0_4_2_2(n143_I0_4_2_2),
    .I0_5_0_0(n143_I0_5_0_0),
    .I0_5_0_1(n143_I0_5_0_1),
    .I0_5_0_2(n143_I0_5_0_2),
    .I0_5_1_0(n143_I0_5_1_0),
    .I0_5_1_1(n143_I0_5_1_1),
    .I0_5_1_2(n143_I0_5_1_2),
    .I0_5_2_0(n143_I0_5_2_0),
    .I0_5_2_1(n143_I0_5_2_1),
    .I0_5_2_2(n143_I0_5_2_2),
    .I0_6_0_0(n143_I0_6_0_0),
    .I0_6_0_1(n143_I0_6_0_1),
    .I0_6_0_2(n143_I0_6_0_2),
    .I0_6_1_0(n143_I0_6_1_0),
    .I0_6_1_1(n143_I0_6_1_1),
    .I0_6_1_2(n143_I0_6_1_2),
    .I0_6_2_0(n143_I0_6_2_0),
    .I0_6_2_1(n143_I0_6_2_1),
    .I0_6_2_2(n143_I0_6_2_2),
    .I0_7_0_0(n143_I0_7_0_0),
    .I0_7_0_1(n143_I0_7_0_1),
    .I0_7_0_2(n143_I0_7_0_2),
    .I0_7_1_0(n143_I0_7_1_0),
    .I0_7_1_1(n143_I0_7_1_1),
    .I0_7_1_2(n143_I0_7_1_2),
    .I0_7_2_0(n143_I0_7_2_0),
    .I0_7_2_1(n143_I0_7_2_1),
    .I0_7_2_2(n143_I0_7_2_2),
    .I1_0_0_0_t0b(n143_I1_0_0_0_t0b),
    .I1_0_0_0_t1b(n143_I1_0_0_0_t1b),
    .I1_1_0_0_t0b(n143_I1_1_0_0_t0b),
    .I1_1_0_0_t1b(n143_I1_1_0_0_t1b),
    .I1_2_0_0_t0b(n143_I1_2_0_0_t0b),
    .I1_2_0_0_t1b(n143_I1_2_0_0_t1b),
    .I1_3_0_0_t0b(n143_I1_3_0_0_t0b),
    .I1_3_0_0_t1b(n143_I1_3_0_0_t1b),
    .I1_4_0_0_t0b(n143_I1_4_0_0_t0b),
    .I1_4_0_0_t1b(n143_I1_4_0_0_t1b),
    .I1_5_0_0_t0b(n143_I1_5_0_0_t0b),
    .I1_5_0_0_t1b(n143_I1_5_0_0_t1b),
    .I1_6_0_0_t0b(n143_I1_6_0_0_t0b),
    .I1_6_0_0_t1b(n143_I1_6_0_0_t1b),
    .I1_7_0_0_t0b(n143_I1_7_0_0_t0b),
    .I1_7_0_0_t1b(n143_I1_7_0_0_t1b),
    .O_0_0_0_t0b(n143_O_0_0_0_t0b),
    .O_0_0_0_t1b_t0b(n143_O_0_0_0_t1b_t0b),
    .O_0_0_0_t1b_t1b(n143_O_0_0_0_t1b_t1b),
    .O_1_0_0_t0b(n143_O_1_0_0_t0b),
    .O_1_0_0_t1b_t0b(n143_O_1_0_0_t1b_t0b),
    .O_1_0_0_t1b_t1b(n143_O_1_0_0_t1b_t1b),
    .O_2_0_0_t0b(n143_O_2_0_0_t0b),
    .O_2_0_0_t1b_t0b(n143_O_2_0_0_t1b_t0b),
    .O_2_0_0_t1b_t1b(n143_O_2_0_0_t1b_t1b),
    .O_3_0_0_t0b(n143_O_3_0_0_t0b),
    .O_3_0_0_t1b_t0b(n143_O_3_0_0_t1b_t0b),
    .O_3_0_0_t1b_t1b(n143_O_3_0_0_t1b_t1b),
    .O_4_0_0_t0b(n143_O_4_0_0_t0b),
    .O_4_0_0_t1b_t0b(n143_O_4_0_0_t1b_t0b),
    .O_4_0_0_t1b_t1b(n143_O_4_0_0_t1b_t1b),
    .O_5_0_0_t0b(n143_O_5_0_0_t0b),
    .O_5_0_0_t1b_t0b(n143_O_5_0_0_t1b_t0b),
    .O_5_0_0_t1b_t1b(n143_O_5_0_0_t1b_t1b),
    .O_6_0_0_t0b(n143_O_6_0_0_t0b),
    .O_6_0_0_t1b_t0b(n143_O_6_0_0_t1b_t0b),
    .O_6_0_0_t1b_t1b(n143_O_6_0_0_t1b_t1b),
    .O_7_0_0_t0b(n143_O_7_0_0_t0b),
    .O_7_0_0_t1b_t0b(n143_O_7_0_0_t1b_t0b),
    .O_7_0_0_t1b_t1b(n143_O_7_0_0_t1b_t1b)
  );
  assign valid_down = n143_valid_down; // @[Top.scala 351:16]
  assign O_0_0_0_t0b = n143_O_0_0_0_t0b; // @[Top.scala 350:7]
  assign O_0_0_0_t1b_t0b = n143_O_0_0_0_t1b_t0b; // @[Top.scala 350:7]
  assign O_0_0_0_t1b_t1b = n143_O_0_0_0_t1b_t1b; // @[Top.scala 350:7]
  assign O_1_0_0_t0b = n143_O_1_0_0_t0b; // @[Top.scala 350:7]
  assign O_1_0_0_t1b_t0b = n143_O_1_0_0_t1b_t0b; // @[Top.scala 350:7]
  assign O_1_0_0_t1b_t1b = n143_O_1_0_0_t1b_t1b; // @[Top.scala 350:7]
  assign O_2_0_0_t0b = n143_O_2_0_0_t0b; // @[Top.scala 350:7]
  assign O_2_0_0_t1b_t0b = n143_O_2_0_0_t1b_t0b; // @[Top.scala 350:7]
  assign O_2_0_0_t1b_t1b = n143_O_2_0_0_t1b_t1b; // @[Top.scala 350:7]
  assign O_3_0_0_t0b = n143_O_3_0_0_t0b; // @[Top.scala 350:7]
  assign O_3_0_0_t1b_t0b = n143_O_3_0_0_t1b_t0b; // @[Top.scala 350:7]
  assign O_3_0_0_t1b_t1b = n143_O_3_0_0_t1b_t1b; // @[Top.scala 350:7]
  assign O_4_0_0_t0b = n143_O_4_0_0_t0b; // @[Top.scala 350:7]
  assign O_4_0_0_t1b_t0b = n143_O_4_0_0_t1b_t0b; // @[Top.scala 350:7]
  assign O_4_0_0_t1b_t1b = n143_O_4_0_0_t1b_t1b; // @[Top.scala 350:7]
  assign O_5_0_0_t0b = n143_O_5_0_0_t0b; // @[Top.scala 350:7]
  assign O_5_0_0_t1b_t0b = n143_O_5_0_0_t1b_t0b; // @[Top.scala 350:7]
  assign O_5_0_0_t1b_t1b = n143_O_5_0_0_t1b_t1b; // @[Top.scala 350:7]
  assign O_6_0_0_t0b = n143_O_6_0_0_t0b; // @[Top.scala 350:7]
  assign O_6_0_0_t1b_t0b = n143_O_6_0_0_t1b_t0b; // @[Top.scala 350:7]
  assign O_6_0_0_t1b_t1b = n143_O_6_0_0_t1b_t1b; // @[Top.scala 350:7]
  assign O_7_0_0_t0b = n143_O_7_0_0_t0b; // @[Top.scala 350:7]
  assign O_7_0_0_t1b_t0b = n143_O_7_0_0_t1b_t0b; // @[Top.scala 350:7]
  assign O_7_0_0_t1b_t1b = n143_O_7_0_0_t1b_t1b; // @[Top.scala 350:7]
  assign counter108_clock = clock;
  assign counter108_reset = reset;
  assign n116_I_0 = counter108_O_0; // @[Top.scala 328:12]
  assign n116_I_1 = counter108_O_1; // @[Top.scala 328:12]
  assign n116_I_2 = counter108_O_2; // @[Top.scala 328:12]
  assign n116_I_3 = counter108_O_3; // @[Top.scala 328:12]
  assign n116_I_4 = counter108_O_4; // @[Top.scala 328:12]
  assign n116_I_5 = counter108_O_5; // @[Top.scala 328:12]
  assign n116_I_6 = counter108_O_6; // @[Top.scala 328:12]
  assign n116_I_7 = counter108_O_7; // @[Top.scala 328:12]
  assign n128_I_0 = counter108_O_0; // @[Top.scala 331:12]
  assign n128_I_1 = counter108_O_1; // @[Top.scala 331:12]
  assign n128_I_2 = counter108_O_2; // @[Top.scala 331:12]
  assign n128_I_3 = counter108_O_3; // @[Top.scala 331:12]
  assign n128_I_4 = counter108_O_4; // @[Top.scala 331:12]
  assign n128_I_5 = counter108_O_5; // @[Top.scala 331:12]
  assign n128_I_6 = counter108_O_6; // @[Top.scala 331:12]
  assign n128_I_7 = counter108_O_7; // @[Top.scala 331:12]
  assign n129_valid_up = n116_valid_down & n128_valid_down; // @[Top.scala 336:19]
  assign n129_I0_0 = n116_O_0; // @[Top.scala 334:13]
  assign n129_I0_1 = n116_O_1; // @[Top.scala 334:13]
  assign n129_I0_2 = n116_O_2; // @[Top.scala 334:13]
  assign n129_I0_3 = n116_O_3; // @[Top.scala 334:13]
  assign n129_I0_4 = n116_O_4; // @[Top.scala 334:13]
  assign n129_I0_5 = n116_O_5; // @[Top.scala 334:13]
  assign n129_I0_6 = n116_O_6; // @[Top.scala 334:13]
  assign n129_I0_7 = n116_O_7; // @[Top.scala 334:13]
  assign n129_I1_0 = n128_O_0; // @[Top.scala 335:13]
  assign n129_I1_1 = n128_O_1; // @[Top.scala 335:13]
  assign n129_I1_2 = n128_O_2; // @[Top.scala 335:13]
  assign n129_I1_3 = n128_O_3; // @[Top.scala 335:13]
  assign n129_I1_4 = n128_O_4; // @[Top.scala 335:13]
  assign n129_I1_5 = n128_O_5; // @[Top.scala 335:13]
  assign n129_I1_6 = n128_O_6; // @[Top.scala 335:13]
  assign n129_I1_7 = n128_O_7; // @[Top.scala 335:13]
  assign n138_valid_up = n129_valid_down; // @[Top.scala 339:19]
  assign n138_I_0_t0b = n129_O_0_t0b; // @[Top.scala 338:12]
  assign n138_I_0_t1b = n129_O_0_t1b; // @[Top.scala 338:12]
  assign n138_I_1_t0b = n129_O_1_t0b; // @[Top.scala 338:12]
  assign n138_I_1_t1b = n129_O_1_t1b; // @[Top.scala 338:12]
  assign n138_I_2_t0b = n129_O_2_t0b; // @[Top.scala 338:12]
  assign n138_I_2_t1b = n129_O_2_t1b; // @[Top.scala 338:12]
  assign n138_I_3_t0b = n129_O_3_t0b; // @[Top.scala 338:12]
  assign n138_I_3_t1b = n129_O_3_t1b; // @[Top.scala 338:12]
  assign n138_I_4_t0b = n129_O_4_t0b; // @[Top.scala 338:12]
  assign n138_I_4_t1b = n129_O_4_t1b; // @[Top.scala 338:12]
  assign n138_I_5_t0b = n129_O_5_t0b; // @[Top.scala 338:12]
  assign n138_I_5_t1b = n129_O_5_t1b; // @[Top.scala 338:12]
  assign n138_I_6_t0b = n129_O_6_t0b; // @[Top.scala 338:12]
  assign n138_I_6_t1b = n129_O_6_t1b; // @[Top.scala 338:12]
  assign n138_I_7_t0b = n129_O_7_t0b; // @[Top.scala 338:12]
  assign n138_I_7_t1b = n129_O_7_t1b; // @[Top.scala 338:12]
  assign n141_valid_up = n138_valid_down; // @[Top.scala 342:19]
  assign n141_I_0_0_t0b = n138_O_0_0_t0b; // @[Top.scala 341:12]
  assign n141_I_0_0_t1b = n138_O_0_0_t1b; // @[Top.scala 341:12]
  assign n141_I_1_0_t0b = n138_O_1_0_t0b; // @[Top.scala 341:12]
  assign n141_I_1_0_t1b = n138_O_1_0_t1b; // @[Top.scala 341:12]
  assign n141_I_2_0_t0b = n138_O_2_0_t0b; // @[Top.scala 341:12]
  assign n141_I_2_0_t1b = n138_O_2_0_t1b; // @[Top.scala 341:12]
  assign n141_I_3_0_t0b = n138_O_3_0_t0b; // @[Top.scala 341:12]
  assign n141_I_3_0_t1b = n138_O_3_0_t1b; // @[Top.scala 341:12]
  assign n141_I_4_0_t0b = n138_O_4_0_t0b; // @[Top.scala 341:12]
  assign n141_I_4_0_t1b = n138_O_4_0_t1b; // @[Top.scala 341:12]
  assign n141_I_5_0_t0b = n138_O_5_0_t0b; // @[Top.scala 341:12]
  assign n141_I_5_0_t1b = n138_O_5_0_t1b; // @[Top.scala 341:12]
  assign n141_I_6_0_t0b = n138_O_6_0_t0b; // @[Top.scala 341:12]
  assign n141_I_6_0_t1b = n138_O_6_0_t1b; // @[Top.scala 341:12]
  assign n141_I_7_0_t0b = n138_O_7_0_t0b; // @[Top.scala 341:12]
  assign n141_I_7_0_t1b = n138_O_7_0_t1b; // @[Top.scala 341:12]
  assign n142_clock = clock;
  assign n142_reset = reset;
  assign n142_valid_up = n141_valid_down; // @[Top.scala 345:19]
  assign n142_I_0_0_0_t0b = n141_O_0_0_0_t0b; // @[Top.scala 344:12]
  assign n142_I_0_0_0_t1b = n141_O_0_0_0_t1b; // @[Top.scala 344:12]
  assign n142_I_1_0_0_t0b = n141_O_1_0_0_t0b; // @[Top.scala 344:12]
  assign n142_I_1_0_0_t1b = n141_O_1_0_0_t1b; // @[Top.scala 344:12]
  assign n142_I_2_0_0_t0b = n141_O_2_0_0_t0b; // @[Top.scala 344:12]
  assign n142_I_2_0_0_t1b = n141_O_2_0_0_t1b; // @[Top.scala 344:12]
  assign n142_I_3_0_0_t0b = n141_O_3_0_0_t0b; // @[Top.scala 344:12]
  assign n142_I_3_0_0_t1b = n141_O_3_0_0_t1b; // @[Top.scala 344:12]
  assign n142_I_4_0_0_t0b = n141_O_4_0_0_t0b; // @[Top.scala 344:12]
  assign n142_I_4_0_0_t1b = n141_O_4_0_0_t1b; // @[Top.scala 344:12]
  assign n142_I_5_0_0_t0b = n141_O_5_0_0_t0b; // @[Top.scala 344:12]
  assign n142_I_5_0_0_t1b = n141_O_5_0_0_t1b; // @[Top.scala 344:12]
  assign n142_I_6_0_0_t0b = n141_O_6_0_0_t0b; // @[Top.scala 344:12]
  assign n142_I_6_0_0_t1b = n141_O_6_0_0_t1b; // @[Top.scala 344:12]
  assign n142_I_7_0_0_t0b = n141_O_7_0_0_t0b; // @[Top.scala 344:12]
  assign n142_I_7_0_0_t1b = n141_O_7_0_0_t1b; // @[Top.scala 344:12]
  assign n143_clock = clock;
  assign n143_reset = reset;
  assign n143_valid_up = valid_up & n142_valid_down; // @[Top.scala 349:19]
  assign n143_I0_0_0_0 = I_0_0_0; // @[Top.scala 347:13]
  assign n143_I0_0_0_1 = I_0_0_1; // @[Top.scala 347:13]
  assign n143_I0_0_0_2 = I_0_0_2; // @[Top.scala 347:13]
  assign n143_I0_0_1_0 = I_0_1_0; // @[Top.scala 347:13]
  assign n143_I0_0_1_1 = I_0_1_1; // @[Top.scala 347:13]
  assign n143_I0_0_1_2 = I_0_1_2; // @[Top.scala 347:13]
  assign n143_I0_0_2_0 = I_0_2_0; // @[Top.scala 347:13]
  assign n143_I0_0_2_1 = I_0_2_1; // @[Top.scala 347:13]
  assign n143_I0_0_2_2 = I_0_2_2; // @[Top.scala 347:13]
  assign n143_I0_1_0_0 = I_1_0_0; // @[Top.scala 347:13]
  assign n143_I0_1_0_1 = I_1_0_1; // @[Top.scala 347:13]
  assign n143_I0_1_0_2 = I_1_0_2; // @[Top.scala 347:13]
  assign n143_I0_1_1_0 = I_1_1_0; // @[Top.scala 347:13]
  assign n143_I0_1_1_1 = I_1_1_1; // @[Top.scala 347:13]
  assign n143_I0_1_1_2 = I_1_1_2; // @[Top.scala 347:13]
  assign n143_I0_1_2_0 = I_1_2_0; // @[Top.scala 347:13]
  assign n143_I0_1_2_1 = I_1_2_1; // @[Top.scala 347:13]
  assign n143_I0_1_2_2 = I_1_2_2; // @[Top.scala 347:13]
  assign n143_I0_2_0_0 = I_2_0_0; // @[Top.scala 347:13]
  assign n143_I0_2_0_1 = I_2_0_1; // @[Top.scala 347:13]
  assign n143_I0_2_0_2 = I_2_0_2; // @[Top.scala 347:13]
  assign n143_I0_2_1_0 = I_2_1_0; // @[Top.scala 347:13]
  assign n143_I0_2_1_1 = I_2_1_1; // @[Top.scala 347:13]
  assign n143_I0_2_1_2 = I_2_1_2; // @[Top.scala 347:13]
  assign n143_I0_2_2_0 = I_2_2_0; // @[Top.scala 347:13]
  assign n143_I0_2_2_1 = I_2_2_1; // @[Top.scala 347:13]
  assign n143_I0_2_2_2 = I_2_2_2; // @[Top.scala 347:13]
  assign n143_I0_3_0_0 = I_3_0_0; // @[Top.scala 347:13]
  assign n143_I0_3_0_1 = I_3_0_1; // @[Top.scala 347:13]
  assign n143_I0_3_0_2 = I_3_0_2; // @[Top.scala 347:13]
  assign n143_I0_3_1_0 = I_3_1_0; // @[Top.scala 347:13]
  assign n143_I0_3_1_1 = I_3_1_1; // @[Top.scala 347:13]
  assign n143_I0_3_1_2 = I_3_1_2; // @[Top.scala 347:13]
  assign n143_I0_3_2_0 = I_3_2_0; // @[Top.scala 347:13]
  assign n143_I0_3_2_1 = I_3_2_1; // @[Top.scala 347:13]
  assign n143_I0_3_2_2 = I_3_2_2; // @[Top.scala 347:13]
  assign n143_I0_4_0_0 = I_4_0_0; // @[Top.scala 347:13]
  assign n143_I0_4_0_1 = I_4_0_1; // @[Top.scala 347:13]
  assign n143_I0_4_0_2 = I_4_0_2; // @[Top.scala 347:13]
  assign n143_I0_4_1_0 = I_4_1_0; // @[Top.scala 347:13]
  assign n143_I0_4_1_1 = I_4_1_1; // @[Top.scala 347:13]
  assign n143_I0_4_1_2 = I_4_1_2; // @[Top.scala 347:13]
  assign n143_I0_4_2_0 = I_4_2_0; // @[Top.scala 347:13]
  assign n143_I0_4_2_1 = I_4_2_1; // @[Top.scala 347:13]
  assign n143_I0_4_2_2 = I_4_2_2; // @[Top.scala 347:13]
  assign n143_I0_5_0_0 = I_5_0_0; // @[Top.scala 347:13]
  assign n143_I0_5_0_1 = I_5_0_1; // @[Top.scala 347:13]
  assign n143_I0_5_0_2 = I_5_0_2; // @[Top.scala 347:13]
  assign n143_I0_5_1_0 = I_5_1_0; // @[Top.scala 347:13]
  assign n143_I0_5_1_1 = I_5_1_1; // @[Top.scala 347:13]
  assign n143_I0_5_1_2 = I_5_1_2; // @[Top.scala 347:13]
  assign n143_I0_5_2_0 = I_5_2_0; // @[Top.scala 347:13]
  assign n143_I0_5_2_1 = I_5_2_1; // @[Top.scala 347:13]
  assign n143_I0_5_2_2 = I_5_2_2; // @[Top.scala 347:13]
  assign n143_I0_6_0_0 = I_6_0_0; // @[Top.scala 347:13]
  assign n143_I0_6_0_1 = I_6_0_1; // @[Top.scala 347:13]
  assign n143_I0_6_0_2 = I_6_0_2; // @[Top.scala 347:13]
  assign n143_I0_6_1_0 = I_6_1_0; // @[Top.scala 347:13]
  assign n143_I0_6_1_1 = I_6_1_1; // @[Top.scala 347:13]
  assign n143_I0_6_1_2 = I_6_1_2; // @[Top.scala 347:13]
  assign n143_I0_6_2_0 = I_6_2_0; // @[Top.scala 347:13]
  assign n143_I0_6_2_1 = I_6_2_1; // @[Top.scala 347:13]
  assign n143_I0_6_2_2 = I_6_2_2; // @[Top.scala 347:13]
  assign n143_I0_7_0_0 = I_7_0_0; // @[Top.scala 347:13]
  assign n143_I0_7_0_1 = I_7_0_1; // @[Top.scala 347:13]
  assign n143_I0_7_0_2 = I_7_0_2; // @[Top.scala 347:13]
  assign n143_I0_7_1_0 = I_7_1_0; // @[Top.scala 347:13]
  assign n143_I0_7_1_1 = I_7_1_1; // @[Top.scala 347:13]
  assign n143_I0_7_1_2 = I_7_1_2; // @[Top.scala 347:13]
  assign n143_I0_7_2_0 = I_7_2_0; // @[Top.scala 347:13]
  assign n143_I0_7_2_1 = I_7_2_1; // @[Top.scala 347:13]
  assign n143_I0_7_2_2 = I_7_2_2; // @[Top.scala 347:13]
  assign n143_I1_0_0_0_t0b = n142_O_0_0_0_t0b; // @[Top.scala 348:13]
  assign n143_I1_0_0_0_t1b = n142_O_0_0_0_t1b; // @[Top.scala 348:13]
  assign n143_I1_1_0_0_t0b = n142_O_1_0_0_t0b; // @[Top.scala 348:13]
  assign n143_I1_1_0_0_t1b = n142_O_1_0_0_t1b; // @[Top.scala 348:13]
  assign n143_I1_2_0_0_t0b = n142_O_2_0_0_t0b; // @[Top.scala 348:13]
  assign n143_I1_2_0_0_t1b = n142_O_2_0_0_t1b; // @[Top.scala 348:13]
  assign n143_I1_3_0_0_t0b = n142_O_3_0_0_t0b; // @[Top.scala 348:13]
  assign n143_I1_3_0_0_t1b = n142_O_3_0_0_t1b; // @[Top.scala 348:13]
  assign n143_I1_4_0_0_t0b = n142_O_4_0_0_t0b; // @[Top.scala 348:13]
  assign n143_I1_4_0_0_t1b = n142_O_4_0_0_t1b; // @[Top.scala 348:13]
  assign n143_I1_5_0_0_t0b = n142_O_5_0_0_t0b; // @[Top.scala 348:13]
  assign n143_I1_5_0_0_t1b = n142_O_5_0_0_t1b; // @[Top.scala 348:13]
  assign n143_I1_6_0_0_t0b = n142_O_6_0_0_t0b; // @[Top.scala 348:13]
  assign n143_I1_6_0_0_t1b = n142_O_6_0_0_t1b; // @[Top.scala 348:13]
  assign n143_I1_7_0_0_t0b = n142_O_7_0_0_t0b; // @[Top.scala 348:13]
  assign n143_I1_7_0_0_t1b = n142_O_7_0_0_t1b; // @[Top.scala 348:13]
endmodule
module MapT_12(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0_0,
  input  [31:0] I_0_0_1,
  input  [31:0] I_0_0_2,
  input  [31:0] I_0_1_0,
  input  [31:0] I_0_1_1,
  input  [31:0] I_0_1_2,
  input  [31:0] I_0_2_0,
  input  [31:0] I_0_2_1,
  input  [31:0] I_0_2_2,
  input  [31:0] I_1_0_0,
  input  [31:0] I_1_0_1,
  input  [31:0] I_1_0_2,
  input  [31:0] I_1_1_0,
  input  [31:0] I_1_1_1,
  input  [31:0] I_1_1_2,
  input  [31:0] I_1_2_0,
  input  [31:0] I_1_2_1,
  input  [31:0] I_1_2_2,
  input  [31:0] I_2_0_0,
  input  [31:0] I_2_0_1,
  input  [31:0] I_2_0_2,
  input  [31:0] I_2_1_0,
  input  [31:0] I_2_1_1,
  input  [31:0] I_2_1_2,
  input  [31:0] I_2_2_0,
  input  [31:0] I_2_2_1,
  input  [31:0] I_2_2_2,
  input  [31:0] I_3_0_0,
  input  [31:0] I_3_0_1,
  input  [31:0] I_3_0_2,
  input  [31:0] I_3_1_0,
  input  [31:0] I_3_1_1,
  input  [31:0] I_3_1_2,
  input  [31:0] I_3_2_0,
  input  [31:0] I_3_2_1,
  input  [31:0] I_3_2_2,
  input  [31:0] I_4_0_0,
  input  [31:0] I_4_0_1,
  input  [31:0] I_4_0_2,
  input  [31:0] I_4_1_0,
  input  [31:0] I_4_1_1,
  input  [31:0] I_4_1_2,
  input  [31:0] I_4_2_0,
  input  [31:0] I_4_2_1,
  input  [31:0] I_4_2_2,
  input  [31:0] I_5_0_0,
  input  [31:0] I_5_0_1,
  input  [31:0] I_5_0_2,
  input  [31:0] I_5_1_0,
  input  [31:0] I_5_1_1,
  input  [31:0] I_5_1_2,
  input  [31:0] I_5_2_0,
  input  [31:0] I_5_2_1,
  input  [31:0] I_5_2_2,
  input  [31:0] I_6_0_0,
  input  [31:0] I_6_0_1,
  input  [31:0] I_6_0_2,
  input  [31:0] I_6_1_0,
  input  [31:0] I_6_1_1,
  input  [31:0] I_6_1_2,
  input  [31:0] I_6_2_0,
  input  [31:0] I_6_2_1,
  input  [31:0] I_6_2_2,
  input  [31:0] I_7_0_0,
  input  [31:0] I_7_0_1,
  input  [31:0] I_7_0_2,
  input  [31:0] I_7_1_0,
  input  [31:0] I_7_1_1,
  input  [31:0] I_7_1_2,
  input  [31:0] I_7_2_0,
  input  [31:0] I_7_2_1,
  input  [31:0] I_7_2_2,
  output [31:0] O_0_0_0_t0b,
  output [31:0] O_0_0_0_t1b_t0b,
  output [31:0] O_0_0_0_t1b_t1b,
  output [31:0] O_1_0_0_t0b,
  output [31:0] O_1_0_0_t1b_t0b,
  output [31:0] O_1_0_0_t1b_t1b,
  output [31:0] O_2_0_0_t0b,
  output [31:0] O_2_0_0_t1b_t0b,
  output [31:0] O_2_0_0_t1b_t1b,
  output [31:0] O_3_0_0_t0b,
  output [31:0] O_3_0_0_t1b_t0b,
  output [31:0] O_3_0_0_t1b_t1b,
  output [31:0] O_4_0_0_t0b,
  output [31:0] O_4_0_0_t1b_t0b,
  output [31:0] O_4_0_0_t1b_t1b,
  output [31:0] O_5_0_0_t0b,
  output [31:0] O_5_0_0_t1b_t0b,
  output [31:0] O_5_0_0_t1b_t1b,
  output [31:0] O_6_0_0_t0b,
  output [31:0] O_6_0_0_t1b_t0b,
  output [31:0] O_6_0_0_t1b_t1b,
  output [31:0] O_7_0_0_t0b,
  output [31:0] O_7_0_0_t1b_t0b,
  output [31:0] O_7_0_0_t1b_t1b
);
  wire  op_clock; // @[MapT.scala 8:20]
  wire  op_reset; // @[MapT.scala 8:20]
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_0_0_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_0_0_t1b_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_0_0_t1b_t1b; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_0_0_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_0_0_t1b_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_0_0_t1b_t1b; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_0_0_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_0_0_t1b_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_0_0_t1b_t1b; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_0_0_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_0_0_t1b_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_0_0_t1b_t1b; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_0_0_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_0_0_t1b_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_0_0_t1b_t1b; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_0_0_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_0_0_t1b_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_0_0_t1b_t1b; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_0_0_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_0_0_t1b_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_0_0_t1b_t1b; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_0_0_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_0_0_t1b_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_0_0_t1b_t1b; // @[MapT.scala 8:20]
  Module_7 op ( // @[MapT.scala 8:20]
    .clock(op_clock),
    .reset(op_reset),
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0(op_I_0_0_0),
    .I_0_0_1(op_I_0_0_1),
    .I_0_0_2(op_I_0_0_2),
    .I_0_1_0(op_I_0_1_0),
    .I_0_1_1(op_I_0_1_1),
    .I_0_1_2(op_I_0_1_2),
    .I_0_2_0(op_I_0_2_0),
    .I_0_2_1(op_I_0_2_1),
    .I_0_2_2(op_I_0_2_2),
    .I_1_0_0(op_I_1_0_0),
    .I_1_0_1(op_I_1_0_1),
    .I_1_0_2(op_I_1_0_2),
    .I_1_1_0(op_I_1_1_0),
    .I_1_1_1(op_I_1_1_1),
    .I_1_1_2(op_I_1_1_2),
    .I_1_2_0(op_I_1_2_0),
    .I_1_2_1(op_I_1_2_1),
    .I_1_2_2(op_I_1_2_2),
    .I_2_0_0(op_I_2_0_0),
    .I_2_0_1(op_I_2_0_1),
    .I_2_0_2(op_I_2_0_2),
    .I_2_1_0(op_I_2_1_0),
    .I_2_1_1(op_I_2_1_1),
    .I_2_1_2(op_I_2_1_2),
    .I_2_2_0(op_I_2_2_0),
    .I_2_2_1(op_I_2_2_1),
    .I_2_2_2(op_I_2_2_2),
    .I_3_0_0(op_I_3_0_0),
    .I_3_0_1(op_I_3_0_1),
    .I_3_0_2(op_I_3_0_2),
    .I_3_1_0(op_I_3_1_0),
    .I_3_1_1(op_I_3_1_1),
    .I_3_1_2(op_I_3_1_2),
    .I_3_2_0(op_I_3_2_0),
    .I_3_2_1(op_I_3_2_1),
    .I_3_2_2(op_I_3_2_2),
    .I_4_0_0(op_I_4_0_0),
    .I_4_0_1(op_I_4_0_1),
    .I_4_0_2(op_I_4_0_2),
    .I_4_1_0(op_I_4_1_0),
    .I_4_1_1(op_I_4_1_1),
    .I_4_1_2(op_I_4_1_2),
    .I_4_2_0(op_I_4_2_0),
    .I_4_2_1(op_I_4_2_1),
    .I_4_2_2(op_I_4_2_2),
    .I_5_0_0(op_I_5_0_0),
    .I_5_0_1(op_I_5_0_1),
    .I_5_0_2(op_I_5_0_2),
    .I_5_1_0(op_I_5_1_0),
    .I_5_1_1(op_I_5_1_1),
    .I_5_1_2(op_I_5_1_2),
    .I_5_2_0(op_I_5_2_0),
    .I_5_2_1(op_I_5_2_1),
    .I_5_2_2(op_I_5_2_2),
    .I_6_0_0(op_I_6_0_0),
    .I_6_0_1(op_I_6_0_1),
    .I_6_0_2(op_I_6_0_2),
    .I_6_1_0(op_I_6_1_0),
    .I_6_1_1(op_I_6_1_1),
    .I_6_1_2(op_I_6_1_2),
    .I_6_2_0(op_I_6_2_0),
    .I_6_2_1(op_I_6_2_1),
    .I_6_2_2(op_I_6_2_2),
    .I_7_0_0(op_I_7_0_0),
    .I_7_0_1(op_I_7_0_1),
    .I_7_0_2(op_I_7_0_2),
    .I_7_1_0(op_I_7_1_0),
    .I_7_1_1(op_I_7_1_1),
    .I_7_1_2(op_I_7_1_2),
    .I_7_2_0(op_I_7_2_0),
    .I_7_2_1(op_I_7_2_1),
    .I_7_2_2(op_I_7_2_2),
    .O_0_0_0_t0b(op_O_0_0_0_t0b),
    .O_0_0_0_t1b_t0b(op_O_0_0_0_t1b_t0b),
    .O_0_0_0_t1b_t1b(op_O_0_0_0_t1b_t1b),
    .O_1_0_0_t0b(op_O_1_0_0_t0b),
    .O_1_0_0_t1b_t0b(op_O_1_0_0_t1b_t0b),
    .O_1_0_0_t1b_t1b(op_O_1_0_0_t1b_t1b),
    .O_2_0_0_t0b(op_O_2_0_0_t0b),
    .O_2_0_0_t1b_t0b(op_O_2_0_0_t1b_t0b),
    .O_2_0_0_t1b_t1b(op_O_2_0_0_t1b_t1b),
    .O_3_0_0_t0b(op_O_3_0_0_t0b),
    .O_3_0_0_t1b_t0b(op_O_3_0_0_t1b_t0b),
    .O_3_0_0_t1b_t1b(op_O_3_0_0_t1b_t1b),
    .O_4_0_0_t0b(op_O_4_0_0_t0b),
    .O_4_0_0_t1b_t0b(op_O_4_0_0_t1b_t0b),
    .O_4_0_0_t1b_t1b(op_O_4_0_0_t1b_t1b),
    .O_5_0_0_t0b(op_O_5_0_0_t0b),
    .O_5_0_0_t1b_t0b(op_O_5_0_0_t1b_t0b),
    .O_5_0_0_t1b_t1b(op_O_5_0_0_t1b_t1b),
    .O_6_0_0_t0b(op_O_6_0_0_t0b),
    .O_6_0_0_t1b_t0b(op_O_6_0_0_t1b_t0b),
    .O_6_0_0_t1b_t1b(op_O_6_0_0_t1b_t1b),
    .O_7_0_0_t0b(op_O_7_0_0_t0b),
    .O_7_0_0_t1b_t0b(op_O_7_0_0_t1b_t0b),
    .O_7_0_0_t1b_t1b(op_O_7_0_0_t1b_t1b)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0_t0b = op_O_0_0_0_t0b; // @[MapT.scala 15:7]
  assign O_0_0_0_t1b_t0b = op_O_0_0_0_t1b_t0b; // @[MapT.scala 15:7]
  assign O_0_0_0_t1b_t1b = op_O_0_0_0_t1b_t1b; // @[MapT.scala 15:7]
  assign O_1_0_0_t0b = op_O_1_0_0_t0b; // @[MapT.scala 15:7]
  assign O_1_0_0_t1b_t0b = op_O_1_0_0_t1b_t0b; // @[MapT.scala 15:7]
  assign O_1_0_0_t1b_t1b = op_O_1_0_0_t1b_t1b; // @[MapT.scala 15:7]
  assign O_2_0_0_t0b = op_O_2_0_0_t0b; // @[MapT.scala 15:7]
  assign O_2_0_0_t1b_t0b = op_O_2_0_0_t1b_t0b; // @[MapT.scala 15:7]
  assign O_2_0_0_t1b_t1b = op_O_2_0_0_t1b_t1b; // @[MapT.scala 15:7]
  assign O_3_0_0_t0b = op_O_3_0_0_t0b; // @[MapT.scala 15:7]
  assign O_3_0_0_t1b_t0b = op_O_3_0_0_t1b_t0b; // @[MapT.scala 15:7]
  assign O_3_0_0_t1b_t1b = op_O_3_0_0_t1b_t1b; // @[MapT.scala 15:7]
  assign O_4_0_0_t0b = op_O_4_0_0_t0b; // @[MapT.scala 15:7]
  assign O_4_0_0_t1b_t0b = op_O_4_0_0_t1b_t0b; // @[MapT.scala 15:7]
  assign O_4_0_0_t1b_t1b = op_O_4_0_0_t1b_t1b; // @[MapT.scala 15:7]
  assign O_5_0_0_t0b = op_O_5_0_0_t0b; // @[MapT.scala 15:7]
  assign O_5_0_0_t1b_t0b = op_O_5_0_0_t1b_t0b; // @[MapT.scala 15:7]
  assign O_5_0_0_t1b_t1b = op_O_5_0_0_t1b_t1b; // @[MapT.scala 15:7]
  assign O_6_0_0_t0b = op_O_6_0_0_t0b; // @[MapT.scala 15:7]
  assign O_6_0_0_t1b_t0b = op_O_6_0_0_t1b_t0b; // @[MapT.scala 15:7]
  assign O_6_0_0_t1b_t1b = op_O_6_0_0_t1b_t1b; // @[MapT.scala 15:7]
  assign O_7_0_0_t0b = op_O_7_0_0_t0b; // @[MapT.scala 15:7]
  assign O_7_0_0_t1b_t0b = op_O_7_0_0_t1b_t0b; // @[MapT.scala 15:7]
  assign O_7_0_0_t1b_t1b = op_O_7_0_0_t1b_t1b; // @[MapT.scala 15:7]
  assign op_clock = clock;
  assign op_reset = reset;
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0 = I_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_1 = I_0_0_1; // @[MapT.scala 14:10]
  assign op_I_0_0_2 = I_0_0_2; // @[MapT.scala 14:10]
  assign op_I_0_1_0 = I_0_1_0; // @[MapT.scala 14:10]
  assign op_I_0_1_1 = I_0_1_1; // @[MapT.scala 14:10]
  assign op_I_0_1_2 = I_0_1_2; // @[MapT.scala 14:10]
  assign op_I_0_2_0 = I_0_2_0; // @[MapT.scala 14:10]
  assign op_I_0_2_1 = I_0_2_1; // @[MapT.scala 14:10]
  assign op_I_0_2_2 = I_0_2_2; // @[MapT.scala 14:10]
  assign op_I_1_0_0 = I_1_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_1 = I_1_0_1; // @[MapT.scala 14:10]
  assign op_I_1_0_2 = I_1_0_2; // @[MapT.scala 14:10]
  assign op_I_1_1_0 = I_1_1_0; // @[MapT.scala 14:10]
  assign op_I_1_1_1 = I_1_1_1; // @[MapT.scala 14:10]
  assign op_I_1_1_2 = I_1_1_2; // @[MapT.scala 14:10]
  assign op_I_1_2_0 = I_1_2_0; // @[MapT.scala 14:10]
  assign op_I_1_2_1 = I_1_2_1; // @[MapT.scala 14:10]
  assign op_I_1_2_2 = I_1_2_2; // @[MapT.scala 14:10]
  assign op_I_2_0_0 = I_2_0_0; // @[MapT.scala 14:10]
  assign op_I_2_0_1 = I_2_0_1; // @[MapT.scala 14:10]
  assign op_I_2_0_2 = I_2_0_2; // @[MapT.scala 14:10]
  assign op_I_2_1_0 = I_2_1_0; // @[MapT.scala 14:10]
  assign op_I_2_1_1 = I_2_1_1; // @[MapT.scala 14:10]
  assign op_I_2_1_2 = I_2_1_2; // @[MapT.scala 14:10]
  assign op_I_2_2_0 = I_2_2_0; // @[MapT.scala 14:10]
  assign op_I_2_2_1 = I_2_2_1; // @[MapT.scala 14:10]
  assign op_I_2_2_2 = I_2_2_2; // @[MapT.scala 14:10]
  assign op_I_3_0_0 = I_3_0_0; // @[MapT.scala 14:10]
  assign op_I_3_0_1 = I_3_0_1; // @[MapT.scala 14:10]
  assign op_I_3_0_2 = I_3_0_2; // @[MapT.scala 14:10]
  assign op_I_3_1_0 = I_3_1_0; // @[MapT.scala 14:10]
  assign op_I_3_1_1 = I_3_1_1; // @[MapT.scala 14:10]
  assign op_I_3_1_2 = I_3_1_2; // @[MapT.scala 14:10]
  assign op_I_3_2_0 = I_3_2_0; // @[MapT.scala 14:10]
  assign op_I_3_2_1 = I_3_2_1; // @[MapT.scala 14:10]
  assign op_I_3_2_2 = I_3_2_2; // @[MapT.scala 14:10]
  assign op_I_4_0_0 = I_4_0_0; // @[MapT.scala 14:10]
  assign op_I_4_0_1 = I_4_0_1; // @[MapT.scala 14:10]
  assign op_I_4_0_2 = I_4_0_2; // @[MapT.scala 14:10]
  assign op_I_4_1_0 = I_4_1_0; // @[MapT.scala 14:10]
  assign op_I_4_1_1 = I_4_1_1; // @[MapT.scala 14:10]
  assign op_I_4_1_2 = I_4_1_2; // @[MapT.scala 14:10]
  assign op_I_4_2_0 = I_4_2_0; // @[MapT.scala 14:10]
  assign op_I_4_2_1 = I_4_2_1; // @[MapT.scala 14:10]
  assign op_I_4_2_2 = I_4_2_2; // @[MapT.scala 14:10]
  assign op_I_5_0_0 = I_5_0_0; // @[MapT.scala 14:10]
  assign op_I_5_0_1 = I_5_0_1; // @[MapT.scala 14:10]
  assign op_I_5_0_2 = I_5_0_2; // @[MapT.scala 14:10]
  assign op_I_5_1_0 = I_5_1_0; // @[MapT.scala 14:10]
  assign op_I_5_1_1 = I_5_1_1; // @[MapT.scala 14:10]
  assign op_I_5_1_2 = I_5_1_2; // @[MapT.scala 14:10]
  assign op_I_5_2_0 = I_5_2_0; // @[MapT.scala 14:10]
  assign op_I_5_2_1 = I_5_2_1; // @[MapT.scala 14:10]
  assign op_I_5_2_2 = I_5_2_2; // @[MapT.scala 14:10]
  assign op_I_6_0_0 = I_6_0_0; // @[MapT.scala 14:10]
  assign op_I_6_0_1 = I_6_0_1; // @[MapT.scala 14:10]
  assign op_I_6_0_2 = I_6_0_2; // @[MapT.scala 14:10]
  assign op_I_6_1_0 = I_6_1_0; // @[MapT.scala 14:10]
  assign op_I_6_1_1 = I_6_1_1; // @[MapT.scala 14:10]
  assign op_I_6_1_2 = I_6_1_2; // @[MapT.scala 14:10]
  assign op_I_6_2_0 = I_6_2_0; // @[MapT.scala 14:10]
  assign op_I_6_2_1 = I_6_2_1; // @[MapT.scala 14:10]
  assign op_I_6_2_2 = I_6_2_2; // @[MapT.scala 14:10]
  assign op_I_7_0_0 = I_7_0_0; // @[MapT.scala 14:10]
  assign op_I_7_0_1 = I_7_0_1; // @[MapT.scala 14:10]
  assign op_I_7_0_2 = I_7_0_2; // @[MapT.scala 14:10]
  assign op_I_7_1_0 = I_7_1_0; // @[MapT.scala 14:10]
  assign op_I_7_1_1 = I_7_1_1; // @[MapT.scala 14:10]
  assign op_I_7_1_2 = I_7_1_2; // @[MapT.scala 14:10]
  assign op_I_7_2_0 = I_7_2_0; // @[MapT.scala 14:10]
  assign op_I_7_2_1 = I_7_2_1; // @[MapT.scala 14:10]
  assign op_I_7_2_2 = I_7_2_2; // @[MapT.scala 14:10]
endmodule
module Passthrough_1(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0_0_t0b,
  input  [31:0] I_0_0_0_t1b_t0b,
  input  [31:0] I_0_0_0_t1b_t1b,
  input  [31:0] I_1_0_0_t0b,
  input  [31:0] I_1_0_0_t1b_t0b,
  input  [31:0] I_1_0_0_t1b_t1b,
  input  [31:0] I_2_0_0_t0b,
  input  [31:0] I_2_0_0_t1b_t0b,
  input  [31:0] I_2_0_0_t1b_t1b,
  input  [31:0] I_3_0_0_t0b,
  input  [31:0] I_3_0_0_t1b_t0b,
  input  [31:0] I_3_0_0_t1b_t1b,
  input  [31:0] I_4_0_0_t0b,
  input  [31:0] I_4_0_0_t1b_t0b,
  input  [31:0] I_4_0_0_t1b_t1b,
  input  [31:0] I_5_0_0_t0b,
  input  [31:0] I_5_0_0_t1b_t0b,
  input  [31:0] I_5_0_0_t1b_t1b,
  input  [31:0] I_6_0_0_t0b,
  input  [31:0] I_6_0_0_t1b_t0b,
  input  [31:0] I_6_0_0_t1b_t1b,
  input  [31:0] I_7_0_0_t0b,
  input  [31:0] I_7_0_0_t1b_t0b,
  input  [31:0] I_7_0_0_t1b_t1b,
  output [31:0] O_0_0_0_t0b,
  output [31:0] O_0_0_0_t1b_t0b,
  output [31:0] O_0_0_0_t1b_t1b,
  output [31:0] O_1_0_0_t0b,
  output [31:0] O_1_0_0_t1b_t0b,
  output [31:0] O_1_0_0_t1b_t1b,
  output [31:0] O_2_0_0_t0b,
  output [31:0] O_2_0_0_t1b_t0b,
  output [31:0] O_2_0_0_t1b_t1b,
  output [31:0] O_3_0_0_t0b,
  output [31:0] O_3_0_0_t1b_t0b,
  output [31:0] O_3_0_0_t1b_t1b,
  output [31:0] O_4_0_0_t0b,
  output [31:0] O_4_0_0_t1b_t0b,
  output [31:0] O_4_0_0_t1b_t1b,
  output [31:0] O_5_0_0_t0b,
  output [31:0] O_5_0_0_t1b_t0b,
  output [31:0] O_5_0_0_t1b_t1b,
  output [31:0] O_6_0_0_t0b,
  output [31:0] O_6_0_0_t1b_t0b,
  output [31:0] O_6_0_0_t1b_t1b,
  output [31:0] O_7_0_0_t0b,
  output [31:0] O_7_0_0_t1b_t0b,
  output [31:0] O_7_0_0_t1b_t1b
);
  assign valid_down = valid_up; // @[Passthrough.scala 18:14]
  assign O_0_0_0_t0b = I_0_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_0_0_0_t1b_t0b = I_0_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_0_0_0_t1b_t1b = I_0_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_1_0_0_t0b = I_1_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_1_0_0_t1b_t0b = I_1_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_1_0_0_t1b_t1b = I_1_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_2_0_0_t0b = I_2_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_2_0_0_t1b_t0b = I_2_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_2_0_0_t1b_t1b = I_2_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_3_0_0_t0b = I_3_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_3_0_0_t1b_t0b = I_3_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_3_0_0_t1b_t1b = I_3_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_4_0_0_t0b = I_4_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_4_0_0_t1b_t0b = I_4_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_4_0_0_t1b_t1b = I_4_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_5_0_0_t0b = I_5_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_5_0_0_t1b_t0b = I_5_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_5_0_0_t1b_t1b = I_5_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_6_0_0_t0b = I_6_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_6_0_0_t1b_t0b = I_6_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_6_0_0_t1b_t1b = I_6_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_7_0_0_t0b = I_7_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_7_0_0_t1b_t0b = I_7_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_7_0_0_t1b_t1b = I_7_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
endmodule
module Passthrough_2(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0_0_t0b,
  input  [31:0] I_0_0_0_t1b_t0b,
  input  [31:0] I_0_0_0_t1b_t1b,
  input  [31:0] I_1_0_0_t0b,
  input  [31:0] I_1_0_0_t1b_t0b,
  input  [31:0] I_1_0_0_t1b_t1b,
  input  [31:0] I_2_0_0_t0b,
  input  [31:0] I_2_0_0_t1b_t0b,
  input  [31:0] I_2_0_0_t1b_t1b,
  input  [31:0] I_3_0_0_t0b,
  input  [31:0] I_3_0_0_t1b_t0b,
  input  [31:0] I_3_0_0_t1b_t1b,
  input  [31:0] I_4_0_0_t0b,
  input  [31:0] I_4_0_0_t1b_t0b,
  input  [31:0] I_4_0_0_t1b_t1b,
  input  [31:0] I_5_0_0_t0b,
  input  [31:0] I_5_0_0_t1b_t0b,
  input  [31:0] I_5_0_0_t1b_t1b,
  input  [31:0] I_6_0_0_t0b,
  input  [31:0] I_6_0_0_t1b_t0b,
  input  [31:0] I_6_0_0_t1b_t1b,
  input  [31:0] I_7_0_0_t0b,
  input  [31:0] I_7_0_0_t1b_t0b,
  input  [31:0] I_7_0_0_t1b_t1b,
  output [31:0] O_0_0_t0b,
  output [31:0] O_0_0_t1b_t0b,
  output [31:0] O_0_0_t1b_t1b,
  output [31:0] O_1_0_t0b,
  output [31:0] O_1_0_t1b_t0b,
  output [31:0] O_1_0_t1b_t1b,
  output [31:0] O_2_0_t0b,
  output [31:0] O_2_0_t1b_t0b,
  output [31:0] O_2_0_t1b_t1b,
  output [31:0] O_3_0_t0b,
  output [31:0] O_3_0_t1b_t0b,
  output [31:0] O_3_0_t1b_t1b,
  output [31:0] O_4_0_t0b,
  output [31:0] O_4_0_t1b_t0b,
  output [31:0] O_4_0_t1b_t1b,
  output [31:0] O_5_0_t0b,
  output [31:0] O_5_0_t1b_t0b,
  output [31:0] O_5_0_t1b_t1b,
  output [31:0] O_6_0_t0b,
  output [31:0] O_6_0_t1b_t0b,
  output [31:0] O_6_0_t1b_t1b,
  output [31:0] O_7_0_t0b,
  output [31:0] O_7_0_t1b_t0b,
  output [31:0] O_7_0_t1b_t1b
);
  assign valid_down = valid_up; // @[Passthrough.scala 18:14]
  assign O_0_0_t0b = I_0_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_0_0_t1b_t0b = I_0_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_0_0_t1b_t1b = I_0_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_1_0_t0b = I_1_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_1_0_t1b_t0b = I_1_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_1_0_t1b_t1b = I_1_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_2_0_t0b = I_2_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_2_0_t1b_t0b = I_2_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_2_0_t1b_t1b = I_2_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_3_0_t0b = I_3_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_3_0_t1b_t0b = I_3_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_3_0_t1b_t1b = I_3_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_4_0_t0b = I_4_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_4_0_t1b_t0b = I_4_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_4_0_t1b_t1b = I_4_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_5_0_t0b = I_5_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_5_0_t1b_t0b = I_5_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_5_0_t1b_t1b = I_5_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_6_0_t0b = I_6_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_6_0_t1b_t0b = I_6_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_6_0_t1b_t1b = I_6_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_7_0_t0b = I_7_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_7_0_t1b_t0b = I_7_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_7_0_t1b_t1b = I_7_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
endmodule
module Passthrough_3(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0_t0b,
  input  [31:0] I_0_0_t1b_t0b,
  input  [31:0] I_0_0_t1b_t1b,
  input  [31:0] I_1_0_t0b,
  input  [31:0] I_1_0_t1b_t0b,
  input  [31:0] I_1_0_t1b_t1b,
  input  [31:0] I_2_0_t0b,
  input  [31:0] I_2_0_t1b_t0b,
  input  [31:0] I_2_0_t1b_t1b,
  input  [31:0] I_3_0_t0b,
  input  [31:0] I_3_0_t1b_t0b,
  input  [31:0] I_3_0_t1b_t1b,
  input  [31:0] I_4_0_t0b,
  input  [31:0] I_4_0_t1b_t0b,
  input  [31:0] I_4_0_t1b_t1b,
  input  [31:0] I_5_0_t0b,
  input  [31:0] I_5_0_t1b_t0b,
  input  [31:0] I_5_0_t1b_t1b,
  input  [31:0] I_6_0_t0b,
  input  [31:0] I_6_0_t1b_t0b,
  input  [31:0] I_6_0_t1b_t1b,
  input  [31:0] I_7_0_t0b,
  input  [31:0] I_7_0_t1b_t0b,
  input  [31:0] I_7_0_t1b_t1b,
  output [31:0] O_0_t0b,
  output [31:0] O_0_t1b_t0b,
  output [31:0] O_0_t1b_t1b,
  output [31:0] O_1_t0b,
  output [31:0] O_1_t1b_t0b,
  output [31:0] O_1_t1b_t1b,
  output [31:0] O_2_t0b,
  output [31:0] O_2_t1b_t0b,
  output [31:0] O_2_t1b_t1b,
  output [31:0] O_3_t0b,
  output [31:0] O_3_t1b_t0b,
  output [31:0] O_3_t1b_t1b,
  output [31:0] O_4_t0b,
  output [31:0] O_4_t1b_t0b,
  output [31:0] O_4_t1b_t1b,
  output [31:0] O_5_t0b,
  output [31:0] O_5_t1b_t0b,
  output [31:0] O_5_t1b_t1b,
  output [31:0] O_6_t0b,
  output [31:0] O_6_t1b_t0b,
  output [31:0] O_6_t1b_t1b,
  output [31:0] O_7_t0b,
  output [31:0] O_7_t1b_t0b,
  output [31:0] O_7_t1b_t1b
);
  assign valid_down = valid_up; // @[Passthrough.scala 18:14]
  assign O_0_t0b = I_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_0_t1b_t0b = I_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_0_t1b_t1b = I_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_1_t0b = I_1_0_t0b; // @[Passthrough.scala 17:68]
  assign O_1_t1b_t0b = I_1_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_1_t1b_t1b = I_1_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_2_t0b = I_2_0_t0b; // @[Passthrough.scala 17:68]
  assign O_2_t1b_t0b = I_2_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_2_t1b_t1b = I_2_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_3_t0b = I_3_0_t0b; // @[Passthrough.scala 17:68]
  assign O_3_t1b_t0b = I_3_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_3_t1b_t1b = I_3_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_4_t0b = I_4_0_t0b; // @[Passthrough.scala 17:68]
  assign O_4_t1b_t0b = I_4_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_4_t1b_t1b = I_4_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_5_t0b = I_5_0_t0b; // @[Passthrough.scala 17:68]
  assign O_5_t1b_t0b = I_5_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_5_t1b_t1b = I_5_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_6_t0b = I_6_0_t0b; // @[Passthrough.scala 17:68]
  assign O_6_t1b_t0b = I_6_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_6_t1b_t1b = I_6_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_7_t0b = I_7_0_t0b; // @[Passthrough.scala 17:68]
  assign O_7_t1b_t0b = I_7_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_7_t1b_t1b = I_7_0_t1b_t1b; // @[Passthrough.scala 17:68]
endmodule
module Fst_1(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_t0b,
  output [31:0] O
);
  assign valid_down = valid_up; // @[Tuple.scala 59:14]
  assign O = I_t0b; // @[Tuple.scala 58:5]
endmodule
module MapS_49(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_t0b,
  input  [31:0] I_1_t0b,
  input  [31:0] I_2_t0b,
  input  [31:0] I_3_t0b,
  input  [31:0] I_4_t0b,
  input  [31:0] I_5_t0b,
  input  [31:0] I_6_t0b,
  input  [31:0] I_7_t0b,
  output [31:0] O_0,
  output [31:0] O_1,
  output [31:0] O_2,
  output [31:0] O_3,
  output [31:0] O_4,
  output [31:0] O_5,
  output [31:0] O_6,
  output [31:0] O_7
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_t0b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_t0b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_O; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_t0b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_O; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_t0b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_O; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_t0b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_O; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_t0b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_O; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_t0b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_O; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_t0b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_O; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  wire  _T_1; // @[MapS.scala 23:83]
  wire  _T_2; // @[MapS.scala 23:83]
  wire  _T_3; // @[MapS.scala 23:83]
  wire  _T_4; // @[MapS.scala 23:83]
  wire  _T_5; // @[MapS.scala 23:83]
  Fst_1 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_t0b(fst_op_I_t0b),
    .O(fst_op_O)
  );
  Fst_1 other_ops_0 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_t0b(other_ops_0_I_t0b),
    .O(other_ops_0_O)
  );
  Fst_1 other_ops_1 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_t0b(other_ops_1_I_t0b),
    .O(other_ops_1_O)
  );
  Fst_1 other_ops_2 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I_t0b(other_ops_2_I_t0b),
    .O(other_ops_2_O)
  );
  Fst_1 other_ops_3 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I_t0b(other_ops_3_I_t0b),
    .O(other_ops_3_O)
  );
  Fst_1 other_ops_4 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I_t0b(other_ops_4_I_t0b),
    .O(other_ops_4_O)
  );
  Fst_1 other_ops_5 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I_t0b(other_ops_5_I_t0b),
    .O(other_ops_5_O)
  );
  Fst_1 other_ops_6 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I_t0b(other_ops_6_I_t0b),
    .O(other_ops_6_O)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[MapS.scala 23:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[MapS.scala 23:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[MapS.scala 23:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[MapS.scala 23:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T_5 & other_ops_6_valid_down; // @[MapS.scala 23:14]
  assign O_0 = fst_op_O; // @[MapS.scala 17:8]
  assign O_1 = other_ops_0_O; // @[MapS.scala 21:12]
  assign O_2 = other_ops_1_O; // @[MapS.scala 21:12]
  assign O_3 = other_ops_2_O; // @[MapS.scala 21:12]
  assign O_4 = other_ops_3_O; // @[MapS.scala 21:12]
  assign O_5 = other_ops_4_O; // @[MapS.scala 21:12]
  assign O_6 = other_ops_5_O; // @[MapS.scala 21:12]
  assign O_7 = other_ops_6_O; // @[MapS.scala 21:12]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_t0b = I_0_t0b; // @[MapS.scala 16:12]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_t0b = I_1_t0b; // @[MapS.scala 20:41]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_t0b = I_2_t0b; // @[MapS.scala 20:41]
  assign other_ops_2_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_2_I_t0b = I_3_t0b; // @[MapS.scala 20:41]
  assign other_ops_3_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_3_I_t0b = I_4_t0b; // @[MapS.scala 20:41]
  assign other_ops_4_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_4_I_t0b = I_5_t0b; // @[MapS.scala 20:41]
  assign other_ops_5_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_5_I_t0b = I_6_t0b; // @[MapS.scala 20:41]
  assign other_ops_6_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_6_I_t0b = I_7_t0b; // @[MapS.scala 20:41]
endmodule
module MapT_13(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_t0b,
  input  [31:0] I_1_t0b,
  input  [31:0] I_2_t0b,
  input  [31:0] I_3_t0b,
  input  [31:0] I_4_t0b,
  input  [31:0] I_5_t0b,
  input  [31:0] I_6_t0b,
  input  [31:0] I_7_t0b,
  output [31:0] O_0,
  output [31:0] O_1,
  output [31:0] O_2,
  output [31:0] O_3,
  output [31:0] O_4,
  output [31:0] O_5,
  output [31:0] O_6,
  output [31:0] O_7
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_3; // @[MapT.scala 8:20]
  wire [31:0] op_O_4; // @[MapT.scala 8:20]
  wire [31:0] op_O_5; // @[MapT.scala 8:20]
  wire [31:0] op_O_6; // @[MapT.scala 8:20]
  wire [31:0] op_O_7; // @[MapT.scala 8:20]
  MapS_49 op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_t0b(op_I_0_t0b),
    .I_1_t0b(op_I_1_t0b),
    .I_2_t0b(op_I_2_t0b),
    .I_3_t0b(op_I_3_t0b),
    .I_4_t0b(op_I_4_t0b),
    .I_5_t0b(op_I_5_t0b),
    .I_6_t0b(op_I_6_t0b),
    .I_7_t0b(op_I_7_t0b),
    .O_0(op_O_0),
    .O_1(op_O_1),
    .O_2(op_O_2),
    .O_3(op_O_3),
    .O_4(op_O_4),
    .O_5(op_O_5),
    .O_6(op_O_6),
    .O_7(op_O_7)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0 = op_O_0; // @[MapT.scala 15:7]
  assign O_1 = op_O_1; // @[MapT.scala 15:7]
  assign O_2 = op_O_2; // @[MapT.scala 15:7]
  assign O_3 = op_O_3; // @[MapT.scala 15:7]
  assign O_4 = op_O_4; // @[MapT.scala 15:7]
  assign O_5 = op_O_5; // @[MapT.scala 15:7]
  assign O_6 = op_O_6; // @[MapT.scala 15:7]
  assign O_7 = op_O_7; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_t0b = I_0_t0b; // @[MapT.scala 14:10]
  assign op_I_1_t0b = I_1_t0b; // @[MapT.scala 14:10]
  assign op_I_2_t0b = I_2_t0b; // @[MapT.scala 14:10]
  assign op_I_3_t0b = I_3_t0b; // @[MapT.scala 14:10]
  assign op_I_4_t0b = I_4_t0b; // @[MapT.scala 14:10]
  assign op_I_5_t0b = I_5_t0b; // @[MapT.scala 14:10]
  assign op_I_6_t0b = I_6_t0b; // @[MapT.scala 14:10]
  assign op_I_7_t0b = I_7_t0b; // @[MapT.scala 14:10]
endmodule
module Map2S_62(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0,
  input  [31:0] I0_1,
  input  [31:0] I0_2,
  input  [31:0] I1_0,
  input  [31:0] I1_1,
  input  [31:0] I1_2,
  output [31:0] O_0_t0b,
  output [31:0] O_0_t1b,
  output [31:0] O_1_t0b,
  output [31:0] O_1_t1b,
  output [31:0] O_2_t0b,
  output [31:0] O_2_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_t1b; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_t1b; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  AtomTuple fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1(fst_op_I1),
    .O_t0b(fst_op_O_t0b),
    .O_t1b(fst_op_O_t1b)
  );
  AtomTuple other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0(other_ops_0_I0),
    .I1(other_ops_0_I1),
    .O_t0b(other_ops_0_O_t0b),
    .O_t1b(other_ops_0_O_t1b)
  );
  AtomTuple other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0(other_ops_1_I0),
    .I1(other_ops_1_I1),
    .O_t0b(other_ops_1_O_t0b),
    .O_t1b(other_ops_1_O_t1b)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[Map2S.scala 26:14]
  assign O_0_t0b = fst_op_O_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b = fst_op_O_t1b; // @[Map2S.scala 19:8]
  assign O_1_t0b = other_ops_0_O_t0b; // @[Map2S.scala 24:12]
  assign O_1_t1b = other_ops_0_O_t1b; // @[Map2S.scala 24:12]
  assign O_2_t0b = other_ops_1_O_t0b; // @[Map2S.scala 24:12]
  assign O_2_t1b = other_ops_1_O_t1b; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0 = I0_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I1 = I1_1; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0 = I0_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1 = I1_2; // @[Map2S.scala 23:43]
endmodule
module Map2S_63(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0_0,
  input  [31:0] I0_0_1,
  input  [31:0] I0_0_2,
  input  [31:0] I0_1_0,
  input  [31:0] I0_1_1,
  input  [31:0] I0_1_2,
  input  [31:0] I0_2_0,
  input  [31:0] I0_2_1,
  input  [31:0] I0_2_2,
  output [31:0] O_0_0_t0b,
  output [31:0] O_0_0_t1b,
  output [31:0] O_0_1_t0b,
  output [31:0] O_0_1_t1b,
  output [31:0] O_0_2_t0b,
  output [31:0] O_0_2_t1b,
  output [31:0] O_1_0_t0b,
  output [31:0] O_1_0_t1b,
  output [31:0] O_1_1_t0b,
  output [31:0] O_1_1_t1b,
  output [31:0] O_1_2_t0b,
  output [31:0] O_1_2_t1b,
  output [31:0] O_2_0_t0b,
  output [31:0] O_2_0_t1b,
  output [31:0] O_2_1_t0b,
  output [31:0] O_2_1_t1b,
  output [31:0] O_2_2_t0b,
  output [31:0] O_2_2_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_2; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_2; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_t1b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_1_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_1_t1b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_2_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_2_t1b; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_0_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_0_t1b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_1_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_1_t1b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_2_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_2_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_0_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_0_t1b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_1_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_1_t1b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_2_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_2_t1b; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  Map2S_62 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I0_1(fst_op_I0_1),
    .I0_2(fst_op_I0_2),
    .I1_0(fst_op_I1_0),
    .I1_1(fst_op_I1_1),
    .I1_2(fst_op_I1_2),
    .O_0_t0b(fst_op_O_0_t0b),
    .O_0_t1b(fst_op_O_0_t1b),
    .O_1_t0b(fst_op_O_1_t0b),
    .O_1_t1b(fst_op_O_1_t1b),
    .O_2_t0b(fst_op_O_2_t0b),
    .O_2_t1b(fst_op_O_2_t1b)
  );
  Map2S_62 other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0(other_ops_0_I0_0),
    .I0_1(other_ops_0_I0_1),
    .I0_2(other_ops_0_I0_2),
    .I1_0(other_ops_0_I1_0),
    .I1_1(other_ops_0_I1_1),
    .I1_2(other_ops_0_I1_2),
    .O_0_t0b(other_ops_0_O_0_t0b),
    .O_0_t1b(other_ops_0_O_0_t1b),
    .O_1_t0b(other_ops_0_O_1_t0b),
    .O_1_t1b(other_ops_0_O_1_t1b),
    .O_2_t0b(other_ops_0_O_2_t0b),
    .O_2_t1b(other_ops_0_O_2_t1b)
  );
  Map2S_62 other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0_0(other_ops_1_I0_0),
    .I0_1(other_ops_1_I0_1),
    .I0_2(other_ops_1_I0_2),
    .I1_0(other_ops_1_I1_0),
    .I1_1(other_ops_1_I1_1),
    .I1_2(other_ops_1_I1_2),
    .O_0_t0b(other_ops_1_O_0_t0b),
    .O_0_t1b(other_ops_1_O_0_t1b),
    .O_1_t0b(other_ops_1_O_1_t0b),
    .O_1_t1b(other_ops_1_O_1_t1b),
    .O_2_t0b(other_ops_1_O_2_t0b),
    .O_2_t1b(other_ops_1_O_2_t1b)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_t0b = fst_op_O_0_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_t1b = fst_op_O_0_t1b; // @[Map2S.scala 19:8]
  assign O_0_1_t0b = fst_op_O_1_t0b; // @[Map2S.scala 19:8]
  assign O_0_1_t1b = fst_op_O_1_t1b; // @[Map2S.scala 19:8]
  assign O_0_2_t0b = fst_op_O_2_t0b; // @[Map2S.scala 19:8]
  assign O_0_2_t1b = fst_op_O_2_t1b; // @[Map2S.scala 19:8]
  assign O_1_0_t0b = other_ops_0_O_0_t0b; // @[Map2S.scala 24:12]
  assign O_1_0_t1b = other_ops_0_O_0_t1b; // @[Map2S.scala 24:12]
  assign O_1_1_t0b = other_ops_0_O_1_t0b; // @[Map2S.scala 24:12]
  assign O_1_1_t1b = other_ops_0_O_1_t1b; // @[Map2S.scala 24:12]
  assign O_1_2_t0b = other_ops_0_O_2_t0b; // @[Map2S.scala 24:12]
  assign O_1_2_t1b = other_ops_0_O_2_t1b; // @[Map2S.scala 24:12]
  assign O_2_0_t0b = other_ops_1_O_0_t0b; // @[Map2S.scala 24:12]
  assign O_2_0_t1b = other_ops_1_O_0_t1b; // @[Map2S.scala 24:12]
  assign O_2_1_t0b = other_ops_1_O_1_t0b; // @[Map2S.scala 24:12]
  assign O_2_1_t1b = other_ops_1_O_1_t1b; // @[Map2S.scala 24:12]
  assign O_2_2_t0b = other_ops_1_O_2_t0b; // @[Map2S.scala 24:12]
  assign O_2_2_t1b = other_ops_1_O_2_t1b; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1 = I0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_2 = I0_0_2; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = 32'h1; // @[Map2S.scala 18:13]
  assign fst_op_I1_1 = 32'h2; // @[Map2S.scala 18:13]
  assign fst_op_I1_2 = 32'h1; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0 = I0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1 = I0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_2 = I0_1_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I1_0 = 32'h2; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_1 = 32'h4; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_2 = 32'h2; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0_0 = I0_2_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1 = I0_2_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_2 = I0_2_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1_0 = 32'h1; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_1 = 32'h2; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_2 = 32'h1; // @[Map2S.scala 23:43]
endmodule
module Mul(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_t0b,
  input  [31:0] I_t1b,
  output [31:0] O
);
  wire [31:0] BlackBoxMulUInt32_I0; // @[Arithmetic.scala 195:27]
  wire [31:0] BlackBoxMulUInt32_I1; // @[Arithmetic.scala 195:27]
  wire [63:0] BlackBoxMulUInt32_O; // @[Arithmetic.scala 195:27]
  wire  BlackBoxMulUInt32_clock; // @[Arithmetic.scala 195:27]
  reg  _T_1; // @[Arithmetic.scala 214:66]
  reg [31:0] _RAND_0;
  reg  _T_2; // @[Arithmetic.scala 214:58]
  reg [31:0] _RAND_1;
  reg  _T_3; // @[Arithmetic.scala 214:50]
  reg [31:0] _RAND_2;
  reg  _T_4; // @[Arithmetic.scala 214:42]
  reg [31:0] _RAND_3;
  reg  _T_5; // @[Arithmetic.scala 214:34]
  reg [31:0] _RAND_4;
  reg  _T_6; // @[Arithmetic.scala 214:26]
  reg [31:0] _RAND_5;
  BlackBoxMulUInt32 BlackBoxMulUInt32 ( // @[Arithmetic.scala 195:27]
    .I0(BlackBoxMulUInt32_I0),
    .I1(BlackBoxMulUInt32_I1),
    .O(BlackBoxMulUInt32_O),
    .clock(BlackBoxMulUInt32_clock)
  );
  assign valid_down = _T_6; // @[Arithmetic.scala 214:16]
  assign O = BlackBoxMulUInt32_O[31:0]; // @[Arithmetic.scala 198:7]
  assign BlackBoxMulUInt32_I0 = I_t0b; // @[Arithmetic.scala 196:21]
  assign BlackBoxMulUInt32_I1 = I_t1b; // @[Arithmetic.scala 197:21]
  assign BlackBoxMulUInt32_clock = clock; // @[Arithmetic.scala 199:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_2 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_3 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_4 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_5 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_6 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      _T_1 <= valid_up;
    end
    if (reset) begin
      _T_2 <= 1'h0;
    end else begin
      _T_2 <= _T_1;
    end
    if (reset) begin
      _T_3 <= 1'h0;
    end else begin
      _T_3 <= _T_2;
    end
    _T_4 <= _T_3;
    _T_5 <= _T_4;
    _T_6 <= _T_5;
  end
endmodule
module MapS_54(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_t0b,
  input  [31:0] I_0_t1b,
  input  [31:0] I_1_t0b,
  input  [31:0] I_1_t1b,
  input  [31:0] I_2_t0b,
  input  [31:0] I_2_t1b,
  output [31:0] O_0,
  output [31:0] O_1,
  output [31:0] O_2
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_t0b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_t1b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O; // @[MapS.scala 9:22]
  wire  other_ops_0_clock; // @[MapS.scala 10:86]
  wire  other_ops_0_reset; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_t0b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_t1b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_O; // @[MapS.scala 10:86]
  wire  other_ops_1_clock; // @[MapS.scala 10:86]
  wire  other_ops_1_reset; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_t0b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_t1b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_O; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  Mul fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_t0b(fst_op_I_t0b),
    .I_t1b(fst_op_I_t1b),
    .O(fst_op_O)
  );
  Mul other_ops_0 ( // @[MapS.scala 10:86]
    .clock(other_ops_0_clock),
    .reset(other_ops_0_reset),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_t0b(other_ops_0_I_t0b),
    .I_t1b(other_ops_0_I_t1b),
    .O(other_ops_0_O)
  );
  Mul other_ops_1 ( // @[MapS.scala 10:86]
    .clock(other_ops_1_clock),
    .reset(other_ops_1_reset),
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_t0b(other_ops_1_I_t0b),
    .I_t1b(other_ops_1_I_t1b),
    .O(other_ops_1_O)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[MapS.scala 23:14]
  assign O_0 = fst_op_O; // @[MapS.scala 17:8]
  assign O_1 = other_ops_0_O; // @[MapS.scala 21:12]
  assign O_2 = other_ops_1_O; // @[MapS.scala 21:12]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_t0b = I_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_t1b = I_0_t1b; // @[MapS.scala 16:12]
  assign other_ops_0_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_0_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_t0b = I_1_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_t1b = I_1_t1b; // @[MapS.scala 20:41]
  assign other_ops_1_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_1_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_t0b = I_2_t0b; // @[MapS.scala 20:41]
  assign other_ops_1_I_t1b = I_2_t1b; // @[MapS.scala 20:41]
endmodule
module MapS_55(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0_t0b,
  input  [31:0] I_0_0_t1b,
  input  [31:0] I_0_1_t0b,
  input  [31:0] I_0_1_t1b,
  input  [31:0] I_0_2_t0b,
  input  [31:0] I_0_2_t1b,
  input  [31:0] I_1_0_t0b,
  input  [31:0] I_1_0_t1b,
  input  [31:0] I_1_1_t0b,
  input  [31:0] I_1_1_t1b,
  input  [31:0] I_1_2_t0b,
  input  [31:0] I_1_2_t1b,
  input  [31:0] I_2_0_t0b,
  input  [31:0] I_2_0_t1b,
  input  [31:0] I_2_1_t0b,
  input  [31:0] I_2_1_t1b,
  input  [31:0] I_2_2_t0b,
  input  [31:0] I_2_2_t1b,
  output [31:0] O_0_0,
  output [31:0] O_0_1,
  output [31:0] O_0_2,
  output [31:0] O_1_0,
  output [31:0] O_1_1,
  output [31:0] O_1_2,
  output [31:0] O_2_0,
  output [31:0] O_2_1,
  output [31:0] O_2_2
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_t0b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_t1b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_1_t0b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_1_t1b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_2_t0b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_2_t1b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_0; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_1; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_2; // @[MapS.scala 9:22]
  wire  other_ops_0_clock; // @[MapS.scala 10:86]
  wire  other_ops_0_reset; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_0_t0b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_0_t1b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_1_t0b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_1_t1b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_2_t0b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_2_t1b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_O_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_O_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_O_2; // @[MapS.scala 10:86]
  wire  other_ops_1_clock; // @[MapS.scala 10:86]
  wire  other_ops_1_reset; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_0_t0b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_0_t1b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_1_t0b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_1_t1b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_2_t0b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_2_t1b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_O_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_O_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_O_2; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  MapS_54 fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_t0b(fst_op_I_0_t0b),
    .I_0_t1b(fst_op_I_0_t1b),
    .I_1_t0b(fst_op_I_1_t0b),
    .I_1_t1b(fst_op_I_1_t1b),
    .I_2_t0b(fst_op_I_2_t0b),
    .I_2_t1b(fst_op_I_2_t1b),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1),
    .O_2(fst_op_O_2)
  );
  MapS_54 other_ops_0 ( // @[MapS.scala 10:86]
    .clock(other_ops_0_clock),
    .reset(other_ops_0_reset),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_t0b(other_ops_0_I_0_t0b),
    .I_0_t1b(other_ops_0_I_0_t1b),
    .I_1_t0b(other_ops_0_I_1_t0b),
    .I_1_t1b(other_ops_0_I_1_t1b),
    .I_2_t0b(other_ops_0_I_2_t0b),
    .I_2_t1b(other_ops_0_I_2_t1b),
    .O_0(other_ops_0_O_0),
    .O_1(other_ops_0_O_1),
    .O_2(other_ops_0_O_2)
  );
  MapS_54 other_ops_1 ( // @[MapS.scala 10:86]
    .clock(other_ops_1_clock),
    .reset(other_ops_1_reset),
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0_t0b(other_ops_1_I_0_t0b),
    .I_0_t1b(other_ops_1_I_0_t1b),
    .I_1_t0b(other_ops_1_I_1_t0b),
    .I_1_t1b(other_ops_1_I_1_t1b),
    .I_2_t0b(other_ops_1_I_2_t0b),
    .I_2_t1b(other_ops_1_I_2_t1b),
    .O_0(other_ops_1_O_0),
    .O_1(other_ops_1_O_1),
    .O_2(other_ops_1_O_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign O_0_1 = fst_op_O_1; // @[MapS.scala 17:8]
  assign O_0_2 = fst_op_O_2; // @[MapS.scala 17:8]
  assign O_1_0 = other_ops_0_O_0; // @[MapS.scala 21:12]
  assign O_1_1 = other_ops_0_O_1; // @[MapS.scala 21:12]
  assign O_1_2 = other_ops_0_O_2; // @[MapS.scala 21:12]
  assign O_2_0 = other_ops_1_O_0; // @[MapS.scala 21:12]
  assign O_2_1 = other_ops_1_O_1; // @[MapS.scala 21:12]
  assign O_2_2 = other_ops_1_O_2; // @[MapS.scala 21:12]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_t0b = I_0_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_0_t1b = I_0_0_t1b; // @[MapS.scala 16:12]
  assign fst_op_I_1_t0b = I_0_1_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_1_t1b = I_0_1_t1b; // @[MapS.scala 16:12]
  assign fst_op_I_2_t0b = I_0_2_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_2_t1b = I_0_2_t1b; // @[MapS.scala 16:12]
  assign other_ops_0_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_0_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_t0b = I_1_0_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_t1b = I_1_0_t1b; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_t0b = I_1_1_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_t1b = I_1_1_t1b; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_t0b = I_1_2_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_t1b = I_1_2_t1b; // @[MapS.scala 20:41]
  assign other_ops_1_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_1_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0_t0b = I_2_0_t0b; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_t1b = I_2_0_t1b; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_t0b = I_2_1_t0b; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_t1b = I_2_1_t1b; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_t0b = I_2_2_t0b; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_t1b = I_2_2_t1b; // @[MapS.scala 20:41]
endmodule
module ReduceS_2(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0,
  input  [31:0] I_1,
  input  [31:0] I_2,
  output [31:0] O_0
);
  wire [31:0] AddNoValid_I_t0b; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_I_t1b; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_O; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_1_I_t0b; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_1_I_t1b; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_1_O; // @[ReduceS.scala 20:43]
  reg [31:0] _T; // @[ReduceS.scala 27:24]
  reg [31:0] _RAND_0;
  reg [31:0] _T_1; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_1;
  reg [31:0] _T_2; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_2;
  reg [31:0] _T_3; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_3;
  reg  _T_4; // @[ReduceS.scala 47:32]
  reg [31:0] _RAND_4;
  reg  _T_5; // @[ReduceS.scala 47:24]
  reg [31:0] _RAND_5;
  AddNoValid AddNoValid ( // @[ReduceS.scala 20:43]
    .I_t0b(AddNoValid_I_t0b),
    .I_t1b(AddNoValid_I_t1b),
    .O(AddNoValid_O)
  );
  AddNoValid AddNoValid_1 ( // @[ReduceS.scala 20:43]
    .I_t0b(AddNoValid_1_I_t0b),
    .I_t1b(AddNoValid_1_I_t1b),
    .O(AddNoValid_1_O)
  );
  assign valid_down = _T_5; // @[ReduceS.scala 47:14]
  assign O_0 = _T; // @[ReduceS.scala 27:14]
  assign AddNoValid_I_t0b = _T_2; // @[ReduceS.scala 43:18]
  assign AddNoValid_I_t1b = AddNoValid_1_O; // @[ReduceS.scala 36:18]
  assign AddNoValid_1_I_t0b = _T_3; // @[ReduceS.scala 43:18]
  assign AddNoValid_1_I_t1b = _T_1; // @[ReduceS.scala 43:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_2 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_3 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T <= AddNoValid_O;
    _T_1 <= I_0;
    _T_2 <= I_1;
    _T_3 <= I_2;
    if (reset) begin
      _T_4 <= 1'h0;
    end else begin
      _T_4 <= valid_up;
    end
    _T_5 <= _T_4;
  end
endmodule
module MapS_56(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0,
  input  [31:0] I_0_1,
  input  [31:0] I_0_2,
  input  [31:0] I_1_0,
  input  [31:0] I_1_1,
  input  [31:0] I_1_2,
  input  [31:0] I_2_0,
  input  [31:0] I_2_1,
  input  [31:0] I_2_2,
  output [31:0] O_0_0,
  output [31:0] O_1_0,
  output [31:0] O_2_0
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_1; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_2; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_0; // @[MapS.scala 9:22]
  wire  other_ops_0_clock; // @[MapS.scala 10:86]
  wire  other_ops_0_reset; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_O_0; // @[MapS.scala 10:86]
  wire  other_ops_1_clock; // @[MapS.scala 10:86]
  wire  other_ops_1_reset; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_O_0; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  ReduceS_2 fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0(fst_op_I_0),
    .I_1(fst_op_I_1),
    .I_2(fst_op_I_2),
    .O_0(fst_op_O_0)
  );
  ReduceS_2 other_ops_0 ( // @[MapS.scala 10:86]
    .clock(other_ops_0_clock),
    .reset(other_ops_0_reset),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0(other_ops_0_I_0),
    .I_1(other_ops_0_I_1),
    .I_2(other_ops_0_I_2),
    .O_0(other_ops_0_O_0)
  );
  ReduceS_2 other_ops_1 ( // @[MapS.scala 10:86]
    .clock(other_ops_1_clock),
    .reset(other_ops_1_reset),
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0(other_ops_1_I_0),
    .I_1(other_ops_1_I_1),
    .I_2(other_ops_1_I_2),
    .O_0(other_ops_1_O_0)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign O_1_0 = other_ops_0_O_0; // @[MapS.scala 21:12]
  assign O_2_0 = other_ops_1_O_0; // @[MapS.scala 21:12]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0 = I_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_1 = I_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_2 = I_0_2; // @[MapS.scala 16:12]
  assign other_ops_0_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_0_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0 = I_1_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_1 = I_1_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_2 = I_1_2; // @[MapS.scala 20:41]
  assign other_ops_1_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_1_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0 = I_2_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_1 = I_2_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_2 = I_2_2; // @[MapS.scala 20:41]
endmodule
module MapSNoValid(
  input  [31:0] I_0_t0b,
  input  [31:0] I_0_t1b,
  output [31:0] O_0
);
  wire [31:0] fst_op_I_t0b; // @[MapS.scala 28:22]
  wire [31:0] fst_op_I_t1b; // @[MapS.scala 28:22]
  wire [31:0] fst_op_O; // @[MapS.scala 28:22]
  AddNoValid fst_op ( // @[MapS.scala 28:22]
    .I_t0b(fst_op_I_t0b),
    .I_t1b(fst_op_I_t1b),
    .O(fst_op_O)
  );
  assign O_0 = fst_op_O; // @[MapS.scala 35:8]
  assign fst_op_I_t0b = I_0_t0b; // @[MapS.scala 34:12]
  assign fst_op_I_t1b = I_0_t1b; // @[MapS.scala 34:12]
endmodule
module ReduceS_3(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0,
  input  [31:0] I_1_0,
  input  [31:0] I_2_0,
  output [31:0] O_0_0
);
  wire [31:0] MapSNoValid_I_0_t0b; // @[ReduceS.scala 20:43]
  wire [31:0] MapSNoValid_I_0_t1b; // @[ReduceS.scala 20:43]
  wire [31:0] MapSNoValid_O_0; // @[ReduceS.scala 20:43]
  wire [31:0] MapSNoValid_1_I_0_t0b; // @[ReduceS.scala 20:43]
  wire [31:0] MapSNoValid_1_I_0_t1b; // @[ReduceS.scala 20:43]
  wire [31:0] MapSNoValid_1_O_0; // @[ReduceS.scala 20:43]
  reg [31:0] _T_0; // @[ReduceS.scala 27:24]
  reg [31:0] _RAND_0;
  reg [31:0] _T_1_0; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_1;
  reg [31:0] _T_2_0; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_2;
  reg [31:0] _T_3_0; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_3;
  reg  _T_4; // @[ReduceS.scala 47:32]
  reg [31:0] _RAND_4;
  reg  _T_5; // @[ReduceS.scala 47:24]
  reg [31:0] _RAND_5;
  MapSNoValid MapSNoValid ( // @[ReduceS.scala 20:43]
    .I_0_t0b(MapSNoValid_I_0_t0b),
    .I_0_t1b(MapSNoValid_I_0_t1b),
    .O_0(MapSNoValid_O_0)
  );
  MapSNoValid MapSNoValid_1 ( // @[ReduceS.scala 20:43]
    .I_0_t0b(MapSNoValid_1_I_0_t0b),
    .I_0_t1b(MapSNoValid_1_I_0_t1b),
    .O_0(MapSNoValid_1_O_0)
  );
  assign valid_down = _T_5; // @[ReduceS.scala 47:14]
  assign O_0_0 = _T_0; // @[ReduceS.scala 27:14]
  assign MapSNoValid_I_0_t0b = _T_1_0; // @[ReduceS.scala 43:18]
  assign MapSNoValid_I_0_t1b = MapSNoValid_1_O_0; // @[ReduceS.scala 36:18]
  assign MapSNoValid_1_I_0_t0b = _T_2_0; // @[ReduceS.scala 43:18]
  assign MapSNoValid_1_I_0_t1b = _T_3_0; // @[ReduceS.scala 43:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1_0 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_2_0 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_3_0 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_0 <= MapSNoValid_O_0;
    _T_1_0 <= I_0_0;
    _T_2_0 <= I_1_0;
    _T_3_0 <= I_2_0;
    if (reset) begin
      _T_4 <= 1'h0;
    end else begin
      _T_4 <= valid_up;
    end
    _T_5 <= _T_4;
  end
endmodule
module InitialDelayCounter_5(
  input   clock,
  input   reset,
  output  valid_down
);
  reg [3:0] value; // @[InitialDelayCounter.scala 8:34]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[InitialDelayCounter.scala 17:17]
  wire [3:0] _T_4; // @[InitialDelayCounter.scala 17:53]
  assign _T_1 = value < 4'hd; // @[InitialDelayCounter.scala 17:17]
  assign _T_4 = value + 4'h1; // @[InitialDelayCounter.scala 17:53]
  assign valid_down = value == 4'hd; // @[InitialDelayCounter.scala 16:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 4'h0;
    end else if (_T_1) begin
      value <= _T_4;
    end
  end
endmodule
module AtomTuple_26(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0,
  input  [7:0]  I1,
  output [31:0] O_t0b,
  output [7:0]  O_t1b
);
  assign valid_down = valid_up; // @[Tuple.scala 51:14]
  assign O_t0b = I0; // @[Tuple.scala 49:9]
  assign O_t1b = I1; // @[Tuple.scala 50:9]
endmodule
module Map2S_64(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0,
  output [31:0] O_0_t0b,
  output [7:0]  O_0_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_t0b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_t1b; // @[Map2S.scala 9:22]
  AtomTuple_26 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1(fst_op_I1),
    .O_t0b(fst_op_O_t0b),
    .O_t1b(fst_op_O_t1b)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_t0b = fst_op_O_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b = fst_op_O_t1b; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1 = 8'sh8; // @[Map2S.scala 18:13]
endmodule
module Map2S_65(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0_0,
  output [31:0] O_0_0_t0b,
  output [7:0]  O_0_0_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_t0b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_t1b; // @[Map2S.scala 9:22]
  Map2S_64 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .O_0_t0b(fst_op_O_0_t0b),
    .O_0_t1b(fst_op_O_0_t1b)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_t0b = fst_op_O_0_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_t1b = fst_op_O_0_t1b; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
endmodule
module Div(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_t0b,
  input  [7:0]  I_t1b,
  output [31:0] O
);
  wire [31:0] BlackBoxMulUInt32_I0; // @[Arithmetic.scala 356:27]
  wire [31:0] BlackBoxMulUInt32_I1; // @[Arithmetic.scala 356:27]
  wire [63:0] BlackBoxMulUInt32_O; // @[Arithmetic.scala 356:27]
  wire  BlackBoxMulUInt32_clock; // @[Arithmetic.scala 356:27]
  wire [8:0] _T_1; // @[Cat.scala 29:58]
  reg  _T_3; // @[Arithmetic.scala 367:66]
  reg [31:0] _RAND_0;
  reg  _T_4; // @[Arithmetic.scala 367:58]
  reg [31:0] _RAND_1;
  reg  _T_5; // @[Arithmetic.scala 367:50]
  reg [31:0] _RAND_2;
  reg  _T_6; // @[Arithmetic.scala 367:42]
  reg [31:0] _RAND_3;
  reg  _T_7; // @[Arithmetic.scala 367:34]
  reg [31:0] _RAND_4;
  reg  _T_8; // @[Arithmetic.scala 367:26]
  reg [31:0] _RAND_5;
  BlackBoxMulUInt32 BlackBoxMulUInt32 ( // @[Arithmetic.scala 356:27]
    .I0(BlackBoxMulUInt32_I0),
    .I1(BlackBoxMulUInt32_I1),
    .O(BlackBoxMulUInt32_O),
    .clock(BlackBoxMulUInt32_clock)
  );
  assign _T_1 = {1'h0,I_t1b}; // @[Cat.scala 29:58]
  assign valid_down = _T_8; // @[Arithmetic.scala 367:16]
  assign O = BlackBoxMulUInt32_O[38:7]; // @[Arithmetic.scala 359:7]
  assign BlackBoxMulUInt32_I0 = I_t0b; // @[Arithmetic.scala 357:21]
  assign BlackBoxMulUInt32_I1 = {{23'd0}, _T_1}; // @[Arithmetic.scala 358:21]
  assign BlackBoxMulUInt32_clock = clock; // @[Arithmetic.scala 360:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_3 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_4 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_5 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_6 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_7 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_8 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_3 <= 1'h0;
    end else begin
      _T_3 <= valid_up;
    end
    if (reset) begin
      _T_4 <= 1'h0;
    end else begin
      _T_4 <= _T_3;
    end
    if (reset) begin
      _T_5 <= 1'h0;
    end else begin
      _T_5 <= _T_4;
    end
    _T_6 <= _T_5;
    _T_7 <= _T_6;
    _T_8 <= _T_7;
  end
endmodule
module MapS_57(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_t0b,
  input  [7:0]  I_0_t1b,
  output [31:0] O_0
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_t1b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O; // @[MapS.scala 9:22]
  Div fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_t0b(fst_op_I_t0b),
    .I_t1b(fst_op_I_t1b),
    .O(fst_op_O)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0 = fst_op_O; // @[MapS.scala 17:8]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_t0b = I_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_t1b = I_0_t1b; // @[MapS.scala 16:12]
endmodule
module MapS_58(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0_t0b,
  input  [7:0]  I_0_0_t1b,
  output [31:0] O_0_0
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_t1b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_0; // @[MapS.scala 9:22]
  MapS_57 fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_t0b(fst_op_I_0_t0b),
    .I_0_t1b(fst_op_I_0_t1b),
    .O_0(fst_op_O_0)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_t0b = I_0_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_0_t1b = I_0_0_t1b; // @[MapS.scala 16:12]
endmodule
module Module_8(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0,
  input  [31:0] I_0_1,
  input  [31:0] I_0_2,
  input  [31:0] I_1_0,
  input  [31:0] I_1_1,
  input  [31:0] I_1_2,
  input  [31:0] I_2_0,
  input  [31:0] I_2_1,
  input  [31:0] I_2_2,
  output [31:0] O_0_0
);
  wire  InitialDelayCounter_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_valid_down; // @[Const.scala 11:33]
  wire  n560_valid_up; // @[Top.scala 358:22]
  wire  n560_valid_down; // @[Top.scala 358:22]
  wire [31:0] n560_I0_0_0; // @[Top.scala 358:22]
  wire [31:0] n560_I0_0_1; // @[Top.scala 358:22]
  wire [31:0] n560_I0_0_2; // @[Top.scala 358:22]
  wire [31:0] n560_I0_1_0; // @[Top.scala 358:22]
  wire [31:0] n560_I0_1_1; // @[Top.scala 358:22]
  wire [31:0] n560_I0_1_2; // @[Top.scala 358:22]
  wire [31:0] n560_I0_2_0; // @[Top.scala 358:22]
  wire [31:0] n560_I0_2_1; // @[Top.scala 358:22]
  wire [31:0] n560_I0_2_2; // @[Top.scala 358:22]
  wire [31:0] n560_O_0_0_t0b; // @[Top.scala 358:22]
  wire [31:0] n560_O_0_0_t1b; // @[Top.scala 358:22]
  wire [31:0] n560_O_0_1_t0b; // @[Top.scala 358:22]
  wire [31:0] n560_O_0_1_t1b; // @[Top.scala 358:22]
  wire [31:0] n560_O_0_2_t0b; // @[Top.scala 358:22]
  wire [31:0] n560_O_0_2_t1b; // @[Top.scala 358:22]
  wire [31:0] n560_O_1_0_t0b; // @[Top.scala 358:22]
  wire [31:0] n560_O_1_0_t1b; // @[Top.scala 358:22]
  wire [31:0] n560_O_1_1_t0b; // @[Top.scala 358:22]
  wire [31:0] n560_O_1_1_t1b; // @[Top.scala 358:22]
  wire [31:0] n560_O_1_2_t0b; // @[Top.scala 358:22]
  wire [31:0] n560_O_1_2_t1b; // @[Top.scala 358:22]
  wire [31:0] n560_O_2_0_t0b; // @[Top.scala 358:22]
  wire [31:0] n560_O_2_0_t1b; // @[Top.scala 358:22]
  wire [31:0] n560_O_2_1_t0b; // @[Top.scala 358:22]
  wire [31:0] n560_O_2_1_t1b; // @[Top.scala 358:22]
  wire [31:0] n560_O_2_2_t0b; // @[Top.scala 358:22]
  wire [31:0] n560_O_2_2_t1b; // @[Top.scala 358:22]
  wire  n571_clock; // @[Top.scala 362:22]
  wire  n571_reset; // @[Top.scala 362:22]
  wire  n571_valid_up; // @[Top.scala 362:22]
  wire  n571_valid_down; // @[Top.scala 362:22]
  wire [31:0] n571_I_0_0_t0b; // @[Top.scala 362:22]
  wire [31:0] n571_I_0_0_t1b; // @[Top.scala 362:22]
  wire [31:0] n571_I_0_1_t0b; // @[Top.scala 362:22]
  wire [31:0] n571_I_0_1_t1b; // @[Top.scala 362:22]
  wire [31:0] n571_I_0_2_t0b; // @[Top.scala 362:22]
  wire [31:0] n571_I_0_2_t1b; // @[Top.scala 362:22]
  wire [31:0] n571_I_1_0_t0b; // @[Top.scala 362:22]
  wire [31:0] n571_I_1_0_t1b; // @[Top.scala 362:22]
  wire [31:0] n571_I_1_1_t0b; // @[Top.scala 362:22]
  wire [31:0] n571_I_1_1_t1b; // @[Top.scala 362:22]
  wire [31:0] n571_I_1_2_t0b; // @[Top.scala 362:22]
  wire [31:0] n571_I_1_2_t1b; // @[Top.scala 362:22]
  wire [31:0] n571_I_2_0_t0b; // @[Top.scala 362:22]
  wire [31:0] n571_I_2_0_t1b; // @[Top.scala 362:22]
  wire [31:0] n571_I_2_1_t0b; // @[Top.scala 362:22]
  wire [31:0] n571_I_2_1_t1b; // @[Top.scala 362:22]
  wire [31:0] n571_I_2_2_t0b; // @[Top.scala 362:22]
  wire [31:0] n571_I_2_2_t1b; // @[Top.scala 362:22]
  wire [31:0] n571_O_0_0; // @[Top.scala 362:22]
  wire [31:0] n571_O_0_1; // @[Top.scala 362:22]
  wire [31:0] n571_O_0_2; // @[Top.scala 362:22]
  wire [31:0] n571_O_1_0; // @[Top.scala 362:22]
  wire [31:0] n571_O_1_1; // @[Top.scala 362:22]
  wire [31:0] n571_O_1_2; // @[Top.scala 362:22]
  wire [31:0] n571_O_2_0; // @[Top.scala 362:22]
  wire [31:0] n571_O_2_1; // @[Top.scala 362:22]
  wire [31:0] n571_O_2_2; // @[Top.scala 362:22]
  wire  n576_clock; // @[Top.scala 365:22]
  wire  n576_reset; // @[Top.scala 365:22]
  wire  n576_valid_up; // @[Top.scala 365:22]
  wire  n576_valid_down; // @[Top.scala 365:22]
  wire [31:0] n576_I_0_0; // @[Top.scala 365:22]
  wire [31:0] n576_I_0_1; // @[Top.scala 365:22]
  wire [31:0] n576_I_0_2; // @[Top.scala 365:22]
  wire [31:0] n576_I_1_0; // @[Top.scala 365:22]
  wire [31:0] n576_I_1_1; // @[Top.scala 365:22]
  wire [31:0] n576_I_1_2; // @[Top.scala 365:22]
  wire [31:0] n576_I_2_0; // @[Top.scala 365:22]
  wire [31:0] n576_I_2_1; // @[Top.scala 365:22]
  wire [31:0] n576_I_2_2; // @[Top.scala 365:22]
  wire [31:0] n576_O_0_0; // @[Top.scala 365:22]
  wire [31:0] n576_O_1_0; // @[Top.scala 365:22]
  wire [31:0] n576_O_2_0; // @[Top.scala 365:22]
  wire  n581_clock; // @[Top.scala 368:22]
  wire  n581_reset; // @[Top.scala 368:22]
  wire  n581_valid_up; // @[Top.scala 368:22]
  wire  n581_valid_down; // @[Top.scala 368:22]
  wire [31:0] n581_I_0_0; // @[Top.scala 368:22]
  wire [31:0] n581_I_1_0; // @[Top.scala 368:22]
  wire [31:0] n581_I_2_0; // @[Top.scala 368:22]
  wire [31:0] n581_O_0_0; // @[Top.scala 368:22]
  wire  InitialDelayCounter_1_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_1_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_1_valid_down; // @[Const.scala 11:33]
  wire  n584_valid_up; // @[Top.scala 372:22]
  wire  n584_valid_down; // @[Top.scala 372:22]
  wire [31:0] n584_I0_0_0; // @[Top.scala 372:22]
  wire [31:0] n584_O_0_0_t0b; // @[Top.scala 372:22]
  wire [7:0] n584_O_0_0_t1b; // @[Top.scala 372:22]
  wire  n595_clock; // @[Top.scala 376:22]
  wire  n595_reset; // @[Top.scala 376:22]
  wire  n595_valid_up; // @[Top.scala 376:22]
  wire  n595_valid_down; // @[Top.scala 376:22]
  wire [31:0] n595_I_0_0_t0b; // @[Top.scala 376:22]
  wire [7:0] n595_I_0_0_t1b; // @[Top.scala 376:22]
  wire [31:0] n595_O_0_0; // @[Top.scala 376:22]
  InitialDelayCounter_2 InitialDelayCounter ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_clock),
    .reset(InitialDelayCounter_reset),
    .valid_down(InitialDelayCounter_valid_down)
  );
  Map2S_63 n560 ( // @[Top.scala 358:22]
    .valid_up(n560_valid_up),
    .valid_down(n560_valid_down),
    .I0_0_0(n560_I0_0_0),
    .I0_0_1(n560_I0_0_1),
    .I0_0_2(n560_I0_0_2),
    .I0_1_0(n560_I0_1_0),
    .I0_1_1(n560_I0_1_1),
    .I0_1_2(n560_I0_1_2),
    .I0_2_0(n560_I0_2_0),
    .I0_2_1(n560_I0_2_1),
    .I0_2_2(n560_I0_2_2),
    .O_0_0_t0b(n560_O_0_0_t0b),
    .O_0_0_t1b(n560_O_0_0_t1b),
    .O_0_1_t0b(n560_O_0_1_t0b),
    .O_0_1_t1b(n560_O_0_1_t1b),
    .O_0_2_t0b(n560_O_0_2_t0b),
    .O_0_2_t1b(n560_O_0_2_t1b),
    .O_1_0_t0b(n560_O_1_0_t0b),
    .O_1_0_t1b(n560_O_1_0_t1b),
    .O_1_1_t0b(n560_O_1_1_t0b),
    .O_1_1_t1b(n560_O_1_1_t1b),
    .O_1_2_t0b(n560_O_1_2_t0b),
    .O_1_2_t1b(n560_O_1_2_t1b),
    .O_2_0_t0b(n560_O_2_0_t0b),
    .O_2_0_t1b(n560_O_2_0_t1b),
    .O_2_1_t0b(n560_O_2_1_t0b),
    .O_2_1_t1b(n560_O_2_1_t1b),
    .O_2_2_t0b(n560_O_2_2_t0b),
    .O_2_2_t1b(n560_O_2_2_t1b)
  );
  MapS_55 n571 ( // @[Top.scala 362:22]
    .clock(n571_clock),
    .reset(n571_reset),
    .valid_up(n571_valid_up),
    .valid_down(n571_valid_down),
    .I_0_0_t0b(n571_I_0_0_t0b),
    .I_0_0_t1b(n571_I_0_0_t1b),
    .I_0_1_t0b(n571_I_0_1_t0b),
    .I_0_1_t1b(n571_I_0_1_t1b),
    .I_0_2_t0b(n571_I_0_2_t0b),
    .I_0_2_t1b(n571_I_0_2_t1b),
    .I_1_0_t0b(n571_I_1_0_t0b),
    .I_1_0_t1b(n571_I_1_0_t1b),
    .I_1_1_t0b(n571_I_1_1_t0b),
    .I_1_1_t1b(n571_I_1_1_t1b),
    .I_1_2_t0b(n571_I_1_2_t0b),
    .I_1_2_t1b(n571_I_1_2_t1b),
    .I_2_0_t0b(n571_I_2_0_t0b),
    .I_2_0_t1b(n571_I_2_0_t1b),
    .I_2_1_t0b(n571_I_2_1_t0b),
    .I_2_1_t1b(n571_I_2_1_t1b),
    .I_2_2_t0b(n571_I_2_2_t0b),
    .I_2_2_t1b(n571_I_2_2_t1b),
    .O_0_0(n571_O_0_0),
    .O_0_1(n571_O_0_1),
    .O_0_2(n571_O_0_2),
    .O_1_0(n571_O_1_0),
    .O_1_1(n571_O_1_1),
    .O_1_2(n571_O_1_2),
    .O_2_0(n571_O_2_0),
    .O_2_1(n571_O_2_1),
    .O_2_2(n571_O_2_2)
  );
  MapS_56 n576 ( // @[Top.scala 365:22]
    .clock(n576_clock),
    .reset(n576_reset),
    .valid_up(n576_valid_up),
    .valid_down(n576_valid_down),
    .I_0_0(n576_I_0_0),
    .I_0_1(n576_I_0_1),
    .I_0_2(n576_I_0_2),
    .I_1_0(n576_I_1_0),
    .I_1_1(n576_I_1_1),
    .I_1_2(n576_I_1_2),
    .I_2_0(n576_I_2_0),
    .I_2_1(n576_I_2_1),
    .I_2_2(n576_I_2_2),
    .O_0_0(n576_O_0_0),
    .O_1_0(n576_O_1_0),
    .O_2_0(n576_O_2_0)
  );
  ReduceS_3 n581 ( // @[Top.scala 368:22]
    .clock(n581_clock),
    .reset(n581_reset),
    .valid_up(n581_valid_up),
    .valid_down(n581_valid_down),
    .I_0_0(n581_I_0_0),
    .I_1_0(n581_I_1_0),
    .I_2_0(n581_I_2_0),
    .O_0_0(n581_O_0_0)
  );
  InitialDelayCounter_5 InitialDelayCounter_1 ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_1_clock),
    .reset(InitialDelayCounter_1_reset),
    .valid_down(InitialDelayCounter_1_valid_down)
  );
  Map2S_65 n584 ( // @[Top.scala 372:22]
    .valid_up(n584_valid_up),
    .valid_down(n584_valid_down),
    .I0_0_0(n584_I0_0_0),
    .O_0_0_t0b(n584_O_0_0_t0b),
    .O_0_0_t1b(n584_O_0_0_t1b)
  );
  MapS_58 n595 ( // @[Top.scala 376:22]
    .clock(n595_clock),
    .reset(n595_reset),
    .valid_up(n595_valid_up),
    .valid_down(n595_valid_down),
    .I_0_0_t0b(n595_I_0_0_t0b),
    .I_0_0_t1b(n595_I_0_0_t1b),
    .O_0_0(n595_O_0_0)
  );
  assign valid_down = n595_valid_down; // @[Top.scala 380:16]
  assign O_0_0 = n595_O_0_0; // @[Top.scala 379:7]
  assign InitialDelayCounter_clock = clock;
  assign InitialDelayCounter_reset = reset;
  assign n560_valid_up = valid_up & InitialDelayCounter_valid_down; // @[Top.scala 361:19]
  assign n560_I0_0_0 = I_0_0; // @[Top.scala 359:13]
  assign n560_I0_0_1 = I_0_1; // @[Top.scala 359:13]
  assign n560_I0_0_2 = I_0_2; // @[Top.scala 359:13]
  assign n560_I0_1_0 = I_1_0; // @[Top.scala 359:13]
  assign n560_I0_1_1 = I_1_1; // @[Top.scala 359:13]
  assign n560_I0_1_2 = I_1_2; // @[Top.scala 359:13]
  assign n560_I0_2_0 = I_2_0; // @[Top.scala 359:13]
  assign n560_I0_2_1 = I_2_1; // @[Top.scala 359:13]
  assign n560_I0_2_2 = I_2_2; // @[Top.scala 359:13]
  assign n571_clock = clock;
  assign n571_reset = reset;
  assign n571_valid_up = n560_valid_down; // @[Top.scala 364:19]
  assign n571_I_0_0_t0b = n560_O_0_0_t0b; // @[Top.scala 363:12]
  assign n571_I_0_0_t1b = n560_O_0_0_t1b; // @[Top.scala 363:12]
  assign n571_I_0_1_t0b = n560_O_0_1_t0b; // @[Top.scala 363:12]
  assign n571_I_0_1_t1b = n560_O_0_1_t1b; // @[Top.scala 363:12]
  assign n571_I_0_2_t0b = n560_O_0_2_t0b; // @[Top.scala 363:12]
  assign n571_I_0_2_t1b = n560_O_0_2_t1b; // @[Top.scala 363:12]
  assign n571_I_1_0_t0b = n560_O_1_0_t0b; // @[Top.scala 363:12]
  assign n571_I_1_0_t1b = n560_O_1_0_t1b; // @[Top.scala 363:12]
  assign n571_I_1_1_t0b = n560_O_1_1_t0b; // @[Top.scala 363:12]
  assign n571_I_1_1_t1b = n560_O_1_1_t1b; // @[Top.scala 363:12]
  assign n571_I_1_2_t0b = n560_O_1_2_t0b; // @[Top.scala 363:12]
  assign n571_I_1_2_t1b = n560_O_1_2_t1b; // @[Top.scala 363:12]
  assign n571_I_2_0_t0b = n560_O_2_0_t0b; // @[Top.scala 363:12]
  assign n571_I_2_0_t1b = n560_O_2_0_t1b; // @[Top.scala 363:12]
  assign n571_I_2_1_t0b = n560_O_2_1_t0b; // @[Top.scala 363:12]
  assign n571_I_2_1_t1b = n560_O_2_1_t1b; // @[Top.scala 363:12]
  assign n571_I_2_2_t0b = n560_O_2_2_t0b; // @[Top.scala 363:12]
  assign n571_I_2_2_t1b = n560_O_2_2_t1b; // @[Top.scala 363:12]
  assign n576_clock = clock;
  assign n576_reset = reset;
  assign n576_valid_up = n571_valid_down; // @[Top.scala 367:19]
  assign n576_I_0_0 = n571_O_0_0; // @[Top.scala 366:12]
  assign n576_I_0_1 = n571_O_0_1; // @[Top.scala 366:12]
  assign n576_I_0_2 = n571_O_0_2; // @[Top.scala 366:12]
  assign n576_I_1_0 = n571_O_1_0; // @[Top.scala 366:12]
  assign n576_I_1_1 = n571_O_1_1; // @[Top.scala 366:12]
  assign n576_I_1_2 = n571_O_1_2; // @[Top.scala 366:12]
  assign n576_I_2_0 = n571_O_2_0; // @[Top.scala 366:12]
  assign n576_I_2_1 = n571_O_2_1; // @[Top.scala 366:12]
  assign n576_I_2_2 = n571_O_2_2; // @[Top.scala 366:12]
  assign n581_clock = clock;
  assign n581_reset = reset;
  assign n581_valid_up = n576_valid_down; // @[Top.scala 370:19]
  assign n581_I_0_0 = n576_O_0_0; // @[Top.scala 369:12]
  assign n581_I_1_0 = n576_O_1_0; // @[Top.scala 369:12]
  assign n581_I_2_0 = n576_O_2_0; // @[Top.scala 369:12]
  assign InitialDelayCounter_1_clock = clock;
  assign InitialDelayCounter_1_reset = reset;
  assign n584_valid_up = n581_valid_down & InitialDelayCounter_1_valid_down; // @[Top.scala 375:19]
  assign n584_I0_0_0 = n581_O_0_0; // @[Top.scala 373:13]
  assign n595_clock = clock;
  assign n595_reset = reset;
  assign n595_valid_up = n584_valid_down; // @[Top.scala 378:19]
  assign n595_I_0_0_t0b = n584_O_0_0_t0b; // @[Top.scala 377:12]
  assign n595_I_0_0_t1b = n584_O_0_0_t1b; // @[Top.scala 377:12]
endmodule
module MapS_59(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0_0,
  input  [31:0] I_0_0_1,
  input  [31:0] I_0_0_2,
  input  [31:0] I_0_1_0,
  input  [31:0] I_0_1_1,
  input  [31:0] I_0_1_2,
  input  [31:0] I_0_2_0,
  input  [31:0] I_0_2_1,
  input  [31:0] I_0_2_2,
  input  [31:0] I_1_0_0,
  input  [31:0] I_1_0_1,
  input  [31:0] I_1_0_2,
  input  [31:0] I_1_1_0,
  input  [31:0] I_1_1_1,
  input  [31:0] I_1_1_2,
  input  [31:0] I_1_2_0,
  input  [31:0] I_1_2_1,
  input  [31:0] I_1_2_2,
  input  [31:0] I_2_0_0,
  input  [31:0] I_2_0_1,
  input  [31:0] I_2_0_2,
  input  [31:0] I_2_1_0,
  input  [31:0] I_2_1_1,
  input  [31:0] I_2_1_2,
  input  [31:0] I_2_2_0,
  input  [31:0] I_2_2_1,
  input  [31:0] I_2_2_2,
  input  [31:0] I_3_0_0,
  input  [31:0] I_3_0_1,
  input  [31:0] I_3_0_2,
  input  [31:0] I_3_1_0,
  input  [31:0] I_3_1_1,
  input  [31:0] I_3_1_2,
  input  [31:0] I_3_2_0,
  input  [31:0] I_3_2_1,
  input  [31:0] I_3_2_2,
  input  [31:0] I_4_0_0,
  input  [31:0] I_4_0_1,
  input  [31:0] I_4_0_2,
  input  [31:0] I_4_1_0,
  input  [31:0] I_4_1_1,
  input  [31:0] I_4_1_2,
  input  [31:0] I_4_2_0,
  input  [31:0] I_4_2_1,
  input  [31:0] I_4_2_2,
  input  [31:0] I_5_0_0,
  input  [31:0] I_5_0_1,
  input  [31:0] I_5_0_2,
  input  [31:0] I_5_1_0,
  input  [31:0] I_5_1_1,
  input  [31:0] I_5_1_2,
  input  [31:0] I_5_2_0,
  input  [31:0] I_5_2_1,
  input  [31:0] I_5_2_2,
  input  [31:0] I_6_0_0,
  input  [31:0] I_6_0_1,
  input  [31:0] I_6_0_2,
  input  [31:0] I_6_1_0,
  input  [31:0] I_6_1_1,
  input  [31:0] I_6_1_2,
  input  [31:0] I_6_2_0,
  input  [31:0] I_6_2_1,
  input  [31:0] I_6_2_2,
  input  [31:0] I_7_0_0,
  input  [31:0] I_7_0_1,
  input  [31:0] I_7_0_2,
  input  [31:0] I_7_1_0,
  input  [31:0] I_7_1_1,
  input  [31:0] I_7_1_2,
  input  [31:0] I_7_2_0,
  input  [31:0] I_7_2_1,
  input  [31:0] I_7_2_2,
  output [31:0] O_0_0_0,
  output [31:0] O_1_0_0,
  output [31:0] O_2_0_0,
  output [31:0] O_3_0_0,
  output [31:0] O_4_0_0,
  output [31:0] O_5_0_0,
  output [31:0] O_6_0_0,
  output [31:0] O_7_0_0
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_0; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_1; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_2; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_1_0; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_1_1; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_1_2; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_2_0; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_2_1; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_2_2; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_0_0; // @[MapS.scala 9:22]
  wire  other_ops_0_clock; // @[MapS.scala 10:86]
  wire  other_ops_0_reset; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_2_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_1_clock; // @[MapS.scala 10:86]
  wire  other_ops_1_reset; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_2_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_2_clock; // @[MapS.scala 10:86]
  wire  other_ops_2_reset; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_2_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_3_clock; // @[MapS.scala 10:86]
  wire  other_ops_3_reset; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_2_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_4_clock; // @[MapS.scala 10:86]
  wire  other_ops_4_reset; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_2_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_5_clock; // @[MapS.scala 10:86]
  wire  other_ops_5_reset; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_2_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_6_clock; // @[MapS.scala 10:86]
  wire  other_ops_6_reset; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_2_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_O_0_0; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  wire  _T_1; // @[MapS.scala 23:83]
  wire  _T_2; // @[MapS.scala 23:83]
  wire  _T_3; // @[MapS.scala 23:83]
  wire  _T_4; // @[MapS.scala 23:83]
  wire  _T_5; // @[MapS.scala 23:83]
  Module_8 fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_0(fst_op_I_0_0),
    .I_0_1(fst_op_I_0_1),
    .I_0_2(fst_op_I_0_2),
    .I_1_0(fst_op_I_1_0),
    .I_1_1(fst_op_I_1_1),
    .I_1_2(fst_op_I_1_2),
    .I_2_0(fst_op_I_2_0),
    .I_2_1(fst_op_I_2_1),
    .I_2_2(fst_op_I_2_2),
    .O_0_0(fst_op_O_0_0)
  );
  Module_8 other_ops_0 ( // @[MapS.scala 10:86]
    .clock(other_ops_0_clock),
    .reset(other_ops_0_reset),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_0(other_ops_0_I_0_0),
    .I_0_1(other_ops_0_I_0_1),
    .I_0_2(other_ops_0_I_0_2),
    .I_1_0(other_ops_0_I_1_0),
    .I_1_1(other_ops_0_I_1_1),
    .I_1_2(other_ops_0_I_1_2),
    .I_2_0(other_ops_0_I_2_0),
    .I_2_1(other_ops_0_I_2_1),
    .I_2_2(other_ops_0_I_2_2),
    .O_0_0(other_ops_0_O_0_0)
  );
  Module_8 other_ops_1 ( // @[MapS.scala 10:86]
    .clock(other_ops_1_clock),
    .reset(other_ops_1_reset),
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0_0(other_ops_1_I_0_0),
    .I_0_1(other_ops_1_I_0_1),
    .I_0_2(other_ops_1_I_0_2),
    .I_1_0(other_ops_1_I_1_0),
    .I_1_1(other_ops_1_I_1_1),
    .I_1_2(other_ops_1_I_1_2),
    .I_2_0(other_ops_1_I_2_0),
    .I_2_1(other_ops_1_I_2_1),
    .I_2_2(other_ops_1_I_2_2),
    .O_0_0(other_ops_1_O_0_0)
  );
  Module_8 other_ops_2 ( // @[MapS.scala 10:86]
    .clock(other_ops_2_clock),
    .reset(other_ops_2_reset),
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I_0_0(other_ops_2_I_0_0),
    .I_0_1(other_ops_2_I_0_1),
    .I_0_2(other_ops_2_I_0_2),
    .I_1_0(other_ops_2_I_1_0),
    .I_1_1(other_ops_2_I_1_1),
    .I_1_2(other_ops_2_I_1_2),
    .I_2_0(other_ops_2_I_2_0),
    .I_2_1(other_ops_2_I_2_1),
    .I_2_2(other_ops_2_I_2_2),
    .O_0_0(other_ops_2_O_0_0)
  );
  Module_8 other_ops_3 ( // @[MapS.scala 10:86]
    .clock(other_ops_3_clock),
    .reset(other_ops_3_reset),
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I_0_0(other_ops_3_I_0_0),
    .I_0_1(other_ops_3_I_0_1),
    .I_0_2(other_ops_3_I_0_2),
    .I_1_0(other_ops_3_I_1_0),
    .I_1_1(other_ops_3_I_1_1),
    .I_1_2(other_ops_3_I_1_2),
    .I_2_0(other_ops_3_I_2_0),
    .I_2_1(other_ops_3_I_2_1),
    .I_2_2(other_ops_3_I_2_2),
    .O_0_0(other_ops_3_O_0_0)
  );
  Module_8 other_ops_4 ( // @[MapS.scala 10:86]
    .clock(other_ops_4_clock),
    .reset(other_ops_4_reset),
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I_0_0(other_ops_4_I_0_0),
    .I_0_1(other_ops_4_I_0_1),
    .I_0_2(other_ops_4_I_0_2),
    .I_1_0(other_ops_4_I_1_0),
    .I_1_1(other_ops_4_I_1_1),
    .I_1_2(other_ops_4_I_1_2),
    .I_2_0(other_ops_4_I_2_0),
    .I_2_1(other_ops_4_I_2_1),
    .I_2_2(other_ops_4_I_2_2),
    .O_0_0(other_ops_4_O_0_0)
  );
  Module_8 other_ops_5 ( // @[MapS.scala 10:86]
    .clock(other_ops_5_clock),
    .reset(other_ops_5_reset),
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I_0_0(other_ops_5_I_0_0),
    .I_0_1(other_ops_5_I_0_1),
    .I_0_2(other_ops_5_I_0_2),
    .I_1_0(other_ops_5_I_1_0),
    .I_1_1(other_ops_5_I_1_1),
    .I_1_2(other_ops_5_I_1_2),
    .I_2_0(other_ops_5_I_2_0),
    .I_2_1(other_ops_5_I_2_1),
    .I_2_2(other_ops_5_I_2_2),
    .O_0_0(other_ops_5_O_0_0)
  );
  Module_8 other_ops_6 ( // @[MapS.scala 10:86]
    .clock(other_ops_6_clock),
    .reset(other_ops_6_reset),
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I_0_0(other_ops_6_I_0_0),
    .I_0_1(other_ops_6_I_0_1),
    .I_0_2(other_ops_6_I_0_2),
    .I_1_0(other_ops_6_I_1_0),
    .I_1_1(other_ops_6_I_1_1),
    .I_1_2(other_ops_6_I_1_2),
    .I_2_0(other_ops_6_I_2_0),
    .I_2_1(other_ops_6_I_2_1),
    .I_2_2(other_ops_6_I_2_2),
    .O_0_0(other_ops_6_O_0_0)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[MapS.scala 23:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[MapS.scala 23:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[MapS.scala 23:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[MapS.scala 23:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T_5 & other_ops_6_valid_down; // @[MapS.scala 23:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[MapS.scala 17:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[MapS.scala 21:12]
  assign O_2_0_0 = other_ops_1_O_0_0; // @[MapS.scala 21:12]
  assign O_3_0_0 = other_ops_2_O_0_0; // @[MapS.scala 21:12]
  assign O_4_0_0 = other_ops_3_O_0_0; // @[MapS.scala 21:12]
  assign O_5_0_0 = other_ops_4_O_0_0; // @[MapS.scala 21:12]
  assign O_6_0_0 = other_ops_5_O_0_0; // @[MapS.scala 21:12]
  assign O_7_0_0 = other_ops_6_O_0_0; // @[MapS.scala 21:12]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_0 = I_0_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_1 = I_0_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_2 = I_0_0_2; // @[MapS.scala 16:12]
  assign fst_op_I_1_0 = I_0_1_0; // @[MapS.scala 16:12]
  assign fst_op_I_1_1 = I_0_1_1; // @[MapS.scala 16:12]
  assign fst_op_I_1_2 = I_0_1_2; // @[MapS.scala 16:12]
  assign fst_op_I_2_0 = I_0_2_0; // @[MapS.scala 16:12]
  assign fst_op_I_2_1 = I_0_2_1; // @[MapS.scala 16:12]
  assign fst_op_I_2_2 = I_0_2_2; // @[MapS.scala 16:12]
  assign other_ops_0_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_0_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_0 = I_1_0_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1 = I_1_0_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2 = I_1_0_2; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_0 = I_1_1_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_1 = I_1_1_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_2 = I_1_1_2; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_0 = I_1_2_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_1 = I_1_2_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_2 = I_1_2_2; // @[MapS.scala 20:41]
  assign other_ops_1_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_1_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0_0 = I_2_0_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1 = I_2_0_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2 = I_2_0_2; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_0 = I_2_1_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_1 = I_2_1_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_2 = I_2_1_2; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_0 = I_2_2_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_1 = I_2_2_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_2 = I_2_2_2; // @[MapS.scala 20:41]
  assign other_ops_2_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_2_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_2_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_2_I_0_0 = I_3_0_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1 = I_3_0_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2 = I_3_0_2; // @[MapS.scala 20:41]
  assign other_ops_2_I_1_0 = I_3_1_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_1_1 = I_3_1_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_1_2 = I_3_1_2; // @[MapS.scala 20:41]
  assign other_ops_2_I_2_0 = I_3_2_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_2_1 = I_3_2_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_2_2 = I_3_2_2; // @[MapS.scala 20:41]
  assign other_ops_3_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_3_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_3_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_3_I_0_0 = I_4_0_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_1 = I_4_0_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_2 = I_4_0_2; // @[MapS.scala 20:41]
  assign other_ops_3_I_1_0 = I_4_1_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_1_1 = I_4_1_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_1_2 = I_4_1_2; // @[MapS.scala 20:41]
  assign other_ops_3_I_2_0 = I_4_2_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_2_1 = I_4_2_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_2_2 = I_4_2_2; // @[MapS.scala 20:41]
  assign other_ops_4_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_4_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_4_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_4_I_0_0 = I_5_0_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_1 = I_5_0_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_2 = I_5_0_2; // @[MapS.scala 20:41]
  assign other_ops_4_I_1_0 = I_5_1_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_1_1 = I_5_1_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_1_2 = I_5_1_2; // @[MapS.scala 20:41]
  assign other_ops_4_I_2_0 = I_5_2_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_2_1 = I_5_2_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_2_2 = I_5_2_2; // @[MapS.scala 20:41]
  assign other_ops_5_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_5_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_5_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_5_I_0_0 = I_6_0_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_1 = I_6_0_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_2 = I_6_0_2; // @[MapS.scala 20:41]
  assign other_ops_5_I_1_0 = I_6_1_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_1_1 = I_6_1_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_1_2 = I_6_1_2; // @[MapS.scala 20:41]
  assign other_ops_5_I_2_0 = I_6_2_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_2_1 = I_6_2_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_2_2 = I_6_2_2; // @[MapS.scala 20:41]
  assign other_ops_6_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_6_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_6_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_6_I_0_0 = I_7_0_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_1 = I_7_0_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_2 = I_7_0_2; // @[MapS.scala 20:41]
  assign other_ops_6_I_1_0 = I_7_1_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_1_1 = I_7_1_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_1_2 = I_7_1_2; // @[MapS.scala 20:41]
  assign other_ops_6_I_2_0 = I_7_2_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_2_1 = I_7_2_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_2_2 = I_7_2_2; // @[MapS.scala 20:41]
endmodule
module MapT_22(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0_0,
  input  [31:0] I_0_0_1,
  input  [31:0] I_0_0_2,
  input  [31:0] I_0_1_0,
  input  [31:0] I_0_1_1,
  input  [31:0] I_0_1_2,
  input  [31:0] I_0_2_0,
  input  [31:0] I_0_2_1,
  input  [31:0] I_0_2_2,
  input  [31:0] I_1_0_0,
  input  [31:0] I_1_0_1,
  input  [31:0] I_1_0_2,
  input  [31:0] I_1_1_0,
  input  [31:0] I_1_1_1,
  input  [31:0] I_1_1_2,
  input  [31:0] I_1_2_0,
  input  [31:0] I_1_2_1,
  input  [31:0] I_1_2_2,
  input  [31:0] I_2_0_0,
  input  [31:0] I_2_0_1,
  input  [31:0] I_2_0_2,
  input  [31:0] I_2_1_0,
  input  [31:0] I_2_1_1,
  input  [31:0] I_2_1_2,
  input  [31:0] I_2_2_0,
  input  [31:0] I_2_2_1,
  input  [31:0] I_2_2_2,
  input  [31:0] I_3_0_0,
  input  [31:0] I_3_0_1,
  input  [31:0] I_3_0_2,
  input  [31:0] I_3_1_0,
  input  [31:0] I_3_1_1,
  input  [31:0] I_3_1_2,
  input  [31:0] I_3_2_0,
  input  [31:0] I_3_2_1,
  input  [31:0] I_3_2_2,
  input  [31:0] I_4_0_0,
  input  [31:0] I_4_0_1,
  input  [31:0] I_4_0_2,
  input  [31:0] I_4_1_0,
  input  [31:0] I_4_1_1,
  input  [31:0] I_4_1_2,
  input  [31:0] I_4_2_0,
  input  [31:0] I_4_2_1,
  input  [31:0] I_4_2_2,
  input  [31:0] I_5_0_0,
  input  [31:0] I_5_0_1,
  input  [31:0] I_5_0_2,
  input  [31:0] I_5_1_0,
  input  [31:0] I_5_1_1,
  input  [31:0] I_5_1_2,
  input  [31:0] I_5_2_0,
  input  [31:0] I_5_2_1,
  input  [31:0] I_5_2_2,
  input  [31:0] I_6_0_0,
  input  [31:0] I_6_0_1,
  input  [31:0] I_6_0_2,
  input  [31:0] I_6_1_0,
  input  [31:0] I_6_1_1,
  input  [31:0] I_6_1_2,
  input  [31:0] I_6_2_0,
  input  [31:0] I_6_2_1,
  input  [31:0] I_6_2_2,
  input  [31:0] I_7_0_0,
  input  [31:0] I_7_0_1,
  input  [31:0] I_7_0_2,
  input  [31:0] I_7_1_0,
  input  [31:0] I_7_1_1,
  input  [31:0] I_7_1_2,
  input  [31:0] I_7_2_0,
  input  [31:0] I_7_2_1,
  input  [31:0] I_7_2_2,
  output [31:0] O_0_0_0,
  output [31:0] O_1_0_0,
  output [31:0] O_2_0_0,
  output [31:0] O_3_0_0,
  output [31:0] O_4_0_0,
  output [31:0] O_5_0_0,
  output [31:0] O_6_0_0,
  output [31:0] O_7_0_0
);
  wire  op_clock; // @[MapT.scala 8:20]
  wire  op_reset; // @[MapT.scala 8:20]
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_0_0; // @[MapT.scala 8:20]
  MapS_59 op ( // @[MapT.scala 8:20]
    .clock(op_clock),
    .reset(op_reset),
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0(op_I_0_0_0),
    .I_0_0_1(op_I_0_0_1),
    .I_0_0_2(op_I_0_0_2),
    .I_0_1_0(op_I_0_1_0),
    .I_0_1_1(op_I_0_1_1),
    .I_0_1_2(op_I_0_1_2),
    .I_0_2_0(op_I_0_2_0),
    .I_0_2_1(op_I_0_2_1),
    .I_0_2_2(op_I_0_2_2),
    .I_1_0_0(op_I_1_0_0),
    .I_1_0_1(op_I_1_0_1),
    .I_1_0_2(op_I_1_0_2),
    .I_1_1_0(op_I_1_1_0),
    .I_1_1_1(op_I_1_1_1),
    .I_1_1_2(op_I_1_1_2),
    .I_1_2_0(op_I_1_2_0),
    .I_1_2_1(op_I_1_2_1),
    .I_1_2_2(op_I_1_2_2),
    .I_2_0_0(op_I_2_0_0),
    .I_2_0_1(op_I_2_0_1),
    .I_2_0_2(op_I_2_0_2),
    .I_2_1_0(op_I_2_1_0),
    .I_2_1_1(op_I_2_1_1),
    .I_2_1_2(op_I_2_1_2),
    .I_2_2_0(op_I_2_2_0),
    .I_2_2_1(op_I_2_2_1),
    .I_2_2_2(op_I_2_2_2),
    .I_3_0_0(op_I_3_0_0),
    .I_3_0_1(op_I_3_0_1),
    .I_3_0_2(op_I_3_0_2),
    .I_3_1_0(op_I_3_1_0),
    .I_3_1_1(op_I_3_1_1),
    .I_3_1_2(op_I_3_1_2),
    .I_3_2_0(op_I_3_2_0),
    .I_3_2_1(op_I_3_2_1),
    .I_3_2_2(op_I_3_2_2),
    .I_4_0_0(op_I_4_0_0),
    .I_4_0_1(op_I_4_0_1),
    .I_4_0_2(op_I_4_0_2),
    .I_4_1_0(op_I_4_1_0),
    .I_4_1_1(op_I_4_1_1),
    .I_4_1_2(op_I_4_1_2),
    .I_4_2_0(op_I_4_2_0),
    .I_4_2_1(op_I_4_2_1),
    .I_4_2_2(op_I_4_2_2),
    .I_5_0_0(op_I_5_0_0),
    .I_5_0_1(op_I_5_0_1),
    .I_5_0_2(op_I_5_0_2),
    .I_5_1_0(op_I_5_1_0),
    .I_5_1_1(op_I_5_1_1),
    .I_5_1_2(op_I_5_1_2),
    .I_5_2_0(op_I_5_2_0),
    .I_5_2_1(op_I_5_2_1),
    .I_5_2_2(op_I_5_2_2),
    .I_6_0_0(op_I_6_0_0),
    .I_6_0_1(op_I_6_0_1),
    .I_6_0_2(op_I_6_0_2),
    .I_6_1_0(op_I_6_1_0),
    .I_6_1_1(op_I_6_1_1),
    .I_6_1_2(op_I_6_1_2),
    .I_6_2_0(op_I_6_2_0),
    .I_6_2_1(op_I_6_2_1),
    .I_6_2_2(op_I_6_2_2),
    .I_7_0_0(op_I_7_0_0),
    .I_7_0_1(op_I_7_0_1),
    .I_7_0_2(op_I_7_0_2),
    .I_7_1_0(op_I_7_1_0),
    .I_7_1_1(op_I_7_1_1),
    .I_7_1_2(op_I_7_1_2),
    .I_7_2_0(op_I_7_2_0),
    .I_7_2_1(op_I_7_2_1),
    .I_7_2_2(op_I_7_2_2),
    .O_0_0_0(op_O_0_0_0),
    .O_1_0_0(op_O_1_0_0),
    .O_2_0_0(op_O_2_0_0),
    .O_3_0_0(op_O_3_0_0),
    .O_4_0_0(op_O_4_0_0),
    .O_5_0_0(op_O_5_0_0),
    .O_6_0_0(op_O_6_0_0),
    .O_7_0_0(op_O_7_0_0)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0 = op_O_0_0_0; // @[MapT.scala 15:7]
  assign O_1_0_0 = op_O_1_0_0; // @[MapT.scala 15:7]
  assign O_2_0_0 = op_O_2_0_0; // @[MapT.scala 15:7]
  assign O_3_0_0 = op_O_3_0_0; // @[MapT.scala 15:7]
  assign O_4_0_0 = op_O_4_0_0; // @[MapT.scala 15:7]
  assign O_5_0_0 = op_O_5_0_0; // @[MapT.scala 15:7]
  assign O_6_0_0 = op_O_6_0_0; // @[MapT.scala 15:7]
  assign O_7_0_0 = op_O_7_0_0; // @[MapT.scala 15:7]
  assign op_clock = clock;
  assign op_reset = reset;
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0 = I_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_1 = I_0_0_1; // @[MapT.scala 14:10]
  assign op_I_0_0_2 = I_0_0_2; // @[MapT.scala 14:10]
  assign op_I_0_1_0 = I_0_1_0; // @[MapT.scala 14:10]
  assign op_I_0_1_1 = I_0_1_1; // @[MapT.scala 14:10]
  assign op_I_0_1_2 = I_0_1_2; // @[MapT.scala 14:10]
  assign op_I_0_2_0 = I_0_2_0; // @[MapT.scala 14:10]
  assign op_I_0_2_1 = I_0_2_1; // @[MapT.scala 14:10]
  assign op_I_0_2_2 = I_0_2_2; // @[MapT.scala 14:10]
  assign op_I_1_0_0 = I_1_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_1 = I_1_0_1; // @[MapT.scala 14:10]
  assign op_I_1_0_2 = I_1_0_2; // @[MapT.scala 14:10]
  assign op_I_1_1_0 = I_1_1_0; // @[MapT.scala 14:10]
  assign op_I_1_1_1 = I_1_1_1; // @[MapT.scala 14:10]
  assign op_I_1_1_2 = I_1_1_2; // @[MapT.scala 14:10]
  assign op_I_1_2_0 = I_1_2_0; // @[MapT.scala 14:10]
  assign op_I_1_2_1 = I_1_2_1; // @[MapT.scala 14:10]
  assign op_I_1_2_2 = I_1_2_2; // @[MapT.scala 14:10]
  assign op_I_2_0_0 = I_2_0_0; // @[MapT.scala 14:10]
  assign op_I_2_0_1 = I_2_0_1; // @[MapT.scala 14:10]
  assign op_I_2_0_2 = I_2_0_2; // @[MapT.scala 14:10]
  assign op_I_2_1_0 = I_2_1_0; // @[MapT.scala 14:10]
  assign op_I_2_1_1 = I_2_1_1; // @[MapT.scala 14:10]
  assign op_I_2_1_2 = I_2_1_2; // @[MapT.scala 14:10]
  assign op_I_2_2_0 = I_2_2_0; // @[MapT.scala 14:10]
  assign op_I_2_2_1 = I_2_2_1; // @[MapT.scala 14:10]
  assign op_I_2_2_2 = I_2_2_2; // @[MapT.scala 14:10]
  assign op_I_3_0_0 = I_3_0_0; // @[MapT.scala 14:10]
  assign op_I_3_0_1 = I_3_0_1; // @[MapT.scala 14:10]
  assign op_I_3_0_2 = I_3_0_2; // @[MapT.scala 14:10]
  assign op_I_3_1_0 = I_3_1_0; // @[MapT.scala 14:10]
  assign op_I_3_1_1 = I_3_1_1; // @[MapT.scala 14:10]
  assign op_I_3_1_2 = I_3_1_2; // @[MapT.scala 14:10]
  assign op_I_3_2_0 = I_3_2_0; // @[MapT.scala 14:10]
  assign op_I_3_2_1 = I_3_2_1; // @[MapT.scala 14:10]
  assign op_I_3_2_2 = I_3_2_2; // @[MapT.scala 14:10]
  assign op_I_4_0_0 = I_4_0_0; // @[MapT.scala 14:10]
  assign op_I_4_0_1 = I_4_0_1; // @[MapT.scala 14:10]
  assign op_I_4_0_2 = I_4_0_2; // @[MapT.scala 14:10]
  assign op_I_4_1_0 = I_4_1_0; // @[MapT.scala 14:10]
  assign op_I_4_1_1 = I_4_1_1; // @[MapT.scala 14:10]
  assign op_I_4_1_2 = I_4_1_2; // @[MapT.scala 14:10]
  assign op_I_4_2_0 = I_4_2_0; // @[MapT.scala 14:10]
  assign op_I_4_2_1 = I_4_2_1; // @[MapT.scala 14:10]
  assign op_I_4_2_2 = I_4_2_2; // @[MapT.scala 14:10]
  assign op_I_5_0_0 = I_5_0_0; // @[MapT.scala 14:10]
  assign op_I_5_0_1 = I_5_0_1; // @[MapT.scala 14:10]
  assign op_I_5_0_2 = I_5_0_2; // @[MapT.scala 14:10]
  assign op_I_5_1_0 = I_5_1_0; // @[MapT.scala 14:10]
  assign op_I_5_1_1 = I_5_1_1; // @[MapT.scala 14:10]
  assign op_I_5_1_2 = I_5_1_2; // @[MapT.scala 14:10]
  assign op_I_5_2_0 = I_5_2_0; // @[MapT.scala 14:10]
  assign op_I_5_2_1 = I_5_2_1; // @[MapT.scala 14:10]
  assign op_I_5_2_2 = I_5_2_2; // @[MapT.scala 14:10]
  assign op_I_6_0_0 = I_6_0_0; // @[MapT.scala 14:10]
  assign op_I_6_0_1 = I_6_0_1; // @[MapT.scala 14:10]
  assign op_I_6_0_2 = I_6_0_2; // @[MapT.scala 14:10]
  assign op_I_6_1_0 = I_6_1_0; // @[MapT.scala 14:10]
  assign op_I_6_1_1 = I_6_1_1; // @[MapT.scala 14:10]
  assign op_I_6_1_2 = I_6_1_2; // @[MapT.scala 14:10]
  assign op_I_6_2_0 = I_6_2_0; // @[MapT.scala 14:10]
  assign op_I_6_2_1 = I_6_2_1; // @[MapT.scala 14:10]
  assign op_I_6_2_2 = I_6_2_2; // @[MapT.scala 14:10]
  assign op_I_7_0_0 = I_7_0_0; // @[MapT.scala 14:10]
  assign op_I_7_0_1 = I_7_0_1; // @[MapT.scala 14:10]
  assign op_I_7_0_2 = I_7_0_2; // @[MapT.scala 14:10]
  assign op_I_7_1_0 = I_7_1_0; // @[MapT.scala 14:10]
  assign op_I_7_1_1 = I_7_1_1; // @[MapT.scala 14:10]
  assign op_I_7_1_2 = I_7_1_2; // @[MapT.scala 14:10]
  assign op_I_7_2_0 = I_7_2_0; // @[MapT.scala 14:10]
  assign op_I_7_2_1 = I_7_2_1; // @[MapT.scala 14:10]
  assign op_I_7_2_2 = I_7_2_2; // @[MapT.scala 14:10]
endmodule
module Passthrough_4(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0_0,
  input  [31:0] I_1_0_0,
  input  [31:0] I_2_0_0,
  input  [31:0] I_3_0_0,
  input  [31:0] I_4_0_0,
  input  [31:0] I_5_0_0,
  input  [31:0] I_6_0_0,
  input  [31:0] I_7_0_0,
  output [31:0] O_0_0,
  output [31:0] O_1_0,
  output [31:0] O_2_0,
  output [31:0] O_3_0,
  output [31:0] O_4_0,
  output [31:0] O_5_0,
  output [31:0] O_6_0,
  output [31:0] O_7_0
);
  assign valid_down = valid_up; // @[Passthrough.scala 18:14]
  assign O_0_0 = I_0_0_0; // @[Passthrough.scala 17:68]
  assign O_1_0 = I_1_0_0; // @[Passthrough.scala 17:68]
  assign O_2_0 = I_2_0_0; // @[Passthrough.scala 17:68]
  assign O_3_0 = I_3_0_0; // @[Passthrough.scala 17:68]
  assign O_4_0 = I_4_0_0; // @[Passthrough.scala 17:68]
  assign O_5_0 = I_5_0_0; // @[Passthrough.scala 17:68]
  assign O_6_0 = I_6_0_0; // @[Passthrough.scala 17:68]
  assign O_7_0 = I_7_0_0; // @[Passthrough.scala 17:68]
endmodule
module Passthrough_5(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0,
  input  [31:0] I_1_0,
  input  [31:0] I_2_0,
  input  [31:0] I_3_0,
  input  [31:0] I_4_0,
  input  [31:0] I_5_0,
  input  [31:0] I_6_0,
  input  [31:0] I_7_0,
  output [31:0] O_0,
  output [31:0] O_1,
  output [31:0] O_2,
  output [31:0] O_3,
  output [31:0] O_4,
  output [31:0] O_5,
  output [31:0] O_6,
  output [31:0] O_7
);
  assign valid_down = valid_up; // @[Passthrough.scala 18:14]
  assign O_0 = I_0_0; // @[Passthrough.scala 17:68]
  assign O_1 = I_1_0; // @[Passthrough.scala 17:68]
  assign O_2 = I_2_0; // @[Passthrough.scala 17:68]
  assign O_3 = I_3_0; // @[Passthrough.scala 17:68]
  assign O_4 = I_4_0; // @[Passthrough.scala 17:68]
  assign O_5 = I_5_0; // @[Passthrough.scala 17:68]
  assign O_6 = I_6_0; // @[Passthrough.scala 17:68]
  assign O_7 = I_7_0; // @[Passthrough.scala 17:68]
endmodule
module FIFO_9(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0,
  input  [31:0] I_1,
  input  [31:0] I_2,
  input  [31:0] I_3,
  input  [31:0] I_4,
  input  [31:0] I_5,
  input  [31:0] I_6,
  input  [31:0] I_7,
  output [31:0] O_0,
  output [31:0] O_1,
  output [31:0] O_2,
  output [31:0] O_3,
  output [31:0] O_4,
  output [31:0] O_5,
  output [31:0] O_6,
  output [31:0] O_7
);
  reg [31:0] _T__0 [0:16]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_0;
  wire [31:0] _T__0__T_15_data; // @[FIFO.scala 23:33]
  wire [4:0] _T__0__T_15_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_1;
  wire [31:0] _T__0__T_5_data; // @[FIFO.scala 23:33]
  wire [4:0] _T__0__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__0__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__0__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__0__T_15_en_pipe_0;
  reg [31:0] _RAND_2;
  reg [4:0] _T__0__T_15_addr_pipe_0;
  reg [31:0] _RAND_3;
  reg [31:0] _T__1 [0:16]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_4;
  wire [31:0] _T__1__T_15_data; // @[FIFO.scala 23:33]
  wire [4:0] _T__1__T_15_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_5;
  wire [31:0] _T__1__T_5_data; // @[FIFO.scala 23:33]
  wire [4:0] _T__1__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__1__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__1__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__1__T_15_en_pipe_0;
  reg [31:0] _RAND_6;
  reg [4:0] _T__1__T_15_addr_pipe_0;
  reg [31:0] _RAND_7;
  reg [31:0] _T__2 [0:16]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_8;
  wire [31:0] _T__2__T_15_data; // @[FIFO.scala 23:33]
  wire [4:0] _T__2__T_15_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_9;
  wire [31:0] _T__2__T_5_data; // @[FIFO.scala 23:33]
  wire [4:0] _T__2__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__2__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__2__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__2__T_15_en_pipe_0;
  reg [31:0] _RAND_10;
  reg [4:0] _T__2__T_15_addr_pipe_0;
  reg [31:0] _RAND_11;
  reg [31:0] _T__3 [0:16]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_12;
  wire [31:0] _T__3__T_15_data; // @[FIFO.scala 23:33]
  wire [4:0] _T__3__T_15_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_13;
  wire [31:0] _T__3__T_5_data; // @[FIFO.scala 23:33]
  wire [4:0] _T__3__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__3__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__3__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__3__T_15_en_pipe_0;
  reg [31:0] _RAND_14;
  reg [4:0] _T__3__T_15_addr_pipe_0;
  reg [31:0] _RAND_15;
  reg [31:0] _T__4 [0:16]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_16;
  wire [31:0] _T__4__T_15_data; // @[FIFO.scala 23:33]
  wire [4:0] _T__4__T_15_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_17;
  wire [31:0] _T__4__T_5_data; // @[FIFO.scala 23:33]
  wire [4:0] _T__4__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__4__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__4__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__4__T_15_en_pipe_0;
  reg [31:0] _RAND_18;
  reg [4:0] _T__4__T_15_addr_pipe_0;
  reg [31:0] _RAND_19;
  reg [31:0] _T__5 [0:16]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_20;
  wire [31:0] _T__5__T_15_data; // @[FIFO.scala 23:33]
  wire [4:0] _T__5__T_15_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_21;
  wire [31:0] _T__5__T_5_data; // @[FIFO.scala 23:33]
  wire [4:0] _T__5__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__5__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__5__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__5__T_15_en_pipe_0;
  reg [31:0] _RAND_22;
  reg [4:0] _T__5__T_15_addr_pipe_0;
  reg [31:0] _RAND_23;
  reg [31:0] _T__6 [0:16]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_24;
  wire [31:0] _T__6__T_15_data; // @[FIFO.scala 23:33]
  wire [4:0] _T__6__T_15_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_25;
  wire [31:0] _T__6__T_5_data; // @[FIFO.scala 23:33]
  wire [4:0] _T__6__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__6__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__6__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__6__T_15_en_pipe_0;
  reg [31:0] _RAND_26;
  reg [4:0] _T__6__T_15_addr_pipe_0;
  reg [31:0] _RAND_27;
  reg [31:0] _T__7 [0:16]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_28;
  wire [31:0] _T__7__T_15_data; // @[FIFO.scala 23:33]
  wire [4:0] _T__7__T_15_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_29;
  wire [31:0] _T__7__T_5_data; // @[FIFO.scala 23:33]
  wire [4:0] _T__7__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__7__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__7__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__7__T_15_en_pipe_0;
  reg [31:0] _RAND_30;
  reg [4:0] _T__7__T_15_addr_pipe_0;
  reg [31:0] _RAND_31;
  reg [4:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_32;
  reg [4:0] value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_33;
  reg [4:0] value_2; // @[Counter.scala 29:33]
  reg [31:0] _RAND_34;
  wire  _T_1; // @[FIFO.scala 33:46]
  wire  _T_2; // @[Counter.scala 37:24]
  wire [4:0] _T_4; // @[Counter.scala 38:22]
  wire  _T_6; // @[FIFO.scala 38:39]
  wire [4:0] _T_9; // @[Counter.scala 38:22]
  wire  _T_10; // @[FIFO.scala 42:39]
  wire  _T_16; // @[Counter.scala 37:24]
  wire [4:0] _T_18; // @[Counter.scala 38:22]
  wire  _GEN_8; // @[FIFO.scala 42:57]
  assign _T__0__T_15_addr = _T__0__T_15_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__0__T_15_data = _T__0[_T__0__T_15_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__0__T_15_data = _T__0__T_15_addr >= 5'h11 ? _RAND_1[31:0] : _T__0[_T__0__T_15_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__0__T_5_data = I_0;
  assign _T__0__T_5_addr = value_2;
  assign _T__0__T_5_mask = 1'h1;
  assign _T__0__T_5_en = valid_up;
  assign _T__1__T_15_addr = _T__1__T_15_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__1__T_15_data = _T__1[_T__1__T_15_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__1__T_15_data = _T__1__T_15_addr >= 5'h11 ? _RAND_5[31:0] : _T__1[_T__1__T_15_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__1__T_5_data = I_1;
  assign _T__1__T_5_addr = value_2;
  assign _T__1__T_5_mask = 1'h1;
  assign _T__1__T_5_en = valid_up;
  assign _T__2__T_15_addr = _T__2__T_15_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__2__T_15_data = _T__2[_T__2__T_15_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__2__T_15_data = _T__2__T_15_addr >= 5'h11 ? _RAND_9[31:0] : _T__2[_T__2__T_15_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__2__T_5_data = I_2;
  assign _T__2__T_5_addr = value_2;
  assign _T__2__T_5_mask = 1'h1;
  assign _T__2__T_5_en = valid_up;
  assign _T__3__T_15_addr = _T__3__T_15_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__3__T_15_data = _T__3[_T__3__T_15_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__3__T_15_data = _T__3__T_15_addr >= 5'h11 ? _RAND_13[31:0] : _T__3[_T__3__T_15_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__3__T_5_data = I_3;
  assign _T__3__T_5_addr = value_2;
  assign _T__3__T_5_mask = 1'h1;
  assign _T__3__T_5_en = valid_up;
  assign _T__4__T_15_addr = _T__4__T_15_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__4__T_15_data = _T__4[_T__4__T_15_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__4__T_15_data = _T__4__T_15_addr >= 5'h11 ? _RAND_17[31:0] : _T__4[_T__4__T_15_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__4__T_5_data = I_4;
  assign _T__4__T_5_addr = value_2;
  assign _T__4__T_5_mask = 1'h1;
  assign _T__4__T_5_en = valid_up;
  assign _T__5__T_15_addr = _T__5__T_15_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__5__T_15_data = _T__5[_T__5__T_15_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__5__T_15_data = _T__5__T_15_addr >= 5'h11 ? _RAND_21[31:0] : _T__5[_T__5__T_15_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__5__T_5_data = I_5;
  assign _T__5__T_5_addr = value_2;
  assign _T__5__T_5_mask = 1'h1;
  assign _T__5__T_5_en = valid_up;
  assign _T__6__T_15_addr = _T__6__T_15_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__6__T_15_data = _T__6[_T__6__T_15_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__6__T_15_data = _T__6__T_15_addr >= 5'h11 ? _RAND_25[31:0] : _T__6[_T__6__T_15_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__6__T_5_data = I_6;
  assign _T__6__T_5_addr = value_2;
  assign _T__6__T_5_mask = 1'h1;
  assign _T__6__T_5_en = valid_up;
  assign _T__7__T_15_addr = _T__7__T_15_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__7__T_15_data = _T__7[_T__7__T_15_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__7__T_15_data = _T__7__T_15_addr >= 5'h11 ? _RAND_29[31:0] : _T__7[_T__7__T_15_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__7__T_5_data = I_7;
  assign _T__7__T_5_addr = value_2;
  assign _T__7__T_5_mask = 1'h1;
  assign _T__7__T_5_en = valid_up;
  assign _T_1 = value == 5'h10; // @[FIFO.scala 33:46]
  assign _T_2 = value_2 == 5'h10; // @[Counter.scala 37:24]
  assign _T_4 = value_2 + 5'h1; // @[Counter.scala 38:22]
  assign _T_6 = value < 5'h10; // @[FIFO.scala 38:39]
  assign _T_9 = value + 5'h1; // @[Counter.scala 38:22]
  assign _T_10 = value >= 5'hf; // @[FIFO.scala 42:39]
  assign _T_16 = value_1 == 5'h10; // @[Counter.scala 37:24]
  assign _T_18 = value_1 + 5'h1; // @[Counter.scala 38:22]
  assign _GEN_8 = _T_10 & _T_10; // @[FIFO.scala 42:57]
  assign valid_down = value == 5'h10; // @[FIFO.scala 33:16]
  assign O_0 = _T__0__T_15_data; // @[FIFO.scala 43:11]
  assign O_1 = _T__1__T_15_data; // @[FIFO.scala 43:11]
  assign O_2 = _T__2__T_15_data; // @[FIFO.scala 43:11]
  assign O_3 = _T__3__T_15_data; // @[FIFO.scala 43:11]
  assign O_4 = _T__4__T_15_data; // @[FIFO.scala 43:11]
  assign O_5 = _T__5__T_15_data; // @[FIFO.scala 43:11]
  assign O_6 = _T__6__T_15_data; // @[FIFO.scala 43:11]
  assign O_7 = _T__7__T_15_data; // @[FIFO.scala 43:11]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 17; initvar = initvar+1)
    _T__0[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T__0__T_15_en_pipe_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T__0__T_15_addr_pipe_0 = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 17; initvar = initvar+1)
    _T__1[initvar] = _RAND_4[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T__1__T_15_en_pipe_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T__1__T_15_addr_pipe_0 = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 17; initvar = initvar+1)
    _T__2[initvar] = _RAND_8[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_9 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T__2__T_15_en_pipe_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T__2__T_15_addr_pipe_0 = _RAND_11[4:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 17; initvar = initvar+1)
    _T__3[initvar] = _RAND_12[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_13 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T__3__T_15_en_pipe_0 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T__3__T_15_addr_pipe_0 = _RAND_15[4:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 17; initvar = initvar+1)
    _T__4[initvar] = _RAND_16[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_17 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T__4__T_15_en_pipe_0 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T__4__T_15_addr_pipe_0 = _RAND_19[4:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 17; initvar = initvar+1)
    _T__5[initvar] = _RAND_20[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_21 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T__5__T_15_en_pipe_0 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T__5__T_15_addr_pipe_0 = _RAND_23[4:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 17; initvar = initvar+1)
    _T__6[initvar] = _RAND_24[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_25 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T__6__T_15_en_pipe_0 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T__6__T_15_addr_pipe_0 = _RAND_27[4:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 17; initvar = initvar+1)
    _T__7[initvar] = _RAND_28[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_29 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T__7__T_15_en_pipe_0 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T__7__T_15_addr_pipe_0 = _RAND_31[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  value = _RAND_32[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  value_1 = _RAND_33[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  value_2 = _RAND_34[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T__0__T_5_en & _T__0__T_5_mask) begin
      _T__0[_T__0__T_5_addr] <= _T__0__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__0__T_15_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__0__T_15_addr_pipe_0 <= value_1;
    end
    if(_T__1__T_5_en & _T__1__T_5_mask) begin
      _T__1[_T__1__T_5_addr] <= _T__1__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__1__T_15_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__1__T_15_addr_pipe_0 <= value_1;
    end
    if(_T__2__T_5_en & _T__2__T_5_mask) begin
      _T__2[_T__2__T_5_addr] <= _T__2__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__2__T_15_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__2__T_15_addr_pipe_0 <= value_1;
    end
    if(_T__3__T_5_en & _T__3__T_5_mask) begin
      _T__3[_T__3__T_5_addr] <= _T__3__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__3__T_15_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__3__T_15_addr_pipe_0 <= value_1;
    end
    if(_T__4__T_5_en & _T__4__T_5_mask) begin
      _T__4[_T__4__T_5_addr] <= _T__4__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__4__T_15_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__4__T_15_addr_pipe_0 <= value_1;
    end
    if(_T__5__T_5_en & _T__5__T_5_mask) begin
      _T__5[_T__5__T_5_addr] <= _T__5__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__5__T_15_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__5__T_15_addr_pipe_0 <= value_1;
    end
    if(_T__6__T_5_en & _T__6__T_5_mask) begin
      _T__6[_T__6__T_5_addr] <= _T__6__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__6__T_15_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__6__T_15_addr_pipe_0 <= value_1;
    end
    if(_T__7__T_5_en & _T__7__T_5_mask) begin
      _T__7[_T__7__T_5_addr] <= _T__7__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__7__T_15_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__7__T_15_addr_pipe_0 <= value_1;
    end
    if (reset) begin
      value <= 5'h0;
    end else if (valid_up) begin
      if (_T_6) begin
        if (_T_1) begin
          value <= 5'h0;
        end else begin
          value <= _T_9;
        end
      end
    end
    if (reset) begin
      value_1 <= 5'h0;
    end else if (valid_up) begin
      if (_T_10) begin
        if (_T_16) begin
          value_1 <= 5'h0;
        end else begin
          value_1 <= _T_18;
        end
      end
    end
    if (reset) begin
      value_2 <= 5'h0;
    end else if (valid_up) begin
      if (_T_2) begin
        value_2 <= 5'h0;
      end else begin
        value_2 <= _T_4;
      end
    end
  end
endmodule
module FIFO_10(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I,
  output [31:0] O
);
  reg [31:0] _T [0:6]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_0;
  wire [31:0] _T__T_15_data; // @[FIFO.scala 23:33]
  wire [2:0] _T__T_15_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_1;
  wire [31:0] _T__T_5_data; // @[FIFO.scala 23:33]
  wire [2:0] _T__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__T_15_en_pipe_0;
  reg [31:0] _RAND_2;
  reg [2:0] _T__T_15_addr_pipe_0;
  reg [31:0] _RAND_3;
  reg [2:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_4;
  reg [2:0] value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  reg [2:0] value_2; // @[Counter.scala 29:33]
  reg [31:0] _RAND_6;
  wire  _T_1; // @[FIFO.scala 33:46]
  wire  _T_2; // @[Counter.scala 37:24]
  wire [2:0] _T_4; // @[Counter.scala 38:22]
  wire  _T_6; // @[FIFO.scala 38:39]
  wire [2:0] _T_9; // @[Counter.scala 38:22]
  wire  _T_10; // @[FIFO.scala 42:39]
  wire  _T_16; // @[Counter.scala 37:24]
  wire [2:0] _T_18; // @[Counter.scala 38:22]
  wire  _GEN_8; // @[FIFO.scala 42:57]
  assign _T__T_15_addr = _T__T_15_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__T_15_data = _T[_T__T_15_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__T_15_data = _T__T_15_addr >= 3'h7 ? _RAND_1[31:0] : _T[_T__T_15_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__T_5_data = I;
  assign _T__T_5_addr = value_2;
  assign _T__T_5_mask = 1'h1;
  assign _T__T_5_en = valid_up;
  assign _T_1 = value == 3'h6; // @[FIFO.scala 33:46]
  assign _T_2 = value_2 == 3'h6; // @[Counter.scala 37:24]
  assign _T_4 = value_2 + 3'h1; // @[Counter.scala 38:22]
  assign _T_6 = value < 3'h6; // @[FIFO.scala 38:39]
  assign _T_9 = value + 3'h1; // @[Counter.scala 38:22]
  assign _T_10 = value >= 3'h5; // @[FIFO.scala 42:39]
  assign _T_16 = value_1 == 3'h6; // @[Counter.scala 37:24]
  assign _T_18 = value_1 + 3'h1; // @[Counter.scala 38:22]
  assign _GEN_8 = _T_10 & _T_10; // @[FIFO.scala 42:57]
  assign valid_down = value == 3'h6; // @[FIFO.scala 33:16]
  assign O = _T__T_15_data; // @[FIFO.scala 43:11]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 7; initvar = initvar+1)
    _T[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T__T_15_en_pipe_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T__T_15_addr_pipe_0 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  value = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value_1 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  value_2 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T__T_5_en & _T__T_5_mask) begin
      _T[_T__T_5_addr] <= _T__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__T_15_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__T_15_addr_pipe_0 <= value_1;
    end
    if (reset) begin
      value <= 3'h0;
    end else if (valid_up) begin
      if (_T_6) begin
        if (_T_1) begin
          value <= 3'h0;
        end else begin
          value <= _T_9;
        end
      end
    end
    if (reset) begin
      value_1 <= 3'h0;
    end else if (valid_up) begin
      if (_T_10) begin
        if (_T_16) begin
          value_1 <= 3'h0;
        end else begin
          value_1 <= _T_18;
        end
      end
    end
    if (reset) begin
      value_2 <= 3'h0;
    end else if (valid_up) begin
      if (_T_2) begin
        value_2 <= 3'h0;
      end else begin
        value_2 <= _T_4;
      end
    end
  end
endmodule
module InitialDelayCounter_6(
  input   clock,
  input   reset,
  output  valid_down
);
  reg [4:0] value; // @[InitialDelayCounter.scala 8:34]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[InitialDelayCounter.scala 17:17]
  wire [4:0] _T_4; // @[InitialDelayCounter.scala 17:53]
  assign _T_1 = value < 5'h13; // @[InitialDelayCounter.scala 17:17]
  assign _T_4 = value + 5'h1; // @[InitialDelayCounter.scala 17:53]
  assign valid_down = value == 5'h13; // @[InitialDelayCounter.scala 16:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 5'h0;
    end else if (_T_1) begin
      value <= _T_4;
    end
  end
endmodule
module Sub(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_t0b,
  input  [31:0] I_t1b,
  output [31:0] O
);
  assign valid_down = valid_up; // @[Arithmetic.scala 139:14]
  assign O = I_t0b - I_t1b; // @[Arithmetic.scala 137:7]
endmodule
module Or(
  input   valid_up,
  output  valid_down,
  input   I_t0b,
  input   I_t1b,
  output  O
);
  assign valid_down = valid_up; // @[Arithmetic.scala 83:14]
  assign O = I_t0b | I_t1b; // @[Arithmetic.scala 82:5]
endmodule
module AtomTuple_33(
  input         valid_up,
  output        valid_down,
  input         I0,
  input  [31:0] I1_t0b,
  input  [31:0] I1_t1b,
  output        O_t0b,
  output [31:0] O_t1b_t0b,
  output [31:0] O_t1b_t1b
);
  assign valid_down = valid_up; // @[Tuple.scala 51:14]
  assign O_t0b = I0; // @[Tuple.scala 49:9]
  assign O_t1b_t0b = I1_t0b; // @[Tuple.scala 50:9]
  assign O_t1b_t1b = I1_t1b; // @[Tuple.scala 50:9]
endmodule
module If_3(
  input         valid_up,
  output        valid_down,
  input         I_t0b,
  input  [31:0] I_t1b_t0b,
  input  [31:0] I_t1b_t1b,
  output [31:0] O
);
  assign valid_down = valid_up; // @[Arithmetic.scala 525:14]
  assign O = I_t0b ? I_t1b_t0b : I_t1b_t1b; // @[Arithmetic.scala 523:9 Arithmetic.scala 524:20]
endmodule
module Module_9(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I0,
  input  [31:0] I1,
  output [31:0] O
);
  wire  n629_clock; // @[Top.scala 387:22]
  wire  n629_reset; // @[Top.scala 387:22]
  wire  n629_valid_up; // @[Top.scala 387:22]
  wire  n629_valid_down; // @[Top.scala 387:22]
  wire [31:0] n629_I; // @[Top.scala 387:22]
  wire [31:0] n629_O; // @[Top.scala 387:22]
  wire  InitialDelayCounter_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_valid_down; // @[Const.scala 11:33]
  wire  n608_valid_up; // @[Top.scala 391:22]
  wire  n608_valid_down; // @[Top.scala 391:22]
  wire [31:0] n608_I0; // @[Top.scala 391:22]
  wire [31:0] n608_I1; // @[Top.scala 391:22]
  wire [31:0] n608_O_t0b; // @[Top.scala 391:22]
  wire [31:0] n608_O_t1b; // @[Top.scala 391:22]
  wire  n609_valid_up; // @[Top.scala 395:22]
  wire  n609_valid_down; // @[Top.scala 395:22]
  wire [31:0] n609_I_t0b; // @[Top.scala 395:22]
  wire [31:0] n609_I_t1b; // @[Top.scala 395:22]
  wire [31:0] n609_O; // @[Top.scala 395:22]
  wire  n611_valid_up; // @[Top.scala 398:22]
  wire  n611_valid_down; // @[Top.scala 398:22]
  wire [31:0] n611_I0; // @[Top.scala 398:22]
  wire [31:0] n611_I1; // @[Top.scala 398:22]
  wire [31:0] n611_O_t0b; // @[Top.scala 398:22]
  wire [31:0] n611_O_t1b; // @[Top.scala 398:22]
  wire  n612_valid_up; // @[Top.scala 402:22]
  wire  n612_valid_down; // @[Top.scala 402:22]
  wire [31:0] n612_I_t0b; // @[Top.scala 402:22]
  wire [31:0] n612_I_t1b; // @[Top.scala 402:22]
  wire [31:0] n612_O; // @[Top.scala 402:22]
  wire  InitialDelayCounter_1_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_1_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_1_valid_down; // @[Const.scala 11:33]
  wire  n613_valid_up; // @[Top.scala 406:22]
  wire  n613_valid_down; // @[Top.scala 406:22]
  wire [31:0] n613_I0; // @[Top.scala 406:22]
  wire [31:0] n613_I1; // @[Top.scala 406:22]
  wire [31:0] n613_O_t0b; // @[Top.scala 406:22]
  wire [31:0] n613_O_t1b; // @[Top.scala 406:22]
  wire  n614_valid_up; // @[Top.scala 410:22]
  wire  n614_valid_down; // @[Top.scala 410:22]
  wire [31:0] n614_I_t0b; // @[Top.scala 410:22]
  wire [31:0] n614_I_t1b; // @[Top.scala 410:22]
  wire [31:0] n614_O; // @[Top.scala 410:22]
  wire  n616_valid_up; // @[Top.scala 413:22]
  wire  n616_valid_down; // @[Top.scala 413:22]
  wire [31:0] n616_I0; // @[Top.scala 413:22]
  wire [31:0] n616_I1; // @[Top.scala 413:22]
  wire [31:0] n616_O_t0b; // @[Top.scala 413:22]
  wire [31:0] n616_O_t1b; // @[Top.scala 413:22]
  wire  n617_valid_up; // @[Top.scala 417:22]
  wire  n617_valid_down; // @[Top.scala 417:22]
  wire [31:0] n617_I_t0b; // @[Top.scala 417:22]
  wire [31:0] n617_I_t1b; // @[Top.scala 417:22]
  wire [31:0] n617_O; // @[Top.scala 417:22]
  wire  n618_valid_up; // @[Top.scala 420:22]
  wire  n618_valid_down; // @[Top.scala 420:22]
  wire  n618_I0; // @[Top.scala 420:22]
  wire  n618_I1; // @[Top.scala 420:22]
  wire  n618_O_t0b; // @[Top.scala 420:22]
  wire  n618_O_t1b; // @[Top.scala 420:22]
  wire  n619_valid_up; // @[Top.scala 424:22]
  wire  n619_valid_down; // @[Top.scala 424:22]
  wire  n619_I_t0b; // @[Top.scala 424:22]
  wire  n619_I_t1b; // @[Top.scala 424:22]
  wire  n619_O; // @[Top.scala 424:22]
  wire  InitialDelayCounter_2_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_2_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_2_valid_down; // @[Const.scala 11:33]
  wire  n622_valid_up; // @[Top.scala 428:22]
  wire  n622_valid_down; // @[Top.scala 428:22]
  wire [31:0] n622_I0; // @[Top.scala 428:22]
  wire [31:0] n622_I1; // @[Top.scala 428:22]
  wire [31:0] n622_O_t0b; // @[Top.scala 428:22]
  wire [31:0] n622_O_t1b; // @[Top.scala 428:22]
  wire  n623_valid_up; // @[Top.scala 432:22]
  wire  n623_valid_down; // @[Top.scala 432:22]
  wire  n623_I0; // @[Top.scala 432:22]
  wire [31:0] n623_I1_t0b; // @[Top.scala 432:22]
  wire [31:0] n623_I1_t1b; // @[Top.scala 432:22]
  wire  n623_O_t0b; // @[Top.scala 432:22]
  wire [31:0] n623_O_t1b_t0b; // @[Top.scala 432:22]
  wire [31:0] n623_O_t1b_t1b; // @[Top.scala 432:22]
  wire  n624_valid_up; // @[Top.scala 436:22]
  wire  n624_valid_down; // @[Top.scala 436:22]
  wire  n624_I_t0b; // @[Top.scala 436:22]
  wire [31:0] n624_I_t1b_t0b; // @[Top.scala 436:22]
  wire [31:0] n624_I_t1b_t1b; // @[Top.scala 436:22]
  wire [31:0] n624_O; // @[Top.scala 436:22]
  wire  InitialDelayCounter_3_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_3_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_3_valid_down; // @[Const.scala 11:33]
  wire  n627_valid_up; // @[Top.scala 440:22]
  wire  n627_valid_down; // @[Top.scala 440:22]
  wire [31:0] n627_I0; // @[Top.scala 440:22]
  wire [7:0] n627_I1; // @[Top.scala 440:22]
  wire [31:0] n627_O_t0b; // @[Top.scala 440:22]
  wire [7:0] n627_O_t1b; // @[Top.scala 440:22]
  wire  n628_clock; // @[Top.scala 444:22]
  wire  n628_reset; // @[Top.scala 444:22]
  wire  n628_valid_up; // @[Top.scala 444:22]
  wire  n628_valid_down; // @[Top.scala 444:22]
  wire [31:0] n628_I_t0b; // @[Top.scala 444:22]
  wire [7:0] n628_I_t1b; // @[Top.scala 444:22]
  wire [31:0] n628_O; // @[Top.scala 444:22]
  wire  n630_valid_up; // @[Top.scala 447:22]
  wire  n630_valid_down; // @[Top.scala 447:22]
  wire [31:0] n630_I0; // @[Top.scala 447:22]
  wire [31:0] n630_I1; // @[Top.scala 447:22]
  wire [31:0] n630_O_t0b; // @[Top.scala 447:22]
  wire [31:0] n630_O_t1b; // @[Top.scala 447:22]
  wire  n631_valid_up; // @[Top.scala 451:22]
  wire  n631_valid_down; // @[Top.scala 451:22]
  wire [31:0] n631_I_t0b; // @[Top.scala 451:22]
  wire [31:0] n631_I_t1b; // @[Top.scala 451:22]
  wire [31:0] n631_O; // @[Top.scala 451:22]
  FIFO_10 n629 ( // @[Top.scala 387:22]
    .clock(n629_clock),
    .reset(n629_reset),
    .valid_up(n629_valid_up),
    .valid_down(n629_valid_down),
    .I(n629_I),
    .O(n629_O)
  );
  InitialDelayCounter_6 InitialDelayCounter ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_clock),
    .reset(InitialDelayCounter_reset),
    .valid_down(InitialDelayCounter_valid_down)
  );
  AtomTuple n608 ( // @[Top.scala 391:22]
    .valid_up(n608_valid_up),
    .valid_down(n608_valid_down),
    .I0(n608_I0),
    .I1(n608_I1),
    .O_t0b(n608_O_t0b),
    .O_t1b(n608_O_t1b)
  );
  Sub n609 ( // @[Top.scala 395:22]
    .valid_up(n609_valid_up),
    .valid_down(n609_valid_down),
    .I_t0b(n609_I_t0b),
    .I_t1b(n609_I_t1b),
    .O(n609_O)
  );
  AtomTuple n611 ( // @[Top.scala 398:22]
    .valid_up(n611_valid_up),
    .valid_down(n611_valid_down),
    .I0(n611_I0),
    .I1(n611_I1),
    .O_t0b(n611_O_t0b),
    .O_t1b(n611_O_t1b)
  );
  Lt n612 ( // @[Top.scala 402:22]
    .valid_up(n612_valid_up),
    .valid_down(n612_valid_down),
    .I_t0b(n612_I_t0b),
    .I_t1b(n612_I_t1b),
    .O(n612_O)
  );
  InitialDelayCounter_6 InitialDelayCounter_1 ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_1_clock),
    .reset(InitialDelayCounter_1_reset),
    .valid_down(InitialDelayCounter_1_valid_down)
  );
  AtomTuple n613 ( // @[Top.scala 406:22]
    .valid_up(n613_valid_up),
    .valid_down(n613_valid_down),
    .I0(n613_I0),
    .I1(n613_I1),
    .O_t0b(n613_O_t0b),
    .O_t1b(n613_O_t1b)
  );
  Sub n614 ( // @[Top.scala 410:22]
    .valid_up(n614_valid_up),
    .valid_down(n614_valid_down),
    .I_t0b(n614_I_t0b),
    .I_t1b(n614_I_t1b),
    .O(n614_O)
  );
  AtomTuple n616 ( // @[Top.scala 413:22]
    .valid_up(n616_valid_up),
    .valid_down(n616_valid_down),
    .I0(n616_I0),
    .I1(n616_I1),
    .O_t0b(n616_O_t0b),
    .O_t1b(n616_O_t1b)
  );
  Lt n617 ( // @[Top.scala 417:22]
    .valid_up(n617_valid_up),
    .valid_down(n617_valid_down),
    .I_t0b(n617_I_t0b),
    .I_t1b(n617_I_t1b),
    .O(n617_O)
  );
  AtomTuple_4 n618 ( // @[Top.scala 420:22]
    .valid_up(n618_valid_up),
    .valid_down(n618_valid_down),
    .I0(n618_I0),
    .I1(n618_I1),
    .O_t0b(n618_O_t0b),
    .O_t1b(n618_O_t1b)
  );
  Or n619 ( // @[Top.scala 424:22]
    .valid_up(n619_valid_up),
    .valid_down(n619_valid_down),
    .I_t0b(n619_I_t0b),
    .I_t1b(n619_I_t1b),
    .O(n619_O)
  );
  InitialDelayCounter_6 InitialDelayCounter_2 ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_2_clock),
    .reset(InitialDelayCounter_2_reset),
    .valid_down(InitialDelayCounter_2_valid_down)
  );
  AtomTuple n622 ( // @[Top.scala 428:22]
    .valid_up(n622_valid_up),
    .valid_down(n622_valid_down),
    .I0(n622_I0),
    .I1(n622_I1),
    .O_t0b(n622_O_t0b),
    .O_t1b(n622_O_t1b)
  );
  AtomTuple_33 n623 ( // @[Top.scala 432:22]
    .valid_up(n623_valid_up),
    .valid_down(n623_valid_down),
    .I0(n623_I0),
    .I1_t0b(n623_I1_t0b),
    .I1_t1b(n623_I1_t1b),
    .O_t0b(n623_O_t0b),
    .O_t1b_t0b(n623_O_t1b_t0b),
    .O_t1b_t1b(n623_O_t1b_t1b)
  );
  If_3 n624 ( // @[Top.scala 436:22]
    .valid_up(n624_valid_up),
    .valid_down(n624_valid_down),
    .I_t0b(n624_I_t0b),
    .I_t1b_t0b(n624_I_t1b_t0b),
    .I_t1b_t1b(n624_I_t1b_t1b),
    .O(n624_O)
  );
  InitialDelayCounter_6 InitialDelayCounter_3 ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_3_clock),
    .reset(InitialDelayCounter_3_reset),
    .valid_down(InitialDelayCounter_3_valid_down)
  );
  AtomTuple_26 n627 ( // @[Top.scala 440:22]
    .valid_up(n627_valid_up),
    .valid_down(n627_valid_down),
    .I0(n627_I0),
    .I1(n627_I1),
    .O_t0b(n627_O_t0b),
    .O_t1b(n627_O_t1b)
  );
  Div n628 ( // @[Top.scala 444:22]
    .clock(n628_clock),
    .reset(n628_reset),
    .valid_up(n628_valid_up),
    .valid_down(n628_valid_down),
    .I_t0b(n628_I_t0b),
    .I_t1b(n628_I_t1b),
    .O(n628_O)
  );
  AtomTuple n630 ( // @[Top.scala 447:22]
    .valid_up(n630_valid_up),
    .valid_down(n630_valid_down),
    .I0(n630_I0),
    .I1(n630_I1),
    .O_t0b(n630_O_t0b),
    .O_t1b(n630_O_t1b)
  );
  Add n631 ( // @[Top.scala 451:22]
    .valid_up(n631_valid_up),
    .valid_down(n631_valid_down),
    .I_t0b(n631_I_t0b),
    .I_t1b(n631_I_t1b),
    .O(n631_O)
  );
  assign valid_down = n631_valid_down; // @[Top.scala 455:16]
  assign O = n631_O; // @[Top.scala 454:7]
  assign n629_clock = clock;
  assign n629_reset = reset;
  assign n629_valid_up = valid_up; // @[Top.scala 389:19]
  assign n629_I = I1; // @[Top.scala 388:12]
  assign InitialDelayCounter_clock = clock;
  assign InitialDelayCounter_reset = reset;
  assign n608_valid_up = valid_up; // @[Top.scala 394:19]
  assign n608_I0 = I0; // @[Top.scala 392:13]
  assign n608_I1 = I1; // @[Top.scala 393:13]
  assign n609_valid_up = n608_valid_down; // @[Top.scala 397:19]
  assign n609_I_t0b = n608_O_t0b; // @[Top.scala 396:12]
  assign n609_I_t1b = n608_O_t1b; // @[Top.scala 396:12]
  assign n611_valid_up = InitialDelayCounter_valid_down & n609_valid_down; // @[Top.scala 401:19]
  assign n611_I0 = 32'hf; // @[Top.scala 399:13]
  assign n611_I1 = n609_O; // @[Top.scala 400:13]
  assign n612_valid_up = n611_valid_down; // @[Top.scala 404:19]
  assign n612_I_t0b = n611_O_t0b; // @[Top.scala 403:12]
  assign n612_I_t1b = n611_O_t1b; // @[Top.scala 403:12]
  assign InitialDelayCounter_1_clock = clock;
  assign InitialDelayCounter_1_reset = reset;
  assign n613_valid_up = valid_up; // @[Top.scala 409:19]
  assign n613_I0 = I1; // @[Top.scala 407:13]
  assign n613_I1 = I0; // @[Top.scala 408:13]
  assign n614_valid_up = n613_valid_down; // @[Top.scala 412:19]
  assign n614_I_t0b = n613_O_t0b; // @[Top.scala 411:12]
  assign n614_I_t1b = n613_O_t1b; // @[Top.scala 411:12]
  assign n616_valid_up = InitialDelayCounter_1_valid_down & n614_valid_down; // @[Top.scala 416:19]
  assign n616_I0 = 32'hf; // @[Top.scala 414:13]
  assign n616_I1 = n614_O; // @[Top.scala 415:13]
  assign n617_valid_up = n616_valid_down; // @[Top.scala 419:19]
  assign n617_I_t0b = n616_O_t0b; // @[Top.scala 418:12]
  assign n617_I_t1b = n616_O_t1b; // @[Top.scala 418:12]
  assign n618_valid_up = n612_valid_down & n617_valid_down; // @[Top.scala 423:19]
  assign n618_I0 = n612_O[0]; // @[Top.scala 421:13]
  assign n618_I1 = n617_O[0]; // @[Top.scala 422:13]
  assign n619_valid_up = n618_valid_down; // @[Top.scala 426:19]
  assign n619_I_t0b = n618_O_t0b; // @[Top.scala 425:12]
  assign n619_I_t1b = n618_O_t1b; // @[Top.scala 425:12]
  assign InitialDelayCounter_2_clock = clock;
  assign InitialDelayCounter_2_reset = reset;
  assign n622_valid_up = n614_valid_down & InitialDelayCounter_2_valid_down; // @[Top.scala 431:19]
  assign n622_I0 = n614_O; // @[Top.scala 429:13]
  assign n622_I1 = 32'h0; // @[Top.scala 430:13]
  assign n623_valid_up = n619_valid_down & n622_valid_down; // @[Top.scala 435:19]
  assign n623_I0 = n619_O; // @[Top.scala 433:13]
  assign n623_I1_t0b = n622_O_t0b; // @[Top.scala 434:13]
  assign n623_I1_t1b = n622_O_t1b; // @[Top.scala 434:13]
  assign n624_valid_up = n623_valid_down; // @[Top.scala 438:19]
  assign n624_I_t0b = n623_O_t0b; // @[Top.scala 437:12]
  assign n624_I_t1b_t0b = n623_O_t1b_t0b; // @[Top.scala 437:12]
  assign n624_I_t1b_t1b = n623_O_t1b_t1b; // @[Top.scala 437:12]
  assign InitialDelayCounter_3_clock = clock;
  assign InitialDelayCounter_3_reset = reset;
  assign n627_valid_up = n624_valid_down & InitialDelayCounter_3_valid_down; // @[Top.scala 443:19]
  assign n627_I0 = n624_O; // @[Top.scala 441:13]
  assign n627_I1 = 8'sh20; // @[Top.scala 442:13]
  assign n628_clock = clock;
  assign n628_reset = reset;
  assign n628_valid_up = n627_valid_down; // @[Top.scala 446:19]
  assign n628_I_t0b = n627_O_t0b; // @[Top.scala 445:12]
  assign n628_I_t1b = n627_O_t1b; // @[Top.scala 445:12]
  assign n630_valid_up = n629_valid_down & n628_valid_down; // @[Top.scala 450:19]
  assign n630_I0 = n629_O; // @[Top.scala 448:13]
  assign n630_I1 = n628_O; // @[Top.scala 449:13]
  assign n631_valid_up = n630_valid_down; // @[Top.scala 453:19]
  assign n631_I_t0b = n630_O_t0b; // @[Top.scala 452:12]
  assign n631_I_t1b = n630_O_t1b; // @[Top.scala 452:12]
endmodule
module Map2S_66(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0,
  input  [31:0] I0_1,
  input  [31:0] I0_2,
  input  [31:0] I0_3,
  input  [31:0] I0_4,
  input  [31:0] I0_5,
  input  [31:0] I0_6,
  input  [31:0] I0_7,
  input  [31:0] I1_0,
  input  [31:0] I1_1,
  input  [31:0] I1_2,
  input  [31:0] I1_3,
  input  [31:0] I1_4,
  input  [31:0] I1_5,
  input  [31:0] I1_6,
  input  [31:0] I1_7,
  output [31:0] O_0,
  output [31:0] O_1,
  output [31:0] O_2,
  output [31:0] O_3,
  output [31:0] O_4,
  output [31:0] O_5,
  output [31:0] O_6,
  output [31:0] O_7
);
  wire  fst_op_clock; // @[Map2S.scala 9:22]
  wire  fst_op_reset; // @[Map2S.scala 9:22]
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O; // @[Map2S.scala 9:22]
  wire  other_ops_0_clock; // @[Map2S.scala 10:86]
  wire  other_ops_0_reset; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O; // @[Map2S.scala 10:86]
  wire  other_ops_1_clock; // @[Map2S.scala 10:86]
  wire  other_ops_1_reset; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O; // @[Map2S.scala 10:86]
  wire  other_ops_2_clock; // @[Map2S.scala 10:86]
  wire  other_ops_2_reset; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O; // @[Map2S.scala 10:86]
  wire  other_ops_3_clock; // @[Map2S.scala 10:86]
  wire  other_ops_3_reset; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O; // @[Map2S.scala 10:86]
  wire  other_ops_4_clock; // @[Map2S.scala 10:86]
  wire  other_ops_4_reset; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O; // @[Map2S.scala 10:86]
  wire  other_ops_5_clock; // @[Map2S.scala 10:86]
  wire  other_ops_5_reset; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O; // @[Map2S.scala 10:86]
  wire  other_ops_6_clock; // @[Map2S.scala 10:86]
  wire  other_ops_6_reset; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  wire  _T_2; // @[Map2S.scala 26:83]
  wire  _T_3; // @[Map2S.scala 26:83]
  wire  _T_4; // @[Map2S.scala 26:83]
  wire  _T_5; // @[Map2S.scala 26:83]
  Module_9 fst_op ( // @[Map2S.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1(fst_op_I1),
    .O(fst_op_O)
  );
  Module_9 other_ops_0 ( // @[Map2S.scala 10:86]
    .clock(other_ops_0_clock),
    .reset(other_ops_0_reset),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0(other_ops_0_I0),
    .I1(other_ops_0_I1),
    .O(other_ops_0_O)
  );
  Module_9 other_ops_1 ( // @[Map2S.scala 10:86]
    .clock(other_ops_1_clock),
    .reset(other_ops_1_reset),
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0(other_ops_1_I0),
    .I1(other_ops_1_I1),
    .O(other_ops_1_O)
  );
  Module_9 other_ops_2 ( // @[Map2S.scala 10:86]
    .clock(other_ops_2_clock),
    .reset(other_ops_2_reset),
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0(other_ops_2_I0),
    .I1(other_ops_2_I1),
    .O(other_ops_2_O)
  );
  Module_9 other_ops_3 ( // @[Map2S.scala 10:86]
    .clock(other_ops_3_clock),
    .reset(other_ops_3_reset),
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I0(other_ops_3_I0),
    .I1(other_ops_3_I1),
    .O(other_ops_3_O)
  );
  Module_9 other_ops_4 ( // @[Map2S.scala 10:86]
    .clock(other_ops_4_clock),
    .reset(other_ops_4_reset),
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I0(other_ops_4_I0),
    .I1(other_ops_4_I1),
    .O(other_ops_4_O)
  );
  Module_9 other_ops_5 ( // @[Map2S.scala 10:86]
    .clock(other_ops_5_clock),
    .reset(other_ops_5_reset),
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I0(other_ops_5_I0),
    .I1(other_ops_5_I1),
    .O(other_ops_5_O)
  );
  Module_9 other_ops_6 ( // @[Map2S.scala 10:86]
    .clock(other_ops_6_clock),
    .reset(other_ops_6_reset),
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I0(other_ops_6_I0),
    .I1(other_ops_6_I1),
    .O(other_ops_6_O)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[Map2S.scala 26:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[Map2S.scala 26:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_5 & other_ops_6_valid_down; // @[Map2S.scala 26:14]
  assign O_0 = fst_op_O; // @[Map2S.scala 19:8]
  assign O_1 = other_ops_0_O; // @[Map2S.scala 24:12]
  assign O_2 = other_ops_1_O; // @[Map2S.scala 24:12]
  assign O_3 = other_ops_2_O; // @[Map2S.scala 24:12]
  assign O_4 = other_ops_3_O; // @[Map2S.scala 24:12]
  assign O_5 = other_ops_4_O; // @[Map2S.scala 24:12]
  assign O_6 = other_ops_5_O; // @[Map2S.scala 24:12]
  assign O_7 = other_ops_6_O; // @[Map2S.scala 24:12]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
  assign other_ops_0_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_0_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0 = I0_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I1 = I1_1; // @[Map2S.scala 23:43]
  assign other_ops_1_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_1_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0 = I0_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1 = I1_2; // @[Map2S.scala 23:43]
  assign other_ops_2_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_2_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0 = I0_3; // @[Map2S.scala 22:43]
  assign other_ops_2_I1 = I1_3; // @[Map2S.scala 23:43]
  assign other_ops_3_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_3_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_3_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_3_I0 = I0_4; // @[Map2S.scala 22:43]
  assign other_ops_3_I1 = I1_4; // @[Map2S.scala 23:43]
  assign other_ops_4_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_4_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_4_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_4_I0 = I0_5; // @[Map2S.scala 22:43]
  assign other_ops_4_I1 = I1_5; // @[Map2S.scala 23:43]
  assign other_ops_5_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_5_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_5_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_5_I0 = I0_6; // @[Map2S.scala 22:43]
  assign other_ops_5_I1 = I1_6; // @[Map2S.scala 23:43]
  assign other_ops_6_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_6_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_6_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_6_I0 = I0_7; // @[Map2S.scala 22:43]
  assign other_ops_6_I1 = I1_7; // @[Map2S.scala 23:43]
endmodule
module Map2T_18(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0,
  input  [31:0] I0_1,
  input  [31:0] I0_2,
  input  [31:0] I0_3,
  input  [31:0] I0_4,
  input  [31:0] I0_5,
  input  [31:0] I0_6,
  input  [31:0] I0_7,
  input  [31:0] I1_0,
  input  [31:0] I1_1,
  input  [31:0] I1_2,
  input  [31:0] I1_3,
  input  [31:0] I1_4,
  input  [31:0] I1_5,
  input  [31:0] I1_6,
  input  [31:0] I1_7,
  output [31:0] O_0,
  output [31:0] O_1,
  output [31:0] O_2,
  output [31:0] O_3,
  output [31:0] O_4,
  output [31:0] O_5,
  output [31:0] O_6,
  output [31:0] O_7
);
  wire  op_clock; // @[Map2T.scala 8:20]
  wire  op_reset; // @[Map2T.scala 8:20]
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_3; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_4; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_5; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_6; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_7; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7; // @[Map2T.scala 8:20]
  Map2S_66 op ( // @[Map2T.scala 8:20]
    .clock(op_clock),
    .reset(op_reset),
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0(op_I0_0),
    .I0_1(op_I0_1),
    .I0_2(op_I0_2),
    .I0_3(op_I0_3),
    .I0_4(op_I0_4),
    .I0_5(op_I0_5),
    .I0_6(op_I0_6),
    .I0_7(op_I0_7),
    .I1_0(op_I1_0),
    .I1_1(op_I1_1),
    .I1_2(op_I1_2),
    .I1_3(op_I1_3),
    .I1_4(op_I1_4),
    .I1_5(op_I1_5),
    .I1_6(op_I1_6),
    .I1_7(op_I1_7),
    .O_0(op_O_0),
    .O_1(op_O_1),
    .O_2(op_O_2),
    .O_3(op_O_3),
    .O_4(op_O_4),
    .O_5(op_O_5),
    .O_6(op_O_6),
    .O_7(op_O_7)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0 = op_O_0; // @[Map2T.scala 17:7]
  assign O_1 = op_O_1; // @[Map2T.scala 17:7]
  assign O_2 = op_O_2; // @[Map2T.scala 17:7]
  assign O_3 = op_O_3; // @[Map2T.scala 17:7]
  assign O_4 = op_O_4; // @[Map2T.scala 17:7]
  assign O_5 = op_O_5; // @[Map2T.scala 17:7]
  assign O_6 = op_O_6; // @[Map2T.scala 17:7]
  assign O_7 = op_O_7; // @[Map2T.scala 17:7]
  assign op_clock = clock;
  assign op_reset = reset;
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0 = I0_0; // @[Map2T.scala 15:11]
  assign op_I0_1 = I0_1; // @[Map2T.scala 15:11]
  assign op_I0_2 = I0_2; // @[Map2T.scala 15:11]
  assign op_I0_3 = I0_3; // @[Map2T.scala 15:11]
  assign op_I0_4 = I0_4; // @[Map2T.scala 15:11]
  assign op_I0_5 = I0_5; // @[Map2T.scala 15:11]
  assign op_I0_6 = I0_6; // @[Map2T.scala 15:11]
  assign op_I0_7 = I0_7; // @[Map2T.scala 15:11]
  assign op_I1_0 = I1_0; // @[Map2T.scala 16:11]
  assign op_I1_1 = I1_1; // @[Map2T.scala 16:11]
  assign op_I1_2 = I1_2; // @[Map2T.scala 16:11]
  assign op_I1_3 = I1_3; // @[Map2T.scala 16:11]
  assign op_I1_4 = I1_4; // @[Map2T.scala 16:11]
  assign op_I1_5 = I1_5; // @[Map2T.scala 16:11]
  assign op_I1_6 = I1_6; // @[Map2T.scala 16:11]
  assign op_I1_7 = I1_7; // @[Map2T.scala 16:11]
endmodule
module Snd_1(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_t1b_t0b,
  input  [31:0] I_t1b_t1b,
  output [31:0] O_t0b,
  output [31:0] O_t1b
);
  assign valid_down = valid_up; // @[Tuple.scala 67:14]
  assign O_t0b = I_t1b_t0b; // @[Tuple.scala 66:5]
  assign O_t1b = I_t1b_t1b; // @[Tuple.scala 66:5]
endmodule
module Fst_2(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_t0b,
  output [31:0] O
);
  assign valid_down = valid_up; // @[Tuple.scala 59:14]
  assign O = I_t0b; // @[Tuple.scala 58:5]
endmodule
module Module_10(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_t1b_t0b,
  input  [31:0] I_t1b_t1b,
  output [31:0] O
);
  wire  n634_valid_up; // @[Top.scala 461:22]
  wire  n634_valid_down; // @[Top.scala 461:22]
  wire [31:0] n634_I_t1b_t0b; // @[Top.scala 461:22]
  wire [31:0] n634_I_t1b_t1b; // @[Top.scala 461:22]
  wire [31:0] n634_O_t0b; // @[Top.scala 461:22]
  wire [31:0] n634_O_t1b; // @[Top.scala 461:22]
  wire  n635_valid_up; // @[Top.scala 464:22]
  wire  n635_valid_down; // @[Top.scala 464:22]
  wire [31:0] n635_I_t0b; // @[Top.scala 464:22]
  wire [31:0] n635_O; // @[Top.scala 464:22]
  Snd_1 n634 ( // @[Top.scala 461:22]
    .valid_up(n634_valid_up),
    .valid_down(n634_valid_down),
    .I_t1b_t0b(n634_I_t1b_t0b),
    .I_t1b_t1b(n634_I_t1b_t1b),
    .O_t0b(n634_O_t0b),
    .O_t1b(n634_O_t1b)
  );
  Fst_2 n635 ( // @[Top.scala 464:22]
    .valid_up(n635_valid_up),
    .valid_down(n635_valid_down),
    .I_t0b(n635_I_t0b),
    .O(n635_O)
  );
  assign valid_down = n635_valid_down; // @[Top.scala 468:16]
  assign O = n635_O; // @[Top.scala 467:7]
  assign n634_valid_up = valid_up; // @[Top.scala 463:19]
  assign n634_I_t1b_t0b = I_t1b_t0b; // @[Top.scala 462:12]
  assign n634_I_t1b_t1b = I_t1b_t1b; // @[Top.scala 462:12]
  assign n635_valid_up = n634_valid_down; // @[Top.scala 466:19]
  assign n635_I_t0b = n634_O_t0b; // @[Top.scala 465:12]
endmodule
module MapS_60(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_t1b_t0b,
  input  [31:0] I_0_t1b_t1b,
  input  [31:0] I_1_t1b_t0b,
  input  [31:0] I_1_t1b_t1b,
  input  [31:0] I_2_t1b_t0b,
  input  [31:0] I_2_t1b_t1b,
  input  [31:0] I_3_t1b_t0b,
  input  [31:0] I_3_t1b_t1b,
  input  [31:0] I_4_t1b_t0b,
  input  [31:0] I_4_t1b_t1b,
  input  [31:0] I_5_t1b_t0b,
  input  [31:0] I_5_t1b_t1b,
  input  [31:0] I_6_t1b_t0b,
  input  [31:0] I_6_t1b_t1b,
  input  [31:0] I_7_t1b_t0b,
  input  [31:0] I_7_t1b_t1b,
  output [31:0] O_0,
  output [31:0] O_1,
  output [31:0] O_2,
  output [31:0] O_3,
  output [31:0] O_4,
  output [31:0] O_5,
  output [31:0] O_6,
  output [31:0] O_7
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_t1b_t0b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_t1b_t1b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_t1b_t0b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_t1b_t1b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_O; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_t1b_t0b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_t1b_t1b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_O; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_t1b_t0b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_t1b_t1b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_O; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_t1b_t0b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_t1b_t1b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_O; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_t1b_t0b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_t1b_t1b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_O; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_t1b_t0b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_t1b_t1b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_O; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_t1b_t0b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_t1b_t1b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_O; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  wire  _T_1; // @[MapS.scala 23:83]
  wire  _T_2; // @[MapS.scala 23:83]
  wire  _T_3; // @[MapS.scala 23:83]
  wire  _T_4; // @[MapS.scala 23:83]
  wire  _T_5; // @[MapS.scala 23:83]
  Module_10 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_t1b_t0b(fst_op_I_t1b_t0b),
    .I_t1b_t1b(fst_op_I_t1b_t1b),
    .O(fst_op_O)
  );
  Module_10 other_ops_0 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_t1b_t0b(other_ops_0_I_t1b_t0b),
    .I_t1b_t1b(other_ops_0_I_t1b_t1b),
    .O(other_ops_0_O)
  );
  Module_10 other_ops_1 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_t1b_t0b(other_ops_1_I_t1b_t0b),
    .I_t1b_t1b(other_ops_1_I_t1b_t1b),
    .O(other_ops_1_O)
  );
  Module_10 other_ops_2 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I_t1b_t0b(other_ops_2_I_t1b_t0b),
    .I_t1b_t1b(other_ops_2_I_t1b_t1b),
    .O(other_ops_2_O)
  );
  Module_10 other_ops_3 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I_t1b_t0b(other_ops_3_I_t1b_t0b),
    .I_t1b_t1b(other_ops_3_I_t1b_t1b),
    .O(other_ops_3_O)
  );
  Module_10 other_ops_4 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I_t1b_t0b(other_ops_4_I_t1b_t0b),
    .I_t1b_t1b(other_ops_4_I_t1b_t1b),
    .O(other_ops_4_O)
  );
  Module_10 other_ops_5 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I_t1b_t0b(other_ops_5_I_t1b_t0b),
    .I_t1b_t1b(other_ops_5_I_t1b_t1b),
    .O(other_ops_5_O)
  );
  Module_10 other_ops_6 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I_t1b_t0b(other_ops_6_I_t1b_t0b),
    .I_t1b_t1b(other_ops_6_I_t1b_t1b),
    .O(other_ops_6_O)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[MapS.scala 23:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[MapS.scala 23:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[MapS.scala 23:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[MapS.scala 23:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T_5 & other_ops_6_valid_down; // @[MapS.scala 23:14]
  assign O_0 = fst_op_O; // @[MapS.scala 17:8]
  assign O_1 = other_ops_0_O; // @[MapS.scala 21:12]
  assign O_2 = other_ops_1_O; // @[MapS.scala 21:12]
  assign O_3 = other_ops_2_O; // @[MapS.scala 21:12]
  assign O_4 = other_ops_3_O; // @[MapS.scala 21:12]
  assign O_5 = other_ops_4_O; // @[MapS.scala 21:12]
  assign O_6 = other_ops_5_O; // @[MapS.scala 21:12]
  assign O_7 = other_ops_6_O; // @[MapS.scala 21:12]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_t1b_t0b = I_0_t1b_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_t1b_t1b = I_0_t1b_t1b; // @[MapS.scala 16:12]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_t1b_t0b = I_1_t1b_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_t1b_t1b = I_1_t1b_t1b; // @[MapS.scala 20:41]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_t1b_t0b = I_2_t1b_t0b; // @[MapS.scala 20:41]
  assign other_ops_1_I_t1b_t1b = I_2_t1b_t1b; // @[MapS.scala 20:41]
  assign other_ops_2_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_2_I_t1b_t0b = I_3_t1b_t0b; // @[MapS.scala 20:41]
  assign other_ops_2_I_t1b_t1b = I_3_t1b_t1b; // @[MapS.scala 20:41]
  assign other_ops_3_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_3_I_t1b_t0b = I_4_t1b_t0b; // @[MapS.scala 20:41]
  assign other_ops_3_I_t1b_t1b = I_4_t1b_t1b; // @[MapS.scala 20:41]
  assign other_ops_4_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_4_I_t1b_t0b = I_5_t1b_t0b; // @[MapS.scala 20:41]
  assign other_ops_4_I_t1b_t1b = I_5_t1b_t1b; // @[MapS.scala 20:41]
  assign other_ops_5_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_5_I_t1b_t0b = I_6_t1b_t0b; // @[MapS.scala 20:41]
  assign other_ops_5_I_t1b_t1b = I_6_t1b_t1b; // @[MapS.scala 20:41]
  assign other_ops_6_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_6_I_t1b_t0b = I_7_t1b_t0b; // @[MapS.scala 20:41]
  assign other_ops_6_I_t1b_t1b = I_7_t1b_t1b; // @[MapS.scala 20:41]
endmodule
module MapT_23(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_t1b_t0b,
  input  [31:0] I_0_t1b_t1b,
  input  [31:0] I_1_t1b_t0b,
  input  [31:0] I_1_t1b_t1b,
  input  [31:0] I_2_t1b_t0b,
  input  [31:0] I_2_t1b_t1b,
  input  [31:0] I_3_t1b_t0b,
  input  [31:0] I_3_t1b_t1b,
  input  [31:0] I_4_t1b_t0b,
  input  [31:0] I_4_t1b_t1b,
  input  [31:0] I_5_t1b_t0b,
  input  [31:0] I_5_t1b_t1b,
  input  [31:0] I_6_t1b_t0b,
  input  [31:0] I_6_t1b_t1b,
  input  [31:0] I_7_t1b_t0b,
  input  [31:0] I_7_t1b_t1b,
  output [31:0] O_0,
  output [31:0] O_1,
  output [31:0] O_2,
  output [31:0] O_3,
  output [31:0] O_4,
  output [31:0] O_5,
  output [31:0] O_6,
  output [31:0] O_7
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_t1b_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_t1b_t1b; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_t1b_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_t1b_t1b; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_t1b_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_t1b_t1b; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_t1b_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_t1b_t1b; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_t1b_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_t1b_t1b; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_t1b_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_t1b_t1b; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_t1b_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_t1b_t1b; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_t1b_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_t1b_t1b; // @[MapT.scala 8:20]
  wire [31:0] op_O_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_3; // @[MapT.scala 8:20]
  wire [31:0] op_O_4; // @[MapT.scala 8:20]
  wire [31:0] op_O_5; // @[MapT.scala 8:20]
  wire [31:0] op_O_6; // @[MapT.scala 8:20]
  wire [31:0] op_O_7; // @[MapT.scala 8:20]
  MapS_60 op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_t1b_t0b(op_I_0_t1b_t0b),
    .I_0_t1b_t1b(op_I_0_t1b_t1b),
    .I_1_t1b_t0b(op_I_1_t1b_t0b),
    .I_1_t1b_t1b(op_I_1_t1b_t1b),
    .I_2_t1b_t0b(op_I_2_t1b_t0b),
    .I_2_t1b_t1b(op_I_2_t1b_t1b),
    .I_3_t1b_t0b(op_I_3_t1b_t0b),
    .I_3_t1b_t1b(op_I_3_t1b_t1b),
    .I_4_t1b_t0b(op_I_4_t1b_t0b),
    .I_4_t1b_t1b(op_I_4_t1b_t1b),
    .I_5_t1b_t0b(op_I_5_t1b_t0b),
    .I_5_t1b_t1b(op_I_5_t1b_t1b),
    .I_6_t1b_t0b(op_I_6_t1b_t0b),
    .I_6_t1b_t1b(op_I_6_t1b_t1b),
    .I_7_t1b_t0b(op_I_7_t1b_t0b),
    .I_7_t1b_t1b(op_I_7_t1b_t1b),
    .O_0(op_O_0),
    .O_1(op_O_1),
    .O_2(op_O_2),
    .O_3(op_O_3),
    .O_4(op_O_4),
    .O_5(op_O_5),
    .O_6(op_O_6),
    .O_7(op_O_7)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0 = op_O_0; // @[MapT.scala 15:7]
  assign O_1 = op_O_1; // @[MapT.scala 15:7]
  assign O_2 = op_O_2; // @[MapT.scala 15:7]
  assign O_3 = op_O_3; // @[MapT.scala 15:7]
  assign O_4 = op_O_4; // @[MapT.scala 15:7]
  assign O_5 = op_O_5; // @[MapT.scala 15:7]
  assign O_6 = op_O_6; // @[MapT.scala 15:7]
  assign O_7 = op_O_7; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_t1b_t0b = I_0_t1b_t0b; // @[MapT.scala 14:10]
  assign op_I_0_t1b_t1b = I_0_t1b_t1b; // @[MapT.scala 14:10]
  assign op_I_1_t1b_t0b = I_1_t1b_t0b; // @[MapT.scala 14:10]
  assign op_I_1_t1b_t1b = I_1_t1b_t1b; // @[MapT.scala 14:10]
  assign op_I_2_t1b_t0b = I_2_t1b_t0b; // @[MapT.scala 14:10]
  assign op_I_2_t1b_t1b = I_2_t1b_t1b; // @[MapT.scala 14:10]
  assign op_I_3_t1b_t0b = I_3_t1b_t0b; // @[MapT.scala 14:10]
  assign op_I_3_t1b_t1b = I_3_t1b_t1b; // @[MapT.scala 14:10]
  assign op_I_4_t1b_t0b = I_4_t1b_t0b; // @[MapT.scala 14:10]
  assign op_I_4_t1b_t1b = I_4_t1b_t1b; // @[MapT.scala 14:10]
  assign op_I_5_t1b_t0b = I_5_t1b_t0b; // @[MapT.scala 14:10]
  assign op_I_5_t1b_t1b = I_5_t1b_t1b; // @[MapT.scala 14:10]
  assign op_I_6_t1b_t0b = I_6_t1b_t0b; // @[MapT.scala 14:10]
  assign op_I_6_t1b_t1b = I_6_t1b_t1b; // @[MapT.scala 14:10]
  assign op_I_7_t1b_t0b = I_7_t1b_t0b; // @[MapT.scala 14:10]
  assign op_I_7_t1b_t1b = I_7_t1b_t1b; // @[MapT.scala 14:10]
endmodule
module ReduceS_4(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0,
  input  [31:0] I_1,
  input  [31:0] I_2,
  output [31:0] O_0
);
  wire [31:0] AddNoValid_I_t0b; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_I_t1b; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_O; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_1_I_t0b; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_1_I_t1b; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_1_O; // @[ReduceS.scala 20:43]
  reg [31:0] _T; // @[ReduceS.scala 27:24]
  reg [31:0] _RAND_0;
  reg [31:0] _T_1; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_1;
  reg [31:0] _T_2; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_2;
  reg [31:0] _T_3; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_3;
  reg  _T_4; // @[ReduceS.scala 47:32]
  reg [31:0] _RAND_4;
  reg  _T_5; // @[ReduceS.scala 47:24]
  reg [31:0] _RAND_5;
  AddNoValid AddNoValid ( // @[ReduceS.scala 20:43]
    .I_t0b(AddNoValid_I_t0b),
    .I_t1b(AddNoValid_I_t1b),
    .O(AddNoValid_O)
  );
  AddNoValid AddNoValid_1 ( // @[ReduceS.scala 20:43]
    .I_t0b(AddNoValid_1_I_t0b),
    .I_t1b(AddNoValid_1_I_t1b),
    .O(AddNoValid_1_O)
  );
  assign valid_down = _T_5; // @[ReduceS.scala 47:14]
  assign O_0 = _T; // @[ReduceS.scala 27:14]
  assign AddNoValid_I_t0b = _T_3; // @[ReduceS.scala 43:18]
  assign AddNoValid_I_t1b = AddNoValid_1_O; // @[ReduceS.scala 36:18]
  assign AddNoValid_1_I_t0b = _T_2; // @[ReduceS.scala 43:18]
  assign AddNoValid_1_I_t1b = _T_1; // @[ReduceS.scala 43:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_2 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_3 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T <= AddNoValid_O;
    _T_1 <= I_0;
    _T_2 <= I_1;
    _T_3 <= I_2;
    if (reset) begin
      _T_4 <= 1'h0;
    end else begin
      _T_4 <= valid_up;
    end
    _T_5 <= _T_4;
  end
endmodule
module MapS_67(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0,
  input  [31:0] I_0_1,
  input  [31:0] I_0_2,
  input  [31:0] I_1_0,
  input  [31:0] I_1_1,
  input  [31:0] I_1_2,
  input  [31:0] I_2_0,
  input  [31:0] I_2_1,
  input  [31:0] I_2_2,
  output [31:0] O_0_0,
  output [31:0] O_1_0,
  output [31:0] O_2_0
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_1; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_2; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_0; // @[MapS.scala 9:22]
  wire  other_ops_0_clock; // @[MapS.scala 10:86]
  wire  other_ops_0_reset; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_O_0; // @[MapS.scala 10:86]
  wire  other_ops_1_clock; // @[MapS.scala 10:86]
  wire  other_ops_1_reset; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_O_0; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  ReduceS_4 fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0(fst_op_I_0),
    .I_1(fst_op_I_1),
    .I_2(fst_op_I_2),
    .O_0(fst_op_O_0)
  );
  ReduceS_4 other_ops_0 ( // @[MapS.scala 10:86]
    .clock(other_ops_0_clock),
    .reset(other_ops_0_reset),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0(other_ops_0_I_0),
    .I_1(other_ops_0_I_1),
    .I_2(other_ops_0_I_2),
    .O_0(other_ops_0_O_0)
  );
  ReduceS_4 other_ops_1 ( // @[MapS.scala 10:86]
    .clock(other_ops_1_clock),
    .reset(other_ops_1_reset),
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0(other_ops_1_I_0),
    .I_1(other_ops_1_I_1),
    .I_2(other_ops_1_I_2),
    .O_0(other_ops_1_O_0)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign O_1_0 = other_ops_0_O_0; // @[MapS.scala 21:12]
  assign O_2_0 = other_ops_1_O_0; // @[MapS.scala 21:12]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0 = I_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_1 = I_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_2 = I_0_2; // @[MapS.scala 16:12]
  assign other_ops_0_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_0_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0 = I_1_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_1 = I_1_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_2 = I_1_2; // @[MapS.scala 20:41]
  assign other_ops_1_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_1_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0 = I_2_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_1 = I_2_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_2 = I_2_2; // @[MapS.scala 20:41]
endmodule
module ReduceS_5(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0,
  input  [31:0] I_1_0,
  input  [31:0] I_2_0,
  output [31:0] O_0_0
);
  wire [31:0] MapSNoValid_I_0_t0b; // @[ReduceS.scala 20:43]
  wire [31:0] MapSNoValid_I_0_t1b; // @[ReduceS.scala 20:43]
  wire [31:0] MapSNoValid_O_0; // @[ReduceS.scala 20:43]
  wire [31:0] MapSNoValid_1_I_0_t0b; // @[ReduceS.scala 20:43]
  wire [31:0] MapSNoValid_1_I_0_t1b; // @[ReduceS.scala 20:43]
  wire [31:0] MapSNoValid_1_O_0; // @[ReduceS.scala 20:43]
  reg [31:0] _T_0; // @[ReduceS.scala 27:24]
  reg [31:0] _RAND_0;
  reg [31:0] _T_1_0; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_1;
  reg [31:0] _T_2_0; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_2;
  reg [31:0] _T_3_0; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_3;
  reg  _T_4; // @[ReduceS.scala 47:32]
  reg [31:0] _RAND_4;
  reg  _T_5; // @[ReduceS.scala 47:24]
  reg [31:0] _RAND_5;
  MapSNoValid MapSNoValid ( // @[ReduceS.scala 20:43]
    .I_0_t0b(MapSNoValid_I_0_t0b),
    .I_0_t1b(MapSNoValid_I_0_t1b),
    .O_0(MapSNoValid_O_0)
  );
  MapSNoValid MapSNoValid_1 ( // @[ReduceS.scala 20:43]
    .I_0_t0b(MapSNoValid_1_I_0_t0b),
    .I_0_t1b(MapSNoValid_1_I_0_t1b),
    .O_0(MapSNoValid_1_O_0)
  );
  assign valid_down = _T_5; // @[ReduceS.scala 47:14]
  assign O_0_0 = _T_0; // @[ReduceS.scala 27:14]
  assign MapSNoValid_I_0_t0b = _T_1_0; // @[ReduceS.scala 43:18]
  assign MapSNoValid_I_0_t1b = MapSNoValid_1_O_0; // @[ReduceS.scala 36:18]
  assign MapSNoValid_1_I_0_t0b = _T_3_0; // @[ReduceS.scala 43:18]
  assign MapSNoValid_1_I_0_t1b = _T_2_0; // @[ReduceS.scala 43:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1_0 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_2_0 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_3_0 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_0 <= MapSNoValid_O_0;
    _T_1_0 <= I_0_0;
    _T_2_0 <= I_1_0;
    _T_3_0 <= I_2_0;
    if (reset) begin
      _T_4 <= 1'h0;
    end else begin
      _T_4 <= valid_up;
    end
    _T_5 <= _T_4;
  end
endmodule
module Module_11(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0,
  input  [31:0] I_0_1,
  input  [31:0] I_0_2,
  input  [31:0] I_1_0,
  input  [31:0] I_1_1,
  input  [31:0] I_1_2,
  input  [31:0] I_2_0,
  input  [31:0] I_2_1,
  input  [31:0] I_2_2,
  output [31:0] O_0_0
);
  wire  InitialDelayCounter_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_valid_down; // @[Const.scala 11:33]
  wire  n746_valid_up; // @[Top.scala 475:22]
  wire  n746_valid_down; // @[Top.scala 475:22]
  wire [31:0] n746_I0_0_0; // @[Top.scala 475:22]
  wire [31:0] n746_I0_0_1; // @[Top.scala 475:22]
  wire [31:0] n746_I0_0_2; // @[Top.scala 475:22]
  wire [31:0] n746_I0_1_0; // @[Top.scala 475:22]
  wire [31:0] n746_I0_1_1; // @[Top.scala 475:22]
  wire [31:0] n746_I0_1_2; // @[Top.scala 475:22]
  wire [31:0] n746_I0_2_0; // @[Top.scala 475:22]
  wire [31:0] n746_I0_2_1; // @[Top.scala 475:22]
  wire [31:0] n746_I0_2_2; // @[Top.scala 475:22]
  wire [31:0] n746_O_0_0_t0b; // @[Top.scala 475:22]
  wire [31:0] n746_O_0_0_t1b; // @[Top.scala 475:22]
  wire [31:0] n746_O_0_1_t0b; // @[Top.scala 475:22]
  wire [31:0] n746_O_0_1_t1b; // @[Top.scala 475:22]
  wire [31:0] n746_O_0_2_t0b; // @[Top.scala 475:22]
  wire [31:0] n746_O_0_2_t1b; // @[Top.scala 475:22]
  wire [31:0] n746_O_1_0_t0b; // @[Top.scala 475:22]
  wire [31:0] n746_O_1_0_t1b; // @[Top.scala 475:22]
  wire [31:0] n746_O_1_1_t0b; // @[Top.scala 475:22]
  wire [31:0] n746_O_1_1_t1b; // @[Top.scala 475:22]
  wire [31:0] n746_O_1_2_t0b; // @[Top.scala 475:22]
  wire [31:0] n746_O_1_2_t1b; // @[Top.scala 475:22]
  wire [31:0] n746_O_2_0_t0b; // @[Top.scala 475:22]
  wire [31:0] n746_O_2_0_t1b; // @[Top.scala 475:22]
  wire [31:0] n746_O_2_1_t0b; // @[Top.scala 475:22]
  wire [31:0] n746_O_2_1_t1b; // @[Top.scala 475:22]
  wire [31:0] n746_O_2_2_t0b; // @[Top.scala 475:22]
  wire [31:0] n746_O_2_2_t1b; // @[Top.scala 475:22]
  wire  n757_clock; // @[Top.scala 479:22]
  wire  n757_reset; // @[Top.scala 479:22]
  wire  n757_valid_up; // @[Top.scala 479:22]
  wire  n757_valid_down; // @[Top.scala 479:22]
  wire [31:0] n757_I_0_0_t0b; // @[Top.scala 479:22]
  wire [31:0] n757_I_0_0_t1b; // @[Top.scala 479:22]
  wire [31:0] n757_I_0_1_t0b; // @[Top.scala 479:22]
  wire [31:0] n757_I_0_1_t1b; // @[Top.scala 479:22]
  wire [31:0] n757_I_0_2_t0b; // @[Top.scala 479:22]
  wire [31:0] n757_I_0_2_t1b; // @[Top.scala 479:22]
  wire [31:0] n757_I_1_0_t0b; // @[Top.scala 479:22]
  wire [31:0] n757_I_1_0_t1b; // @[Top.scala 479:22]
  wire [31:0] n757_I_1_1_t0b; // @[Top.scala 479:22]
  wire [31:0] n757_I_1_1_t1b; // @[Top.scala 479:22]
  wire [31:0] n757_I_1_2_t0b; // @[Top.scala 479:22]
  wire [31:0] n757_I_1_2_t1b; // @[Top.scala 479:22]
  wire [31:0] n757_I_2_0_t0b; // @[Top.scala 479:22]
  wire [31:0] n757_I_2_0_t1b; // @[Top.scala 479:22]
  wire [31:0] n757_I_2_1_t0b; // @[Top.scala 479:22]
  wire [31:0] n757_I_2_1_t1b; // @[Top.scala 479:22]
  wire [31:0] n757_I_2_2_t0b; // @[Top.scala 479:22]
  wire [31:0] n757_I_2_2_t1b; // @[Top.scala 479:22]
  wire [31:0] n757_O_0_0; // @[Top.scala 479:22]
  wire [31:0] n757_O_0_1; // @[Top.scala 479:22]
  wire [31:0] n757_O_0_2; // @[Top.scala 479:22]
  wire [31:0] n757_O_1_0; // @[Top.scala 479:22]
  wire [31:0] n757_O_1_1; // @[Top.scala 479:22]
  wire [31:0] n757_O_1_2; // @[Top.scala 479:22]
  wire [31:0] n757_O_2_0; // @[Top.scala 479:22]
  wire [31:0] n757_O_2_1; // @[Top.scala 479:22]
  wire [31:0] n757_O_2_2; // @[Top.scala 479:22]
  wire  n762_clock; // @[Top.scala 482:22]
  wire  n762_reset; // @[Top.scala 482:22]
  wire  n762_valid_up; // @[Top.scala 482:22]
  wire  n762_valid_down; // @[Top.scala 482:22]
  wire [31:0] n762_I_0_0; // @[Top.scala 482:22]
  wire [31:0] n762_I_0_1; // @[Top.scala 482:22]
  wire [31:0] n762_I_0_2; // @[Top.scala 482:22]
  wire [31:0] n762_I_1_0; // @[Top.scala 482:22]
  wire [31:0] n762_I_1_1; // @[Top.scala 482:22]
  wire [31:0] n762_I_1_2; // @[Top.scala 482:22]
  wire [31:0] n762_I_2_0; // @[Top.scala 482:22]
  wire [31:0] n762_I_2_1; // @[Top.scala 482:22]
  wire [31:0] n762_I_2_2; // @[Top.scala 482:22]
  wire [31:0] n762_O_0_0; // @[Top.scala 482:22]
  wire [31:0] n762_O_1_0; // @[Top.scala 482:22]
  wire [31:0] n762_O_2_0; // @[Top.scala 482:22]
  wire  n767_clock; // @[Top.scala 485:22]
  wire  n767_reset; // @[Top.scala 485:22]
  wire  n767_valid_up; // @[Top.scala 485:22]
  wire  n767_valid_down; // @[Top.scala 485:22]
  wire [31:0] n767_I_0_0; // @[Top.scala 485:22]
  wire [31:0] n767_I_1_0; // @[Top.scala 485:22]
  wire [31:0] n767_I_2_0; // @[Top.scala 485:22]
  wire [31:0] n767_O_0_0; // @[Top.scala 485:22]
  wire  InitialDelayCounter_1_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_1_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_1_valid_down; // @[Const.scala 11:33]
  wire  n770_valid_up; // @[Top.scala 489:22]
  wire  n770_valid_down; // @[Top.scala 489:22]
  wire [31:0] n770_I0_0_0; // @[Top.scala 489:22]
  wire [31:0] n770_O_0_0_t0b; // @[Top.scala 489:22]
  wire [7:0] n770_O_0_0_t1b; // @[Top.scala 489:22]
  wire  n781_clock; // @[Top.scala 493:22]
  wire  n781_reset; // @[Top.scala 493:22]
  wire  n781_valid_up; // @[Top.scala 493:22]
  wire  n781_valid_down; // @[Top.scala 493:22]
  wire [31:0] n781_I_0_0_t0b; // @[Top.scala 493:22]
  wire [7:0] n781_I_0_0_t1b; // @[Top.scala 493:22]
  wire [31:0] n781_O_0_0; // @[Top.scala 493:22]
  InitialDelayCounter_2 InitialDelayCounter ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_clock),
    .reset(InitialDelayCounter_reset),
    .valid_down(InitialDelayCounter_valid_down)
  );
  Map2S_63 n746 ( // @[Top.scala 475:22]
    .valid_up(n746_valid_up),
    .valid_down(n746_valid_down),
    .I0_0_0(n746_I0_0_0),
    .I0_0_1(n746_I0_0_1),
    .I0_0_2(n746_I0_0_2),
    .I0_1_0(n746_I0_1_0),
    .I0_1_1(n746_I0_1_1),
    .I0_1_2(n746_I0_1_2),
    .I0_2_0(n746_I0_2_0),
    .I0_2_1(n746_I0_2_1),
    .I0_2_2(n746_I0_2_2),
    .O_0_0_t0b(n746_O_0_0_t0b),
    .O_0_0_t1b(n746_O_0_0_t1b),
    .O_0_1_t0b(n746_O_0_1_t0b),
    .O_0_1_t1b(n746_O_0_1_t1b),
    .O_0_2_t0b(n746_O_0_2_t0b),
    .O_0_2_t1b(n746_O_0_2_t1b),
    .O_1_0_t0b(n746_O_1_0_t0b),
    .O_1_0_t1b(n746_O_1_0_t1b),
    .O_1_1_t0b(n746_O_1_1_t0b),
    .O_1_1_t1b(n746_O_1_1_t1b),
    .O_1_2_t0b(n746_O_1_2_t0b),
    .O_1_2_t1b(n746_O_1_2_t1b),
    .O_2_0_t0b(n746_O_2_0_t0b),
    .O_2_0_t1b(n746_O_2_0_t1b),
    .O_2_1_t0b(n746_O_2_1_t0b),
    .O_2_1_t1b(n746_O_2_1_t1b),
    .O_2_2_t0b(n746_O_2_2_t0b),
    .O_2_2_t1b(n746_O_2_2_t1b)
  );
  MapS_55 n757 ( // @[Top.scala 479:22]
    .clock(n757_clock),
    .reset(n757_reset),
    .valid_up(n757_valid_up),
    .valid_down(n757_valid_down),
    .I_0_0_t0b(n757_I_0_0_t0b),
    .I_0_0_t1b(n757_I_0_0_t1b),
    .I_0_1_t0b(n757_I_0_1_t0b),
    .I_0_1_t1b(n757_I_0_1_t1b),
    .I_0_2_t0b(n757_I_0_2_t0b),
    .I_0_2_t1b(n757_I_0_2_t1b),
    .I_1_0_t0b(n757_I_1_0_t0b),
    .I_1_0_t1b(n757_I_1_0_t1b),
    .I_1_1_t0b(n757_I_1_1_t0b),
    .I_1_1_t1b(n757_I_1_1_t1b),
    .I_1_2_t0b(n757_I_1_2_t0b),
    .I_1_2_t1b(n757_I_1_2_t1b),
    .I_2_0_t0b(n757_I_2_0_t0b),
    .I_2_0_t1b(n757_I_2_0_t1b),
    .I_2_1_t0b(n757_I_2_1_t0b),
    .I_2_1_t1b(n757_I_2_1_t1b),
    .I_2_2_t0b(n757_I_2_2_t0b),
    .I_2_2_t1b(n757_I_2_2_t1b),
    .O_0_0(n757_O_0_0),
    .O_0_1(n757_O_0_1),
    .O_0_2(n757_O_0_2),
    .O_1_0(n757_O_1_0),
    .O_1_1(n757_O_1_1),
    .O_1_2(n757_O_1_2),
    .O_2_0(n757_O_2_0),
    .O_2_1(n757_O_2_1),
    .O_2_2(n757_O_2_2)
  );
  MapS_67 n762 ( // @[Top.scala 482:22]
    .clock(n762_clock),
    .reset(n762_reset),
    .valid_up(n762_valid_up),
    .valid_down(n762_valid_down),
    .I_0_0(n762_I_0_0),
    .I_0_1(n762_I_0_1),
    .I_0_2(n762_I_0_2),
    .I_1_0(n762_I_1_0),
    .I_1_1(n762_I_1_1),
    .I_1_2(n762_I_1_2),
    .I_2_0(n762_I_2_0),
    .I_2_1(n762_I_2_1),
    .I_2_2(n762_I_2_2),
    .O_0_0(n762_O_0_0),
    .O_1_0(n762_O_1_0),
    .O_2_0(n762_O_2_0)
  );
  ReduceS_5 n767 ( // @[Top.scala 485:22]
    .clock(n767_clock),
    .reset(n767_reset),
    .valid_up(n767_valid_up),
    .valid_down(n767_valid_down),
    .I_0_0(n767_I_0_0),
    .I_1_0(n767_I_1_0),
    .I_2_0(n767_I_2_0),
    .O_0_0(n767_O_0_0)
  );
  InitialDelayCounter_5 InitialDelayCounter_1 ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_1_clock),
    .reset(InitialDelayCounter_1_reset),
    .valid_down(InitialDelayCounter_1_valid_down)
  );
  Map2S_65 n770 ( // @[Top.scala 489:22]
    .valid_up(n770_valid_up),
    .valid_down(n770_valid_down),
    .I0_0_0(n770_I0_0_0),
    .O_0_0_t0b(n770_O_0_0_t0b),
    .O_0_0_t1b(n770_O_0_0_t1b)
  );
  MapS_58 n781 ( // @[Top.scala 493:22]
    .clock(n781_clock),
    .reset(n781_reset),
    .valid_up(n781_valid_up),
    .valid_down(n781_valid_down),
    .I_0_0_t0b(n781_I_0_0_t0b),
    .I_0_0_t1b(n781_I_0_0_t1b),
    .O_0_0(n781_O_0_0)
  );
  assign valid_down = n781_valid_down; // @[Top.scala 497:16]
  assign O_0_0 = n781_O_0_0; // @[Top.scala 496:7]
  assign InitialDelayCounter_clock = clock;
  assign InitialDelayCounter_reset = reset;
  assign n746_valid_up = valid_up & InitialDelayCounter_valid_down; // @[Top.scala 478:19]
  assign n746_I0_0_0 = I_0_0; // @[Top.scala 476:13]
  assign n746_I0_0_1 = I_0_1; // @[Top.scala 476:13]
  assign n746_I0_0_2 = I_0_2; // @[Top.scala 476:13]
  assign n746_I0_1_0 = I_1_0; // @[Top.scala 476:13]
  assign n746_I0_1_1 = I_1_1; // @[Top.scala 476:13]
  assign n746_I0_1_2 = I_1_2; // @[Top.scala 476:13]
  assign n746_I0_2_0 = I_2_0; // @[Top.scala 476:13]
  assign n746_I0_2_1 = I_2_1; // @[Top.scala 476:13]
  assign n746_I0_2_2 = I_2_2; // @[Top.scala 476:13]
  assign n757_clock = clock;
  assign n757_reset = reset;
  assign n757_valid_up = n746_valid_down; // @[Top.scala 481:19]
  assign n757_I_0_0_t0b = n746_O_0_0_t0b; // @[Top.scala 480:12]
  assign n757_I_0_0_t1b = n746_O_0_0_t1b; // @[Top.scala 480:12]
  assign n757_I_0_1_t0b = n746_O_0_1_t0b; // @[Top.scala 480:12]
  assign n757_I_0_1_t1b = n746_O_0_1_t1b; // @[Top.scala 480:12]
  assign n757_I_0_2_t0b = n746_O_0_2_t0b; // @[Top.scala 480:12]
  assign n757_I_0_2_t1b = n746_O_0_2_t1b; // @[Top.scala 480:12]
  assign n757_I_1_0_t0b = n746_O_1_0_t0b; // @[Top.scala 480:12]
  assign n757_I_1_0_t1b = n746_O_1_0_t1b; // @[Top.scala 480:12]
  assign n757_I_1_1_t0b = n746_O_1_1_t0b; // @[Top.scala 480:12]
  assign n757_I_1_1_t1b = n746_O_1_1_t1b; // @[Top.scala 480:12]
  assign n757_I_1_2_t0b = n746_O_1_2_t0b; // @[Top.scala 480:12]
  assign n757_I_1_2_t1b = n746_O_1_2_t1b; // @[Top.scala 480:12]
  assign n757_I_2_0_t0b = n746_O_2_0_t0b; // @[Top.scala 480:12]
  assign n757_I_2_0_t1b = n746_O_2_0_t1b; // @[Top.scala 480:12]
  assign n757_I_2_1_t0b = n746_O_2_1_t0b; // @[Top.scala 480:12]
  assign n757_I_2_1_t1b = n746_O_2_1_t1b; // @[Top.scala 480:12]
  assign n757_I_2_2_t0b = n746_O_2_2_t0b; // @[Top.scala 480:12]
  assign n757_I_2_2_t1b = n746_O_2_2_t1b; // @[Top.scala 480:12]
  assign n762_clock = clock;
  assign n762_reset = reset;
  assign n762_valid_up = n757_valid_down; // @[Top.scala 484:19]
  assign n762_I_0_0 = n757_O_0_0; // @[Top.scala 483:12]
  assign n762_I_0_1 = n757_O_0_1; // @[Top.scala 483:12]
  assign n762_I_0_2 = n757_O_0_2; // @[Top.scala 483:12]
  assign n762_I_1_0 = n757_O_1_0; // @[Top.scala 483:12]
  assign n762_I_1_1 = n757_O_1_1; // @[Top.scala 483:12]
  assign n762_I_1_2 = n757_O_1_2; // @[Top.scala 483:12]
  assign n762_I_2_0 = n757_O_2_0; // @[Top.scala 483:12]
  assign n762_I_2_1 = n757_O_2_1; // @[Top.scala 483:12]
  assign n762_I_2_2 = n757_O_2_2; // @[Top.scala 483:12]
  assign n767_clock = clock;
  assign n767_reset = reset;
  assign n767_valid_up = n762_valid_down; // @[Top.scala 487:19]
  assign n767_I_0_0 = n762_O_0_0; // @[Top.scala 486:12]
  assign n767_I_1_0 = n762_O_1_0; // @[Top.scala 486:12]
  assign n767_I_2_0 = n762_O_2_0; // @[Top.scala 486:12]
  assign InitialDelayCounter_1_clock = clock;
  assign InitialDelayCounter_1_reset = reset;
  assign n770_valid_up = n767_valid_down & InitialDelayCounter_1_valid_down; // @[Top.scala 492:19]
  assign n770_I0_0_0 = n767_O_0_0; // @[Top.scala 490:13]
  assign n781_clock = clock;
  assign n781_reset = reset;
  assign n781_valid_up = n770_valid_down; // @[Top.scala 495:19]
  assign n781_I_0_0_t0b = n770_O_0_0_t0b; // @[Top.scala 494:12]
  assign n781_I_0_0_t1b = n770_O_0_0_t1b; // @[Top.scala 494:12]
endmodule
module MapS_70(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0_0,
  input  [31:0] I_0_0_1,
  input  [31:0] I_0_0_2,
  input  [31:0] I_0_1_0,
  input  [31:0] I_0_1_1,
  input  [31:0] I_0_1_2,
  input  [31:0] I_0_2_0,
  input  [31:0] I_0_2_1,
  input  [31:0] I_0_2_2,
  input  [31:0] I_1_0_0,
  input  [31:0] I_1_0_1,
  input  [31:0] I_1_0_2,
  input  [31:0] I_1_1_0,
  input  [31:0] I_1_1_1,
  input  [31:0] I_1_1_2,
  input  [31:0] I_1_2_0,
  input  [31:0] I_1_2_1,
  input  [31:0] I_1_2_2,
  input  [31:0] I_2_0_0,
  input  [31:0] I_2_0_1,
  input  [31:0] I_2_0_2,
  input  [31:0] I_2_1_0,
  input  [31:0] I_2_1_1,
  input  [31:0] I_2_1_2,
  input  [31:0] I_2_2_0,
  input  [31:0] I_2_2_1,
  input  [31:0] I_2_2_2,
  input  [31:0] I_3_0_0,
  input  [31:0] I_3_0_1,
  input  [31:0] I_3_0_2,
  input  [31:0] I_3_1_0,
  input  [31:0] I_3_1_1,
  input  [31:0] I_3_1_2,
  input  [31:0] I_3_2_0,
  input  [31:0] I_3_2_1,
  input  [31:0] I_3_2_2,
  input  [31:0] I_4_0_0,
  input  [31:0] I_4_0_1,
  input  [31:0] I_4_0_2,
  input  [31:0] I_4_1_0,
  input  [31:0] I_4_1_1,
  input  [31:0] I_4_1_2,
  input  [31:0] I_4_2_0,
  input  [31:0] I_4_2_1,
  input  [31:0] I_4_2_2,
  input  [31:0] I_5_0_0,
  input  [31:0] I_5_0_1,
  input  [31:0] I_5_0_2,
  input  [31:0] I_5_1_0,
  input  [31:0] I_5_1_1,
  input  [31:0] I_5_1_2,
  input  [31:0] I_5_2_0,
  input  [31:0] I_5_2_1,
  input  [31:0] I_5_2_2,
  input  [31:0] I_6_0_0,
  input  [31:0] I_6_0_1,
  input  [31:0] I_6_0_2,
  input  [31:0] I_6_1_0,
  input  [31:0] I_6_1_1,
  input  [31:0] I_6_1_2,
  input  [31:0] I_6_2_0,
  input  [31:0] I_6_2_1,
  input  [31:0] I_6_2_2,
  input  [31:0] I_7_0_0,
  input  [31:0] I_7_0_1,
  input  [31:0] I_7_0_2,
  input  [31:0] I_7_1_0,
  input  [31:0] I_7_1_1,
  input  [31:0] I_7_1_2,
  input  [31:0] I_7_2_0,
  input  [31:0] I_7_2_1,
  input  [31:0] I_7_2_2,
  output [31:0] O_0_0_0,
  output [31:0] O_1_0_0,
  output [31:0] O_2_0_0,
  output [31:0] O_3_0_0,
  output [31:0] O_4_0_0,
  output [31:0] O_5_0_0,
  output [31:0] O_6_0_0,
  output [31:0] O_7_0_0
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_0; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_1; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_2; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_1_0; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_1_1; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_1_2; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_2_0; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_2_1; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_2_2; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_0_0; // @[MapS.scala 9:22]
  wire  other_ops_0_clock; // @[MapS.scala 10:86]
  wire  other_ops_0_reset; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_2_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_1_clock; // @[MapS.scala 10:86]
  wire  other_ops_1_reset; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_2_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_2_clock; // @[MapS.scala 10:86]
  wire  other_ops_2_reset; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_2_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_3_clock; // @[MapS.scala 10:86]
  wire  other_ops_3_reset; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_2_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_4_clock; // @[MapS.scala 10:86]
  wire  other_ops_4_reset; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_2_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_5_clock; // @[MapS.scala 10:86]
  wire  other_ops_5_reset; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_2_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_6_clock; // @[MapS.scala 10:86]
  wire  other_ops_6_reset; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_2_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_O_0_0; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  wire  _T_1; // @[MapS.scala 23:83]
  wire  _T_2; // @[MapS.scala 23:83]
  wire  _T_3; // @[MapS.scala 23:83]
  wire  _T_4; // @[MapS.scala 23:83]
  wire  _T_5; // @[MapS.scala 23:83]
  Module_11 fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_0(fst_op_I_0_0),
    .I_0_1(fst_op_I_0_1),
    .I_0_2(fst_op_I_0_2),
    .I_1_0(fst_op_I_1_0),
    .I_1_1(fst_op_I_1_1),
    .I_1_2(fst_op_I_1_2),
    .I_2_0(fst_op_I_2_0),
    .I_2_1(fst_op_I_2_1),
    .I_2_2(fst_op_I_2_2),
    .O_0_0(fst_op_O_0_0)
  );
  Module_11 other_ops_0 ( // @[MapS.scala 10:86]
    .clock(other_ops_0_clock),
    .reset(other_ops_0_reset),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_0(other_ops_0_I_0_0),
    .I_0_1(other_ops_0_I_0_1),
    .I_0_2(other_ops_0_I_0_2),
    .I_1_0(other_ops_0_I_1_0),
    .I_1_1(other_ops_0_I_1_1),
    .I_1_2(other_ops_0_I_1_2),
    .I_2_0(other_ops_0_I_2_0),
    .I_2_1(other_ops_0_I_2_1),
    .I_2_2(other_ops_0_I_2_2),
    .O_0_0(other_ops_0_O_0_0)
  );
  Module_11 other_ops_1 ( // @[MapS.scala 10:86]
    .clock(other_ops_1_clock),
    .reset(other_ops_1_reset),
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0_0(other_ops_1_I_0_0),
    .I_0_1(other_ops_1_I_0_1),
    .I_0_2(other_ops_1_I_0_2),
    .I_1_0(other_ops_1_I_1_0),
    .I_1_1(other_ops_1_I_1_1),
    .I_1_2(other_ops_1_I_1_2),
    .I_2_0(other_ops_1_I_2_0),
    .I_2_1(other_ops_1_I_2_1),
    .I_2_2(other_ops_1_I_2_2),
    .O_0_0(other_ops_1_O_0_0)
  );
  Module_11 other_ops_2 ( // @[MapS.scala 10:86]
    .clock(other_ops_2_clock),
    .reset(other_ops_2_reset),
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I_0_0(other_ops_2_I_0_0),
    .I_0_1(other_ops_2_I_0_1),
    .I_0_2(other_ops_2_I_0_2),
    .I_1_0(other_ops_2_I_1_0),
    .I_1_1(other_ops_2_I_1_1),
    .I_1_2(other_ops_2_I_1_2),
    .I_2_0(other_ops_2_I_2_0),
    .I_2_1(other_ops_2_I_2_1),
    .I_2_2(other_ops_2_I_2_2),
    .O_0_0(other_ops_2_O_0_0)
  );
  Module_11 other_ops_3 ( // @[MapS.scala 10:86]
    .clock(other_ops_3_clock),
    .reset(other_ops_3_reset),
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I_0_0(other_ops_3_I_0_0),
    .I_0_1(other_ops_3_I_0_1),
    .I_0_2(other_ops_3_I_0_2),
    .I_1_0(other_ops_3_I_1_0),
    .I_1_1(other_ops_3_I_1_1),
    .I_1_2(other_ops_3_I_1_2),
    .I_2_0(other_ops_3_I_2_0),
    .I_2_1(other_ops_3_I_2_1),
    .I_2_2(other_ops_3_I_2_2),
    .O_0_0(other_ops_3_O_0_0)
  );
  Module_11 other_ops_4 ( // @[MapS.scala 10:86]
    .clock(other_ops_4_clock),
    .reset(other_ops_4_reset),
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I_0_0(other_ops_4_I_0_0),
    .I_0_1(other_ops_4_I_0_1),
    .I_0_2(other_ops_4_I_0_2),
    .I_1_0(other_ops_4_I_1_0),
    .I_1_1(other_ops_4_I_1_1),
    .I_1_2(other_ops_4_I_1_2),
    .I_2_0(other_ops_4_I_2_0),
    .I_2_1(other_ops_4_I_2_1),
    .I_2_2(other_ops_4_I_2_2),
    .O_0_0(other_ops_4_O_0_0)
  );
  Module_11 other_ops_5 ( // @[MapS.scala 10:86]
    .clock(other_ops_5_clock),
    .reset(other_ops_5_reset),
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I_0_0(other_ops_5_I_0_0),
    .I_0_1(other_ops_5_I_0_1),
    .I_0_2(other_ops_5_I_0_2),
    .I_1_0(other_ops_5_I_1_0),
    .I_1_1(other_ops_5_I_1_1),
    .I_1_2(other_ops_5_I_1_2),
    .I_2_0(other_ops_5_I_2_0),
    .I_2_1(other_ops_5_I_2_1),
    .I_2_2(other_ops_5_I_2_2),
    .O_0_0(other_ops_5_O_0_0)
  );
  Module_11 other_ops_6 ( // @[MapS.scala 10:86]
    .clock(other_ops_6_clock),
    .reset(other_ops_6_reset),
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I_0_0(other_ops_6_I_0_0),
    .I_0_1(other_ops_6_I_0_1),
    .I_0_2(other_ops_6_I_0_2),
    .I_1_0(other_ops_6_I_1_0),
    .I_1_1(other_ops_6_I_1_1),
    .I_1_2(other_ops_6_I_1_2),
    .I_2_0(other_ops_6_I_2_0),
    .I_2_1(other_ops_6_I_2_1),
    .I_2_2(other_ops_6_I_2_2),
    .O_0_0(other_ops_6_O_0_0)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[MapS.scala 23:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[MapS.scala 23:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[MapS.scala 23:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[MapS.scala 23:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T_5 & other_ops_6_valid_down; // @[MapS.scala 23:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[MapS.scala 17:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[MapS.scala 21:12]
  assign O_2_0_0 = other_ops_1_O_0_0; // @[MapS.scala 21:12]
  assign O_3_0_0 = other_ops_2_O_0_0; // @[MapS.scala 21:12]
  assign O_4_0_0 = other_ops_3_O_0_0; // @[MapS.scala 21:12]
  assign O_5_0_0 = other_ops_4_O_0_0; // @[MapS.scala 21:12]
  assign O_6_0_0 = other_ops_5_O_0_0; // @[MapS.scala 21:12]
  assign O_7_0_0 = other_ops_6_O_0_0; // @[MapS.scala 21:12]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_0 = I_0_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_1 = I_0_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_2 = I_0_0_2; // @[MapS.scala 16:12]
  assign fst_op_I_1_0 = I_0_1_0; // @[MapS.scala 16:12]
  assign fst_op_I_1_1 = I_0_1_1; // @[MapS.scala 16:12]
  assign fst_op_I_1_2 = I_0_1_2; // @[MapS.scala 16:12]
  assign fst_op_I_2_0 = I_0_2_0; // @[MapS.scala 16:12]
  assign fst_op_I_2_1 = I_0_2_1; // @[MapS.scala 16:12]
  assign fst_op_I_2_2 = I_0_2_2; // @[MapS.scala 16:12]
  assign other_ops_0_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_0_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_0 = I_1_0_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1 = I_1_0_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2 = I_1_0_2; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_0 = I_1_1_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_1 = I_1_1_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_2 = I_1_1_2; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_0 = I_1_2_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_1 = I_1_2_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_2 = I_1_2_2; // @[MapS.scala 20:41]
  assign other_ops_1_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_1_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0_0 = I_2_0_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1 = I_2_0_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2 = I_2_0_2; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_0 = I_2_1_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_1 = I_2_1_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_2 = I_2_1_2; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_0 = I_2_2_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_1 = I_2_2_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_2 = I_2_2_2; // @[MapS.scala 20:41]
  assign other_ops_2_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_2_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_2_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_2_I_0_0 = I_3_0_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1 = I_3_0_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2 = I_3_0_2; // @[MapS.scala 20:41]
  assign other_ops_2_I_1_0 = I_3_1_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_1_1 = I_3_1_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_1_2 = I_3_1_2; // @[MapS.scala 20:41]
  assign other_ops_2_I_2_0 = I_3_2_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_2_1 = I_3_2_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_2_2 = I_3_2_2; // @[MapS.scala 20:41]
  assign other_ops_3_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_3_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_3_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_3_I_0_0 = I_4_0_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_1 = I_4_0_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_2 = I_4_0_2; // @[MapS.scala 20:41]
  assign other_ops_3_I_1_0 = I_4_1_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_1_1 = I_4_1_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_1_2 = I_4_1_2; // @[MapS.scala 20:41]
  assign other_ops_3_I_2_0 = I_4_2_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_2_1 = I_4_2_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_2_2 = I_4_2_2; // @[MapS.scala 20:41]
  assign other_ops_4_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_4_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_4_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_4_I_0_0 = I_5_0_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_1 = I_5_0_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_2 = I_5_0_2; // @[MapS.scala 20:41]
  assign other_ops_4_I_1_0 = I_5_1_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_1_1 = I_5_1_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_1_2 = I_5_1_2; // @[MapS.scala 20:41]
  assign other_ops_4_I_2_0 = I_5_2_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_2_1 = I_5_2_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_2_2 = I_5_2_2; // @[MapS.scala 20:41]
  assign other_ops_5_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_5_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_5_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_5_I_0_0 = I_6_0_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_1 = I_6_0_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_2 = I_6_0_2; // @[MapS.scala 20:41]
  assign other_ops_5_I_1_0 = I_6_1_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_1_1 = I_6_1_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_1_2 = I_6_1_2; // @[MapS.scala 20:41]
  assign other_ops_5_I_2_0 = I_6_2_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_2_1 = I_6_2_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_2_2 = I_6_2_2; // @[MapS.scala 20:41]
  assign other_ops_6_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_6_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_6_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_6_I_0_0 = I_7_0_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_1 = I_7_0_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_2 = I_7_0_2; // @[MapS.scala 20:41]
  assign other_ops_6_I_1_0 = I_7_1_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_1_1 = I_7_1_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_1_2 = I_7_1_2; // @[MapS.scala 20:41]
  assign other_ops_6_I_2_0 = I_7_2_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_2_1 = I_7_2_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_2_2 = I_7_2_2; // @[MapS.scala 20:41]
endmodule
module MapT_32(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0_0,
  input  [31:0] I_0_0_1,
  input  [31:0] I_0_0_2,
  input  [31:0] I_0_1_0,
  input  [31:0] I_0_1_1,
  input  [31:0] I_0_1_2,
  input  [31:0] I_0_2_0,
  input  [31:0] I_0_2_1,
  input  [31:0] I_0_2_2,
  input  [31:0] I_1_0_0,
  input  [31:0] I_1_0_1,
  input  [31:0] I_1_0_2,
  input  [31:0] I_1_1_0,
  input  [31:0] I_1_1_1,
  input  [31:0] I_1_1_2,
  input  [31:0] I_1_2_0,
  input  [31:0] I_1_2_1,
  input  [31:0] I_1_2_2,
  input  [31:0] I_2_0_0,
  input  [31:0] I_2_0_1,
  input  [31:0] I_2_0_2,
  input  [31:0] I_2_1_0,
  input  [31:0] I_2_1_1,
  input  [31:0] I_2_1_2,
  input  [31:0] I_2_2_0,
  input  [31:0] I_2_2_1,
  input  [31:0] I_2_2_2,
  input  [31:0] I_3_0_0,
  input  [31:0] I_3_0_1,
  input  [31:0] I_3_0_2,
  input  [31:0] I_3_1_0,
  input  [31:0] I_3_1_1,
  input  [31:0] I_3_1_2,
  input  [31:0] I_3_2_0,
  input  [31:0] I_3_2_1,
  input  [31:0] I_3_2_2,
  input  [31:0] I_4_0_0,
  input  [31:0] I_4_0_1,
  input  [31:0] I_4_0_2,
  input  [31:0] I_4_1_0,
  input  [31:0] I_4_1_1,
  input  [31:0] I_4_1_2,
  input  [31:0] I_4_2_0,
  input  [31:0] I_4_2_1,
  input  [31:0] I_4_2_2,
  input  [31:0] I_5_0_0,
  input  [31:0] I_5_0_1,
  input  [31:0] I_5_0_2,
  input  [31:0] I_5_1_0,
  input  [31:0] I_5_1_1,
  input  [31:0] I_5_1_2,
  input  [31:0] I_5_2_0,
  input  [31:0] I_5_2_1,
  input  [31:0] I_5_2_2,
  input  [31:0] I_6_0_0,
  input  [31:0] I_6_0_1,
  input  [31:0] I_6_0_2,
  input  [31:0] I_6_1_0,
  input  [31:0] I_6_1_1,
  input  [31:0] I_6_1_2,
  input  [31:0] I_6_2_0,
  input  [31:0] I_6_2_1,
  input  [31:0] I_6_2_2,
  input  [31:0] I_7_0_0,
  input  [31:0] I_7_0_1,
  input  [31:0] I_7_0_2,
  input  [31:0] I_7_1_0,
  input  [31:0] I_7_1_1,
  input  [31:0] I_7_1_2,
  input  [31:0] I_7_2_0,
  input  [31:0] I_7_2_1,
  input  [31:0] I_7_2_2,
  output [31:0] O_0_0_0,
  output [31:0] O_1_0_0,
  output [31:0] O_2_0_0,
  output [31:0] O_3_0_0,
  output [31:0] O_4_0_0,
  output [31:0] O_5_0_0,
  output [31:0] O_6_0_0,
  output [31:0] O_7_0_0
);
  wire  op_clock; // @[MapT.scala 8:20]
  wire  op_reset; // @[MapT.scala 8:20]
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_0_0; // @[MapT.scala 8:20]
  MapS_70 op ( // @[MapT.scala 8:20]
    .clock(op_clock),
    .reset(op_reset),
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0(op_I_0_0_0),
    .I_0_0_1(op_I_0_0_1),
    .I_0_0_2(op_I_0_0_2),
    .I_0_1_0(op_I_0_1_0),
    .I_0_1_1(op_I_0_1_1),
    .I_0_1_2(op_I_0_1_2),
    .I_0_2_0(op_I_0_2_0),
    .I_0_2_1(op_I_0_2_1),
    .I_0_2_2(op_I_0_2_2),
    .I_1_0_0(op_I_1_0_0),
    .I_1_0_1(op_I_1_0_1),
    .I_1_0_2(op_I_1_0_2),
    .I_1_1_0(op_I_1_1_0),
    .I_1_1_1(op_I_1_1_1),
    .I_1_1_2(op_I_1_1_2),
    .I_1_2_0(op_I_1_2_0),
    .I_1_2_1(op_I_1_2_1),
    .I_1_2_2(op_I_1_2_2),
    .I_2_0_0(op_I_2_0_0),
    .I_2_0_1(op_I_2_0_1),
    .I_2_0_2(op_I_2_0_2),
    .I_2_1_0(op_I_2_1_0),
    .I_2_1_1(op_I_2_1_1),
    .I_2_1_2(op_I_2_1_2),
    .I_2_2_0(op_I_2_2_0),
    .I_2_2_1(op_I_2_2_1),
    .I_2_2_2(op_I_2_2_2),
    .I_3_0_0(op_I_3_0_0),
    .I_3_0_1(op_I_3_0_1),
    .I_3_0_2(op_I_3_0_2),
    .I_3_1_0(op_I_3_1_0),
    .I_3_1_1(op_I_3_1_1),
    .I_3_1_2(op_I_3_1_2),
    .I_3_2_0(op_I_3_2_0),
    .I_3_2_1(op_I_3_2_1),
    .I_3_2_2(op_I_3_2_2),
    .I_4_0_0(op_I_4_0_0),
    .I_4_0_1(op_I_4_0_1),
    .I_4_0_2(op_I_4_0_2),
    .I_4_1_0(op_I_4_1_0),
    .I_4_1_1(op_I_4_1_1),
    .I_4_1_2(op_I_4_1_2),
    .I_4_2_0(op_I_4_2_0),
    .I_4_2_1(op_I_4_2_1),
    .I_4_2_2(op_I_4_2_2),
    .I_5_0_0(op_I_5_0_0),
    .I_5_0_1(op_I_5_0_1),
    .I_5_0_2(op_I_5_0_2),
    .I_5_1_0(op_I_5_1_0),
    .I_5_1_1(op_I_5_1_1),
    .I_5_1_2(op_I_5_1_2),
    .I_5_2_0(op_I_5_2_0),
    .I_5_2_1(op_I_5_2_1),
    .I_5_2_2(op_I_5_2_2),
    .I_6_0_0(op_I_6_0_0),
    .I_6_0_1(op_I_6_0_1),
    .I_6_0_2(op_I_6_0_2),
    .I_6_1_0(op_I_6_1_0),
    .I_6_1_1(op_I_6_1_1),
    .I_6_1_2(op_I_6_1_2),
    .I_6_2_0(op_I_6_2_0),
    .I_6_2_1(op_I_6_2_1),
    .I_6_2_2(op_I_6_2_2),
    .I_7_0_0(op_I_7_0_0),
    .I_7_0_1(op_I_7_0_1),
    .I_7_0_2(op_I_7_0_2),
    .I_7_1_0(op_I_7_1_0),
    .I_7_1_1(op_I_7_1_1),
    .I_7_1_2(op_I_7_1_2),
    .I_7_2_0(op_I_7_2_0),
    .I_7_2_1(op_I_7_2_1),
    .I_7_2_2(op_I_7_2_2),
    .O_0_0_0(op_O_0_0_0),
    .O_1_0_0(op_O_1_0_0),
    .O_2_0_0(op_O_2_0_0),
    .O_3_0_0(op_O_3_0_0),
    .O_4_0_0(op_O_4_0_0),
    .O_5_0_0(op_O_5_0_0),
    .O_6_0_0(op_O_6_0_0),
    .O_7_0_0(op_O_7_0_0)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0 = op_O_0_0_0; // @[MapT.scala 15:7]
  assign O_1_0_0 = op_O_1_0_0; // @[MapT.scala 15:7]
  assign O_2_0_0 = op_O_2_0_0; // @[MapT.scala 15:7]
  assign O_3_0_0 = op_O_3_0_0; // @[MapT.scala 15:7]
  assign O_4_0_0 = op_O_4_0_0; // @[MapT.scala 15:7]
  assign O_5_0_0 = op_O_5_0_0; // @[MapT.scala 15:7]
  assign O_6_0_0 = op_O_6_0_0; // @[MapT.scala 15:7]
  assign O_7_0_0 = op_O_7_0_0; // @[MapT.scala 15:7]
  assign op_clock = clock;
  assign op_reset = reset;
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0 = I_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_1 = I_0_0_1; // @[MapT.scala 14:10]
  assign op_I_0_0_2 = I_0_0_2; // @[MapT.scala 14:10]
  assign op_I_0_1_0 = I_0_1_0; // @[MapT.scala 14:10]
  assign op_I_0_1_1 = I_0_1_1; // @[MapT.scala 14:10]
  assign op_I_0_1_2 = I_0_1_2; // @[MapT.scala 14:10]
  assign op_I_0_2_0 = I_0_2_0; // @[MapT.scala 14:10]
  assign op_I_0_2_1 = I_0_2_1; // @[MapT.scala 14:10]
  assign op_I_0_2_2 = I_0_2_2; // @[MapT.scala 14:10]
  assign op_I_1_0_0 = I_1_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_1 = I_1_0_1; // @[MapT.scala 14:10]
  assign op_I_1_0_2 = I_1_0_2; // @[MapT.scala 14:10]
  assign op_I_1_1_0 = I_1_1_0; // @[MapT.scala 14:10]
  assign op_I_1_1_1 = I_1_1_1; // @[MapT.scala 14:10]
  assign op_I_1_1_2 = I_1_1_2; // @[MapT.scala 14:10]
  assign op_I_1_2_0 = I_1_2_0; // @[MapT.scala 14:10]
  assign op_I_1_2_1 = I_1_2_1; // @[MapT.scala 14:10]
  assign op_I_1_2_2 = I_1_2_2; // @[MapT.scala 14:10]
  assign op_I_2_0_0 = I_2_0_0; // @[MapT.scala 14:10]
  assign op_I_2_0_1 = I_2_0_1; // @[MapT.scala 14:10]
  assign op_I_2_0_2 = I_2_0_2; // @[MapT.scala 14:10]
  assign op_I_2_1_0 = I_2_1_0; // @[MapT.scala 14:10]
  assign op_I_2_1_1 = I_2_1_1; // @[MapT.scala 14:10]
  assign op_I_2_1_2 = I_2_1_2; // @[MapT.scala 14:10]
  assign op_I_2_2_0 = I_2_2_0; // @[MapT.scala 14:10]
  assign op_I_2_2_1 = I_2_2_1; // @[MapT.scala 14:10]
  assign op_I_2_2_2 = I_2_2_2; // @[MapT.scala 14:10]
  assign op_I_3_0_0 = I_3_0_0; // @[MapT.scala 14:10]
  assign op_I_3_0_1 = I_3_0_1; // @[MapT.scala 14:10]
  assign op_I_3_0_2 = I_3_0_2; // @[MapT.scala 14:10]
  assign op_I_3_1_0 = I_3_1_0; // @[MapT.scala 14:10]
  assign op_I_3_1_1 = I_3_1_1; // @[MapT.scala 14:10]
  assign op_I_3_1_2 = I_3_1_2; // @[MapT.scala 14:10]
  assign op_I_3_2_0 = I_3_2_0; // @[MapT.scala 14:10]
  assign op_I_3_2_1 = I_3_2_1; // @[MapT.scala 14:10]
  assign op_I_3_2_2 = I_3_2_2; // @[MapT.scala 14:10]
  assign op_I_4_0_0 = I_4_0_0; // @[MapT.scala 14:10]
  assign op_I_4_0_1 = I_4_0_1; // @[MapT.scala 14:10]
  assign op_I_4_0_2 = I_4_0_2; // @[MapT.scala 14:10]
  assign op_I_4_1_0 = I_4_1_0; // @[MapT.scala 14:10]
  assign op_I_4_1_1 = I_4_1_1; // @[MapT.scala 14:10]
  assign op_I_4_1_2 = I_4_1_2; // @[MapT.scala 14:10]
  assign op_I_4_2_0 = I_4_2_0; // @[MapT.scala 14:10]
  assign op_I_4_2_1 = I_4_2_1; // @[MapT.scala 14:10]
  assign op_I_4_2_2 = I_4_2_2; // @[MapT.scala 14:10]
  assign op_I_5_0_0 = I_5_0_0; // @[MapT.scala 14:10]
  assign op_I_5_0_1 = I_5_0_1; // @[MapT.scala 14:10]
  assign op_I_5_0_2 = I_5_0_2; // @[MapT.scala 14:10]
  assign op_I_5_1_0 = I_5_1_0; // @[MapT.scala 14:10]
  assign op_I_5_1_1 = I_5_1_1; // @[MapT.scala 14:10]
  assign op_I_5_1_2 = I_5_1_2; // @[MapT.scala 14:10]
  assign op_I_5_2_0 = I_5_2_0; // @[MapT.scala 14:10]
  assign op_I_5_2_1 = I_5_2_1; // @[MapT.scala 14:10]
  assign op_I_5_2_2 = I_5_2_2; // @[MapT.scala 14:10]
  assign op_I_6_0_0 = I_6_0_0; // @[MapT.scala 14:10]
  assign op_I_6_0_1 = I_6_0_1; // @[MapT.scala 14:10]
  assign op_I_6_0_2 = I_6_0_2; // @[MapT.scala 14:10]
  assign op_I_6_1_0 = I_6_1_0; // @[MapT.scala 14:10]
  assign op_I_6_1_1 = I_6_1_1; // @[MapT.scala 14:10]
  assign op_I_6_1_2 = I_6_1_2; // @[MapT.scala 14:10]
  assign op_I_6_2_0 = I_6_2_0; // @[MapT.scala 14:10]
  assign op_I_6_2_1 = I_6_2_1; // @[MapT.scala 14:10]
  assign op_I_6_2_2 = I_6_2_2; // @[MapT.scala 14:10]
  assign op_I_7_0_0 = I_7_0_0; // @[MapT.scala 14:10]
  assign op_I_7_0_1 = I_7_0_1; // @[MapT.scala 14:10]
  assign op_I_7_0_2 = I_7_0_2; // @[MapT.scala 14:10]
  assign op_I_7_1_0 = I_7_1_0; // @[MapT.scala 14:10]
  assign op_I_7_1_1 = I_7_1_1; // @[MapT.scala 14:10]
  assign op_I_7_1_2 = I_7_1_2; // @[MapT.scala 14:10]
  assign op_I_7_2_0 = I_7_2_0; // @[MapT.scala 14:10]
  assign op_I_7_2_1 = I_7_2_1; // @[MapT.scala 14:10]
  assign op_I_7_2_2 = I_7_2_2; // @[MapT.scala 14:10]
endmodule
module Snd_3(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_t1b,
  output [31:0] O
);
  assign valid_down = valid_up; // @[Tuple.scala 67:14]
  assign O = I_t1b; // @[Tuple.scala 66:5]
endmodule
module Module_13(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_t1b_t0b,
  input  [31:0] I_t1b_t1b,
  output [31:0] O
);
  wire  n820_valid_up; // @[Top.scala 578:22]
  wire  n820_valid_down; // @[Top.scala 578:22]
  wire [31:0] n820_I_t1b_t0b; // @[Top.scala 578:22]
  wire [31:0] n820_I_t1b_t1b; // @[Top.scala 578:22]
  wire [31:0] n820_O_t0b; // @[Top.scala 578:22]
  wire [31:0] n820_O_t1b; // @[Top.scala 578:22]
  wire  n821_valid_up; // @[Top.scala 581:22]
  wire  n821_valid_down; // @[Top.scala 581:22]
  wire [31:0] n821_I_t1b; // @[Top.scala 581:22]
  wire [31:0] n821_O; // @[Top.scala 581:22]
  Snd_1 n820 ( // @[Top.scala 578:22]
    .valid_up(n820_valid_up),
    .valid_down(n820_valid_down),
    .I_t1b_t0b(n820_I_t1b_t0b),
    .I_t1b_t1b(n820_I_t1b_t1b),
    .O_t0b(n820_O_t0b),
    .O_t1b(n820_O_t1b)
  );
  Snd_3 n821 ( // @[Top.scala 581:22]
    .valid_up(n821_valid_up),
    .valid_down(n821_valid_down),
    .I_t1b(n821_I_t1b),
    .O(n821_O)
  );
  assign valid_down = n821_valid_down; // @[Top.scala 585:16]
  assign O = n821_O; // @[Top.scala 584:7]
  assign n820_valid_up = valid_up; // @[Top.scala 580:19]
  assign n820_I_t1b_t0b = I_t1b_t0b; // @[Top.scala 579:12]
  assign n820_I_t1b_t1b = I_t1b_t1b; // @[Top.scala 579:12]
  assign n821_valid_up = n820_valid_down; // @[Top.scala 583:19]
  assign n821_I_t1b = n820_O_t1b; // @[Top.scala 582:12]
endmodule
module MapS_71(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_t1b_t0b,
  input  [31:0] I_0_t1b_t1b,
  input  [31:0] I_1_t1b_t0b,
  input  [31:0] I_1_t1b_t1b,
  input  [31:0] I_2_t1b_t0b,
  input  [31:0] I_2_t1b_t1b,
  input  [31:0] I_3_t1b_t0b,
  input  [31:0] I_3_t1b_t1b,
  input  [31:0] I_4_t1b_t0b,
  input  [31:0] I_4_t1b_t1b,
  input  [31:0] I_5_t1b_t0b,
  input  [31:0] I_5_t1b_t1b,
  input  [31:0] I_6_t1b_t0b,
  input  [31:0] I_6_t1b_t1b,
  input  [31:0] I_7_t1b_t0b,
  input  [31:0] I_7_t1b_t1b,
  output [31:0] O_0,
  output [31:0] O_1,
  output [31:0] O_2,
  output [31:0] O_3,
  output [31:0] O_4,
  output [31:0] O_5,
  output [31:0] O_6,
  output [31:0] O_7
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_t1b_t0b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_t1b_t1b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_t1b_t0b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_t1b_t1b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_O; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_t1b_t0b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_t1b_t1b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_O; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_t1b_t0b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_t1b_t1b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_O; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_t1b_t0b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_t1b_t1b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_O; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_t1b_t0b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_t1b_t1b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_O; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_t1b_t0b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_t1b_t1b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_O; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_t1b_t0b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_t1b_t1b; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_O; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  wire  _T_1; // @[MapS.scala 23:83]
  wire  _T_2; // @[MapS.scala 23:83]
  wire  _T_3; // @[MapS.scala 23:83]
  wire  _T_4; // @[MapS.scala 23:83]
  wire  _T_5; // @[MapS.scala 23:83]
  Module_13 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_t1b_t0b(fst_op_I_t1b_t0b),
    .I_t1b_t1b(fst_op_I_t1b_t1b),
    .O(fst_op_O)
  );
  Module_13 other_ops_0 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_t1b_t0b(other_ops_0_I_t1b_t0b),
    .I_t1b_t1b(other_ops_0_I_t1b_t1b),
    .O(other_ops_0_O)
  );
  Module_13 other_ops_1 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_t1b_t0b(other_ops_1_I_t1b_t0b),
    .I_t1b_t1b(other_ops_1_I_t1b_t1b),
    .O(other_ops_1_O)
  );
  Module_13 other_ops_2 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I_t1b_t0b(other_ops_2_I_t1b_t0b),
    .I_t1b_t1b(other_ops_2_I_t1b_t1b),
    .O(other_ops_2_O)
  );
  Module_13 other_ops_3 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I_t1b_t0b(other_ops_3_I_t1b_t0b),
    .I_t1b_t1b(other_ops_3_I_t1b_t1b),
    .O(other_ops_3_O)
  );
  Module_13 other_ops_4 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I_t1b_t0b(other_ops_4_I_t1b_t0b),
    .I_t1b_t1b(other_ops_4_I_t1b_t1b),
    .O(other_ops_4_O)
  );
  Module_13 other_ops_5 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I_t1b_t0b(other_ops_5_I_t1b_t0b),
    .I_t1b_t1b(other_ops_5_I_t1b_t1b),
    .O(other_ops_5_O)
  );
  Module_13 other_ops_6 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I_t1b_t0b(other_ops_6_I_t1b_t0b),
    .I_t1b_t1b(other_ops_6_I_t1b_t1b),
    .O(other_ops_6_O)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[MapS.scala 23:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[MapS.scala 23:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[MapS.scala 23:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[MapS.scala 23:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T_5 & other_ops_6_valid_down; // @[MapS.scala 23:14]
  assign O_0 = fst_op_O; // @[MapS.scala 17:8]
  assign O_1 = other_ops_0_O; // @[MapS.scala 21:12]
  assign O_2 = other_ops_1_O; // @[MapS.scala 21:12]
  assign O_3 = other_ops_2_O; // @[MapS.scala 21:12]
  assign O_4 = other_ops_3_O; // @[MapS.scala 21:12]
  assign O_5 = other_ops_4_O; // @[MapS.scala 21:12]
  assign O_6 = other_ops_5_O; // @[MapS.scala 21:12]
  assign O_7 = other_ops_6_O; // @[MapS.scala 21:12]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_t1b_t0b = I_0_t1b_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_t1b_t1b = I_0_t1b_t1b; // @[MapS.scala 16:12]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_t1b_t0b = I_1_t1b_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_t1b_t1b = I_1_t1b_t1b; // @[MapS.scala 20:41]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_t1b_t0b = I_2_t1b_t0b; // @[MapS.scala 20:41]
  assign other_ops_1_I_t1b_t1b = I_2_t1b_t1b; // @[MapS.scala 20:41]
  assign other_ops_2_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_2_I_t1b_t0b = I_3_t1b_t0b; // @[MapS.scala 20:41]
  assign other_ops_2_I_t1b_t1b = I_3_t1b_t1b; // @[MapS.scala 20:41]
  assign other_ops_3_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_3_I_t1b_t0b = I_4_t1b_t0b; // @[MapS.scala 20:41]
  assign other_ops_3_I_t1b_t1b = I_4_t1b_t1b; // @[MapS.scala 20:41]
  assign other_ops_4_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_4_I_t1b_t0b = I_5_t1b_t0b; // @[MapS.scala 20:41]
  assign other_ops_4_I_t1b_t1b = I_5_t1b_t1b; // @[MapS.scala 20:41]
  assign other_ops_5_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_5_I_t1b_t0b = I_6_t1b_t0b; // @[MapS.scala 20:41]
  assign other_ops_5_I_t1b_t1b = I_6_t1b_t1b; // @[MapS.scala 20:41]
  assign other_ops_6_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_6_I_t1b_t0b = I_7_t1b_t0b; // @[MapS.scala 20:41]
  assign other_ops_6_I_t1b_t1b = I_7_t1b_t1b; // @[MapS.scala 20:41]
endmodule
module MapT_33(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_t1b_t0b,
  input  [31:0] I_0_t1b_t1b,
  input  [31:0] I_1_t1b_t0b,
  input  [31:0] I_1_t1b_t1b,
  input  [31:0] I_2_t1b_t0b,
  input  [31:0] I_2_t1b_t1b,
  input  [31:0] I_3_t1b_t0b,
  input  [31:0] I_3_t1b_t1b,
  input  [31:0] I_4_t1b_t0b,
  input  [31:0] I_4_t1b_t1b,
  input  [31:0] I_5_t1b_t0b,
  input  [31:0] I_5_t1b_t1b,
  input  [31:0] I_6_t1b_t0b,
  input  [31:0] I_6_t1b_t1b,
  input  [31:0] I_7_t1b_t0b,
  input  [31:0] I_7_t1b_t1b,
  output [31:0] O_0,
  output [31:0] O_1,
  output [31:0] O_2,
  output [31:0] O_3,
  output [31:0] O_4,
  output [31:0] O_5,
  output [31:0] O_6,
  output [31:0] O_7
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_t1b_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_t1b_t1b; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_t1b_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_t1b_t1b; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_t1b_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_t1b_t1b; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_t1b_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_t1b_t1b; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_t1b_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_t1b_t1b; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_t1b_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_t1b_t1b; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_t1b_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_t1b_t1b; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_t1b_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_t1b_t1b; // @[MapT.scala 8:20]
  wire [31:0] op_O_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_3; // @[MapT.scala 8:20]
  wire [31:0] op_O_4; // @[MapT.scala 8:20]
  wire [31:0] op_O_5; // @[MapT.scala 8:20]
  wire [31:0] op_O_6; // @[MapT.scala 8:20]
  wire [31:0] op_O_7; // @[MapT.scala 8:20]
  MapS_71 op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_t1b_t0b(op_I_0_t1b_t0b),
    .I_0_t1b_t1b(op_I_0_t1b_t1b),
    .I_1_t1b_t0b(op_I_1_t1b_t0b),
    .I_1_t1b_t1b(op_I_1_t1b_t1b),
    .I_2_t1b_t0b(op_I_2_t1b_t0b),
    .I_2_t1b_t1b(op_I_2_t1b_t1b),
    .I_3_t1b_t0b(op_I_3_t1b_t0b),
    .I_3_t1b_t1b(op_I_3_t1b_t1b),
    .I_4_t1b_t0b(op_I_4_t1b_t0b),
    .I_4_t1b_t1b(op_I_4_t1b_t1b),
    .I_5_t1b_t0b(op_I_5_t1b_t0b),
    .I_5_t1b_t1b(op_I_5_t1b_t1b),
    .I_6_t1b_t0b(op_I_6_t1b_t0b),
    .I_6_t1b_t1b(op_I_6_t1b_t1b),
    .I_7_t1b_t0b(op_I_7_t1b_t0b),
    .I_7_t1b_t1b(op_I_7_t1b_t1b),
    .O_0(op_O_0),
    .O_1(op_O_1),
    .O_2(op_O_2),
    .O_3(op_O_3),
    .O_4(op_O_4),
    .O_5(op_O_5),
    .O_6(op_O_6),
    .O_7(op_O_7)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0 = op_O_0; // @[MapT.scala 15:7]
  assign O_1 = op_O_1; // @[MapT.scala 15:7]
  assign O_2 = op_O_2; // @[MapT.scala 15:7]
  assign O_3 = op_O_3; // @[MapT.scala 15:7]
  assign O_4 = op_O_4; // @[MapT.scala 15:7]
  assign O_5 = op_O_5; // @[MapT.scala 15:7]
  assign O_6 = op_O_6; // @[MapT.scala 15:7]
  assign O_7 = op_O_7; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_t1b_t0b = I_0_t1b_t0b; // @[MapT.scala 14:10]
  assign op_I_0_t1b_t1b = I_0_t1b_t1b; // @[MapT.scala 14:10]
  assign op_I_1_t1b_t0b = I_1_t1b_t0b; // @[MapT.scala 14:10]
  assign op_I_1_t1b_t1b = I_1_t1b_t1b; // @[MapT.scala 14:10]
  assign op_I_2_t1b_t0b = I_2_t1b_t0b; // @[MapT.scala 14:10]
  assign op_I_2_t1b_t1b = I_2_t1b_t1b; // @[MapT.scala 14:10]
  assign op_I_3_t1b_t0b = I_3_t1b_t0b; // @[MapT.scala 14:10]
  assign op_I_3_t1b_t1b = I_3_t1b_t1b; // @[MapT.scala 14:10]
  assign op_I_4_t1b_t0b = I_4_t1b_t0b; // @[MapT.scala 14:10]
  assign op_I_4_t1b_t1b = I_4_t1b_t1b; // @[MapT.scala 14:10]
  assign op_I_5_t1b_t0b = I_5_t1b_t0b; // @[MapT.scala 14:10]
  assign op_I_5_t1b_t1b = I_5_t1b_t1b; // @[MapT.scala 14:10]
  assign op_I_6_t1b_t0b = I_6_t1b_t0b; // @[MapT.scala 14:10]
  assign op_I_6_t1b_t1b = I_6_t1b_t1b; // @[MapT.scala 14:10]
  assign op_I_7_t1b_t0b = I_7_t1b_t0b; // @[MapT.scala 14:10]
  assign op_I_7_t1b_t1b = I_7_t1b_t1b; // @[MapT.scala 14:10]
endmodule
module ReduceS_6(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0,
  input  [31:0] I_1,
  input  [31:0] I_2,
  output [31:0] O_0
);
  wire [31:0] AddNoValid_I_t0b; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_I_t1b; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_O; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_1_I_t0b; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_1_I_t1b; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_1_O; // @[ReduceS.scala 20:43]
  reg [31:0] _T; // @[ReduceS.scala 27:24]
  reg [31:0] _RAND_0;
  reg [31:0] _T_1; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_1;
  reg [31:0] _T_2; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_2;
  reg [31:0] _T_3; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_3;
  reg  _T_4; // @[ReduceS.scala 47:32]
  reg [31:0] _RAND_4;
  reg  _T_5; // @[ReduceS.scala 47:24]
  reg [31:0] _RAND_5;
  AddNoValid AddNoValid ( // @[ReduceS.scala 20:43]
    .I_t0b(AddNoValid_I_t0b),
    .I_t1b(AddNoValid_I_t1b),
    .O(AddNoValid_O)
  );
  AddNoValid AddNoValid_1 ( // @[ReduceS.scala 20:43]
    .I_t0b(AddNoValid_1_I_t0b),
    .I_t1b(AddNoValid_1_I_t1b),
    .O(AddNoValid_1_O)
  );
  assign valid_down = _T_5; // @[ReduceS.scala 47:14]
  assign O_0 = _T; // @[ReduceS.scala 27:14]
  assign AddNoValid_I_t0b = _T_2; // @[ReduceS.scala 43:18]
  assign AddNoValid_I_t1b = AddNoValid_1_O; // @[ReduceS.scala 36:18]
  assign AddNoValid_1_I_t0b = _T_1; // @[ReduceS.scala 43:18]
  assign AddNoValid_1_I_t1b = _T_3; // @[ReduceS.scala 43:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_2 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_3 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T <= AddNoValid_O;
    _T_1 <= I_0;
    _T_2 <= I_1;
    _T_3 <= I_2;
    if (reset) begin
      _T_4 <= 1'h0;
    end else begin
      _T_4 <= valid_up;
    end
    _T_5 <= _T_4;
  end
endmodule
module MapS_78(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0,
  input  [31:0] I_0_1,
  input  [31:0] I_0_2,
  input  [31:0] I_1_0,
  input  [31:0] I_1_1,
  input  [31:0] I_1_2,
  input  [31:0] I_2_0,
  input  [31:0] I_2_1,
  input  [31:0] I_2_2,
  output [31:0] O_0_0,
  output [31:0] O_1_0,
  output [31:0] O_2_0
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_1; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_2; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_0; // @[MapS.scala 9:22]
  wire  other_ops_0_clock; // @[MapS.scala 10:86]
  wire  other_ops_0_reset; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_O_0; // @[MapS.scala 10:86]
  wire  other_ops_1_clock; // @[MapS.scala 10:86]
  wire  other_ops_1_reset; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_O_0; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  ReduceS_6 fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0(fst_op_I_0),
    .I_1(fst_op_I_1),
    .I_2(fst_op_I_2),
    .O_0(fst_op_O_0)
  );
  ReduceS_6 other_ops_0 ( // @[MapS.scala 10:86]
    .clock(other_ops_0_clock),
    .reset(other_ops_0_reset),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0(other_ops_0_I_0),
    .I_1(other_ops_0_I_1),
    .I_2(other_ops_0_I_2),
    .O_0(other_ops_0_O_0)
  );
  ReduceS_6 other_ops_1 ( // @[MapS.scala 10:86]
    .clock(other_ops_1_clock),
    .reset(other_ops_1_reset),
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0(other_ops_1_I_0),
    .I_1(other_ops_1_I_1),
    .I_2(other_ops_1_I_2),
    .O_0(other_ops_1_O_0)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign O_1_0 = other_ops_0_O_0; // @[MapS.scala 21:12]
  assign O_2_0 = other_ops_1_O_0; // @[MapS.scala 21:12]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0 = I_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_1 = I_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_2 = I_0_2; // @[MapS.scala 16:12]
  assign other_ops_0_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_0_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0 = I_1_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_1 = I_1_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_2 = I_1_2; // @[MapS.scala 20:41]
  assign other_ops_1_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_1_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0 = I_2_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_1 = I_2_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_2 = I_2_2; // @[MapS.scala 20:41]
endmodule
module ReduceS_7(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0,
  input  [31:0] I_1_0,
  input  [31:0] I_2_0,
  output [31:0] O_0_0
);
  wire [31:0] MapSNoValid_I_0_t0b; // @[ReduceS.scala 20:43]
  wire [31:0] MapSNoValid_I_0_t1b; // @[ReduceS.scala 20:43]
  wire [31:0] MapSNoValid_O_0; // @[ReduceS.scala 20:43]
  wire [31:0] MapSNoValid_1_I_0_t0b; // @[ReduceS.scala 20:43]
  wire [31:0] MapSNoValid_1_I_0_t1b; // @[ReduceS.scala 20:43]
  wire [31:0] MapSNoValid_1_O_0; // @[ReduceS.scala 20:43]
  reg [31:0] _T_0; // @[ReduceS.scala 27:24]
  reg [31:0] _RAND_0;
  reg [31:0] _T_1_0; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_1;
  reg [31:0] _T_2_0; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_2;
  reg [31:0] _T_3_0; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_3;
  reg  _T_4; // @[ReduceS.scala 47:32]
  reg [31:0] _RAND_4;
  reg  _T_5; // @[ReduceS.scala 47:24]
  reg [31:0] _RAND_5;
  MapSNoValid MapSNoValid ( // @[ReduceS.scala 20:43]
    .I_0_t0b(MapSNoValid_I_0_t0b),
    .I_0_t1b(MapSNoValid_I_0_t1b),
    .O_0(MapSNoValid_O_0)
  );
  MapSNoValid MapSNoValid_1 ( // @[ReduceS.scala 20:43]
    .I_0_t0b(MapSNoValid_1_I_0_t0b),
    .I_0_t1b(MapSNoValid_1_I_0_t1b),
    .O_0(MapSNoValid_1_O_0)
  );
  assign valid_down = _T_5; // @[ReduceS.scala 47:14]
  assign O_0_0 = _T_0; // @[ReduceS.scala 27:14]
  assign MapSNoValid_I_0_t0b = _T_3_0; // @[ReduceS.scala 43:18]
  assign MapSNoValid_I_0_t1b = MapSNoValid_1_O_0; // @[ReduceS.scala 36:18]
  assign MapSNoValid_1_I_0_t0b = _T_2_0; // @[ReduceS.scala 43:18]
  assign MapSNoValid_1_I_0_t1b = _T_1_0; // @[ReduceS.scala 43:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1_0 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_2_0 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_3_0 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_0 <= MapSNoValid_O_0;
    _T_1_0 <= I_0_0;
    _T_2_0 <= I_1_0;
    _T_3_0 <= I_2_0;
    if (reset) begin
      _T_4 <= 1'h0;
    end else begin
      _T_4 <= valid_up;
    end
    _T_5 <= _T_4;
  end
endmodule
module Module_14(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0,
  input  [31:0] I_0_1,
  input  [31:0] I_0_2,
  input  [31:0] I_1_0,
  input  [31:0] I_1_1,
  input  [31:0] I_1_2,
  input  [31:0] I_2_0,
  input  [31:0] I_2_1,
  input  [31:0] I_2_2,
  output [31:0] O_0_0
);
  wire  InitialDelayCounter_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_valid_down; // @[Const.scala 11:33]
  wire  n932_valid_up; // @[Top.scala 592:22]
  wire  n932_valid_down; // @[Top.scala 592:22]
  wire [31:0] n932_I0_0_0; // @[Top.scala 592:22]
  wire [31:0] n932_I0_0_1; // @[Top.scala 592:22]
  wire [31:0] n932_I0_0_2; // @[Top.scala 592:22]
  wire [31:0] n932_I0_1_0; // @[Top.scala 592:22]
  wire [31:0] n932_I0_1_1; // @[Top.scala 592:22]
  wire [31:0] n932_I0_1_2; // @[Top.scala 592:22]
  wire [31:0] n932_I0_2_0; // @[Top.scala 592:22]
  wire [31:0] n932_I0_2_1; // @[Top.scala 592:22]
  wire [31:0] n932_I0_2_2; // @[Top.scala 592:22]
  wire [31:0] n932_O_0_0_t0b; // @[Top.scala 592:22]
  wire [31:0] n932_O_0_0_t1b; // @[Top.scala 592:22]
  wire [31:0] n932_O_0_1_t0b; // @[Top.scala 592:22]
  wire [31:0] n932_O_0_1_t1b; // @[Top.scala 592:22]
  wire [31:0] n932_O_0_2_t0b; // @[Top.scala 592:22]
  wire [31:0] n932_O_0_2_t1b; // @[Top.scala 592:22]
  wire [31:0] n932_O_1_0_t0b; // @[Top.scala 592:22]
  wire [31:0] n932_O_1_0_t1b; // @[Top.scala 592:22]
  wire [31:0] n932_O_1_1_t0b; // @[Top.scala 592:22]
  wire [31:0] n932_O_1_1_t1b; // @[Top.scala 592:22]
  wire [31:0] n932_O_1_2_t0b; // @[Top.scala 592:22]
  wire [31:0] n932_O_1_2_t1b; // @[Top.scala 592:22]
  wire [31:0] n932_O_2_0_t0b; // @[Top.scala 592:22]
  wire [31:0] n932_O_2_0_t1b; // @[Top.scala 592:22]
  wire [31:0] n932_O_2_1_t0b; // @[Top.scala 592:22]
  wire [31:0] n932_O_2_1_t1b; // @[Top.scala 592:22]
  wire [31:0] n932_O_2_2_t0b; // @[Top.scala 592:22]
  wire [31:0] n932_O_2_2_t1b; // @[Top.scala 592:22]
  wire  n943_clock; // @[Top.scala 596:22]
  wire  n943_reset; // @[Top.scala 596:22]
  wire  n943_valid_up; // @[Top.scala 596:22]
  wire  n943_valid_down; // @[Top.scala 596:22]
  wire [31:0] n943_I_0_0_t0b; // @[Top.scala 596:22]
  wire [31:0] n943_I_0_0_t1b; // @[Top.scala 596:22]
  wire [31:0] n943_I_0_1_t0b; // @[Top.scala 596:22]
  wire [31:0] n943_I_0_1_t1b; // @[Top.scala 596:22]
  wire [31:0] n943_I_0_2_t0b; // @[Top.scala 596:22]
  wire [31:0] n943_I_0_2_t1b; // @[Top.scala 596:22]
  wire [31:0] n943_I_1_0_t0b; // @[Top.scala 596:22]
  wire [31:0] n943_I_1_0_t1b; // @[Top.scala 596:22]
  wire [31:0] n943_I_1_1_t0b; // @[Top.scala 596:22]
  wire [31:0] n943_I_1_1_t1b; // @[Top.scala 596:22]
  wire [31:0] n943_I_1_2_t0b; // @[Top.scala 596:22]
  wire [31:0] n943_I_1_2_t1b; // @[Top.scala 596:22]
  wire [31:0] n943_I_2_0_t0b; // @[Top.scala 596:22]
  wire [31:0] n943_I_2_0_t1b; // @[Top.scala 596:22]
  wire [31:0] n943_I_2_1_t0b; // @[Top.scala 596:22]
  wire [31:0] n943_I_2_1_t1b; // @[Top.scala 596:22]
  wire [31:0] n943_I_2_2_t0b; // @[Top.scala 596:22]
  wire [31:0] n943_I_2_2_t1b; // @[Top.scala 596:22]
  wire [31:0] n943_O_0_0; // @[Top.scala 596:22]
  wire [31:0] n943_O_0_1; // @[Top.scala 596:22]
  wire [31:0] n943_O_0_2; // @[Top.scala 596:22]
  wire [31:0] n943_O_1_0; // @[Top.scala 596:22]
  wire [31:0] n943_O_1_1; // @[Top.scala 596:22]
  wire [31:0] n943_O_1_2; // @[Top.scala 596:22]
  wire [31:0] n943_O_2_0; // @[Top.scala 596:22]
  wire [31:0] n943_O_2_1; // @[Top.scala 596:22]
  wire [31:0] n943_O_2_2; // @[Top.scala 596:22]
  wire  n948_clock; // @[Top.scala 599:22]
  wire  n948_reset; // @[Top.scala 599:22]
  wire  n948_valid_up; // @[Top.scala 599:22]
  wire  n948_valid_down; // @[Top.scala 599:22]
  wire [31:0] n948_I_0_0; // @[Top.scala 599:22]
  wire [31:0] n948_I_0_1; // @[Top.scala 599:22]
  wire [31:0] n948_I_0_2; // @[Top.scala 599:22]
  wire [31:0] n948_I_1_0; // @[Top.scala 599:22]
  wire [31:0] n948_I_1_1; // @[Top.scala 599:22]
  wire [31:0] n948_I_1_2; // @[Top.scala 599:22]
  wire [31:0] n948_I_2_0; // @[Top.scala 599:22]
  wire [31:0] n948_I_2_1; // @[Top.scala 599:22]
  wire [31:0] n948_I_2_2; // @[Top.scala 599:22]
  wire [31:0] n948_O_0_0; // @[Top.scala 599:22]
  wire [31:0] n948_O_1_0; // @[Top.scala 599:22]
  wire [31:0] n948_O_2_0; // @[Top.scala 599:22]
  wire  n953_clock; // @[Top.scala 602:22]
  wire  n953_reset; // @[Top.scala 602:22]
  wire  n953_valid_up; // @[Top.scala 602:22]
  wire  n953_valid_down; // @[Top.scala 602:22]
  wire [31:0] n953_I_0_0; // @[Top.scala 602:22]
  wire [31:0] n953_I_1_0; // @[Top.scala 602:22]
  wire [31:0] n953_I_2_0; // @[Top.scala 602:22]
  wire [31:0] n953_O_0_0; // @[Top.scala 602:22]
  wire  InitialDelayCounter_1_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_1_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_1_valid_down; // @[Const.scala 11:33]
  wire  n956_valid_up; // @[Top.scala 606:22]
  wire  n956_valid_down; // @[Top.scala 606:22]
  wire [31:0] n956_I0_0_0; // @[Top.scala 606:22]
  wire [31:0] n956_O_0_0_t0b; // @[Top.scala 606:22]
  wire [7:0] n956_O_0_0_t1b; // @[Top.scala 606:22]
  wire  n967_clock; // @[Top.scala 610:22]
  wire  n967_reset; // @[Top.scala 610:22]
  wire  n967_valid_up; // @[Top.scala 610:22]
  wire  n967_valid_down; // @[Top.scala 610:22]
  wire [31:0] n967_I_0_0_t0b; // @[Top.scala 610:22]
  wire [7:0] n967_I_0_0_t1b; // @[Top.scala 610:22]
  wire [31:0] n967_O_0_0; // @[Top.scala 610:22]
  InitialDelayCounter_2 InitialDelayCounter ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_clock),
    .reset(InitialDelayCounter_reset),
    .valid_down(InitialDelayCounter_valid_down)
  );
  Map2S_63 n932 ( // @[Top.scala 592:22]
    .valid_up(n932_valid_up),
    .valid_down(n932_valid_down),
    .I0_0_0(n932_I0_0_0),
    .I0_0_1(n932_I0_0_1),
    .I0_0_2(n932_I0_0_2),
    .I0_1_0(n932_I0_1_0),
    .I0_1_1(n932_I0_1_1),
    .I0_1_2(n932_I0_1_2),
    .I0_2_0(n932_I0_2_0),
    .I0_2_1(n932_I0_2_1),
    .I0_2_2(n932_I0_2_2),
    .O_0_0_t0b(n932_O_0_0_t0b),
    .O_0_0_t1b(n932_O_0_0_t1b),
    .O_0_1_t0b(n932_O_0_1_t0b),
    .O_0_1_t1b(n932_O_0_1_t1b),
    .O_0_2_t0b(n932_O_0_2_t0b),
    .O_0_2_t1b(n932_O_0_2_t1b),
    .O_1_0_t0b(n932_O_1_0_t0b),
    .O_1_0_t1b(n932_O_1_0_t1b),
    .O_1_1_t0b(n932_O_1_1_t0b),
    .O_1_1_t1b(n932_O_1_1_t1b),
    .O_1_2_t0b(n932_O_1_2_t0b),
    .O_1_2_t1b(n932_O_1_2_t1b),
    .O_2_0_t0b(n932_O_2_0_t0b),
    .O_2_0_t1b(n932_O_2_0_t1b),
    .O_2_1_t0b(n932_O_2_1_t0b),
    .O_2_1_t1b(n932_O_2_1_t1b),
    .O_2_2_t0b(n932_O_2_2_t0b),
    .O_2_2_t1b(n932_O_2_2_t1b)
  );
  MapS_55 n943 ( // @[Top.scala 596:22]
    .clock(n943_clock),
    .reset(n943_reset),
    .valid_up(n943_valid_up),
    .valid_down(n943_valid_down),
    .I_0_0_t0b(n943_I_0_0_t0b),
    .I_0_0_t1b(n943_I_0_0_t1b),
    .I_0_1_t0b(n943_I_0_1_t0b),
    .I_0_1_t1b(n943_I_0_1_t1b),
    .I_0_2_t0b(n943_I_0_2_t0b),
    .I_0_2_t1b(n943_I_0_2_t1b),
    .I_1_0_t0b(n943_I_1_0_t0b),
    .I_1_0_t1b(n943_I_1_0_t1b),
    .I_1_1_t0b(n943_I_1_1_t0b),
    .I_1_1_t1b(n943_I_1_1_t1b),
    .I_1_2_t0b(n943_I_1_2_t0b),
    .I_1_2_t1b(n943_I_1_2_t1b),
    .I_2_0_t0b(n943_I_2_0_t0b),
    .I_2_0_t1b(n943_I_2_0_t1b),
    .I_2_1_t0b(n943_I_2_1_t0b),
    .I_2_1_t1b(n943_I_2_1_t1b),
    .I_2_2_t0b(n943_I_2_2_t0b),
    .I_2_2_t1b(n943_I_2_2_t1b),
    .O_0_0(n943_O_0_0),
    .O_0_1(n943_O_0_1),
    .O_0_2(n943_O_0_2),
    .O_1_0(n943_O_1_0),
    .O_1_1(n943_O_1_1),
    .O_1_2(n943_O_1_2),
    .O_2_0(n943_O_2_0),
    .O_2_1(n943_O_2_1),
    .O_2_2(n943_O_2_2)
  );
  MapS_78 n948 ( // @[Top.scala 599:22]
    .clock(n948_clock),
    .reset(n948_reset),
    .valid_up(n948_valid_up),
    .valid_down(n948_valid_down),
    .I_0_0(n948_I_0_0),
    .I_0_1(n948_I_0_1),
    .I_0_2(n948_I_0_2),
    .I_1_0(n948_I_1_0),
    .I_1_1(n948_I_1_1),
    .I_1_2(n948_I_1_2),
    .I_2_0(n948_I_2_0),
    .I_2_1(n948_I_2_1),
    .I_2_2(n948_I_2_2),
    .O_0_0(n948_O_0_0),
    .O_1_0(n948_O_1_0),
    .O_2_0(n948_O_2_0)
  );
  ReduceS_7 n953 ( // @[Top.scala 602:22]
    .clock(n953_clock),
    .reset(n953_reset),
    .valid_up(n953_valid_up),
    .valid_down(n953_valid_down),
    .I_0_0(n953_I_0_0),
    .I_1_0(n953_I_1_0),
    .I_2_0(n953_I_2_0),
    .O_0_0(n953_O_0_0)
  );
  InitialDelayCounter_5 InitialDelayCounter_1 ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_1_clock),
    .reset(InitialDelayCounter_1_reset),
    .valid_down(InitialDelayCounter_1_valid_down)
  );
  Map2S_65 n956 ( // @[Top.scala 606:22]
    .valid_up(n956_valid_up),
    .valid_down(n956_valid_down),
    .I0_0_0(n956_I0_0_0),
    .O_0_0_t0b(n956_O_0_0_t0b),
    .O_0_0_t1b(n956_O_0_0_t1b)
  );
  MapS_58 n967 ( // @[Top.scala 610:22]
    .clock(n967_clock),
    .reset(n967_reset),
    .valid_up(n967_valid_up),
    .valid_down(n967_valid_down),
    .I_0_0_t0b(n967_I_0_0_t0b),
    .I_0_0_t1b(n967_I_0_0_t1b),
    .O_0_0(n967_O_0_0)
  );
  assign valid_down = n967_valid_down; // @[Top.scala 614:16]
  assign O_0_0 = n967_O_0_0; // @[Top.scala 613:7]
  assign InitialDelayCounter_clock = clock;
  assign InitialDelayCounter_reset = reset;
  assign n932_valid_up = valid_up & InitialDelayCounter_valid_down; // @[Top.scala 595:19]
  assign n932_I0_0_0 = I_0_0; // @[Top.scala 593:13]
  assign n932_I0_0_1 = I_0_1; // @[Top.scala 593:13]
  assign n932_I0_0_2 = I_0_2; // @[Top.scala 593:13]
  assign n932_I0_1_0 = I_1_0; // @[Top.scala 593:13]
  assign n932_I0_1_1 = I_1_1; // @[Top.scala 593:13]
  assign n932_I0_1_2 = I_1_2; // @[Top.scala 593:13]
  assign n932_I0_2_0 = I_2_0; // @[Top.scala 593:13]
  assign n932_I0_2_1 = I_2_1; // @[Top.scala 593:13]
  assign n932_I0_2_2 = I_2_2; // @[Top.scala 593:13]
  assign n943_clock = clock;
  assign n943_reset = reset;
  assign n943_valid_up = n932_valid_down; // @[Top.scala 598:19]
  assign n943_I_0_0_t0b = n932_O_0_0_t0b; // @[Top.scala 597:12]
  assign n943_I_0_0_t1b = n932_O_0_0_t1b; // @[Top.scala 597:12]
  assign n943_I_0_1_t0b = n932_O_0_1_t0b; // @[Top.scala 597:12]
  assign n943_I_0_1_t1b = n932_O_0_1_t1b; // @[Top.scala 597:12]
  assign n943_I_0_2_t0b = n932_O_0_2_t0b; // @[Top.scala 597:12]
  assign n943_I_0_2_t1b = n932_O_0_2_t1b; // @[Top.scala 597:12]
  assign n943_I_1_0_t0b = n932_O_1_0_t0b; // @[Top.scala 597:12]
  assign n943_I_1_0_t1b = n932_O_1_0_t1b; // @[Top.scala 597:12]
  assign n943_I_1_1_t0b = n932_O_1_1_t0b; // @[Top.scala 597:12]
  assign n943_I_1_1_t1b = n932_O_1_1_t1b; // @[Top.scala 597:12]
  assign n943_I_1_2_t0b = n932_O_1_2_t0b; // @[Top.scala 597:12]
  assign n943_I_1_2_t1b = n932_O_1_2_t1b; // @[Top.scala 597:12]
  assign n943_I_2_0_t0b = n932_O_2_0_t0b; // @[Top.scala 597:12]
  assign n943_I_2_0_t1b = n932_O_2_0_t1b; // @[Top.scala 597:12]
  assign n943_I_2_1_t0b = n932_O_2_1_t0b; // @[Top.scala 597:12]
  assign n943_I_2_1_t1b = n932_O_2_1_t1b; // @[Top.scala 597:12]
  assign n943_I_2_2_t0b = n932_O_2_2_t0b; // @[Top.scala 597:12]
  assign n943_I_2_2_t1b = n932_O_2_2_t1b; // @[Top.scala 597:12]
  assign n948_clock = clock;
  assign n948_reset = reset;
  assign n948_valid_up = n943_valid_down; // @[Top.scala 601:19]
  assign n948_I_0_0 = n943_O_0_0; // @[Top.scala 600:12]
  assign n948_I_0_1 = n943_O_0_1; // @[Top.scala 600:12]
  assign n948_I_0_2 = n943_O_0_2; // @[Top.scala 600:12]
  assign n948_I_1_0 = n943_O_1_0; // @[Top.scala 600:12]
  assign n948_I_1_1 = n943_O_1_1; // @[Top.scala 600:12]
  assign n948_I_1_2 = n943_O_1_2; // @[Top.scala 600:12]
  assign n948_I_2_0 = n943_O_2_0; // @[Top.scala 600:12]
  assign n948_I_2_1 = n943_O_2_1; // @[Top.scala 600:12]
  assign n948_I_2_2 = n943_O_2_2; // @[Top.scala 600:12]
  assign n953_clock = clock;
  assign n953_reset = reset;
  assign n953_valid_up = n948_valid_down; // @[Top.scala 604:19]
  assign n953_I_0_0 = n948_O_0_0; // @[Top.scala 603:12]
  assign n953_I_1_0 = n948_O_1_0; // @[Top.scala 603:12]
  assign n953_I_2_0 = n948_O_2_0; // @[Top.scala 603:12]
  assign InitialDelayCounter_1_clock = clock;
  assign InitialDelayCounter_1_reset = reset;
  assign n956_valid_up = n953_valid_down & InitialDelayCounter_1_valid_down; // @[Top.scala 609:19]
  assign n956_I0_0_0 = n953_O_0_0; // @[Top.scala 607:13]
  assign n967_clock = clock;
  assign n967_reset = reset;
  assign n967_valid_up = n956_valid_down; // @[Top.scala 612:19]
  assign n967_I_0_0_t0b = n956_O_0_0_t0b; // @[Top.scala 611:12]
  assign n967_I_0_0_t1b = n956_O_0_0_t1b; // @[Top.scala 611:12]
endmodule
module MapS_81(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0_0,
  input  [31:0] I_0_0_1,
  input  [31:0] I_0_0_2,
  input  [31:0] I_0_1_0,
  input  [31:0] I_0_1_1,
  input  [31:0] I_0_1_2,
  input  [31:0] I_0_2_0,
  input  [31:0] I_0_2_1,
  input  [31:0] I_0_2_2,
  input  [31:0] I_1_0_0,
  input  [31:0] I_1_0_1,
  input  [31:0] I_1_0_2,
  input  [31:0] I_1_1_0,
  input  [31:0] I_1_1_1,
  input  [31:0] I_1_1_2,
  input  [31:0] I_1_2_0,
  input  [31:0] I_1_2_1,
  input  [31:0] I_1_2_2,
  input  [31:0] I_2_0_0,
  input  [31:0] I_2_0_1,
  input  [31:0] I_2_0_2,
  input  [31:0] I_2_1_0,
  input  [31:0] I_2_1_1,
  input  [31:0] I_2_1_2,
  input  [31:0] I_2_2_0,
  input  [31:0] I_2_2_1,
  input  [31:0] I_2_2_2,
  input  [31:0] I_3_0_0,
  input  [31:0] I_3_0_1,
  input  [31:0] I_3_0_2,
  input  [31:0] I_3_1_0,
  input  [31:0] I_3_1_1,
  input  [31:0] I_3_1_2,
  input  [31:0] I_3_2_0,
  input  [31:0] I_3_2_1,
  input  [31:0] I_3_2_2,
  input  [31:0] I_4_0_0,
  input  [31:0] I_4_0_1,
  input  [31:0] I_4_0_2,
  input  [31:0] I_4_1_0,
  input  [31:0] I_4_1_1,
  input  [31:0] I_4_1_2,
  input  [31:0] I_4_2_0,
  input  [31:0] I_4_2_1,
  input  [31:0] I_4_2_2,
  input  [31:0] I_5_0_0,
  input  [31:0] I_5_0_1,
  input  [31:0] I_5_0_2,
  input  [31:0] I_5_1_0,
  input  [31:0] I_5_1_1,
  input  [31:0] I_5_1_2,
  input  [31:0] I_5_2_0,
  input  [31:0] I_5_2_1,
  input  [31:0] I_5_2_2,
  input  [31:0] I_6_0_0,
  input  [31:0] I_6_0_1,
  input  [31:0] I_6_0_2,
  input  [31:0] I_6_1_0,
  input  [31:0] I_6_1_1,
  input  [31:0] I_6_1_2,
  input  [31:0] I_6_2_0,
  input  [31:0] I_6_2_1,
  input  [31:0] I_6_2_2,
  input  [31:0] I_7_0_0,
  input  [31:0] I_7_0_1,
  input  [31:0] I_7_0_2,
  input  [31:0] I_7_1_0,
  input  [31:0] I_7_1_1,
  input  [31:0] I_7_1_2,
  input  [31:0] I_7_2_0,
  input  [31:0] I_7_2_1,
  input  [31:0] I_7_2_2,
  output [31:0] O_0_0_0,
  output [31:0] O_1_0_0,
  output [31:0] O_2_0_0,
  output [31:0] O_3_0_0,
  output [31:0] O_4_0_0,
  output [31:0] O_5_0_0,
  output [31:0] O_6_0_0,
  output [31:0] O_7_0_0
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_0; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_1; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_2; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_1_0; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_1_1; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_1_2; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_2_0; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_2_1; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_2_2; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_0_0; // @[MapS.scala 9:22]
  wire  other_ops_0_clock; // @[MapS.scala 10:86]
  wire  other_ops_0_reset; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_2_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_1_clock; // @[MapS.scala 10:86]
  wire  other_ops_1_reset; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_2_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_2_clock; // @[MapS.scala 10:86]
  wire  other_ops_2_reset; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_2_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_3_clock; // @[MapS.scala 10:86]
  wire  other_ops_3_reset; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_2_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_4_clock; // @[MapS.scala 10:86]
  wire  other_ops_4_reset; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_2_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_5_clock; // @[MapS.scala 10:86]
  wire  other_ops_5_reset; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_2_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_6_clock; // @[MapS.scala 10:86]
  wire  other_ops_6_reset; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_2_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_O_0_0; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  wire  _T_1; // @[MapS.scala 23:83]
  wire  _T_2; // @[MapS.scala 23:83]
  wire  _T_3; // @[MapS.scala 23:83]
  wire  _T_4; // @[MapS.scala 23:83]
  wire  _T_5; // @[MapS.scala 23:83]
  Module_14 fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_0(fst_op_I_0_0),
    .I_0_1(fst_op_I_0_1),
    .I_0_2(fst_op_I_0_2),
    .I_1_0(fst_op_I_1_0),
    .I_1_1(fst_op_I_1_1),
    .I_1_2(fst_op_I_1_2),
    .I_2_0(fst_op_I_2_0),
    .I_2_1(fst_op_I_2_1),
    .I_2_2(fst_op_I_2_2),
    .O_0_0(fst_op_O_0_0)
  );
  Module_14 other_ops_0 ( // @[MapS.scala 10:86]
    .clock(other_ops_0_clock),
    .reset(other_ops_0_reset),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_0(other_ops_0_I_0_0),
    .I_0_1(other_ops_0_I_0_1),
    .I_0_2(other_ops_0_I_0_2),
    .I_1_0(other_ops_0_I_1_0),
    .I_1_1(other_ops_0_I_1_1),
    .I_1_2(other_ops_0_I_1_2),
    .I_2_0(other_ops_0_I_2_0),
    .I_2_1(other_ops_0_I_2_1),
    .I_2_2(other_ops_0_I_2_2),
    .O_0_0(other_ops_0_O_0_0)
  );
  Module_14 other_ops_1 ( // @[MapS.scala 10:86]
    .clock(other_ops_1_clock),
    .reset(other_ops_1_reset),
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0_0(other_ops_1_I_0_0),
    .I_0_1(other_ops_1_I_0_1),
    .I_0_2(other_ops_1_I_0_2),
    .I_1_0(other_ops_1_I_1_0),
    .I_1_1(other_ops_1_I_1_1),
    .I_1_2(other_ops_1_I_1_2),
    .I_2_0(other_ops_1_I_2_0),
    .I_2_1(other_ops_1_I_2_1),
    .I_2_2(other_ops_1_I_2_2),
    .O_0_0(other_ops_1_O_0_0)
  );
  Module_14 other_ops_2 ( // @[MapS.scala 10:86]
    .clock(other_ops_2_clock),
    .reset(other_ops_2_reset),
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I_0_0(other_ops_2_I_0_0),
    .I_0_1(other_ops_2_I_0_1),
    .I_0_2(other_ops_2_I_0_2),
    .I_1_0(other_ops_2_I_1_0),
    .I_1_1(other_ops_2_I_1_1),
    .I_1_2(other_ops_2_I_1_2),
    .I_2_0(other_ops_2_I_2_0),
    .I_2_1(other_ops_2_I_2_1),
    .I_2_2(other_ops_2_I_2_2),
    .O_0_0(other_ops_2_O_0_0)
  );
  Module_14 other_ops_3 ( // @[MapS.scala 10:86]
    .clock(other_ops_3_clock),
    .reset(other_ops_3_reset),
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I_0_0(other_ops_3_I_0_0),
    .I_0_1(other_ops_3_I_0_1),
    .I_0_2(other_ops_3_I_0_2),
    .I_1_0(other_ops_3_I_1_0),
    .I_1_1(other_ops_3_I_1_1),
    .I_1_2(other_ops_3_I_1_2),
    .I_2_0(other_ops_3_I_2_0),
    .I_2_1(other_ops_3_I_2_1),
    .I_2_2(other_ops_3_I_2_2),
    .O_0_0(other_ops_3_O_0_0)
  );
  Module_14 other_ops_4 ( // @[MapS.scala 10:86]
    .clock(other_ops_4_clock),
    .reset(other_ops_4_reset),
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I_0_0(other_ops_4_I_0_0),
    .I_0_1(other_ops_4_I_0_1),
    .I_0_2(other_ops_4_I_0_2),
    .I_1_0(other_ops_4_I_1_0),
    .I_1_1(other_ops_4_I_1_1),
    .I_1_2(other_ops_4_I_1_2),
    .I_2_0(other_ops_4_I_2_0),
    .I_2_1(other_ops_4_I_2_1),
    .I_2_2(other_ops_4_I_2_2),
    .O_0_0(other_ops_4_O_0_0)
  );
  Module_14 other_ops_5 ( // @[MapS.scala 10:86]
    .clock(other_ops_5_clock),
    .reset(other_ops_5_reset),
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I_0_0(other_ops_5_I_0_0),
    .I_0_1(other_ops_5_I_0_1),
    .I_0_2(other_ops_5_I_0_2),
    .I_1_0(other_ops_5_I_1_0),
    .I_1_1(other_ops_5_I_1_1),
    .I_1_2(other_ops_5_I_1_2),
    .I_2_0(other_ops_5_I_2_0),
    .I_2_1(other_ops_5_I_2_1),
    .I_2_2(other_ops_5_I_2_2),
    .O_0_0(other_ops_5_O_0_0)
  );
  Module_14 other_ops_6 ( // @[MapS.scala 10:86]
    .clock(other_ops_6_clock),
    .reset(other_ops_6_reset),
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I_0_0(other_ops_6_I_0_0),
    .I_0_1(other_ops_6_I_0_1),
    .I_0_2(other_ops_6_I_0_2),
    .I_1_0(other_ops_6_I_1_0),
    .I_1_1(other_ops_6_I_1_1),
    .I_1_2(other_ops_6_I_1_2),
    .I_2_0(other_ops_6_I_2_0),
    .I_2_1(other_ops_6_I_2_1),
    .I_2_2(other_ops_6_I_2_2),
    .O_0_0(other_ops_6_O_0_0)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[MapS.scala 23:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[MapS.scala 23:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[MapS.scala 23:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[MapS.scala 23:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T_5 & other_ops_6_valid_down; // @[MapS.scala 23:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[MapS.scala 17:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[MapS.scala 21:12]
  assign O_2_0_0 = other_ops_1_O_0_0; // @[MapS.scala 21:12]
  assign O_3_0_0 = other_ops_2_O_0_0; // @[MapS.scala 21:12]
  assign O_4_0_0 = other_ops_3_O_0_0; // @[MapS.scala 21:12]
  assign O_5_0_0 = other_ops_4_O_0_0; // @[MapS.scala 21:12]
  assign O_6_0_0 = other_ops_5_O_0_0; // @[MapS.scala 21:12]
  assign O_7_0_0 = other_ops_6_O_0_0; // @[MapS.scala 21:12]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_0 = I_0_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_1 = I_0_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_2 = I_0_0_2; // @[MapS.scala 16:12]
  assign fst_op_I_1_0 = I_0_1_0; // @[MapS.scala 16:12]
  assign fst_op_I_1_1 = I_0_1_1; // @[MapS.scala 16:12]
  assign fst_op_I_1_2 = I_0_1_2; // @[MapS.scala 16:12]
  assign fst_op_I_2_0 = I_0_2_0; // @[MapS.scala 16:12]
  assign fst_op_I_2_1 = I_0_2_1; // @[MapS.scala 16:12]
  assign fst_op_I_2_2 = I_0_2_2; // @[MapS.scala 16:12]
  assign other_ops_0_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_0_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_0 = I_1_0_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1 = I_1_0_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2 = I_1_0_2; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_0 = I_1_1_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_1 = I_1_1_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_2 = I_1_1_2; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_0 = I_1_2_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_1 = I_1_2_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_2 = I_1_2_2; // @[MapS.scala 20:41]
  assign other_ops_1_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_1_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0_0 = I_2_0_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1 = I_2_0_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2 = I_2_0_2; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_0 = I_2_1_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_1 = I_2_1_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_2 = I_2_1_2; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_0 = I_2_2_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_1 = I_2_2_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_2 = I_2_2_2; // @[MapS.scala 20:41]
  assign other_ops_2_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_2_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_2_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_2_I_0_0 = I_3_0_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1 = I_3_0_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2 = I_3_0_2; // @[MapS.scala 20:41]
  assign other_ops_2_I_1_0 = I_3_1_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_1_1 = I_3_1_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_1_2 = I_3_1_2; // @[MapS.scala 20:41]
  assign other_ops_2_I_2_0 = I_3_2_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_2_1 = I_3_2_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_2_2 = I_3_2_2; // @[MapS.scala 20:41]
  assign other_ops_3_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_3_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_3_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_3_I_0_0 = I_4_0_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_1 = I_4_0_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_2 = I_4_0_2; // @[MapS.scala 20:41]
  assign other_ops_3_I_1_0 = I_4_1_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_1_1 = I_4_1_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_1_2 = I_4_1_2; // @[MapS.scala 20:41]
  assign other_ops_3_I_2_0 = I_4_2_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_2_1 = I_4_2_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_2_2 = I_4_2_2; // @[MapS.scala 20:41]
  assign other_ops_4_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_4_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_4_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_4_I_0_0 = I_5_0_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_1 = I_5_0_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_2 = I_5_0_2; // @[MapS.scala 20:41]
  assign other_ops_4_I_1_0 = I_5_1_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_1_1 = I_5_1_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_1_2 = I_5_1_2; // @[MapS.scala 20:41]
  assign other_ops_4_I_2_0 = I_5_2_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_2_1 = I_5_2_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_2_2 = I_5_2_2; // @[MapS.scala 20:41]
  assign other_ops_5_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_5_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_5_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_5_I_0_0 = I_6_0_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_1 = I_6_0_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_2 = I_6_0_2; // @[MapS.scala 20:41]
  assign other_ops_5_I_1_0 = I_6_1_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_1_1 = I_6_1_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_1_2 = I_6_1_2; // @[MapS.scala 20:41]
  assign other_ops_5_I_2_0 = I_6_2_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_2_1 = I_6_2_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_2_2 = I_6_2_2; // @[MapS.scala 20:41]
  assign other_ops_6_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_6_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_6_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_6_I_0_0 = I_7_0_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_1 = I_7_0_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_2 = I_7_0_2; // @[MapS.scala 20:41]
  assign other_ops_6_I_1_0 = I_7_1_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_1_1 = I_7_1_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_1_2 = I_7_1_2; // @[MapS.scala 20:41]
  assign other_ops_6_I_2_0 = I_7_2_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_2_1 = I_7_2_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_2_2 = I_7_2_2; // @[MapS.scala 20:41]
endmodule
module MapT_42(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0_0,
  input  [31:0] I_0_0_1,
  input  [31:0] I_0_0_2,
  input  [31:0] I_0_1_0,
  input  [31:0] I_0_1_1,
  input  [31:0] I_0_1_2,
  input  [31:0] I_0_2_0,
  input  [31:0] I_0_2_1,
  input  [31:0] I_0_2_2,
  input  [31:0] I_1_0_0,
  input  [31:0] I_1_0_1,
  input  [31:0] I_1_0_2,
  input  [31:0] I_1_1_0,
  input  [31:0] I_1_1_1,
  input  [31:0] I_1_1_2,
  input  [31:0] I_1_2_0,
  input  [31:0] I_1_2_1,
  input  [31:0] I_1_2_2,
  input  [31:0] I_2_0_0,
  input  [31:0] I_2_0_1,
  input  [31:0] I_2_0_2,
  input  [31:0] I_2_1_0,
  input  [31:0] I_2_1_1,
  input  [31:0] I_2_1_2,
  input  [31:0] I_2_2_0,
  input  [31:0] I_2_2_1,
  input  [31:0] I_2_2_2,
  input  [31:0] I_3_0_0,
  input  [31:0] I_3_0_1,
  input  [31:0] I_3_0_2,
  input  [31:0] I_3_1_0,
  input  [31:0] I_3_1_1,
  input  [31:0] I_3_1_2,
  input  [31:0] I_3_2_0,
  input  [31:0] I_3_2_1,
  input  [31:0] I_3_2_2,
  input  [31:0] I_4_0_0,
  input  [31:0] I_4_0_1,
  input  [31:0] I_4_0_2,
  input  [31:0] I_4_1_0,
  input  [31:0] I_4_1_1,
  input  [31:0] I_4_1_2,
  input  [31:0] I_4_2_0,
  input  [31:0] I_4_2_1,
  input  [31:0] I_4_2_2,
  input  [31:0] I_5_0_0,
  input  [31:0] I_5_0_1,
  input  [31:0] I_5_0_2,
  input  [31:0] I_5_1_0,
  input  [31:0] I_5_1_1,
  input  [31:0] I_5_1_2,
  input  [31:0] I_5_2_0,
  input  [31:0] I_5_2_1,
  input  [31:0] I_5_2_2,
  input  [31:0] I_6_0_0,
  input  [31:0] I_6_0_1,
  input  [31:0] I_6_0_2,
  input  [31:0] I_6_1_0,
  input  [31:0] I_6_1_1,
  input  [31:0] I_6_1_2,
  input  [31:0] I_6_2_0,
  input  [31:0] I_6_2_1,
  input  [31:0] I_6_2_2,
  input  [31:0] I_7_0_0,
  input  [31:0] I_7_0_1,
  input  [31:0] I_7_0_2,
  input  [31:0] I_7_1_0,
  input  [31:0] I_7_1_1,
  input  [31:0] I_7_1_2,
  input  [31:0] I_7_2_0,
  input  [31:0] I_7_2_1,
  input  [31:0] I_7_2_2,
  output [31:0] O_0_0_0,
  output [31:0] O_1_0_0,
  output [31:0] O_2_0_0,
  output [31:0] O_3_0_0,
  output [31:0] O_4_0_0,
  output [31:0] O_5_0_0,
  output [31:0] O_6_0_0,
  output [31:0] O_7_0_0
);
  wire  op_clock; // @[MapT.scala 8:20]
  wire  op_reset; // @[MapT.scala 8:20]
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_0_0; // @[MapT.scala 8:20]
  MapS_81 op ( // @[MapT.scala 8:20]
    .clock(op_clock),
    .reset(op_reset),
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0(op_I_0_0_0),
    .I_0_0_1(op_I_0_0_1),
    .I_0_0_2(op_I_0_0_2),
    .I_0_1_0(op_I_0_1_0),
    .I_0_1_1(op_I_0_1_1),
    .I_0_1_2(op_I_0_1_2),
    .I_0_2_0(op_I_0_2_0),
    .I_0_2_1(op_I_0_2_1),
    .I_0_2_2(op_I_0_2_2),
    .I_1_0_0(op_I_1_0_0),
    .I_1_0_1(op_I_1_0_1),
    .I_1_0_2(op_I_1_0_2),
    .I_1_1_0(op_I_1_1_0),
    .I_1_1_1(op_I_1_1_1),
    .I_1_1_2(op_I_1_1_2),
    .I_1_2_0(op_I_1_2_0),
    .I_1_2_1(op_I_1_2_1),
    .I_1_2_2(op_I_1_2_2),
    .I_2_0_0(op_I_2_0_0),
    .I_2_0_1(op_I_2_0_1),
    .I_2_0_2(op_I_2_0_2),
    .I_2_1_0(op_I_2_1_0),
    .I_2_1_1(op_I_2_1_1),
    .I_2_1_2(op_I_2_1_2),
    .I_2_2_0(op_I_2_2_0),
    .I_2_2_1(op_I_2_2_1),
    .I_2_2_2(op_I_2_2_2),
    .I_3_0_0(op_I_3_0_0),
    .I_3_0_1(op_I_3_0_1),
    .I_3_0_2(op_I_3_0_2),
    .I_3_1_0(op_I_3_1_0),
    .I_3_1_1(op_I_3_1_1),
    .I_3_1_2(op_I_3_1_2),
    .I_3_2_0(op_I_3_2_0),
    .I_3_2_1(op_I_3_2_1),
    .I_3_2_2(op_I_3_2_2),
    .I_4_0_0(op_I_4_0_0),
    .I_4_0_1(op_I_4_0_1),
    .I_4_0_2(op_I_4_0_2),
    .I_4_1_0(op_I_4_1_0),
    .I_4_1_1(op_I_4_1_1),
    .I_4_1_2(op_I_4_1_2),
    .I_4_2_0(op_I_4_2_0),
    .I_4_2_1(op_I_4_2_1),
    .I_4_2_2(op_I_4_2_2),
    .I_5_0_0(op_I_5_0_0),
    .I_5_0_1(op_I_5_0_1),
    .I_5_0_2(op_I_5_0_2),
    .I_5_1_0(op_I_5_1_0),
    .I_5_1_1(op_I_5_1_1),
    .I_5_1_2(op_I_5_1_2),
    .I_5_2_0(op_I_5_2_0),
    .I_5_2_1(op_I_5_2_1),
    .I_5_2_2(op_I_5_2_2),
    .I_6_0_0(op_I_6_0_0),
    .I_6_0_1(op_I_6_0_1),
    .I_6_0_2(op_I_6_0_2),
    .I_6_1_0(op_I_6_1_0),
    .I_6_1_1(op_I_6_1_1),
    .I_6_1_2(op_I_6_1_2),
    .I_6_2_0(op_I_6_2_0),
    .I_6_2_1(op_I_6_2_1),
    .I_6_2_2(op_I_6_2_2),
    .I_7_0_0(op_I_7_0_0),
    .I_7_0_1(op_I_7_0_1),
    .I_7_0_2(op_I_7_0_2),
    .I_7_1_0(op_I_7_1_0),
    .I_7_1_1(op_I_7_1_1),
    .I_7_1_2(op_I_7_1_2),
    .I_7_2_0(op_I_7_2_0),
    .I_7_2_1(op_I_7_2_1),
    .I_7_2_2(op_I_7_2_2),
    .O_0_0_0(op_O_0_0_0),
    .O_1_0_0(op_O_1_0_0),
    .O_2_0_0(op_O_2_0_0),
    .O_3_0_0(op_O_3_0_0),
    .O_4_0_0(op_O_4_0_0),
    .O_5_0_0(op_O_5_0_0),
    .O_6_0_0(op_O_6_0_0),
    .O_7_0_0(op_O_7_0_0)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0 = op_O_0_0_0; // @[MapT.scala 15:7]
  assign O_1_0_0 = op_O_1_0_0; // @[MapT.scala 15:7]
  assign O_2_0_0 = op_O_2_0_0; // @[MapT.scala 15:7]
  assign O_3_0_0 = op_O_3_0_0; // @[MapT.scala 15:7]
  assign O_4_0_0 = op_O_4_0_0; // @[MapT.scala 15:7]
  assign O_5_0_0 = op_O_5_0_0; // @[MapT.scala 15:7]
  assign O_6_0_0 = op_O_6_0_0; // @[MapT.scala 15:7]
  assign O_7_0_0 = op_O_7_0_0; // @[MapT.scala 15:7]
  assign op_clock = clock;
  assign op_reset = reset;
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0 = I_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_1 = I_0_0_1; // @[MapT.scala 14:10]
  assign op_I_0_0_2 = I_0_0_2; // @[MapT.scala 14:10]
  assign op_I_0_1_0 = I_0_1_0; // @[MapT.scala 14:10]
  assign op_I_0_1_1 = I_0_1_1; // @[MapT.scala 14:10]
  assign op_I_0_1_2 = I_0_1_2; // @[MapT.scala 14:10]
  assign op_I_0_2_0 = I_0_2_0; // @[MapT.scala 14:10]
  assign op_I_0_2_1 = I_0_2_1; // @[MapT.scala 14:10]
  assign op_I_0_2_2 = I_0_2_2; // @[MapT.scala 14:10]
  assign op_I_1_0_0 = I_1_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_1 = I_1_0_1; // @[MapT.scala 14:10]
  assign op_I_1_0_2 = I_1_0_2; // @[MapT.scala 14:10]
  assign op_I_1_1_0 = I_1_1_0; // @[MapT.scala 14:10]
  assign op_I_1_1_1 = I_1_1_1; // @[MapT.scala 14:10]
  assign op_I_1_1_2 = I_1_1_2; // @[MapT.scala 14:10]
  assign op_I_1_2_0 = I_1_2_0; // @[MapT.scala 14:10]
  assign op_I_1_2_1 = I_1_2_1; // @[MapT.scala 14:10]
  assign op_I_1_2_2 = I_1_2_2; // @[MapT.scala 14:10]
  assign op_I_2_0_0 = I_2_0_0; // @[MapT.scala 14:10]
  assign op_I_2_0_1 = I_2_0_1; // @[MapT.scala 14:10]
  assign op_I_2_0_2 = I_2_0_2; // @[MapT.scala 14:10]
  assign op_I_2_1_0 = I_2_1_0; // @[MapT.scala 14:10]
  assign op_I_2_1_1 = I_2_1_1; // @[MapT.scala 14:10]
  assign op_I_2_1_2 = I_2_1_2; // @[MapT.scala 14:10]
  assign op_I_2_2_0 = I_2_2_0; // @[MapT.scala 14:10]
  assign op_I_2_2_1 = I_2_2_1; // @[MapT.scala 14:10]
  assign op_I_2_2_2 = I_2_2_2; // @[MapT.scala 14:10]
  assign op_I_3_0_0 = I_3_0_0; // @[MapT.scala 14:10]
  assign op_I_3_0_1 = I_3_0_1; // @[MapT.scala 14:10]
  assign op_I_3_0_2 = I_3_0_2; // @[MapT.scala 14:10]
  assign op_I_3_1_0 = I_3_1_0; // @[MapT.scala 14:10]
  assign op_I_3_1_1 = I_3_1_1; // @[MapT.scala 14:10]
  assign op_I_3_1_2 = I_3_1_2; // @[MapT.scala 14:10]
  assign op_I_3_2_0 = I_3_2_0; // @[MapT.scala 14:10]
  assign op_I_3_2_1 = I_3_2_1; // @[MapT.scala 14:10]
  assign op_I_3_2_2 = I_3_2_2; // @[MapT.scala 14:10]
  assign op_I_4_0_0 = I_4_0_0; // @[MapT.scala 14:10]
  assign op_I_4_0_1 = I_4_0_1; // @[MapT.scala 14:10]
  assign op_I_4_0_2 = I_4_0_2; // @[MapT.scala 14:10]
  assign op_I_4_1_0 = I_4_1_0; // @[MapT.scala 14:10]
  assign op_I_4_1_1 = I_4_1_1; // @[MapT.scala 14:10]
  assign op_I_4_1_2 = I_4_1_2; // @[MapT.scala 14:10]
  assign op_I_4_2_0 = I_4_2_0; // @[MapT.scala 14:10]
  assign op_I_4_2_1 = I_4_2_1; // @[MapT.scala 14:10]
  assign op_I_4_2_2 = I_4_2_2; // @[MapT.scala 14:10]
  assign op_I_5_0_0 = I_5_0_0; // @[MapT.scala 14:10]
  assign op_I_5_0_1 = I_5_0_1; // @[MapT.scala 14:10]
  assign op_I_5_0_2 = I_5_0_2; // @[MapT.scala 14:10]
  assign op_I_5_1_0 = I_5_1_0; // @[MapT.scala 14:10]
  assign op_I_5_1_1 = I_5_1_1; // @[MapT.scala 14:10]
  assign op_I_5_1_2 = I_5_1_2; // @[MapT.scala 14:10]
  assign op_I_5_2_0 = I_5_2_0; // @[MapT.scala 14:10]
  assign op_I_5_2_1 = I_5_2_1; // @[MapT.scala 14:10]
  assign op_I_5_2_2 = I_5_2_2; // @[MapT.scala 14:10]
  assign op_I_6_0_0 = I_6_0_0; // @[MapT.scala 14:10]
  assign op_I_6_0_1 = I_6_0_1; // @[MapT.scala 14:10]
  assign op_I_6_0_2 = I_6_0_2; // @[MapT.scala 14:10]
  assign op_I_6_1_0 = I_6_1_0; // @[MapT.scala 14:10]
  assign op_I_6_1_1 = I_6_1_1; // @[MapT.scala 14:10]
  assign op_I_6_1_2 = I_6_1_2; // @[MapT.scala 14:10]
  assign op_I_6_2_0 = I_6_2_0; // @[MapT.scala 14:10]
  assign op_I_6_2_1 = I_6_2_1; // @[MapT.scala 14:10]
  assign op_I_6_2_2 = I_6_2_2; // @[MapT.scala 14:10]
  assign op_I_7_0_0 = I_7_0_0; // @[MapT.scala 14:10]
  assign op_I_7_0_1 = I_7_0_1; // @[MapT.scala 14:10]
  assign op_I_7_0_2 = I_7_0_2; // @[MapT.scala 14:10]
  assign op_I_7_1_0 = I_7_1_0; // @[MapT.scala 14:10]
  assign op_I_7_1_1 = I_7_1_1; // @[MapT.scala 14:10]
  assign op_I_7_1_2 = I_7_1_2; // @[MapT.scala 14:10]
  assign op_I_7_2_0 = I_7_2_0; // @[MapT.scala 14:10]
  assign op_I_7_2_1 = I_7_2_1; // @[MapT.scala 14:10]
  assign op_I_7_2_2 = I_7_2_2; // @[MapT.scala 14:10]
endmodule
module Map2S_93(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0,
  input  [31:0] I0_1,
  input  [31:0] I0_2,
  input  [31:0] I0_3,
  input  [31:0] I0_4,
  input  [31:0] I0_5,
  input  [31:0] I0_6,
  input  [31:0] I0_7,
  input  [31:0] I1_0,
  input  [31:0] I1_1,
  input  [31:0] I1_2,
  input  [31:0] I1_3,
  input  [31:0] I1_4,
  input  [31:0] I1_5,
  input  [31:0] I1_6,
  input  [31:0] I1_7,
  output [31:0] O_0_t0b,
  output [31:0] O_0_t1b,
  output [31:0] O_1_t0b,
  output [31:0] O_1_t1b,
  output [31:0] O_2_t0b,
  output [31:0] O_2_t1b,
  output [31:0] O_3_t0b,
  output [31:0] O_3_t1b,
  output [31:0] O_4_t0b,
  output [31:0] O_4_t1b,
  output [31:0] O_5_t0b,
  output [31:0] O_5_t1b,
  output [31:0] O_6_t0b,
  output [31:0] O_6_t1b,
  output [31:0] O_7_t0b,
  output [31:0] O_7_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_t1b; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_t1b; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  wire  _T_2; // @[Map2S.scala 26:83]
  wire  _T_3; // @[Map2S.scala 26:83]
  wire  _T_4; // @[Map2S.scala 26:83]
  wire  _T_5; // @[Map2S.scala 26:83]
  AtomTuple fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1(fst_op_I1),
    .O_t0b(fst_op_O_t0b),
    .O_t1b(fst_op_O_t1b)
  );
  AtomTuple other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0(other_ops_0_I0),
    .I1(other_ops_0_I1),
    .O_t0b(other_ops_0_O_t0b),
    .O_t1b(other_ops_0_O_t1b)
  );
  AtomTuple other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0(other_ops_1_I0),
    .I1(other_ops_1_I1),
    .O_t0b(other_ops_1_O_t0b),
    .O_t1b(other_ops_1_O_t1b)
  );
  AtomTuple other_ops_2 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0(other_ops_2_I0),
    .I1(other_ops_2_I1),
    .O_t0b(other_ops_2_O_t0b),
    .O_t1b(other_ops_2_O_t1b)
  );
  AtomTuple other_ops_3 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I0(other_ops_3_I0),
    .I1(other_ops_3_I1),
    .O_t0b(other_ops_3_O_t0b),
    .O_t1b(other_ops_3_O_t1b)
  );
  AtomTuple other_ops_4 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I0(other_ops_4_I0),
    .I1(other_ops_4_I1),
    .O_t0b(other_ops_4_O_t0b),
    .O_t1b(other_ops_4_O_t1b)
  );
  AtomTuple other_ops_5 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I0(other_ops_5_I0),
    .I1(other_ops_5_I1),
    .O_t0b(other_ops_5_O_t0b),
    .O_t1b(other_ops_5_O_t1b)
  );
  AtomTuple other_ops_6 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I0(other_ops_6_I0),
    .I1(other_ops_6_I1),
    .O_t0b(other_ops_6_O_t0b),
    .O_t1b(other_ops_6_O_t1b)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[Map2S.scala 26:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[Map2S.scala 26:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_5 & other_ops_6_valid_down; // @[Map2S.scala 26:14]
  assign O_0_t0b = fst_op_O_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b = fst_op_O_t1b; // @[Map2S.scala 19:8]
  assign O_1_t0b = other_ops_0_O_t0b; // @[Map2S.scala 24:12]
  assign O_1_t1b = other_ops_0_O_t1b; // @[Map2S.scala 24:12]
  assign O_2_t0b = other_ops_1_O_t0b; // @[Map2S.scala 24:12]
  assign O_2_t1b = other_ops_1_O_t1b; // @[Map2S.scala 24:12]
  assign O_3_t0b = other_ops_2_O_t0b; // @[Map2S.scala 24:12]
  assign O_3_t1b = other_ops_2_O_t1b; // @[Map2S.scala 24:12]
  assign O_4_t0b = other_ops_3_O_t0b; // @[Map2S.scala 24:12]
  assign O_4_t1b = other_ops_3_O_t1b; // @[Map2S.scala 24:12]
  assign O_5_t0b = other_ops_4_O_t0b; // @[Map2S.scala 24:12]
  assign O_5_t1b = other_ops_4_O_t1b; // @[Map2S.scala 24:12]
  assign O_6_t0b = other_ops_5_O_t0b; // @[Map2S.scala 24:12]
  assign O_6_t1b = other_ops_5_O_t1b; // @[Map2S.scala 24:12]
  assign O_7_t0b = other_ops_6_O_t0b; // @[Map2S.scala 24:12]
  assign O_7_t1b = other_ops_6_O_t1b; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0 = I0_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I1 = I1_1; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0 = I0_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1 = I1_2; // @[Map2S.scala 23:43]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0 = I0_3; // @[Map2S.scala 22:43]
  assign other_ops_2_I1 = I1_3; // @[Map2S.scala 23:43]
  assign other_ops_3_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_3_I0 = I0_4; // @[Map2S.scala 22:43]
  assign other_ops_3_I1 = I1_4; // @[Map2S.scala 23:43]
  assign other_ops_4_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_4_I0 = I0_5; // @[Map2S.scala 22:43]
  assign other_ops_4_I1 = I1_5; // @[Map2S.scala 23:43]
  assign other_ops_5_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_5_I0 = I0_6; // @[Map2S.scala 22:43]
  assign other_ops_5_I1 = I1_6; // @[Map2S.scala 23:43]
  assign other_ops_6_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_6_I0 = I0_7; // @[Map2S.scala 22:43]
  assign other_ops_6_I1 = I1_7; // @[Map2S.scala 23:43]
endmodule
module Map2T_37(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0,
  input  [31:0] I0_1,
  input  [31:0] I0_2,
  input  [31:0] I0_3,
  input  [31:0] I0_4,
  input  [31:0] I0_5,
  input  [31:0] I0_6,
  input  [31:0] I0_7,
  input  [31:0] I1_0,
  input  [31:0] I1_1,
  input  [31:0] I1_2,
  input  [31:0] I1_3,
  input  [31:0] I1_4,
  input  [31:0] I1_5,
  input  [31:0] I1_6,
  input  [31:0] I1_7,
  output [31:0] O_0_t0b,
  output [31:0] O_0_t1b,
  output [31:0] O_1_t0b,
  output [31:0] O_1_t1b,
  output [31:0] O_2_t0b,
  output [31:0] O_2_t1b,
  output [31:0] O_3_t0b,
  output [31:0] O_3_t1b,
  output [31:0] O_4_t0b,
  output [31:0] O_4_t1b,
  output [31:0] O_5_t0b,
  output [31:0] O_5_t1b,
  output [31:0] O_6_t0b,
  output [31:0] O_6_t1b,
  output [31:0] O_7_t0b,
  output [31:0] O_7_t1b
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_3; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_4; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_5; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_6; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_7; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_t1b; // @[Map2T.scala 8:20]
  Map2S_93 op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0(op_I0_0),
    .I0_1(op_I0_1),
    .I0_2(op_I0_2),
    .I0_3(op_I0_3),
    .I0_4(op_I0_4),
    .I0_5(op_I0_5),
    .I0_6(op_I0_6),
    .I0_7(op_I0_7),
    .I1_0(op_I1_0),
    .I1_1(op_I1_1),
    .I1_2(op_I1_2),
    .I1_3(op_I1_3),
    .I1_4(op_I1_4),
    .I1_5(op_I1_5),
    .I1_6(op_I1_6),
    .I1_7(op_I1_7),
    .O_0_t0b(op_O_0_t0b),
    .O_0_t1b(op_O_0_t1b),
    .O_1_t0b(op_O_1_t0b),
    .O_1_t1b(op_O_1_t1b),
    .O_2_t0b(op_O_2_t0b),
    .O_2_t1b(op_O_2_t1b),
    .O_3_t0b(op_O_3_t0b),
    .O_3_t1b(op_O_3_t1b),
    .O_4_t0b(op_O_4_t0b),
    .O_4_t1b(op_O_4_t1b),
    .O_5_t0b(op_O_5_t0b),
    .O_5_t1b(op_O_5_t1b),
    .O_6_t0b(op_O_6_t0b),
    .O_6_t1b(op_O_6_t1b),
    .O_7_t0b(op_O_7_t0b),
    .O_7_t1b(op_O_7_t1b)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_t0b = op_O_0_t0b; // @[Map2T.scala 17:7]
  assign O_0_t1b = op_O_0_t1b; // @[Map2T.scala 17:7]
  assign O_1_t0b = op_O_1_t0b; // @[Map2T.scala 17:7]
  assign O_1_t1b = op_O_1_t1b; // @[Map2T.scala 17:7]
  assign O_2_t0b = op_O_2_t0b; // @[Map2T.scala 17:7]
  assign O_2_t1b = op_O_2_t1b; // @[Map2T.scala 17:7]
  assign O_3_t0b = op_O_3_t0b; // @[Map2T.scala 17:7]
  assign O_3_t1b = op_O_3_t1b; // @[Map2T.scala 17:7]
  assign O_4_t0b = op_O_4_t0b; // @[Map2T.scala 17:7]
  assign O_4_t1b = op_O_4_t1b; // @[Map2T.scala 17:7]
  assign O_5_t0b = op_O_5_t0b; // @[Map2T.scala 17:7]
  assign O_5_t1b = op_O_5_t1b; // @[Map2T.scala 17:7]
  assign O_6_t0b = op_O_6_t0b; // @[Map2T.scala 17:7]
  assign O_6_t1b = op_O_6_t1b; // @[Map2T.scala 17:7]
  assign O_7_t0b = op_O_7_t0b; // @[Map2T.scala 17:7]
  assign O_7_t1b = op_O_7_t1b; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0 = I0_0; // @[Map2T.scala 15:11]
  assign op_I0_1 = I0_1; // @[Map2T.scala 15:11]
  assign op_I0_2 = I0_2; // @[Map2T.scala 15:11]
  assign op_I0_3 = I0_3; // @[Map2T.scala 15:11]
  assign op_I0_4 = I0_4; // @[Map2T.scala 15:11]
  assign op_I0_5 = I0_5; // @[Map2T.scala 15:11]
  assign op_I0_6 = I0_6; // @[Map2T.scala 15:11]
  assign op_I0_7 = I0_7; // @[Map2T.scala 15:11]
  assign op_I1_0 = I1_0; // @[Map2T.scala 16:11]
  assign op_I1_1 = I1_1; // @[Map2T.scala 16:11]
  assign op_I1_2 = I1_2; // @[Map2T.scala 16:11]
  assign op_I1_3 = I1_3; // @[Map2T.scala 16:11]
  assign op_I1_4 = I1_4; // @[Map2T.scala 16:11]
  assign op_I1_5 = I1_5; // @[Map2T.scala 16:11]
  assign op_I1_6 = I1_6; // @[Map2T.scala 16:11]
  assign op_I1_7 = I1_7; // @[Map2T.scala 16:11]
endmodule
module Map2S_94(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0,
  input  [31:0] I0_1,
  input  [31:0] I0_2,
  input  [31:0] I0_3,
  input  [31:0] I0_4,
  input  [31:0] I0_5,
  input  [31:0] I0_6,
  input  [31:0] I0_7,
  input  [31:0] I1_0_t0b,
  input  [31:0] I1_0_t1b,
  input  [31:0] I1_1_t0b,
  input  [31:0] I1_1_t1b,
  input  [31:0] I1_2_t0b,
  input  [31:0] I1_2_t1b,
  input  [31:0] I1_3_t0b,
  input  [31:0] I1_3_t1b,
  input  [31:0] I1_4_t0b,
  input  [31:0] I1_4_t1b,
  input  [31:0] I1_5_t0b,
  input  [31:0] I1_5_t1b,
  input  [31:0] I1_6_t0b,
  input  [31:0] I1_6_t1b,
  input  [31:0] I1_7_t0b,
  input  [31:0] I1_7_t1b,
  output [31:0] O_0_t0b,
  output [31:0] O_0_t1b_t0b,
  output [31:0] O_0_t1b_t1b,
  output [31:0] O_1_t0b,
  output [31:0] O_1_t1b_t0b,
  output [31:0] O_1_t1b_t1b,
  output [31:0] O_2_t0b,
  output [31:0] O_2_t1b_t0b,
  output [31:0] O_2_t1b_t1b,
  output [31:0] O_3_t0b,
  output [31:0] O_3_t1b_t0b,
  output [31:0] O_3_t1b_t1b,
  output [31:0] O_4_t0b,
  output [31:0] O_4_t1b_t0b,
  output [31:0] O_4_t1b_t1b,
  output [31:0] O_5_t0b,
  output [31:0] O_5_t1b_t0b,
  output [31:0] O_5_t1b_t1b,
  output [31:0] O_6_t0b,
  output [31:0] O_6_t1b_t0b,
  output [31:0] O_6_t1b_t1b,
  output [31:0] O_7_t0b,
  output [31:0] O_7_t1b_t0b,
  output [31:0] O_7_t1b_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_t1b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_t1b_t1b; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I1_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I1_t1b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_t1b_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_t1b_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I1_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I1_t1b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_t1b_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_t1b_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I1_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I1_t1b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_t1b_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_t1b_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I1_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I1_t1b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_t1b_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_t1b_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I1_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I1_t1b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_t1b_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_t1b_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I1_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I1_t1b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_t1b_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_t1b_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I1_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I1_t1b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_t1b_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_t1b_t1b; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  wire  _T_2; // @[Map2S.scala 26:83]
  wire  _T_3; // @[Map2S.scala 26:83]
  wire  _T_4; // @[Map2S.scala 26:83]
  wire  _T_5; // @[Map2S.scala 26:83]
  AtomTuple_10 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1_t0b(fst_op_I1_t0b),
    .I1_t1b(fst_op_I1_t1b),
    .O_t0b(fst_op_O_t0b),
    .O_t1b_t0b(fst_op_O_t1b_t0b),
    .O_t1b_t1b(fst_op_O_t1b_t1b)
  );
  AtomTuple_10 other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0(other_ops_0_I0),
    .I1_t0b(other_ops_0_I1_t0b),
    .I1_t1b(other_ops_0_I1_t1b),
    .O_t0b(other_ops_0_O_t0b),
    .O_t1b_t0b(other_ops_0_O_t1b_t0b),
    .O_t1b_t1b(other_ops_0_O_t1b_t1b)
  );
  AtomTuple_10 other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0(other_ops_1_I0),
    .I1_t0b(other_ops_1_I1_t0b),
    .I1_t1b(other_ops_1_I1_t1b),
    .O_t0b(other_ops_1_O_t0b),
    .O_t1b_t0b(other_ops_1_O_t1b_t0b),
    .O_t1b_t1b(other_ops_1_O_t1b_t1b)
  );
  AtomTuple_10 other_ops_2 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0(other_ops_2_I0),
    .I1_t0b(other_ops_2_I1_t0b),
    .I1_t1b(other_ops_2_I1_t1b),
    .O_t0b(other_ops_2_O_t0b),
    .O_t1b_t0b(other_ops_2_O_t1b_t0b),
    .O_t1b_t1b(other_ops_2_O_t1b_t1b)
  );
  AtomTuple_10 other_ops_3 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I0(other_ops_3_I0),
    .I1_t0b(other_ops_3_I1_t0b),
    .I1_t1b(other_ops_3_I1_t1b),
    .O_t0b(other_ops_3_O_t0b),
    .O_t1b_t0b(other_ops_3_O_t1b_t0b),
    .O_t1b_t1b(other_ops_3_O_t1b_t1b)
  );
  AtomTuple_10 other_ops_4 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I0(other_ops_4_I0),
    .I1_t0b(other_ops_4_I1_t0b),
    .I1_t1b(other_ops_4_I1_t1b),
    .O_t0b(other_ops_4_O_t0b),
    .O_t1b_t0b(other_ops_4_O_t1b_t0b),
    .O_t1b_t1b(other_ops_4_O_t1b_t1b)
  );
  AtomTuple_10 other_ops_5 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I0(other_ops_5_I0),
    .I1_t0b(other_ops_5_I1_t0b),
    .I1_t1b(other_ops_5_I1_t1b),
    .O_t0b(other_ops_5_O_t0b),
    .O_t1b_t0b(other_ops_5_O_t1b_t0b),
    .O_t1b_t1b(other_ops_5_O_t1b_t1b)
  );
  AtomTuple_10 other_ops_6 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I0(other_ops_6_I0),
    .I1_t0b(other_ops_6_I1_t0b),
    .I1_t1b(other_ops_6_I1_t1b),
    .O_t0b(other_ops_6_O_t0b),
    .O_t1b_t0b(other_ops_6_O_t1b_t0b),
    .O_t1b_t1b(other_ops_6_O_t1b_t1b)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[Map2S.scala 26:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[Map2S.scala 26:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_5 & other_ops_6_valid_down; // @[Map2S.scala 26:14]
  assign O_0_t0b = fst_op_O_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b_t0b = fst_op_O_t1b_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b_t1b = fst_op_O_t1b_t1b; // @[Map2S.scala 19:8]
  assign O_1_t0b = other_ops_0_O_t0b; // @[Map2S.scala 24:12]
  assign O_1_t1b_t0b = other_ops_0_O_t1b_t0b; // @[Map2S.scala 24:12]
  assign O_1_t1b_t1b = other_ops_0_O_t1b_t1b; // @[Map2S.scala 24:12]
  assign O_2_t0b = other_ops_1_O_t0b; // @[Map2S.scala 24:12]
  assign O_2_t1b_t0b = other_ops_1_O_t1b_t0b; // @[Map2S.scala 24:12]
  assign O_2_t1b_t1b = other_ops_1_O_t1b_t1b; // @[Map2S.scala 24:12]
  assign O_3_t0b = other_ops_2_O_t0b; // @[Map2S.scala 24:12]
  assign O_3_t1b_t0b = other_ops_2_O_t1b_t0b; // @[Map2S.scala 24:12]
  assign O_3_t1b_t1b = other_ops_2_O_t1b_t1b; // @[Map2S.scala 24:12]
  assign O_4_t0b = other_ops_3_O_t0b; // @[Map2S.scala 24:12]
  assign O_4_t1b_t0b = other_ops_3_O_t1b_t0b; // @[Map2S.scala 24:12]
  assign O_4_t1b_t1b = other_ops_3_O_t1b_t1b; // @[Map2S.scala 24:12]
  assign O_5_t0b = other_ops_4_O_t0b; // @[Map2S.scala 24:12]
  assign O_5_t1b_t0b = other_ops_4_O_t1b_t0b; // @[Map2S.scala 24:12]
  assign O_5_t1b_t1b = other_ops_4_O_t1b_t1b; // @[Map2S.scala 24:12]
  assign O_6_t0b = other_ops_5_O_t0b; // @[Map2S.scala 24:12]
  assign O_6_t1b_t0b = other_ops_5_O_t1b_t0b; // @[Map2S.scala 24:12]
  assign O_6_t1b_t1b = other_ops_5_O_t1b_t1b; // @[Map2S.scala 24:12]
  assign O_7_t0b = other_ops_6_O_t0b; // @[Map2S.scala 24:12]
  assign O_7_t1b_t0b = other_ops_6_O_t1b_t0b; // @[Map2S.scala 24:12]
  assign O_7_t1b_t1b = other_ops_6_O_t1b_t1b; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1_t0b = I1_0_t0b; // @[Map2S.scala 18:13]
  assign fst_op_I1_t1b = I1_0_t1b; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0 = I0_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I1_t0b = I1_1_t0b; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_t1b = I1_1_t1b; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0 = I0_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1_t0b = I1_2_t0b; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_t1b = I1_2_t1b; // @[Map2S.scala 23:43]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0 = I0_3; // @[Map2S.scala 22:43]
  assign other_ops_2_I1_t0b = I1_3_t0b; // @[Map2S.scala 23:43]
  assign other_ops_2_I1_t1b = I1_3_t1b; // @[Map2S.scala 23:43]
  assign other_ops_3_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_3_I0 = I0_4; // @[Map2S.scala 22:43]
  assign other_ops_3_I1_t0b = I1_4_t0b; // @[Map2S.scala 23:43]
  assign other_ops_3_I1_t1b = I1_4_t1b; // @[Map2S.scala 23:43]
  assign other_ops_4_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_4_I0 = I0_5; // @[Map2S.scala 22:43]
  assign other_ops_4_I1_t0b = I1_5_t0b; // @[Map2S.scala 23:43]
  assign other_ops_4_I1_t1b = I1_5_t1b; // @[Map2S.scala 23:43]
  assign other_ops_5_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_5_I0 = I0_6; // @[Map2S.scala 22:43]
  assign other_ops_5_I1_t0b = I1_6_t0b; // @[Map2S.scala 23:43]
  assign other_ops_5_I1_t1b = I1_6_t1b; // @[Map2S.scala 23:43]
  assign other_ops_6_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_6_I0 = I0_7; // @[Map2S.scala 22:43]
  assign other_ops_6_I1_t0b = I1_7_t0b; // @[Map2S.scala 23:43]
  assign other_ops_6_I1_t1b = I1_7_t1b; // @[Map2S.scala 23:43]
endmodule
module Map2T_38(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0,
  input  [31:0] I0_1,
  input  [31:0] I0_2,
  input  [31:0] I0_3,
  input  [31:0] I0_4,
  input  [31:0] I0_5,
  input  [31:0] I0_6,
  input  [31:0] I0_7,
  input  [31:0] I1_0_t0b,
  input  [31:0] I1_0_t1b,
  input  [31:0] I1_1_t0b,
  input  [31:0] I1_1_t1b,
  input  [31:0] I1_2_t0b,
  input  [31:0] I1_2_t1b,
  input  [31:0] I1_3_t0b,
  input  [31:0] I1_3_t1b,
  input  [31:0] I1_4_t0b,
  input  [31:0] I1_4_t1b,
  input  [31:0] I1_5_t0b,
  input  [31:0] I1_5_t1b,
  input  [31:0] I1_6_t0b,
  input  [31:0] I1_6_t1b,
  input  [31:0] I1_7_t0b,
  input  [31:0] I1_7_t1b,
  output [31:0] O_0_t0b,
  output [31:0] O_0_t1b_t0b,
  output [31:0] O_0_t1b_t1b,
  output [31:0] O_1_t0b,
  output [31:0] O_1_t1b_t0b,
  output [31:0] O_1_t1b_t1b,
  output [31:0] O_2_t0b,
  output [31:0] O_2_t1b_t0b,
  output [31:0] O_2_t1b_t1b,
  output [31:0] O_3_t0b,
  output [31:0] O_3_t1b_t0b,
  output [31:0] O_3_t1b_t1b,
  output [31:0] O_4_t0b,
  output [31:0] O_4_t1b_t0b,
  output [31:0] O_4_t1b_t1b,
  output [31:0] O_5_t0b,
  output [31:0] O_5_t1b_t0b,
  output [31:0] O_5_t1b_t1b,
  output [31:0] O_6_t0b,
  output [31:0] O_6_t1b_t0b,
  output [31:0] O_6_t1b_t1b,
  output [31:0] O_7_t0b,
  output [31:0] O_7_t1b_t0b,
  output [31:0] O_7_t1b_t1b
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_0_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_0_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_1_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_1_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_2_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_2_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_3_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_3_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_4_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_4_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_5_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_5_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_6_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_6_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_7_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_7_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_t1b_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_t1b_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_t1b_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_t1b_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_t1b_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_t1b_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_t1b_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_t1b_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_t1b_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_t1b_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_t1b_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_t1b_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_t1b_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_t1b_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_t1b_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_t1b_t1b; // @[Map2T.scala 8:20]
  Map2S_94 op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0(op_I0_0),
    .I0_1(op_I0_1),
    .I0_2(op_I0_2),
    .I0_3(op_I0_3),
    .I0_4(op_I0_4),
    .I0_5(op_I0_5),
    .I0_6(op_I0_6),
    .I0_7(op_I0_7),
    .I1_0_t0b(op_I1_0_t0b),
    .I1_0_t1b(op_I1_0_t1b),
    .I1_1_t0b(op_I1_1_t0b),
    .I1_1_t1b(op_I1_1_t1b),
    .I1_2_t0b(op_I1_2_t0b),
    .I1_2_t1b(op_I1_2_t1b),
    .I1_3_t0b(op_I1_3_t0b),
    .I1_3_t1b(op_I1_3_t1b),
    .I1_4_t0b(op_I1_4_t0b),
    .I1_4_t1b(op_I1_4_t1b),
    .I1_5_t0b(op_I1_5_t0b),
    .I1_5_t1b(op_I1_5_t1b),
    .I1_6_t0b(op_I1_6_t0b),
    .I1_6_t1b(op_I1_6_t1b),
    .I1_7_t0b(op_I1_7_t0b),
    .I1_7_t1b(op_I1_7_t1b),
    .O_0_t0b(op_O_0_t0b),
    .O_0_t1b_t0b(op_O_0_t1b_t0b),
    .O_0_t1b_t1b(op_O_0_t1b_t1b),
    .O_1_t0b(op_O_1_t0b),
    .O_1_t1b_t0b(op_O_1_t1b_t0b),
    .O_1_t1b_t1b(op_O_1_t1b_t1b),
    .O_2_t0b(op_O_2_t0b),
    .O_2_t1b_t0b(op_O_2_t1b_t0b),
    .O_2_t1b_t1b(op_O_2_t1b_t1b),
    .O_3_t0b(op_O_3_t0b),
    .O_3_t1b_t0b(op_O_3_t1b_t0b),
    .O_3_t1b_t1b(op_O_3_t1b_t1b),
    .O_4_t0b(op_O_4_t0b),
    .O_4_t1b_t0b(op_O_4_t1b_t0b),
    .O_4_t1b_t1b(op_O_4_t1b_t1b),
    .O_5_t0b(op_O_5_t0b),
    .O_5_t1b_t0b(op_O_5_t1b_t0b),
    .O_5_t1b_t1b(op_O_5_t1b_t1b),
    .O_6_t0b(op_O_6_t0b),
    .O_6_t1b_t0b(op_O_6_t1b_t0b),
    .O_6_t1b_t1b(op_O_6_t1b_t1b),
    .O_7_t0b(op_O_7_t0b),
    .O_7_t1b_t0b(op_O_7_t1b_t0b),
    .O_7_t1b_t1b(op_O_7_t1b_t1b)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_t0b = op_O_0_t0b; // @[Map2T.scala 17:7]
  assign O_0_t1b_t0b = op_O_0_t1b_t0b; // @[Map2T.scala 17:7]
  assign O_0_t1b_t1b = op_O_0_t1b_t1b; // @[Map2T.scala 17:7]
  assign O_1_t0b = op_O_1_t0b; // @[Map2T.scala 17:7]
  assign O_1_t1b_t0b = op_O_1_t1b_t0b; // @[Map2T.scala 17:7]
  assign O_1_t1b_t1b = op_O_1_t1b_t1b; // @[Map2T.scala 17:7]
  assign O_2_t0b = op_O_2_t0b; // @[Map2T.scala 17:7]
  assign O_2_t1b_t0b = op_O_2_t1b_t0b; // @[Map2T.scala 17:7]
  assign O_2_t1b_t1b = op_O_2_t1b_t1b; // @[Map2T.scala 17:7]
  assign O_3_t0b = op_O_3_t0b; // @[Map2T.scala 17:7]
  assign O_3_t1b_t0b = op_O_3_t1b_t0b; // @[Map2T.scala 17:7]
  assign O_3_t1b_t1b = op_O_3_t1b_t1b; // @[Map2T.scala 17:7]
  assign O_4_t0b = op_O_4_t0b; // @[Map2T.scala 17:7]
  assign O_4_t1b_t0b = op_O_4_t1b_t0b; // @[Map2T.scala 17:7]
  assign O_4_t1b_t1b = op_O_4_t1b_t1b; // @[Map2T.scala 17:7]
  assign O_5_t0b = op_O_5_t0b; // @[Map2T.scala 17:7]
  assign O_5_t1b_t0b = op_O_5_t1b_t0b; // @[Map2T.scala 17:7]
  assign O_5_t1b_t1b = op_O_5_t1b_t1b; // @[Map2T.scala 17:7]
  assign O_6_t0b = op_O_6_t0b; // @[Map2T.scala 17:7]
  assign O_6_t1b_t0b = op_O_6_t1b_t0b; // @[Map2T.scala 17:7]
  assign O_6_t1b_t1b = op_O_6_t1b_t1b; // @[Map2T.scala 17:7]
  assign O_7_t0b = op_O_7_t0b; // @[Map2T.scala 17:7]
  assign O_7_t1b_t0b = op_O_7_t1b_t0b; // @[Map2T.scala 17:7]
  assign O_7_t1b_t1b = op_O_7_t1b_t1b; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0 = I0_0; // @[Map2T.scala 15:11]
  assign op_I0_1 = I0_1; // @[Map2T.scala 15:11]
  assign op_I0_2 = I0_2; // @[Map2T.scala 15:11]
  assign op_I0_3 = I0_3; // @[Map2T.scala 15:11]
  assign op_I0_4 = I0_4; // @[Map2T.scala 15:11]
  assign op_I0_5 = I0_5; // @[Map2T.scala 15:11]
  assign op_I0_6 = I0_6; // @[Map2T.scala 15:11]
  assign op_I0_7 = I0_7; // @[Map2T.scala 15:11]
  assign op_I1_0_t0b = I1_0_t0b; // @[Map2T.scala 16:11]
  assign op_I1_0_t1b = I1_0_t1b; // @[Map2T.scala 16:11]
  assign op_I1_1_t0b = I1_1_t0b; // @[Map2T.scala 16:11]
  assign op_I1_1_t1b = I1_1_t1b; // @[Map2T.scala 16:11]
  assign op_I1_2_t0b = I1_2_t0b; // @[Map2T.scala 16:11]
  assign op_I1_2_t1b = I1_2_t1b; // @[Map2T.scala 16:11]
  assign op_I1_3_t0b = I1_3_t0b; // @[Map2T.scala 16:11]
  assign op_I1_3_t1b = I1_3_t1b; // @[Map2T.scala 16:11]
  assign op_I1_4_t0b = I1_4_t0b; // @[Map2T.scala 16:11]
  assign op_I1_4_t1b = I1_4_t1b; // @[Map2T.scala 16:11]
  assign op_I1_5_t0b = I1_5_t0b; // @[Map2T.scala 16:11]
  assign op_I1_5_t1b = I1_5_t1b; // @[Map2T.scala 16:11]
  assign op_I1_6_t0b = I1_6_t0b; // @[Map2T.scala 16:11]
  assign op_I1_6_t1b = I1_6_t1b; // @[Map2T.scala 16:11]
  assign op_I1_7_t0b = I1_7_t0b; // @[Map2T.scala 16:11]
  assign op_I1_7_t1b = I1_7_t1b; // @[Map2T.scala 16:11]
endmodule
module FIFO_15(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_t0b,
  input  [31:0] I_0_t1b_t0b,
  input  [31:0] I_0_t1b_t1b,
  input  [31:0] I_1_t0b,
  input  [31:0] I_1_t1b_t0b,
  input  [31:0] I_1_t1b_t1b,
  input  [31:0] I_2_t0b,
  input  [31:0] I_2_t1b_t0b,
  input  [31:0] I_2_t1b_t1b,
  input  [31:0] I_3_t0b,
  input  [31:0] I_3_t1b_t0b,
  input  [31:0] I_3_t1b_t1b,
  input  [31:0] I_4_t0b,
  input  [31:0] I_4_t1b_t0b,
  input  [31:0] I_4_t1b_t1b,
  input  [31:0] I_5_t0b,
  input  [31:0] I_5_t1b_t0b,
  input  [31:0] I_5_t1b_t1b,
  input  [31:0] I_6_t0b,
  input  [31:0] I_6_t1b_t0b,
  input  [31:0] I_6_t1b_t1b,
  input  [31:0] I_7_t0b,
  input  [31:0] I_7_t1b_t0b,
  input  [31:0] I_7_t1b_t1b,
  output [31:0] O_0_t0b,
  output [31:0] O_0_t1b_t0b,
  output [31:0] O_0_t1b_t1b,
  output [31:0] O_1_t0b,
  output [31:0] O_1_t1b_t0b,
  output [31:0] O_1_t1b_t1b,
  output [31:0] O_2_t0b,
  output [31:0] O_2_t1b_t0b,
  output [31:0] O_2_t1b_t1b,
  output [31:0] O_3_t0b,
  output [31:0] O_3_t1b_t0b,
  output [31:0] O_3_t1b_t1b,
  output [31:0] O_4_t0b,
  output [31:0] O_4_t1b_t0b,
  output [31:0] O_4_t1b_t1b,
  output [31:0] O_5_t0b,
  output [31:0] O_5_t1b_t0b,
  output [31:0] O_5_t1b_t1b,
  output [31:0] O_6_t0b,
  output [31:0] O_6_t1b_t0b,
  output [31:0] O_6_t1b_t1b,
  output [31:0] O_7_t0b,
  output [31:0] O_7_t1b_t0b,
  output [31:0] O_7_t1b_t1b
);
  reg [31:0] _T__0_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_0;
  reg [31:0] _T__0_t1b_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_1;
  reg [31:0] _T__0_t1b_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_2;
  reg [31:0] _T__1_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_3;
  reg [31:0] _T__1_t1b_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_4;
  reg [31:0] _T__1_t1b_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_5;
  reg [31:0] _T__2_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_6;
  reg [31:0] _T__2_t1b_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_7;
  reg [31:0] _T__2_t1b_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_8;
  reg [31:0] _T__3_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_9;
  reg [31:0] _T__3_t1b_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_10;
  reg [31:0] _T__3_t1b_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_11;
  reg [31:0] _T__4_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_12;
  reg [31:0] _T__4_t1b_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_13;
  reg [31:0] _T__4_t1b_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_14;
  reg [31:0] _T__5_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_15;
  reg [31:0] _T__5_t1b_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_16;
  reg [31:0] _T__5_t1b_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_17;
  reg [31:0] _T__6_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_18;
  reg [31:0] _T__6_t1b_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_19;
  reg [31:0] _T__6_t1b_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_20;
  reg [31:0] _T__7_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_21;
  reg [31:0] _T__7_t1b_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_22;
  reg [31:0] _T__7_t1b_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_23;
  reg  _T_1; // @[FIFO.scala 15:27]
  reg [31:0] _RAND_24;
  assign valid_down = _T_1; // @[FIFO.scala 16:16]
  assign O_0_t0b = _T__0_t0b; // @[FIFO.scala 14:7]
  assign O_0_t1b_t0b = _T__0_t1b_t0b; // @[FIFO.scala 14:7]
  assign O_0_t1b_t1b = _T__0_t1b_t1b; // @[FIFO.scala 14:7]
  assign O_1_t0b = _T__1_t0b; // @[FIFO.scala 14:7]
  assign O_1_t1b_t0b = _T__1_t1b_t0b; // @[FIFO.scala 14:7]
  assign O_1_t1b_t1b = _T__1_t1b_t1b; // @[FIFO.scala 14:7]
  assign O_2_t0b = _T__2_t0b; // @[FIFO.scala 14:7]
  assign O_2_t1b_t0b = _T__2_t1b_t0b; // @[FIFO.scala 14:7]
  assign O_2_t1b_t1b = _T__2_t1b_t1b; // @[FIFO.scala 14:7]
  assign O_3_t0b = _T__3_t0b; // @[FIFO.scala 14:7]
  assign O_3_t1b_t0b = _T__3_t1b_t0b; // @[FIFO.scala 14:7]
  assign O_3_t1b_t1b = _T__3_t1b_t1b; // @[FIFO.scala 14:7]
  assign O_4_t0b = _T__4_t0b; // @[FIFO.scala 14:7]
  assign O_4_t1b_t0b = _T__4_t1b_t0b; // @[FIFO.scala 14:7]
  assign O_4_t1b_t1b = _T__4_t1b_t1b; // @[FIFO.scala 14:7]
  assign O_5_t0b = _T__5_t0b; // @[FIFO.scala 14:7]
  assign O_5_t1b_t0b = _T__5_t1b_t0b; // @[FIFO.scala 14:7]
  assign O_5_t1b_t1b = _T__5_t1b_t1b; // @[FIFO.scala 14:7]
  assign O_6_t0b = _T__6_t0b; // @[FIFO.scala 14:7]
  assign O_6_t1b_t0b = _T__6_t1b_t0b; // @[FIFO.scala 14:7]
  assign O_6_t1b_t1b = _T__6_t1b_t1b; // @[FIFO.scala 14:7]
  assign O_7_t0b = _T__7_t0b; // @[FIFO.scala 14:7]
  assign O_7_t1b_t0b = _T__7_t1b_t0b; // @[FIFO.scala 14:7]
  assign O_7_t1b_t1b = _T__7_t1b_t1b; // @[FIFO.scala 14:7]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T__0_t0b = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T__0_t1b_t0b = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T__0_t1b_t1b = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T__1_t0b = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T__1_t1b_t0b = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T__1_t1b_t1b = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T__2_t0b = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T__2_t1b_t0b = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T__2_t1b_t1b = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T__3_t0b = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T__3_t1b_t0b = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T__3_t1b_t1b = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T__4_t0b = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T__4_t1b_t0b = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T__4_t1b_t1b = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T__5_t0b = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T__5_t1b_t0b = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T__5_t1b_t1b = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T__6_t0b = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T__6_t1b_t0b = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T__6_t1b_t1b = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T__7_t0b = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T__7_t1b_t0b = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T__7_t1b_t1b = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_1 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T__0_t0b <= I_0_t0b;
    _T__0_t1b_t0b <= I_0_t1b_t0b;
    _T__0_t1b_t1b <= I_0_t1b_t1b;
    _T__1_t0b <= I_1_t0b;
    _T__1_t1b_t0b <= I_1_t1b_t0b;
    _T__1_t1b_t1b <= I_1_t1b_t1b;
    _T__2_t0b <= I_2_t0b;
    _T__2_t1b_t0b <= I_2_t1b_t0b;
    _T__2_t1b_t1b <= I_2_t1b_t1b;
    _T__3_t0b <= I_3_t0b;
    _T__3_t1b_t0b <= I_3_t1b_t0b;
    _T__3_t1b_t1b <= I_3_t1b_t1b;
    _T__4_t0b <= I_4_t0b;
    _T__4_t1b_t0b <= I_4_t1b_t0b;
    _T__4_t1b_t1b <= I_4_t1b_t1b;
    _T__5_t0b <= I_5_t0b;
    _T__5_t1b_t0b <= I_5_t1b_t0b;
    _T__5_t1b_t1b <= I_5_t1b_t1b;
    _T__6_t0b <= I_6_t0b;
    _T__6_t1b_t0b <= I_6_t1b_t0b;
    _T__6_t1b_t1b <= I_6_t1b_t1b;
    _T__7_t0b <= I_7_t0b;
    _T__7_t1b_t0b <= I_7_t1b_t0b;
    _T__7_t1b_t1b <= I_7_t1b_t1b;
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      _T_1 <= valid_up;
    end
  end
endmodule
module Top(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0,
  input  [31:0] I_1,
  input  [31:0] I_2,
  input  [31:0] I_3,
  input  [31:0] I_4,
  input  [31:0] I_5,
  input  [31:0] I_6,
  input  [31:0] I_7,
  output [31:0] O_0_t0b,
  output [31:0] O_0_t1b_t0b,
  output [31:0] O_0_t1b_t1b,
  output [31:0] O_1_t0b,
  output [31:0] O_1_t1b_t0b,
  output [31:0] O_1_t1b_t1b,
  output [31:0] O_2_t0b,
  output [31:0] O_2_t1b_t0b,
  output [31:0] O_2_t1b_t1b,
  output [31:0] O_3_t0b,
  output [31:0] O_3_t1b_t0b,
  output [31:0] O_3_t1b_t1b,
  output [31:0] O_4_t0b,
  output [31:0] O_4_t1b_t0b,
  output [31:0] O_4_t1b_t1b,
  output [31:0] O_5_t0b,
  output [31:0] O_5_t1b_t0b,
  output [31:0] O_5_t1b_t1b,
  output [31:0] O_6_t0b,
  output [31:0] O_6_t1b_t0b,
  output [31:0] O_6_t1b_t1b,
  output [31:0] O_7_t0b,
  output [31:0] O_7_t1b_t0b,
  output [31:0] O_7_t1b_t1b
);
  wire  n1_clock; // @[Top.scala 695:20]
  wire  n1_reset; // @[Top.scala 695:20]
  wire  n1_valid_up; // @[Top.scala 695:20]
  wire  n1_valid_down; // @[Top.scala 695:20]
  wire [31:0] n1_I_0; // @[Top.scala 695:20]
  wire [31:0] n1_I_1; // @[Top.scala 695:20]
  wire [31:0] n1_I_2; // @[Top.scala 695:20]
  wire [31:0] n1_I_3; // @[Top.scala 695:20]
  wire [31:0] n1_I_4; // @[Top.scala 695:20]
  wire [31:0] n1_I_5; // @[Top.scala 695:20]
  wire [31:0] n1_I_6; // @[Top.scala 695:20]
  wire [31:0] n1_I_7; // @[Top.scala 695:20]
  wire [31:0] n1_O_0; // @[Top.scala 695:20]
  wire [31:0] n1_O_1; // @[Top.scala 695:20]
  wire [31:0] n1_O_2; // @[Top.scala 695:20]
  wire [31:0] n1_O_3; // @[Top.scala 695:20]
  wire [31:0] n1_O_4; // @[Top.scala 695:20]
  wire [31:0] n1_O_5; // @[Top.scala 695:20]
  wire [31:0] n1_O_6; // @[Top.scala 695:20]
  wire [31:0] n1_O_7; // @[Top.scala 695:20]
  wire  n2_clock; // @[Top.scala 698:20]
  wire  n2_reset; // @[Top.scala 698:20]
  wire  n2_valid_up; // @[Top.scala 698:20]
  wire  n2_valid_down; // @[Top.scala 698:20]
  wire [31:0] n2_I_0; // @[Top.scala 698:20]
  wire [31:0] n2_I_1; // @[Top.scala 698:20]
  wire [31:0] n2_I_2; // @[Top.scala 698:20]
  wire [31:0] n2_I_3; // @[Top.scala 698:20]
  wire [31:0] n2_I_4; // @[Top.scala 698:20]
  wire [31:0] n2_I_5; // @[Top.scala 698:20]
  wire [31:0] n2_I_6; // @[Top.scala 698:20]
  wire [31:0] n2_I_7; // @[Top.scala 698:20]
  wire [31:0] n2_O_0; // @[Top.scala 698:20]
  wire [31:0] n2_O_1; // @[Top.scala 698:20]
  wire [31:0] n2_O_2; // @[Top.scala 698:20]
  wire [31:0] n2_O_3; // @[Top.scala 698:20]
  wire [31:0] n2_O_4; // @[Top.scala 698:20]
  wire [31:0] n2_O_5; // @[Top.scala 698:20]
  wire [31:0] n2_O_6; // @[Top.scala 698:20]
  wire [31:0] n2_O_7; // @[Top.scala 698:20]
  wire  n3_clock; // @[Top.scala 701:20]
  wire  n3_reset; // @[Top.scala 701:20]
  wire  n3_valid_up; // @[Top.scala 701:20]
  wire  n3_valid_down; // @[Top.scala 701:20]
  wire [31:0] n3_I_0; // @[Top.scala 701:20]
  wire [31:0] n3_I_1; // @[Top.scala 701:20]
  wire [31:0] n3_I_2; // @[Top.scala 701:20]
  wire [31:0] n3_I_3; // @[Top.scala 701:20]
  wire [31:0] n3_I_4; // @[Top.scala 701:20]
  wire [31:0] n3_I_5; // @[Top.scala 701:20]
  wire [31:0] n3_I_6; // @[Top.scala 701:20]
  wire [31:0] n3_I_7; // @[Top.scala 701:20]
  wire [31:0] n3_O_0; // @[Top.scala 701:20]
  wire [31:0] n3_O_1; // @[Top.scala 701:20]
  wire [31:0] n3_O_2; // @[Top.scala 701:20]
  wire [31:0] n3_O_3; // @[Top.scala 701:20]
  wire [31:0] n3_O_4; // @[Top.scala 701:20]
  wire [31:0] n3_O_5; // @[Top.scala 701:20]
  wire [31:0] n3_O_6; // @[Top.scala 701:20]
  wire [31:0] n3_O_7; // @[Top.scala 701:20]
  wire  n4_clock; // @[Top.scala 704:20]
  wire  n4_valid_up; // @[Top.scala 704:20]
  wire  n4_valid_down; // @[Top.scala 704:20]
  wire [31:0] n4_I_0; // @[Top.scala 704:20]
  wire [31:0] n4_I_1; // @[Top.scala 704:20]
  wire [31:0] n4_I_2; // @[Top.scala 704:20]
  wire [31:0] n4_I_3; // @[Top.scala 704:20]
  wire [31:0] n4_I_4; // @[Top.scala 704:20]
  wire [31:0] n4_I_5; // @[Top.scala 704:20]
  wire [31:0] n4_I_6; // @[Top.scala 704:20]
  wire [31:0] n4_I_7; // @[Top.scala 704:20]
  wire [31:0] n4_O_0; // @[Top.scala 704:20]
  wire [31:0] n4_O_1; // @[Top.scala 704:20]
  wire [31:0] n4_O_2; // @[Top.scala 704:20]
  wire [31:0] n4_O_3; // @[Top.scala 704:20]
  wire [31:0] n4_O_4; // @[Top.scala 704:20]
  wire [31:0] n4_O_5; // @[Top.scala 704:20]
  wire [31:0] n4_O_6; // @[Top.scala 704:20]
  wire [31:0] n4_O_7; // @[Top.scala 704:20]
  wire  n5_clock; // @[Top.scala 707:20]
  wire  n5_valid_up; // @[Top.scala 707:20]
  wire  n5_valid_down; // @[Top.scala 707:20]
  wire [31:0] n5_I_0; // @[Top.scala 707:20]
  wire [31:0] n5_I_1; // @[Top.scala 707:20]
  wire [31:0] n5_I_2; // @[Top.scala 707:20]
  wire [31:0] n5_I_3; // @[Top.scala 707:20]
  wire [31:0] n5_I_4; // @[Top.scala 707:20]
  wire [31:0] n5_I_5; // @[Top.scala 707:20]
  wire [31:0] n5_I_6; // @[Top.scala 707:20]
  wire [31:0] n5_I_7; // @[Top.scala 707:20]
  wire [31:0] n5_O_0; // @[Top.scala 707:20]
  wire [31:0] n5_O_1; // @[Top.scala 707:20]
  wire [31:0] n5_O_2; // @[Top.scala 707:20]
  wire [31:0] n5_O_3; // @[Top.scala 707:20]
  wire [31:0] n5_O_4; // @[Top.scala 707:20]
  wire [31:0] n5_O_5; // @[Top.scala 707:20]
  wire [31:0] n5_O_6; // @[Top.scala 707:20]
  wire [31:0] n5_O_7; // @[Top.scala 707:20]
  wire  n6_valid_up; // @[Top.scala 710:20]
  wire  n6_valid_down; // @[Top.scala 710:20]
  wire [31:0] n6_I0_0; // @[Top.scala 710:20]
  wire [31:0] n6_I0_1; // @[Top.scala 710:20]
  wire [31:0] n6_I0_2; // @[Top.scala 710:20]
  wire [31:0] n6_I0_3; // @[Top.scala 710:20]
  wire [31:0] n6_I0_4; // @[Top.scala 710:20]
  wire [31:0] n6_I0_5; // @[Top.scala 710:20]
  wire [31:0] n6_I0_6; // @[Top.scala 710:20]
  wire [31:0] n6_I0_7; // @[Top.scala 710:20]
  wire [31:0] n6_I1_0; // @[Top.scala 710:20]
  wire [31:0] n6_I1_1; // @[Top.scala 710:20]
  wire [31:0] n6_I1_2; // @[Top.scala 710:20]
  wire [31:0] n6_I1_3; // @[Top.scala 710:20]
  wire [31:0] n6_I1_4; // @[Top.scala 710:20]
  wire [31:0] n6_I1_5; // @[Top.scala 710:20]
  wire [31:0] n6_I1_6; // @[Top.scala 710:20]
  wire [31:0] n6_I1_7; // @[Top.scala 710:20]
  wire [31:0] n6_O_0_0; // @[Top.scala 710:20]
  wire [31:0] n6_O_0_1; // @[Top.scala 710:20]
  wire [31:0] n6_O_1_0; // @[Top.scala 710:20]
  wire [31:0] n6_O_1_1; // @[Top.scala 710:20]
  wire [31:0] n6_O_2_0; // @[Top.scala 710:20]
  wire [31:0] n6_O_2_1; // @[Top.scala 710:20]
  wire [31:0] n6_O_3_0; // @[Top.scala 710:20]
  wire [31:0] n6_O_3_1; // @[Top.scala 710:20]
  wire [31:0] n6_O_4_0; // @[Top.scala 710:20]
  wire [31:0] n6_O_4_1; // @[Top.scala 710:20]
  wire [31:0] n6_O_5_0; // @[Top.scala 710:20]
  wire [31:0] n6_O_5_1; // @[Top.scala 710:20]
  wire [31:0] n6_O_6_0; // @[Top.scala 710:20]
  wire [31:0] n6_O_6_1; // @[Top.scala 710:20]
  wire [31:0] n6_O_7_0; // @[Top.scala 710:20]
  wire [31:0] n6_O_7_1; // @[Top.scala 710:20]
  wire  n13_valid_up; // @[Top.scala 714:21]
  wire  n13_valid_down; // @[Top.scala 714:21]
  wire [31:0] n13_I0_0_0; // @[Top.scala 714:21]
  wire [31:0] n13_I0_0_1; // @[Top.scala 714:21]
  wire [31:0] n13_I0_1_0; // @[Top.scala 714:21]
  wire [31:0] n13_I0_1_1; // @[Top.scala 714:21]
  wire [31:0] n13_I0_2_0; // @[Top.scala 714:21]
  wire [31:0] n13_I0_2_1; // @[Top.scala 714:21]
  wire [31:0] n13_I0_3_0; // @[Top.scala 714:21]
  wire [31:0] n13_I0_3_1; // @[Top.scala 714:21]
  wire [31:0] n13_I0_4_0; // @[Top.scala 714:21]
  wire [31:0] n13_I0_4_1; // @[Top.scala 714:21]
  wire [31:0] n13_I0_5_0; // @[Top.scala 714:21]
  wire [31:0] n13_I0_5_1; // @[Top.scala 714:21]
  wire [31:0] n13_I0_6_0; // @[Top.scala 714:21]
  wire [31:0] n13_I0_6_1; // @[Top.scala 714:21]
  wire [31:0] n13_I0_7_0; // @[Top.scala 714:21]
  wire [31:0] n13_I0_7_1; // @[Top.scala 714:21]
  wire [31:0] n13_I1_0; // @[Top.scala 714:21]
  wire [31:0] n13_I1_1; // @[Top.scala 714:21]
  wire [31:0] n13_I1_2; // @[Top.scala 714:21]
  wire [31:0] n13_I1_3; // @[Top.scala 714:21]
  wire [31:0] n13_I1_4; // @[Top.scala 714:21]
  wire [31:0] n13_I1_5; // @[Top.scala 714:21]
  wire [31:0] n13_I1_6; // @[Top.scala 714:21]
  wire [31:0] n13_I1_7; // @[Top.scala 714:21]
  wire [31:0] n13_O_0_0; // @[Top.scala 714:21]
  wire [31:0] n13_O_0_1; // @[Top.scala 714:21]
  wire [31:0] n13_O_0_2; // @[Top.scala 714:21]
  wire [31:0] n13_O_1_0; // @[Top.scala 714:21]
  wire [31:0] n13_O_1_1; // @[Top.scala 714:21]
  wire [31:0] n13_O_1_2; // @[Top.scala 714:21]
  wire [31:0] n13_O_2_0; // @[Top.scala 714:21]
  wire [31:0] n13_O_2_1; // @[Top.scala 714:21]
  wire [31:0] n13_O_2_2; // @[Top.scala 714:21]
  wire [31:0] n13_O_3_0; // @[Top.scala 714:21]
  wire [31:0] n13_O_3_1; // @[Top.scala 714:21]
  wire [31:0] n13_O_3_2; // @[Top.scala 714:21]
  wire [31:0] n13_O_4_0; // @[Top.scala 714:21]
  wire [31:0] n13_O_4_1; // @[Top.scala 714:21]
  wire [31:0] n13_O_4_2; // @[Top.scala 714:21]
  wire [31:0] n13_O_5_0; // @[Top.scala 714:21]
  wire [31:0] n13_O_5_1; // @[Top.scala 714:21]
  wire [31:0] n13_O_5_2; // @[Top.scala 714:21]
  wire [31:0] n13_O_6_0; // @[Top.scala 714:21]
  wire [31:0] n13_O_6_1; // @[Top.scala 714:21]
  wire [31:0] n13_O_6_2; // @[Top.scala 714:21]
  wire [31:0] n13_O_7_0; // @[Top.scala 714:21]
  wire [31:0] n13_O_7_1; // @[Top.scala 714:21]
  wire [31:0] n13_O_7_2; // @[Top.scala 714:21]
  wire  n22_valid_up; // @[Top.scala 718:21]
  wire  n22_valid_down; // @[Top.scala 718:21]
  wire [31:0] n22_I_0_0; // @[Top.scala 718:21]
  wire [31:0] n22_I_0_1; // @[Top.scala 718:21]
  wire [31:0] n22_I_0_2; // @[Top.scala 718:21]
  wire [31:0] n22_I_1_0; // @[Top.scala 718:21]
  wire [31:0] n22_I_1_1; // @[Top.scala 718:21]
  wire [31:0] n22_I_1_2; // @[Top.scala 718:21]
  wire [31:0] n22_I_2_0; // @[Top.scala 718:21]
  wire [31:0] n22_I_2_1; // @[Top.scala 718:21]
  wire [31:0] n22_I_2_2; // @[Top.scala 718:21]
  wire [31:0] n22_I_3_0; // @[Top.scala 718:21]
  wire [31:0] n22_I_3_1; // @[Top.scala 718:21]
  wire [31:0] n22_I_3_2; // @[Top.scala 718:21]
  wire [31:0] n22_I_4_0; // @[Top.scala 718:21]
  wire [31:0] n22_I_4_1; // @[Top.scala 718:21]
  wire [31:0] n22_I_4_2; // @[Top.scala 718:21]
  wire [31:0] n22_I_5_0; // @[Top.scala 718:21]
  wire [31:0] n22_I_5_1; // @[Top.scala 718:21]
  wire [31:0] n22_I_5_2; // @[Top.scala 718:21]
  wire [31:0] n22_I_6_0; // @[Top.scala 718:21]
  wire [31:0] n22_I_6_1; // @[Top.scala 718:21]
  wire [31:0] n22_I_6_2; // @[Top.scala 718:21]
  wire [31:0] n22_I_7_0; // @[Top.scala 718:21]
  wire [31:0] n22_I_7_1; // @[Top.scala 718:21]
  wire [31:0] n22_I_7_2; // @[Top.scala 718:21]
  wire [31:0] n22_O_0_0_0; // @[Top.scala 718:21]
  wire [31:0] n22_O_0_0_1; // @[Top.scala 718:21]
  wire [31:0] n22_O_0_0_2; // @[Top.scala 718:21]
  wire [31:0] n22_O_1_0_0; // @[Top.scala 718:21]
  wire [31:0] n22_O_1_0_1; // @[Top.scala 718:21]
  wire [31:0] n22_O_1_0_2; // @[Top.scala 718:21]
  wire [31:0] n22_O_2_0_0; // @[Top.scala 718:21]
  wire [31:0] n22_O_2_0_1; // @[Top.scala 718:21]
  wire [31:0] n22_O_2_0_2; // @[Top.scala 718:21]
  wire [31:0] n22_O_3_0_0; // @[Top.scala 718:21]
  wire [31:0] n22_O_3_0_1; // @[Top.scala 718:21]
  wire [31:0] n22_O_3_0_2; // @[Top.scala 718:21]
  wire [31:0] n22_O_4_0_0; // @[Top.scala 718:21]
  wire [31:0] n22_O_4_0_1; // @[Top.scala 718:21]
  wire [31:0] n22_O_4_0_2; // @[Top.scala 718:21]
  wire [31:0] n22_O_5_0_0; // @[Top.scala 718:21]
  wire [31:0] n22_O_5_0_1; // @[Top.scala 718:21]
  wire [31:0] n22_O_5_0_2; // @[Top.scala 718:21]
  wire [31:0] n22_O_6_0_0; // @[Top.scala 718:21]
  wire [31:0] n22_O_6_0_1; // @[Top.scala 718:21]
  wire [31:0] n22_O_6_0_2; // @[Top.scala 718:21]
  wire [31:0] n22_O_7_0_0; // @[Top.scala 718:21]
  wire [31:0] n22_O_7_0_1; // @[Top.scala 718:21]
  wire [31:0] n22_O_7_0_2; // @[Top.scala 718:21]
  wire  n29_valid_up; // @[Top.scala 721:21]
  wire  n29_valid_down; // @[Top.scala 721:21]
  wire [31:0] n29_I_0_0_0; // @[Top.scala 721:21]
  wire [31:0] n29_I_0_0_1; // @[Top.scala 721:21]
  wire [31:0] n29_I_0_0_2; // @[Top.scala 721:21]
  wire [31:0] n29_I_1_0_0; // @[Top.scala 721:21]
  wire [31:0] n29_I_1_0_1; // @[Top.scala 721:21]
  wire [31:0] n29_I_1_0_2; // @[Top.scala 721:21]
  wire [31:0] n29_I_2_0_0; // @[Top.scala 721:21]
  wire [31:0] n29_I_2_0_1; // @[Top.scala 721:21]
  wire [31:0] n29_I_2_0_2; // @[Top.scala 721:21]
  wire [31:0] n29_I_3_0_0; // @[Top.scala 721:21]
  wire [31:0] n29_I_3_0_1; // @[Top.scala 721:21]
  wire [31:0] n29_I_3_0_2; // @[Top.scala 721:21]
  wire [31:0] n29_I_4_0_0; // @[Top.scala 721:21]
  wire [31:0] n29_I_4_0_1; // @[Top.scala 721:21]
  wire [31:0] n29_I_4_0_2; // @[Top.scala 721:21]
  wire [31:0] n29_I_5_0_0; // @[Top.scala 721:21]
  wire [31:0] n29_I_5_0_1; // @[Top.scala 721:21]
  wire [31:0] n29_I_5_0_2; // @[Top.scala 721:21]
  wire [31:0] n29_I_6_0_0; // @[Top.scala 721:21]
  wire [31:0] n29_I_6_0_1; // @[Top.scala 721:21]
  wire [31:0] n29_I_6_0_2; // @[Top.scala 721:21]
  wire [31:0] n29_I_7_0_0; // @[Top.scala 721:21]
  wire [31:0] n29_I_7_0_1; // @[Top.scala 721:21]
  wire [31:0] n29_I_7_0_2; // @[Top.scala 721:21]
  wire [31:0] n29_O_0_0; // @[Top.scala 721:21]
  wire [31:0] n29_O_0_1; // @[Top.scala 721:21]
  wire [31:0] n29_O_0_2; // @[Top.scala 721:21]
  wire [31:0] n29_O_1_0; // @[Top.scala 721:21]
  wire [31:0] n29_O_1_1; // @[Top.scala 721:21]
  wire [31:0] n29_O_1_2; // @[Top.scala 721:21]
  wire [31:0] n29_O_2_0; // @[Top.scala 721:21]
  wire [31:0] n29_O_2_1; // @[Top.scala 721:21]
  wire [31:0] n29_O_2_2; // @[Top.scala 721:21]
  wire [31:0] n29_O_3_0; // @[Top.scala 721:21]
  wire [31:0] n29_O_3_1; // @[Top.scala 721:21]
  wire [31:0] n29_O_3_2; // @[Top.scala 721:21]
  wire [31:0] n29_O_4_0; // @[Top.scala 721:21]
  wire [31:0] n29_O_4_1; // @[Top.scala 721:21]
  wire [31:0] n29_O_4_2; // @[Top.scala 721:21]
  wire [31:0] n29_O_5_0; // @[Top.scala 721:21]
  wire [31:0] n29_O_5_1; // @[Top.scala 721:21]
  wire [31:0] n29_O_5_2; // @[Top.scala 721:21]
  wire [31:0] n29_O_6_0; // @[Top.scala 721:21]
  wire [31:0] n29_O_6_1; // @[Top.scala 721:21]
  wire [31:0] n29_O_6_2; // @[Top.scala 721:21]
  wire [31:0] n29_O_7_0; // @[Top.scala 721:21]
  wire [31:0] n29_O_7_1; // @[Top.scala 721:21]
  wire [31:0] n29_O_7_2; // @[Top.scala 721:21]
  wire  n30_clock; // @[Top.scala 724:21]
  wire  n30_valid_up; // @[Top.scala 724:21]
  wire  n30_valid_down; // @[Top.scala 724:21]
  wire [31:0] n30_I_0; // @[Top.scala 724:21]
  wire [31:0] n30_I_1; // @[Top.scala 724:21]
  wire [31:0] n30_I_2; // @[Top.scala 724:21]
  wire [31:0] n30_I_3; // @[Top.scala 724:21]
  wire [31:0] n30_I_4; // @[Top.scala 724:21]
  wire [31:0] n30_I_5; // @[Top.scala 724:21]
  wire [31:0] n30_I_6; // @[Top.scala 724:21]
  wire [31:0] n30_I_7; // @[Top.scala 724:21]
  wire [31:0] n30_O_0; // @[Top.scala 724:21]
  wire [31:0] n30_O_1; // @[Top.scala 724:21]
  wire [31:0] n30_O_2; // @[Top.scala 724:21]
  wire [31:0] n30_O_3; // @[Top.scala 724:21]
  wire [31:0] n30_O_4; // @[Top.scala 724:21]
  wire [31:0] n30_O_5; // @[Top.scala 724:21]
  wire [31:0] n30_O_6; // @[Top.scala 724:21]
  wire [31:0] n30_O_7; // @[Top.scala 724:21]
  wire  n31_clock; // @[Top.scala 727:21]
  wire  n31_valid_up; // @[Top.scala 727:21]
  wire  n31_valid_down; // @[Top.scala 727:21]
  wire [31:0] n31_I_0; // @[Top.scala 727:21]
  wire [31:0] n31_I_1; // @[Top.scala 727:21]
  wire [31:0] n31_I_2; // @[Top.scala 727:21]
  wire [31:0] n31_I_3; // @[Top.scala 727:21]
  wire [31:0] n31_I_4; // @[Top.scala 727:21]
  wire [31:0] n31_I_5; // @[Top.scala 727:21]
  wire [31:0] n31_I_6; // @[Top.scala 727:21]
  wire [31:0] n31_I_7; // @[Top.scala 727:21]
  wire [31:0] n31_O_0; // @[Top.scala 727:21]
  wire [31:0] n31_O_1; // @[Top.scala 727:21]
  wire [31:0] n31_O_2; // @[Top.scala 727:21]
  wire [31:0] n31_O_3; // @[Top.scala 727:21]
  wire [31:0] n31_O_4; // @[Top.scala 727:21]
  wire [31:0] n31_O_5; // @[Top.scala 727:21]
  wire [31:0] n31_O_6; // @[Top.scala 727:21]
  wire [31:0] n31_O_7; // @[Top.scala 727:21]
  wire  n32_valid_up; // @[Top.scala 730:21]
  wire  n32_valid_down; // @[Top.scala 730:21]
  wire [31:0] n32_I0_0; // @[Top.scala 730:21]
  wire [31:0] n32_I0_1; // @[Top.scala 730:21]
  wire [31:0] n32_I0_2; // @[Top.scala 730:21]
  wire [31:0] n32_I0_3; // @[Top.scala 730:21]
  wire [31:0] n32_I0_4; // @[Top.scala 730:21]
  wire [31:0] n32_I0_5; // @[Top.scala 730:21]
  wire [31:0] n32_I0_6; // @[Top.scala 730:21]
  wire [31:0] n32_I0_7; // @[Top.scala 730:21]
  wire [31:0] n32_I1_0; // @[Top.scala 730:21]
  wire [31:0] n32_I1_1; // @[Top.scala 730:21]
  wire [31:0] n32_I1_2; // @[Top.scala 730:21]
  wire [31:0] n32_I1_3; // @[Top.scala 730:21]
  wire [31:0] n32_I1_4; // @[Top.scala 730:21]
  wire [31:0] n32_I1_5; // @[Top.scala 730:21]
  wire [31:0] n32_I1_6; // @[Top.scala 730:21]
  wire [31:0] n32_I1_7; // @[Top.scala 730:21]
  wire [31:0] n32_O_0_0; // @[Top.scala 730:21]
  wire [31:0] n32_O_0_1; // @[Top.scala 730:21]
  wire [31:0] n32_O_1_0; // @[Top.scala 730:21]
  wire [31:0] n32_O_1_1; // @[Top.scala 730:21]
  wire [31:0] n32_O_2_0; // @[Top.scala 730:21]
  wire [31:0] n32_O_2_1; // @[Top.scala 730:21]
  wire [31:0] n32_O_3_0; // @[Top.scala 730:21]
  wire [31:0] n32_O_3_1; // @[Top.scala 730:21]
  wire [31:0] n32_O_4_0; // @[Top.scala 730:21]
  wire [31:0] n32_O_4_1; // @[Top.scala 730:21]
  wire [31:0] n32_O_5_0; // @[Top.scala 730:21]
  wire [31:0] n32_O_5_1; // @[Top.scala 730:21]
  wire [31:0] n32_O_6_0; // @[Top.scala 730:21]
  wire [31:0] n32_O_6_1; // @[Top.scala 730:21]
  wire [31:0] n32_O_7_0; // @[Top.scala 730:21]
  wire [31:0] n32_O_7_1; // @[Top.scala 730:21]
  wire  n39_valid_up; // @[Top.scala 734:21]
  wire  n39_valid_down; // @[Top.scala 734:21]
  wire [31:0] n39_I0_0_0; // @[Top.scala 734:21]
  wire [31:0] n39_I0_0_1; // @[Top.scala 734:21]
  wire [31:0] n39_I0_1_0; // @[Top.scala 734:21]
  wire [31:0] n39_I0_1_1; // @[Top.scala 734:21]
  wire [31:0] n39_I0_2_0; // @[Top.scala 734:21]
  wire [31:0] n39_I0_2_1; // @[Top.scala 734:21]
  wire [31:0] n39_I0_3_0; // @[Top.scala 734:21]
  wire [31:0] n39_I0_3_1; // @[Top.scala 734:21]
  wire [31:0] n39_I0_4_0; // @[Top.scala 734:21]
  wire [31:0] n39_I0_4_1; // @[Top.scala 734:21]
  wire [31:0] n39_I0_5_0; // @[Top.scala 734:21]
  wire [31:0] n39_I0_5_1; // @[Top.scala 734:21]
  wire [31:0] n39_I0_6_0; // @[Top.scala 734:21]
  wire [31:0] n39_I0_6_1; // @[Top.scala 734:21]
  wire [31:0] n39_I0_7_0; // @[Top.scala 734:21]
  wire [31:0] n39_I0_7_1; // @[Top.scala 734:21]
  wire [31:0] n39_I1_0; // @[Top.scala 734:21]
  wire [31:0] n39_I1_1; // @[Top.scala 734:21]
  wire [31:0] n39_I1_2; // @[Top.scala 734:21]
  wire [31:0] n39_I1_3; // @[Top.scala 734:21]
  wire [31:0] n39_I1_4; // @[Top.scala 734:21]
  wire [31:0] n39_I1_5; // @[Top.scala 734:21]
  wire [31:0] n39_I1_6; // @[Top.scala 734:21]
  wire [31:0] n39_I1_7; // @[Top.scala 734:21]
  wire [31:0] n39_O_0_0; // @[Top.scala 734:21]
  wire [31:0] n39_O_0_1; // @[Top.scala 734:21]
  wire [31:0] n39_O_0_2; // @[Top.scala 734:21]
  wire [31:0] n39_O_1_0; // @[Top.scala 734:21]
  wire [31:0] n39_O_1_1; // @[Top.scala 734:21]
  wire [31:0] n39_O_1_2; // @[Top.scala 734:21]
  wire [31:0] n39_O_2_0; // @[Top.scala 734:21]
  wire [31:0] n39_O_2_1; // @[Top.scala 734:21]
  wire [31:0] n39_O_2_2; // @[Top.scala 734:21]
  wire [31:0] n39_O_3_0; // @[Top.scala 734:21]
  wire [31:0] n39_O_3_1; // @[Top.scala 734:21]
  wire [31:0] n39_O_3_2; // @[Top.scala 734:21]
  wire [31:0] n39_O_4_0; // @[Top.scala 734:21]
  wire [31:0] n39_O_4_1; // @[Top.scala 734:21]
  wire [31:0] n39_O_4_2; // @[Top.scala 734:21]
  wire [31:0] n39_O_5_0; // @[Top.scala 734:21]
  wire [31:0] n39_O_5_1; // @[Top.scala 734:21]
  wire [31:0] n39_O_5_2; // @[Top.scala 734:21]
  wire [31:0] n39_O_6_0; // @[Top.scala 734:21]
  wire [31:0] n39_O_6_1; // @[Top.scala 734:21]
  wire [31:0] n39_O_6_2; // @[Top.scala 734:21]
  wire [31:0] n39_O_7_0; // @[Top.scala 734:21]
  wire [31:0] n39_O_7_1; // @[Top.scala 734:21]
  wire [31:0] n39_O_7_2; // @[Top.scala 734:21]
  wire  n48_valid_up; // @[Top.scala 738:21]
  wire  n48_valid_down; // @[Top.scala 738:21]
  wire [31:0] n48_I_0_0; // @[Top.scala 738:21]
  wire [31:0] n48_I_0_1; // @[Top.scala 738:21]
  wire [31:0] n48_I_0_2; // @[Top.scala 738:21]
  wire [31:0] n48_I_1_0; // @[Top.scala 738:21]
  wire [31:0] n48_I_1_1; // @[Top.scala 738:21]
  wire [31:0] n48_I_1_2; // @[Top.scala 738:21]
  wire [31:0] n48_I_2_0; // @[Top.scala 738:21]
  wire [31:0] n48_I_2_1; // @[Top.scala 738:21]
  wire [31:0] n48_I_2_2; // @[Top.scala 738:21]
  wire [31:0] n48_I_3_0; // @[Top.scala 738:21]
  wire [31:0] n48_I_3_1; // @[Top.scala 738:21]
  wire [31:0] n48_I_3_2; // @[Top.scala 738:21]
  wire [31:0] n48_I_4_0; // @[Top.scala 738:21]
  wire [31:0] n48_I_4_1; // @[Top.scala 738:21]
  wire [31:0] n48_I_4_2; // @[Top.scala 738:21]
  wire [31:0] n48_I_5_0; // @[Top.scala 738:21]
  wire [31:0] n48_I_5_1; // @[Top.scala 738:21]
  wire [31:0] n48_I_5_2; // @[Top.scala 738:21]
  wire [31:0] n48_I_6_0; // @[Top.scala 738:21]
  wire [31:0] n48_I_6_1; // @[Top.scala 738:21]
  wire [31:0] n48_I_6_2; // @[Top.scala 738:21]
  wire [31:0] n48_I_7_0; // @[Top.scala 738:21]
  wire [31:0] n48_I_7_1; // @[Top.scala 738:21]
  wire [31:0] n48_I_7_2; // @[Top.scala 738:21]
  wire [31:0] n48_O_0_0_0; // @[Top.scala 738:21]
  wire [31:0] n48_O_0_0_1; // @[Top.scala 738:21]
  wire [31:0] n48_O_0_0_2; // @[Top.scala 738:21]
  wire [31:0] n48_O_1_0_0; // @[Top.scala 738:21]
  wire [31:0] n48_O_1_0_1; // @[Top.scala 738:21]
  wire [31:0] n48_O_1_0_2; // @[Top.scala 738:21]
  wire [31:0] n48_O_2_0_0; // @[Top.scala 738:21]
  wire [31:0] n48_O_2_0_1; // @[Top.scala 738:21]
  wire [31:0] n48_O_2_0_2; // @[Top.scala 738:21]
  wire [31:0] n48_O_3_0_0; // @[Top.scala 738:21]
  wire [31:0] n48_O_3_0_1; // @[Top.scala 738:21]
  wire [31:0] n48_O_3_0_2; // @[Top.scala 738:21]
  wire [31:0] n48_O_4_0_0; // @[Top.scala 738:21]
  wire [31:0] n48_O_4_0_1; // @[Top.scala 738:21]
  wire [31:0] n48_O_4_0_2; // @[Top.scala 738:21]
  wire [31:0] n48_O_5_0_0; // @[Top.scala 738:21]
  wire [31:0] n48_O_5_0_1; // @[Top.scala 738:21]
  wire [31:0] n48_O_5_0_2; // @[Top.scala 738:21]
  wire [31:0] n48_O_6_0_0; // @[Top.scala 738:21]
  wire [31:0] n48_O_6_0_1; // @[Top.scala 738:21]
  wire [31:0] n48_O_6_0_2; // @[Top.scala 738:21]
  wire [31:0] n48_O_7_0_0; // @[Top.scala 738:21]
  wire [31:0] n48_O_7_0_1; // @[Top.scala 738:21]
  wire [31:0] n48_O_7_0_2; // @[Top.scala 738:21]
  wire  n55_valid_up; // @[Top.scala 741:21]
  wire  n55_valid_down; // @[Top.scala 741:21]
  wire [31:0] n55_I_0_0_0; // @[Top.scala 741:21]
  wire [31:0] n55_I_0_0_1; // @[Top.scala 741:21]
  wire [31:0] n55_I_0_0_2; // @[Top.scala 741:21]
  wire [31:0] n55_I_1_0_0; // @[Top.scala 741:21]
  wire [31:0] n55_I_1_0_1; // @[Top.scala 741:21]
  wire [31:0] n55_I_1_0_2; // @[Top.scala 741:21]
  wire [31:0] n55_I_2_0_0; // @[Top.scala 741:21]
  wire [31:0] n55_I_2_0_1; // @[Top.scala 741:21]
  wire [31:0] n55_I_2_0_2; // @[Top.scala 741:21]
  wire [31:0] n55_I_3_0_0; // @[Top.scala 741:21]
  wire [31:0] n55_I_3_0_1; // @[Top.scala 741:21]
  wire [31:0] n55_I_3_0_2; // @[Top.scala 741:21]
  wire [31:0] n55_I_4_0_0; // @[Top.scala 741:21]
  wire [31:0] n55_I_4_0_1; // @[Top.scala 741:21]
  wire [31:0] n55_I_4_0_2; // @[Top.scala 741:21]
  wire [31:0] n55_I_5_0_0; // @[Top.scala 741:21]
  wire [31:0] n55_I_5_0_1; // @[Top.scala 741:21]
  wire [31:0] n55_I_5_0_2; // @[Top.scala 741:21]
  wire [31:0] n55_I_6_0_0; // @[Top.scala 741:21]
  wire [31:0] n55_I_6_0_1; // @[Top.scala 741:21]
  wire [31:0] n55_I_6_0_2; // @[Top.scala 741:21]
  wire [31:0] n55_I_7_0_0; // @[Top.scala 741:21]
  wire [31:0] n55_I_7_0_1; // @[Top.scala 741:21]
  wire [31:0] n55_I_7_0_2; // @[Top.scala 741:21]
  wire [31:0] n55_O_0_0; // @[Top.scala 741:21]
  wire [31:0] n55_O_0_1; // @[Top.scala 741:21]
  wire [31:0] n55_O_0_2; // @[Top.scala 741:21]
  wire [31:0] n55_O_1_0; // @[Top.scala 741:21]
  wire [31:0] n55_O_1_1; // @[Top.scala 741:21]
  wire [31:0] n55_O_1_2; // @[Top.scala 741:21]
  wire [31:0] n55_O_2_0; // @[Top.scala 741:21]
  wire [31:0] n55_O_2_1; // @[Top.scala 741:21]
  wire [31:0] n55_O_2_2; // @[Top.scala 741:21]
  wire [31:0] n55_O_3_0; // @[Top.scala 741:21]
  wire [31:0] n55_O_3_1; // @[Top.scala 741:21]
  wire [31:0] n55_O_3_2; // @[Top.scala 741:21]
  wire [31:0] n55_O_4_0; // @[Top.scala 741:21]
  wire [31:0] n55_O_4_1; // @[Top.scala 741:21]
  wire [31:0] n55_O_4_2; // @[Top.scala 741:21]
  wire [31:0] n55_O_5_0; // @[Top.scala 741:21]
  wire [31:0] n55_O_5_1; // @[Top.scala 741:21]
  wire [31:0] n55_O_5_2; // @[Top.scala 741:21]
  wire [31:0] n55_O_6_0; // @[Top.scala 741:21]
  wire [31:0] n55_O_6_1; // @[Top.scala 741:21]
  wire [31:0] n55_O_6_2; // @[Top.scala 741:21]
  wire [31:0] n55_O_7_0; // @[Top.scala 741:21]
  wire [31:0] n55_O_7_1; // @[Top.scala 741:21]
  wire [31:0] n55_O_7_2; // @[Top.scala 741:21]
  wire  n56_valid_up; // @[Top.scala 744:21]
  wire  n56_valid_down; // @[Top.scala 744:21]
  wire [31:0] n56_I0_0_0; // @[Top.scala 744:21]
  wire [31:0] n56_I0_0_1; // @[Top.scala 744:21]
  wire [31:0] n56_I0_0_2; // @[Top.scala 744:21]
  wire [31:0] n56_I0_1_0; // @[Top.scala 744:21]
  wire [31:0] n56_I0_1_1; // @[Top.scala 744:21]
  wire [31:0] n56_I0_1_2; // @[Top.scala 744:21]
  wire [31:0] n56_I0_2_0; // @[Top.scala 744:21]
  wire [31:0] n56_I0_2_1; // @[Top.scala 744:21]
  wire [31:0] n56_I0_2_2; // @[Top.scala 744:21]
  wire [31:0] n56_I0_3_0; // @[Top.scala 744:21]
  wire [31:0] n56_I0_3_1; // @[Top.scala 744:21]
  wire [31:0] n56_I0_3_2; // @[Top.scala 744:21]
  wire [31:0] n56_I0_4_0; // @[Top.scala 744:21]
  wire [31:0] n56_I0_4_1; // @[Top.scala 744:21]
  wire [31:0] n56_I0_4_2; // @[Top.scala 744:21]
  wire [31:0] n56_I0_5_0; // @[Top.scala 744:21]
  wire [31:0] n56_I0_5_1; // @[Top.scala 744:21]
  wire [31:0] n56_I0_5_2; // @[Top.scala 744:21]
  wire [31:0] n56_I0_6_0; // @[Top.scala 744:21]
  wire [31:0] n56_I0_6_1; // @[Top.scala 744:21]
  wire [31:0] n56_I0_6_2; // @[Top.scala 744:21]
  wire [31:0] n56_I0_7_0; // @[Top.scala 744:21]
  wire [31:0] n56_I0_7_1; // @[Top.scala 744:21]
  wire [31:0] n56_I0_7_2; // @[Top.scala 744:21]
  wire [31:0] n56_I1_0_0; // @[Top.scala 744:21]
  wire [31:0] n56_I1_0_1; // @[Top.scala 744:21]
  wire [31:0] n56_I1_0_2; // @[Top.scala 744:21]
  wire [31:0] n56_I1_1_0; // @[Top.scala 744:21]
  wire [31:0] n56_I1_1_1; // @[Top.scala 744:21]
  wire [31:0] n56_I1_1_2; // @[Top.scala 744:21]
  wire [31:0] n56_I1_2_0; // @[Top.scala 744:21]
  wire [31:0] n56_I1_2_1; // @[Top.scala 744:21]
  wire [31:0] n56_I1_2_2; // @[Top.scala 744:21]
  wire [31:0] n56_I1_3_0; // @[Top.scala 744:21]
  wire [31:0] n56_I1_3_1; // @[Top.scala 744:21]
  wire [31:0] n56_I1_3_2; // @[Top.scala 744:21]
  wire [31:0] n56_I1_4_0; // @[Top.scala 744:21]
  wire [31:0] n56_I1_4_1; // @[Top.scala 744:21]
  wire [31:0] n56_I1_4_2; // @[Top.scala 744:21]
  wire [31:0] n56_I1_5_0; // @[Top.scala 744:21]
  wire [31:0] n56_I1_5_1; // @[Top.scala 744:21]
  wire [31:0] n56_I1_5_2; // @[Top.scala 744:21]
  wire [31:0] n56_I1_6_0; // @[Top.scala 744:21]
  wire [31:0] n56_I1_6_1; // @[Top.scala 744:21]
  wire [31:0] n56_I1_6_2; // @[Top.scala 744:21]
  wire [31:0] n56_I1_7_0; // @[Top.scala 744:21]
  wire [31:0] n56_I1_7_1; // @[Top.scala 744:21]
  wire [31:0] n56_I1_7_2; // @[Top.scala 744:21]
  wire [31:0] n56_O_0_0_0; // @[Top.scala 744:21]
  wire [31:0] n56_O_0_0_1; // @[Top.scala 744:21]
  wire [31:0] n56_O_0_0_2; // @[Top.scala 744:21]
  wire [31:0] n56_O_0_1_0; // @[Top.scala 744:21]
  wire [31:0] n56_O_0_1_1; // @[Top.scala 744:21]
  wire [31:0] n56_O_0_1_2; // @[Top.scala 744:21]
  wire [31:0] n56_O_1_0_0; // @[Top.scala 744:21]
  wire [31:0] n56_O_1_0_1; // @[Top.scala 744:21]
  wire [31:0] n56_O_1_0_2; // @[Top.scala 744:21]
  wire [31:0] n56_O_1_1_0; // @[Top.scala 744:21]
  wire [31:0] n56_O_1_1_1; // @[Top.scala 744:21]
  wire [31:0] n56_O_1_1_2; // @[Top.scala 744:21]
  wire [31:0] n56_O_2_0_0; // @[Top.scala 744:21]
  wire [31:0] n56_O_2_0_1; // @[Top.scala 744:21]
  wire [31:0] n56_O_2_0_2; // @[Top.scala 744:21]
  wire [31:0] n56_O_2_1_0; // @[Top.scala 744:21]
  wire [31:0] n56_O_2_1_1; // @[Top.scala 744:21]
  wire [31:0] n56_O_2_1_2; // @[Top.scala 744:21]
  wire [31:0] n56_O_3_0_0; // @[Top.scala 744:21]
  wire [31:0] n56_O_3_0_1; // @[Top.scala 744:21]
  wire [31:0] n56_O_3_0_2; // @[Top.scala 744:21]
  wire [31:0] n56_O_3_1_0; // @[Top.scala 744:21]
  wire [31:0] n56_O_3_1_1; // @[Top.scala 744:21]
  wire [31:0] n56_O_3_1_2; // @[Top.scala 744:21]
  wire [31:0] n56_O_4_0_0; // @[Top.scala 744:21]
  wire [31:0] n56_O_4_0_1; // @[Top.scala 744:21]
  wire [31:0] n56_O_4_0_2; // @[Top.scala 744:21]
  wire [31:0] n56_O_4_1_0; // @[Top.scala 744:21]
  wire [31:0] n56_O_4_1_1; // @[Top.scala 744:21]
  wire [31:0] n56_O_4_1_2; // @[Top.scala 744:21]
  wire [31:0] n56_O_5_0_0; // @[Top.scala 744:21]
  wire [31:0] n56_O_5_0_1; // @[Top.scala 744:21]
  wire [31:0] n56_O_5_0_2; // @[Top.scala 744:21]
  wire [31:0] n56_O_5_1_0; // @[Top.scala 744:21]
  wire [31:0] n56_O_5_1_1; // @[Top.scala 744:21]
  wire [31:0] n56_O_5_1_2; // @[Top.scala 744:21]
  wire [31:0] n56_O_6_0_0; // @[Top.scala 744:21]
  wire [31:0] n56_O_6_0_1; // @[Top.scala 744:21]
  wire [31:0] n56_O_6_0_2; // @[Top.scala 744:21]
  wire [31:0] n56_O_6_1_0; // @[Top.scala 744:21]
  wire [31:0] n56_O_6_1_1; // @[Top.scala 744:21]
  wire [31:0] n56_O_6_1_2; // @[Top.scala 744:21]
  wire [31:0] n56_O_7_0_0; // @[Top.scala 744:21]
  wire [31:0] n56_O_7_0_1; // @[Top.scala 744:21]
  wire [31:0] n56_O_7_0_2; // @[Top.scala 744:21]
  wire [31:0] n56_O_7_1_0; // @[Top.scala 744:21]
  wire [31:0] n56_O_7_1_1; // @[Top.scala 744:21]
  wire [31:0] n56_O_7_1_2; // @[Top.scala 744:21]
  wire  n63_clock; // @[Top.scala 748:21]
  wire  n63_valid_up; // @[Top.scala 748:21]
  wire  n63_valid_down; // @[Top.scala 748:21]
  wire [31:0] n63_I_0; // @[Top.scala 748:21]
  wire [31:0] n63_I_1; // @[Top.scala 748:21]
  wire [31:0] n63_I_2; // @[Top.scala 748:21]
  wire [31:0] n63_I_3; // @[Top.scala 748:21]
  wire [31:0] n63_I_4; // @[Top.scala 748:21]
  wire [31:0] n63_I_5; // @[Top.scala 748:21]
  wire [31:0] n63_I_6; // @[Top.scala 748:21]
  wire [31:0] n63_I_7; // @[Top.scala 748:21]
  wire [31:0] n63_O_0; // @[Top.scala 748:21]
  wire [31:0] n63_O_1; // @[Top.scala 748:21]
  wire [31:0] n63_O_2; // @[Top.scala 748:21]
  wire [31:0] n63_O_3; // @[Top.scala 748:21]
  wire [31:0] n63_O_4; // @[Top.scala 748:21]
  wire [31:0] n63_O_5; // @[Top.scala 748:21]
  wire [31:0] n63_O_6; // @[Top.scala 748:21]
  wire [31:0] n63_O_7; // @[Top.scala 748:21]
  wire  n64_clock; // @[Top.scala 751:21]
  wire  n64_valid_up; // @[Top.scala 751:21]
  wire  n64_valid_down; // @[Top.scala 751:21]
  wire [31:0] n64_I_0; // @[Top.scala 751:21]
  wire [31:0] n64_I_1; // @[Top.scala 751:21]
  wire [31:0] n64_I_2; // @[Top.scala 751:21]
  wire [31:0] n64_I_3; // @[Top.scala 751:21]
  wire [31:0] n64_I_4; // @[Top.scala 751:21]
  wire [31:0] n64_I_5; // @[Top.scala 751:21]
  wire [31:0] n64_I_6; // @[Top.scala 751:21]
  wire [31:0] n64_I_7; // @[Top.scala 751:21]
  wire [31:0] n64_O_0; // @[Top.scala 751:21]
  wire [31:0] n64_O_1; // @[Top.scala 751:21]
  wire [31:0] n64_O_2; // @[Top.scala 751:21]
  wire [31:0] n64_O_3; // @[Top.scala 751:21]
  wire [31:0] n64_O_4; // @[Top.scala 751:21]
  wire [31:0] n64_O_5; // @[Top.scala 751:21]
  wire [31:0] n64_O_6; // @[Top.scala 751:21]
  wire [31:0] n64_O_7; // @[Top.scala 751:21]
  wire  n65_valid_up; // @[Top.scala 754:21]
  wire  n65_valid_down; // @[Top.scala 754:21]
  wire [31:0] n65_I0_0; // @[Top.scala 754:21]
  wire [31:0] n65_I0_1; // @[Top.scala 754:21]
  wire [31:0] n65_I0_2; // @[Top.scala 754:21]
  wire [31:0] n65_I0_3; // @[Top.scala 754:21]
  wire [31:0] n65_I0_4; // @[Top.scala 754:21]
  wire [31:0] n65_I0_5; // @[Top.scala 754:21]
  wire [31:0] n65_I0_6; // @[Top.scala 754:21]
  wire [31:0] n65_I0_7; // @[Top.scala 754:21]
  wire [31:0] n65_I1_0; // @[Top.scala 754:21]
  wire [31:0] n65_I1_1; // @[Top.scala 754:21]
  wire [31:0] n65_I1_2; // @[Top.scala 754:21]
  wire [31:0] n65_I1_3; // @[Top.scala 754:21]
  wire [31:0] n65_I1_4; // @[Top.scala 754:21]
  wire [31:0] n65_I1_5; // @[Top.scala 754:21]
  wire [31:0] n65_I1_6; // @[Top.scala 754:21]
  wire [31:0] n65_I1_7; // @[Top.scala 754:21]
  wire [31:0] n65_O_0_0; // @[Top.scala 754:21]
  wire [31:0] n65_O_0_1; // @[Top.scala 754:21]
  wire [31:0] n65_O_1_0; // @[Top.scala 754:21]
  wire [31:0] n65_O_1_1; // @[Top.scala 754:21]
  wire [31:0] n65_O_2_0; // @[Top.scala 754:21]
  wire [31:0] n65_O_2_1; // @[Top.scala 754:21]
  wire [31:0] n65_O_3_0; // @[Top.scala 754:21]
  wire [31:0] n65_O_3_1; // @[Top.scala 754:21]
  wire [31:0] n65_O_4_0; // @[Top.scala 754:21]
  wire [31:0] n65_O_4_1; // @[Top.scala 754:21]
  wire [31:0] n65_O_5_0; // @[Top.scala 754:21]
  wire [31:0] n65_O_5_1; // @[Top.scala 754:21]
  wire [31:0] n65_O_6_0; // @[Top.scala 754:21]
  wire [31:0] n65_O_6_1; // @[Top.scala 754:21]
  wire [31:0] n65_O_7_0; // @[Top.scala 754:21]
  wire [31:0] n65_O_7_1; // @[Top.scala 754:21]
  wire  n72_valid_up; // @[Top.scala 758:21]
  wire  n72_valid_down; // @[Top.scala 758:21]
  wire [31:0] n72_I0_0_0; // @[Top.scala 758:21]
  wire [31:0] n72_I0_0_1; // @[Top.scala 758:21]
  wire [31:0] n72_I0_1_0; // @[Top.scala 758:21]
  wire [31:0] n72_I0_1_1; // @[Top.scala 758:21]
  wire [31:0] n72_I0_2_0; // @[Top.scala 758:21]
  wire [31:0] n72_I0_2_1; // @[Top.scala 758:21]
  wire [31:0] n72_I0_3_0; // @[Top.scala 758:21]
  wire [31:0] n72_I0_3_1; // @[Top.scala 758:21]
  wire [31:0] n72_I0_4_0; // @[Top.scala 758:21]
  wire [31:0] n72_I0_4_1; // @[Top.scala 758:21]
  wire [31:0] n72_I0_5_0; // @[Top.scala 758:21]
  wire [31:0] n72_I0_5_1; // @[Top.scala 758:21]
  wire [31:0] n72_I0_6_0; // @[Top.scala 758:21]
  wire [31:0] n72_I0_6_1; // @[Top.scala 758:21]
  wire [31:0] n72_I0_7_0; // @[Top.scala 758:21]
  wire [31:0] n72_I0_7_1; // @[Top.scala 758:21]
  wire [31:0] n72_I1_0; // @[Top.scala 758:21]
  wire [31:0] n72_I1_1; // @[Top.scala 758:21]
  wire [31:0] n72_I1_2; // @[Top.scala 758:21]
  wire [31:0] n72_I1_3; // @[Top.scala 758:21]
  wire [31:0] n72_I1_4; // @[Top.scala 758:21]
  wire [31:0] n72_I1_5; // @[Top.scala 758:21]
  wire [31:0] n72_I1_6; // @[Top.scala 758:21]
  wire [31:0] n72_I1_7; // @[Top.scala 758:21]
  wire [31:0] n72_O_0_0; // @[Top.scala 758:21]
  wire [31:0] n72_O_0_1; // @[Top.scala 758:21]
  wire [31:0] n72_O_0_2; // @[Top.scala 758:21]
  wire [31:0] n72_O_1_0; // @[Top.scala 758:21]
  wire [31:0] n72_O_1_1; // @[Top.scala 758:21]
  wire [31:0] n72_O_1_2; // @[Top.scala 758:21]
  wire [31:0] n72_O_2_0; // @[Top.scala 758:21]
  wire [31:0] n72_O_2_1; // @[Top.scala 758:21]
  wire [31:0] n72_O_2_2; // @[Top.scala 758:21]
  wire [31:0] n72_O_3_0; // @[Top.scala 758:21]
  wire [31:0] n72_O_3_1; // @[Top.scala 758:21]
  wire [31:0] n72_O_3_2; // @[Top.scala 758:21]
  wire [31:0] n72_O_4_0; // @[Top.scala 758:21]
  wire [31:0] n72_O_4_1; // @[Top.scala 758:21]
  wire [31:0] n72_O_4_2; // @[Top.scala 758:21]
  wire [31:0] n72_O_5_0; // @[Top.scala 758:21]
  wire [31:0] n72_O_5_1; // @[Top.scala 758:21]
  wire [31:0] n72_O_5_2; // @[Top.scala 758:21]
  wire [31:0] n72_O_6_0; // @[Top.scala 758:21]
  wire [31:0] n72_O_6_1; // @[Top.scala 758:21]
  wire [31:0] n72_O_6_2; // @[Top.scala 758:21]
  wire [31:0] n72_O_7_0; // @[Top.scala 758:21]
  wire [31:0] n72_O_7_1; // @[Top.scala 758:21]
  wire [31:0] n72_O_7_2; // @[Top.scala 758:21]
  wire  n81_valid_up; // @[Top.scala 762:21]
  wire  n81_valid_down; // @[Top.scala 762:21]
  wire [31:0] n81_I_0_0; // @[Top.scala 762:21]
  wire [31:0] n81_I_0_1; // @[Top.scala 762:21]
  wire [31:0] n81_I_0_2; // @[Top.scala 762:21]
  wire [31:0] n81_I_1_0; // @[Top.scala 762:21]
  wire [31:0] n81_I_1_1; // @[Top.scala 762:21]
  wire [31:0] n81_I_1_2; // @[Top.scala 762:21]
  wire [31:0] n81_I_2_0; // @[Top.scala 762:21]
  wire [31:0] n81_I_2_1; // @[Top.scala 762:21]
  wire [31:0] n81_I_2_2; // @[Top.scala 762:21]
  wire [31:0] n81_I_3_0; // @[Top.scala 762:21]
  wire [31:0] n81_I_3_1; // @[Top.scala 762:21]
  wire [31:0] n81_I_3_2; // @[Top.scala 762:21]
  wire [31:0] n81_I_4_0; // @[Top.scala 762:21]
  wire [31:0] n81_I_4_1; // @[Top.scala 762:21]
  wire [31:0] n81_I_4_2; // @[Top.scala 762:21]
  wire [31:0] n81_I_5_0; // @[Top.scala 762:21]
  wire [31:0] n81_I_5_1; // @[Top.scala 762:21]
  wire [31:0] n81_I_5_2; // @[Top.scala 762:21]
  wire [31:0] n81_I_6_0; // @[Top.scala 762:21]
  wire [31:0] n81_I_6_1; // @[Top.scala 762:21]
  wire [31:0] n81_I_6_2; // @[Top.scala 762:21]
  wire [31:0] n81_I_7_0; // @[Top.scala 762:21]
  wire [31:0] n81_I_7_1; // @[Top.scala 762:21]
  wire [31:0] n81_I_7_2; // @[Top.scala 762:21]
  wire [31:0] n81_O_0_0_0; // @[Top.scala 762:21]
  wire [31:0] n81_O_0_0_1; // @[Top.scala 762:21]
  wire [31:0] n81_O_0_0_2; // @[Top.scala 762:21]
  wire [31:0] n81_O_1_0_0; // @[Top.scala 762:21]
  wire [31:0] n81_O_1_0_1; // @[Top.scala 762:21]
  wire [31:0] n81_O_1_0_2; // @[Top.scala 762:21]
  wire [31:0] n81_O_2_0_0; // @[Top.scala 762:21]
  wire [31:0] n81_O_2_0_1; // @[Top.scala 762:21]
  wire [31:0] n81_O_2_0_2; // @[Top.scala 762:21]
  wire [31:0] n81_O_3_0_0; // @[Top.scala 762:21]
  wire [31:0] n81_O_3_0_1; // @[Top.scala 762:21]
  wire [31:0] n81_O_3_0_2; // @[Top.scala 762:21]
  wire [31:0] n81_O_4_0_0; // @[Top.scala 762:21]
  wire [31:0] n81_O_4_0_1; // @[Top.scala 762:21]
  wire [31:0] n81_O_4_0_2; // @[Top.scala 762:21]
  wire [31:0] n81_O_5_0_0; // @[Top.scala 762:21]
  wire [31:0] n81_O_5_0_1; // @[Top.scala 762:21]
  wire [31:0] n81_O_5_0_2; // @[Top.scala 762:21]
  wire [31:0] n81_O_6_0_0; // @[Top.scala 762:21]
  wire [31:0] n81_O_6_0_1; // @[Top.scala 762:21]
  wire [31:0] n81_O_6_0_2; // @[Top.scala 762:21]
  wire [31:0] n81_O_7_0_0; // @[Top.scala 762:21]
  wire [31:0] n81_O_7_0_1; // @[Top.scala 762:21]
  wire [31:0] n81_O_7_0_2; // @[Top.scala 762:21]
  wire  n88_valid_up; // @[Top.scala 765:21]
  wire  n88_valid_down; // @[Top.scala 765:21]
  wire [31:0] n88_I_0_0_0; // @[Top.scala 765:21]
  wire [31:0] n88_I_0_0_1; // @[Top.scala 765:21]
  wire [31:0] n88_I_0_0_2; // @[Top.scala 765:21]
  wire [31:0] n88_I_1_0_0; // @[Top.scala 765:21]
  wire [31:0] n88_I_1_0_1; // @[Top.scala 765:21]
  wire [31:0] n88_I_1_0_2; // @[Top.scala 765:21]
  wire [31:0] n88_I_2_0_0; // @[Top.scala 765:21]
  wire [31:0] n88_I_2_0_1; // @[Top.scala 765:21]
  wire [31:0] n88_I_2_0_2; // @[Top.scala 765:21]
  wire [31:0] n88_I_3_0_0; // @[Top.scala 765:21]
  wire [31:0] n88_I_3_0_1; // @[Top.scala 765:21]
  wire [31:0] n88_I_3_0_2; // @[Top.scala 765:21]
  wire [31:0] n88_I_4_0_0; // @[Top.scala 765:21]
  wire [31:0] n88_I_4_0_1; // @[Top.scala 765:21]
  wire [31:0] n88_I_4_0_2; // @[Top.scala 765:21]
  wire [31:0] n88_I_5_0_0; // @[Top.scala 765:21]
  wire [31:0] n88_I_5_0_1; // @[Top.scala 765:21]
  wire [31:0] n88_I_5_0_2; // @[Top.scala 765:21]
  wire [31:0] n88_I_6_0_0; // @[Top.scala 765:21]
  wire [31:0] n88_I_6_0_1; // @[Top.scala 765:21]
  wire [31:0] n88_I_6_0_2; // @[Top.scala 765:21]
  wire [31:0] n88_I_7_0_0; // @[Top.scala 765:21]
  wire [31:0] n88_I_7_0_1; // @[Top.scala 765:21]
  wire [31:0] n88_I_7_0_2; // @[Top.scala 765:21]
  wire [31:0] n88_O_0_0; // @[Top.scala 765:21]
  wire [31:0] n88_O_0_1; // @[Top.scala 765:21]
  wire [31:0] n88_O_0_2; // @[Top.scala 765:21]
  wire [31:0] n88_O_1_0; // @[Top.scala 765:21]
  wire [31:0] n88_O_1_1; // @[Top.scala 765:21]
  wire [31:0] n88_O_1_2; // @[Top.scala 765:21]
  wire [31:0] n88_O_2_0; // @[Top.scala 765:21]
  wire [31:0] n88_O_2_1; // @[Top.scala 765:21]
  wire [31:0] n88_O_2_2; // @[Top.scala 765:21]
  wire [31:0] n88_O_3_0; // @[Top.scala 765:21]
  wire [31:0] n88_O_3_1; // @[Top.scala 765:21]
  wire [31:0] n88_O_3_2; // @[Top.scala 765:21]
  wire [31:0] n88_O_4_0; // @[Top.scala 765:21]
  wire [31:0] n88_O_4_1; // @[Top.scala 765:21]
  wire [31:0] n88_O_4_2; // @[Top.scala 765:21]
  wire [31:0] n88_O_5_0; // @[Top.scala 765:21]
  wire [31:0] n88_O_5_1; // @[Top.scala 765:21]
  wire [31:0] n88_O_5_2; // @[Top.scala 765:21]
  wire [31:0] n88_O_6_0; // @[Top.scala 765:21]
  wire [31:0] n88_O_6_1; // @[Top.scala 765:21]
  wire [31:0] n88_O_6_2; // @[Top.scala 765:21]
  wire [31:0] n88_O_7_0; // @[Top.scala 765:21]
  wire [31:0] n88_O_7_1; // @[Top.scala 765:21]
  wire [31:0] n88_O_7_2; // @[Top.scala 765:21]
  wire  n89_valid_up; // @[Top.scala 768:21]
  wire  n89_valid_down; // @[Top.scala 768:21]
  wire [31:0] n89_I0_0_0_0; // @[Top.scala 768:21]
  wire [31:0] n89_I0_0_0_1; // @[Top.scala 768:21]
  wire [31:0] n89_I0_0_0_2; // @[Top.scala 768:21]
  wire [31:0] n89_I0_0_1_0; // @[Top.scala 768:21]
  wire [31:0] n89_I0_0_1_1; // @[Top.scala 768:21]
  wire [31:0] n89_I0_0_1_2; // @[Top.scala 768:21]
  wire [31:0] n89_I0_1_0_0; // @[Top.scala 768:21]
  wire [31:0] n89_I0_1_0_1; // @[Top.scala 768:21]
  wire [31:0] n89_I0_1_0_2; // @[Top.scala 768:21]
  wire [31:0] n89_I0_1_1_0; // @[Top.scala 768:21]
  wire [31:0] n89_I0_1_1_1; // @[Top.scala 768:21]
  wire [31:0] n89_I0_1_1_2; // @[Top.scala 768:21]
  wire [31:0] n89_I0_2_0_0; // @[Top.scala 768:21]
  wire [31:0] n89_I0_2_0_1; // @[Top.scala 768:21]
  wire [31:0] n89_I0_2_0_2; // @[Top.scala 768:21]
  wire [31:0] n89_I0_2_1_0; // @[Top.scala 768:21]
  wire [31:0] n89_I0_2_1_1; // @[Top.scala 768:21]
  wire [31:0] n89_I0_2_1_2; // @[Top.scala 768:21]
  wire [31:0] n89_I0_3_0_0; // @[Top.scala 768:21]
  wire [31:0] n89_I0_3_0_1; // @[Top.scala 768:21]
  wire [31:0] n89_I0_3_0_2; // @[Top.scala 768:21]
  wire [31:0] n89_I0_3_1_0; // @[Top.scala 768:21]
  wire [31:0] n89_I0_3_1_1; // @[Top.scala 768:21]
  wire [31:0] n89_I0_3_1_2; // @[Top.scala 768:21]
  wire [31:0] n89_I0_4_0_0; // @[Top.scala 768:21]
  wire [31:0] n89_I0_4_0_1; // @[Top.scala 768:21]
  wire [31:0] n89_I0_4_0_2; // @[Top.scala 768:21]
  wire [31:0] n89_I0_4_1_0; // @[Top.scala 768:21]
  wire [31:0] n89_I0_4_1_1; // @[Top.scala 768:21]
  wire [31:0] n89_I0_4_1_2; // @[Top.scala 768:21]
  wire [31:0] n89_I0_5_0_0; // @[Top.scala 768:21]
  wire [31:0] n89_I0_5_0_1; // @[Top.scala 768:21]
  wire [31:0] n89_I0_5_0_2; // @[Top.scala 768:21]
  wire [31:0] n89_I0_5_1_0; // @[Top.scala 768:21]
  wire [31:0] n89_I0_5_1_1; // @[Top.scala 768:21]
  wire [31:0] n89_I0_5_1_2; // @[Top.scala 768:21]
  wire [31:0] n89_I0_6_0_0; // @[Top.scala 768:21]
  wire [31:0] n89_I0_6_0_1; // @[Top.scala 768:21]
  wire [31:0] n89_I0_6_0_2; // @[Top.scala 768:21]
  wire [31:0] n89_I0_6_1_0; // @[Top.scala 768:21]
  wire [31:0] n89_I0_6_1_1; // @[Top.scala 768:21]
  wire [31:0] n89_I0_6_1_2; // @[Top.scala 768:21]
  wire [31:0] n89_I0_7_0_0; // @[Top.scala 768:21]
  wire [31:0] n89_I0_7_0_1; // @[Top.scala 768:21]
  wire [31:0] n89_I0_7_0_2; // @[Top.scala 768:21]
  wire [31:0] n89_I0_7_1_0; // @[Top.scala 768:21]
  wire [31:0] n89_I0_7_1_1; // @[Top.scala 768:21]
  wire [31:0] n89_I0_7_1_2; // @[Top.scala 768:21]
  wire [31:0] n89_I1_0_0; // @[Top.scala 768:21]
  wire [31:0] n89_I1_0_1; // @[Top.scala 768:21]
  wire [31:0] n89_I1_0_2; // @[Top.scala 768:21]
  wire [31:0] n89_I1_1_0; // @[Top.scala 768:21]
  wire [31:0] n89_I1_1_1; // @[Top.scala 768:21]
  wire [31:0] n89_I1_1_2; // @[Top.scala 768:21]
  wire [31:0] n89_I1_2_0; // @[Top.scala 768:21]
  wire [31:0] n89_I1_2_1; // @[Top.scala 768:21]
  wire [31:0] n89_I1_2_2; // @[Top.scala 768:21]
  wire [31:0] n89_I1_3_0; // @[Top.scala 768:21]
  wire [31:0] n89_I1_3_1; // @[Top.scala 768:21]
  wire [31:0] n89_I1_3_2; // @[Top.scala 768:21]
  wire [31:0] n89_I1_4_0; // @[Top.scala 768:21]
  wire [31:0] n89_I1_4_1; // @[Top.scala 768:21]
  wire [31:0] n89_I1_4_2; // @[Top.scala 768:21]
  wire [31:0] n89_I1_5_0; // @[Top.scala 768:21]
  wire [31:0] n89_I1_5_1; // @[Top.scala 768:21]
  wire [31:0] n89_I1_5_2; // @[Top.scala 768:21]
  wire [31:0] n89_I1_6_0; // @[Top.scala 768:21]
  wire [31:0] n89_I1_6_1; // @[Top.scala 768:21]
  wire [31:0] n89_I1_6_2; // @[Top.scala 768:21]
  wire [31:0] n89_I1_7_0; // @[Top.scala 768:21]
  wire [31:0] n89_I1_7_1; // @[Top.scala 768:21]
  wire [31:0] n89_I1_7_2; // @[Top.scala 768:21]
  wire [31:0] n89_O_0_0_0; // @[Top.scala 768:21]
  wire [31:0] n89_O_0_0_1; // @[Top.scala 768:21]
  wire [31:0] n89_O_0_0_2; // @[Top.scala 768:21]
  wire [31:0] n89_O_0_1_0; // @[Top.scala 768:21]
  wire [31:0] n89_O_0_1_1; // @[Top.scala 768:21]
  wire [31:0] n89_O_0_1_2; // @[Top.scala 768:21]
  wire [31:0] n89_O_0_2_0; // @[Top.scala 768:21]
  wire [31:0] n89_O_0_2_1; // @[Top.scala 768:21]
  wire [31:0] n89_O_0_2_2; // @[Top.scala 768:21]
  wire [31:0] n89_O_1_0_0; // @[Top.scala 768:21]
  wire [31:0] n89_O_1_0_1; // @[Top.scala 768:21]
  wire [31:0] n89_O_1_0_2; // @[Top.scala 768:21]
  wire [31:0] n89_O_1_1_0; // @[Top.scala 768:21]
  wire [31:0] n89_O_1_1_1; // @[Top.scala 768:21]
  wire [31:0] n89_O_1_1_2; // @[Top.scala 768:21]
  wire [31:0] n89_O_1_2_0; // @[Top.scala 768:21]
  wire [31:0] n89_O_1_2_1; // @[Top.scala 768:21]
  wire [31:0] n89_O_1_2_2; // @[Top.scala 768:21]
  wire [31:0] n89_O_2_0_0; // @[Top.scala 768:21]
  wire [31:0] n89_O_2_0_1; // @[Top.scala 768:21]
  wire [31:0] n89_O_2_0_2; // @[Top.scala 768:21]
  wire [31:0] n89_O_2_1_0; // @[Top.scala 768:21]
  wire [31:0] n89_O_2_1_1; // @[Top.scala 768:21]
  wire [31:0] n89_O_2_1_2; // @[Top.scala 768:21]
  wire [31:0] n89_O_2_2_0; // @[Top.scala 768:21]
  wire [31:0] n89_O_2_2_1; // @[Top.scala 768:21]
  wire [31:0] n89_O_2_2_2; // @[Top.scala 768:21]
  wire [31:0] n89_O_3_0_0; // @[Top.scala 768:21]
  wire [31:0] n89_O_3_0_1; // @[Top.scala 768:21]
  wire [31:0] n89_O_3_0_2; // @[Top.scala 768:21]
  wire [31:0] n89_O_3_1_0; // @[Top.scala 768:21]
  wire [31:0] n89_O_3_1_1; // @[Top.scala 768:21]
  wire [31:0] n89_O_3_1_2; // @[Top.scala 768:21]
  wire [31:0] n89_O_3_2_0; // @[Top.scala 768:21]
  wire [31:0] n89_O_3_2_1; // @[Top.scala 768:21]
  wire [31:0] n89_O_3_2_2; // @[Top.scala 768:21]
  wire [31:0] n89_O_4_0_0; // @[Top.scala 768:21]
  wire [31:0] n89_O_4_0_1; // @[Top.scala 768:21]
  wire [31:0] n89_O_4_0_2; // @[Top.scala 768:21]
  wire [31:0] n89_O_4_1_0; // @[Top.scala 768:21]
  wire [31:0] n89_O_4_1_1; // @[Top.scala 768:21]
  wire [31:0] n89_O_4_1_2; // @[Top.scala 768:21]
  wire [31:0] n89_O_4_2_0; // @[Top.scala 768:21]
  wire [31:0] n89_O_4_2_1; // @[Top.scala 768:21]
  wire [31:0] n89_O_4_2_2; // @[Top.scala 768:21]
  wire [31:0] n89_O_5_0_0; // @[Top.scala 768:21]
  wire [31:0] n89_O_5_0_1; // @[Top.scala 768:21]
  wire [31:0] n89_O_5_0_2; // @[Top.scala 768:21]
  wire [31:0] n89_O_5_1_0; // @[Top.scala 768:21]
  wire [31:0] n89_O_5_1_1; // @[Top.scala 768:21]
  wire [31:0] n89_O_5_1_2; // @[Top.scala 768:21]
  wire [31:0] n89_O_5_2_0; // @[Top.scala 768:21]
  wire [31:0] n89_O_5_2_1; // @[Top.scala 768:21]
  wire [31:0] n89_O_5_2_2; // @[Top.scala 768:21]
  wire [31:0] n89_O_6_0_0; // @[Top.scala 768:21]
  wire [31:0] n89_O_6_0_1; // @[Top.scala 768:21]
  wire [31:0] n89_O_6_0_2; // @[Top.scala 768:21]
  wire [31:0] n89_O_6_1_0; // @[Top.scala 768:21]
  wire [31:0] n89_O_6_1_1; // @[Top.scala 768:21]
  wire [31:0] n89_O_6_1_2; // @[Top.scala 768:21]
  wire [31:0] n89_O_6_2_0; // @[Top.scala 768:21]
  wire [31:0] n89_O_6_2_1; // @[Top.scala 768:21]
  wire [31:0] n89_O_6_2_2; // @[Top.scala 768:21]
  wire [31:0] n89_O_7_0_0; // @[Top.scala 768:21]
  wire [31:0] n89_O_7_0_1; // @[Top.scala 768:21]
  wire [31:0] n89_O_7_0_2; // @[Top.scala 768:21]
  wire [31:0] n89_O_7_1_0; // @[Top.scala 768:21]
  wire [31:0] n89_O_7_1_1; // @[Top.scala 768:21]
  wire [31:0] n89_O_7_1_2; // @[Top.scala 768:21]
  wire [31:0] n89_O_7_2_0; // @[Top.scala 768:21]
  wire [31:0] n89_O_7_2_1; // @[Top.scala 768:21]
  wire [31:0] n89_O_7_2_2; // @[Top.scala 768:21]
  wire  n98_valid_up; // @[Top.scala 772:21]
  wire  n98_valid_down; // @[Top.scala 772:21]
  wire [31:0] n98_I_0_0_0; // @[Top.scala 772:21]
  wire [31:0] n98_I_0_0_1; // @[Top.scala 772:21]
  wire [31:0] n98_I_0_0_2; // @[Top.scala 772:21]
  wire [31:0] n98_I_0_1_0; // @[Top.scala 772:21]
  wire [31:0] n98_I_0_1_1; // @[Top.scala 772:21]
  wire [31:0] n98_I_0_1_2; // @[Top.scala 772:21]
  wire [31:0] n98_I_0_2_0; // @[Top.scala 772:21]
  wire [31:0] n98_I_0_2_1; // @[Top.scala 772:21]
  wire [31:0] n98_I_0_2_2; // @[Top.scala 772:21]
  wire [31:0] n98_I_1_0_0; // @[Top.scala 772:21]
  wire [31:0] n98_I_1_0_1; // @[Top.scala 772:21]
  wire [31:0] n98_I_1_0_2; // @[Top.scala 772:21]
  wire [31:0] n98_I_1_1_0; // @[Top.scala 772:21]
  wire [31:0] n98_I_1_1_1; // @[Top.scala 772:21]
  wire [31:0] n98_I_1_1_2; // @[Top.scala 772:21]
  wire [31:0] n98_I_1_2_0; // @[Top.scala 772:21]
  wire [31:0] n98_I_1_2_1; // @[Top.scala 772:21]
  wire [31:0] n98_I_1_2_2; // @[Top.scala 772:21]
  wire [31:0] n98_I_2_0_0; // @[Top.scala 772:21]
  wire [31:0] n98_I_2_0_1; // @[Top.scala 772:21]
  wire [31:0] n98_I_2_0_2; // @[Top.scala 772:21]
  wire [31:0] n98_I_2_1_0; // @[Top.scala 772:21]
  wire [31:0] n98_I_2_1_1; // @[Top.scala 772:21]
  wire [31:0] n98_I_2_1_2; // @[Top.scala 772:21]
  wire [31:0] n98_I_2_2_0; // @[Top.scala 772:21]
  wire [31:0] n98_I_2_2_1; // @[Top.scala 772:21]
  wire [31:0] n98_I_2_2_2; // @[Top.scala 772:21]
  wire [31:0] n98_I_3_0_0; // @[Top.scala 772:21]
  wire [31:0] n98_I_3_0_1; // @[Top.scala 772:21]
  wire [31:0] n98_I_3_0_2; // @[Top.scala 772:21]
  wire [31:0] n98_I_3_1_0; // @[Top.scala 772:21]
  wire [31:0] n98_I_3_1_1; // @[Top.scala 772:21]
  wire [31:0] n98_I_3_1_2; // @[Top.scala 772:21]
  wire [31:0] n98_I_3_2_0; // @[Top.scala 772:21]
  wire [31:0] n98_I_3_2_1; // @[Top.scala 772:21]
  wire [31:0] n98_I_3_2_2; // @[Top.scala 772:21]
  wire [31:0] n98_I_4_0_0; // @[Top.scala 772:21]
  wire [31:0] n98_I_4_0_1; // @[Top.scala 772:21]
  wire [31:0] n98_I_4_0_2; // @[Top.scala 772:21]
  wire [31:0] n98_I_4_1_0; // @[Top.scala 772:21]
  wire [31:0] n98_I_4_1_1; // @[Top.scala 772:21]
  wire [31:0] n98_I_4_1_2; // @[Top.scala 772:21]
  wire [31:0] n98_I_4_2_0; // @[Top.scala 772:21]
  wire [31:0] n98_I_4_2_1; // @[Top.scala 772:21]
  wire [31:0] n98_I_4_2_2; // @[Top.scala 772:21]
  wire [31:0] n98_I_5_0_0; // @[Top.scala 772:21]
  wire [31:0] n98_I_5_0_1; // @[Top.scala 772:21]
  wire [31:0] n98_I_5_0_2; // @[Top.scala 772:21]
  wire [31:0] n98_I_5_1_0; // @[Top.scala 772:21]
  wire [31:0] n98_I_5_1_1; // @[Top.scala 772:21]
  wire [31:0] n98_I_5_1_2; // @[Top.scala 772:21]
  wire [31:0] n98_I_5_2_0; // @[Top.scala 772:21]
  wire [31:0] n98_I_5_2_1; // @[Top.scala 772:21]
  wire [31:0] n98_I_5_2_2; // @[Top.scala 772:21]
  wire [31:0] n98_I_6_0_0; // @[Top.scala 772:21]
  wire [31:0] n98_I_6_0_1; // @[Top.scala 772:21]
  wire [31:0] n98_I_6_0_2; // @[Top.scala 772:21]
  wire [31:0] n98_I_6_1_0; // @[Top.scala 772:21]
  wire [31:0] n98_I_6_1_1; // @[Top.scala 772:21]
  wire [31:0] n98_I_6_1_2; // @[Top.scala 772:21]
  wire [31:0] n98_I_6_2_0; // @[Top.scala 772:21]
  wire [31:0] n98_I_6_2_1; // @[Top.scala 772:21]
  wire [31:0] n98_I_6_2_2; // @[Top.scala 772:21]
  wire [31:0] n98_I_7_0_0; // @[Top.scala 772:21]
  wire [31:0] n98_I_7_0_1; // @[Top.scala 772:21]
  wire [31:0] n98_I_7_0_2; // @[Top.scala 772:21]
  wire [31:0] n98_I_7_1_0; // @[Top.scala 772:21]
  wire [31:0] n98_I_7_1_1; // @[Top.scala 772:21]
  wire [31:0] n98_I_7_1_2; // @[Top.scala 772:21]
  wire [31:0] n98_I_7_2_0; // @[Top.scala 772:21]
  wire [31:0] n98_I_7_2_1; // @[Top.scala 772:21]
  wire [31:0] n98_I_7_2_2; // @[Top.scala 772:21]
  wire [31:0] n98_O_0_0_0_0; // @[Top.scala 772:21]
  wire [31:0] n98_O_0_0_0_1; // @[Top.scala 772:21]
  wire [31:0] n98_O_0_0_0_2; // @[Top.scala 772:21]
  wire [31:0] n98_O_0_0_1_0; // @[Top.scala 772:21]
  wire [31:0] n98_O_0_0_1_1; // @[Top.scala 772:21]
  wire [31:0] n98_O_0_0_1_2; // @[Top.scala 772:21]
  wire [31:0] n98_O_0_0_2_0; // @[Top.scala 772:21]
  wire [31:0] n98_O_0_0_2_1; // @[Top.scala 772:21]
  wire [31:0] n98_O_0_0_2_2; // @[Top.scala 772:21]
  wire [31:0] n98_O_1_0_0_0; // @[Top.scala 772:21]
  wire [31:0] n98_O_1_0_0_1; // @[Top.scala 772:21]
  wire [31:0] n98_O_1_0_0_2; // @[Top.scala 772:21]
  wire [31:0] n98_O_1_0_1_0; // @[Top.scala 772:21]
  wire [31:0] n98_O_1_0_1_1; // @[Top.scala 772:21]
  wire [31:0] n98_O_1_0_1_2; // @[Top.scala 772:21]
  wire [31:0] n98_O_1_0_2_0; // @[Top.scala 772:21]
  wire [31:0] n98_O_1_0_2_1; // @[Top.scala 772:21]
  wire [31:0] n98_O_1_0_2_2; // @[Top.scala 772:21]
  wire [31:0] n98_O_2_0_0_0; // @[Top.scala 772:21]
  wire [31:0] n98_O_2_0_0_1; // @[Top.scala 772:21]
  wire [31:0] n98_O_2_0_0_2; // @[Top.scala 772:21]
  wire [31:0] n98_O_2_0_1_0; // @[Top.scala 772:21]
  wire [31:0] n98_O_2_0_1_1; // @[Top.scala 772:21]
  wire [31:0] n98_O_2_0_1_2; // @[Top.scala 772:21]
  wire [31:0] n98_O_2_0_2_0; // @[Top.scala 772:21]
  wire [31:0] n98_O_2_0_2_1; // @[Top.scala 772:21]
  wire [31:0] n98_O_2_0_2_2; // @[Top.scala 772:21]
  wire [31:0] n98_O_3_0_0_0; // @[Top.scala 772:21]
  wire [31:0] n98_O_3_0_0_1; // @[Top.scala 772:21]
  wire [31:0] n98_O_3_0_0_2; // @[Top.scala 772:21]
  wire [31:0] n98_O_3_0_1_0; // @[Top.scala 772:21]
  wire [31:0] n98_O_3_0_1_1; // @[Top.scala 772:21]
  wire [31:0] n98_O_3_0_1_2; // @[Top.scala 772:21]
  wire [31:0] n98_O_3_0_2_0; // @[Top.scala 772:21]
  wire [31:0] n98_O_3_0_2_1; // @[Top.scala 772:21]
  wire [31:0] n98_O_3_0_2_2; // @[Top.scala 772:21]
  wire [31:0] n98_O_4_0_0_0; // @[Top.scala 772:21]
  wire [31:0] n98_O_4_0_0_1; // @[Top.scala 772:21]
  wire [31:0] n98_O_4_0_0_2; // @[Top.scala 772:21]
  wire [31:0] n98_O_4_0_1_0; // @[Top.scala 772:21]
  wire [31:0] n98_O_4_0_1_1; // @[Top.scala 772:21]
  wire [31:0] n98_O_4_0_1_2; // @[Top.scala 772:21]
  wire [31:0] n98_O_4_0_2_0; // @[Top.scala 772:21]
  wire [31:0] n98_O_4_0_2_1; // @[Top.scala 772:21]
  wire [31:0] n98_O_4_0_2_2; // @[Top.scala 772:21]
  wire [31:0] n98_O_5_0_0_0; // @[Top.scala 772:21]
  wire [31:0] n98_O_5_0_0_1; // @[Top.scala 772:21]
  wire [31:0] n98_O_5_0_0_2; // @[Top.scala 772:21]
  wire [31:0] n98_O_5_0_1_0; // @[Top.scala 772:21]
  wire [31:0] n98_O_5_0_1_1; // @[Top.scala 772:21]
  wire [31:0] n98_O_5_0_1_2; // @[Top.scala 772:21]
  wire [31:0] n98_O_5_0_2_0; // @[Top.scala 772:21]
  wire [31:0] n98_O_5_0_2_1; // @[Top.scala 772:21]
  wire [31:0] n98_O_5_0_2_2; // @[Top.scala 772:21]
  wire [31:0] n98_O_6_0_0_0; // @[Top.scala 772:21]
  wire [31:0] n98_O_6_0_0_1; // @[Top.scala 772:21]
  wire [31:0] n98_O_6_0_0_2; // @[Top.scala 772:21]
  wire [31:0] n98_O_6_0_1_0; // @[Top.scala 772:21]
  wire [31:0] n98_O_6_0_1_1; // @[Top.scala 772:21]
  wire [31:0] n98_O_6_0_1_2; // @[Top.scala 772:21]
  wire [31:0] n98_O_6_0_2_0; // @[Top.scala 772:21]
  wire [31:0] n98_O_6_0_2_1; // @[Top.scala 772:21]
  wire [31:0] n98_O_6_0_2_2; // @[Top.scala 772:21]
  wire [31:0] n98_O_7_0_0_0; // @[Top.scala 772:21]
  wire [31:0] n98_O_7_0_0_1; // @[Top.scala 772:21]
  wire [31:0] n98_O_7_0_0_2; // @[Top.scala 772:21]
  wire [31:0] n98_O_7_0_1_0; // @[Top.scala 772:21]
  wire [31:0] n98_O_7_0_1_1; // @[Top.scala 772:21]
  wire [31:0] n98_O_7_0_1_2; // @[Top.scala 772:21]
  wire [31:0] n98_O_7_0_2_0; // @[Top.scala 772:21]
  wire [31:0] n98_O_7_0_2_1; // @[Top.scala 772:21]
  wire [31:0] n98_O_7_0_2_2; // @[Top.scala 772:21]
  wire  n105_valid_up; // @[Top.scala 775:22]
  wire  n105_valid_down; // @[Top.scala 775:22]
  wire [31:0] n105_I_0_0_0_0; // @[Top.scala 775:22]
  wire [31:0] n105_I_0_0_0_1; // @[Top.scala 775:22]
  wire [31:0] n105_I_0_0_0_2; // @[Top.scala 775:22]
  wire [31:0] n105_I_0_0_1_0; // @[Top.scala 775:22]
  wire [31:0] n105_I_0_0_1_1; // @[Top.scala 775:22]
  wire [31:0] n105_I_0_0_1_2; // @[Top.scala 775:22]
  wire [31:0] n105_I_0_0_2_0; // @[Top.scala 775:22]
  wire [31:0] n105_I_0_0_2_1; // @[Top.scala 775:22]
  wire [31:0] n105_I_0_0_2_2; // @[Top.scala 775:22]
  wire [31:0] n105_I_1_0_0_0; // @[Top.scala 775:22]
  wire [31:0] n105_I_1_0_0_1; // @[Top.scala 775:22]
  wire [31:0] n105_I_1_0_0_2; // @[Top.scala 775:22]
  wire [31:0] n105_I_1_0_1_0; // @[Top.scala 775:22]
  wire [31:0] n105_I_1_0_1_1; // @[Top.scala 775:22]
  wire [31:0] n105_I_1_0_1_2; // @[Top.scala 775:22]
  wire [31:0] n105_I_1_0_2_0; // @[Top.scala 775:22]
  wire [31:0] n105_I_1_0_2_1; // @[Top.scala 775:22]
  wire [31:0] n105_I_1_0_2_2; // @[Top.scala 775:22]
  wire [31:0] n105_I_2_0_0_0; // @[Top.scala 775:22]
  wire [31:0] n105_I_2_0_0_1; // @[Top.scala 775:22]
  wire [31:0] n105_I_2_0_0_2; // @[Top.scala 775:22]
  wire [31:0] n105_I_2_0_1_0; // @[Top.scala 775:22]
  wire [31:0] n105_I_2_0_1_1; // @[Top.scala 775:22]
  wire [31:0] n105_I_2_0_1_2; // @[Top.scala 775:22]
  wire [31:0] n105_I_2_0_2_0; // @[Top.scala 775:22]
  wire [31:0] n105_I_2_0_2_1; // @[Top.scala 775:22]
  wire [31:0] n105_I_2_0_2_2; // @[Top.scala 775:22]
  wire [31:0] n105_I_3_0_0_0; // @[Top.scala 775:22]
  wire [31:0] n105_I_3_0_0_1; // @[Top.scala 775:22]
  wire [31:0] n105_I_3_0_0_2; // @[Top.scala 775:22]
  wire [31:0] n105_I_3_0_1_0; // @[Top.scala 775:22]
  wire [31:0] n105_I_3_0_1_1; // @[Top.scala 775:22]
  wire [31:0] n105_I_3_0_1_2; // @[Top.scala 775:22]
  wire [31:0] n105_I_3_0_2_0; // @[Top.scala 775:22]
  wire [31:0] n105_I_3_0_2_1; // @[Top.scala 775:22]
  wire [31:0] n105_I_3_0_2_2; // @[Top.scala 775:22]
  wire [31:0] n105_I_4_0_0_0; // @[Top.scala 775:22]
  wire [31:0] n105_I_4_0_0_1; // @[Top.scala 775:22]
  wire [31:0] n105_I_4_0_0_2; // @[Top.scala 775:22]
  wire [31:0] n105_I_4_0_1_0; // @[Top.scala 775:22]
  wire [31:0] n105_I_4_0_1_1; // @[Top.scala 775:22]
  wire [31:0] n105_I_4_0_1_2; // @[Top.scala 775:22]
  wire [31:0] n105_I_4_0_2_0; // @[Top.scala 775:22]
  wire [31:0] n105_I_4_0_2_1; // @[Top.scala 775:22]
  wire [31:0] n105_I_4_0_2_2; // @[Top.scala 775:22]
  wire [31:0] n105_I_5_0_0_0; // @[Top.scala 775:22]
  wire [31:0] n105_I_5_0_0_1; // @[Top.scala 775:22]
  wire [31:0] n105_I_5_0_0_2; // @[Top.scala 775:22]
  wire [31:0] n105_I_5_0_1_0; // @[Top.scala 775:22]
  wire [31:0] n105_I_5_0_1_1; // @[Top.scala 775:22]
  wire [31:0] n105_I_5_0_1_2; // @[Top.scala 775:22]
  wire [31:0] n105_I_5_0_2_0; // @[Top.scala 775:22]
  wire [31:0] n105_I_5_0_2_1; // @[Top.scala 775:22]
  wire [31:0] n105_I_5_0_2_2; // @[Top.scala 775:22]
  wire [31:0] n105_I_6_0_0_0; // @[Top.scala 775:22]
  wire [31:0] n105_I_6_0_0_1; // @[Top.scala 775:22]
  wire [31:0] n105_I_6_0_0_2; // @[Top.scala 775:22]
  wire [31:0] n105_I_6_0_1_0; // @[Top.scala 775:22]
  wire [31:0] n105_I_6_0_1_1; // @[Top.scala 775:22]
  wire [31:0] n105_I_6_0_1_2; // @[Top.scala 775:22]
  wire [31:0] n105_I_6_0_2_0; // @[Top.scala 775:22]
  wire [31:0] n105_I_6_0_2_1; // @[Top.scala 775:22]
  wire [31:0] n105_I_6_0_2_2; // @[Top.scala 775:22]
  wire [31:0] n105_I_7_0_0_0; // @[Top.scala 775:22]
  wire [31:0] n105_I_7_0_0_1; // @[Top.scala 775:22]
  wire [31:0] n105_I_7_0_0_2; // @[Top.scala 775:22]
  wire [31:0] n105_I_7_0_1_0; // @[Top.scala 775:22]
  wire [31:0] n105_I_7_0_1_1; // @[Top.scala 775:22]
  wire [31:0] n105_I_7_0_1_2; // @[Top.scala 775:22]
  wire [31:0] n105_I_7_0_2_0; // @[Top.scala 775:22]
  wire [31:0] n105_I_7_0_2_1; // @[Top.scala 775:22]
  wire [31:0] n105_I_7_0_2_2; // @[Top.scala 775:22]
  wire [31:0] n105_O_0_0_0; // @[Top.scala 775:22]
  wire [31:0] n105_O_0_0_1; // @[Top.scala 775:22]
  wire [31:0] n105_O_0_0_2; // @[Top.scala 775:22]
  wire [31:0] n105_O_0_1_0; // @[Top.scala 775:22]
  wire [31:0] n105_O_0_1_1; // @[Top.scala 775:22]
  wire [31:0] n105_O_0_1_2; // @[Top.scala 775:22]
  wire [31:0] n105_O_0_2_0; // @[Top.scala 775:22]
  wire [31:0] n105_O_0_2_1; // @[Top.scala 775:22]
  wire [31:0] n105_O_0_2_2; // @[Top.scala 775:22]
  wire [31:0] n105_O_1_0_0; // @[Top.scala 775:22]
  wire [31:0] n105_O_1_0_1; // @[Top.scala 775:22]
  wire [31:0] n105_O_1_0_2; // @[Top.scala 775:22]
  wire [31:0] n105_O_1_1_0; // @[Top.scala 775:22]
  wire [31:0] n105_O_1_1_1; // @[Top.scala 775:22]
  wire [31:0] n105_O_1_1_2; // @[Top.scala 775:22]
  wire [31:0] n105_O_1_2_0; // @[Top.scala 775:22]
  wire [31:0] n105_O_1_2_1; // @[Top.scala 775:22]
  wire [31:0] n105_O_1_2_2; // @[Top.scala 775:22]
  wire [31:0] n105_O_2_0_0; // @[Top.scala 775:22]
  wire [31:0] n105_O_2_0_1; // @[Top.scala 775:22]
  wire [31:0] n105_O_2_0_2; // @[Top.scala 775:22]
  wire [31:0] n105_O_2_1_0; // @[Top.scala 775:22]
  wire [31:0] n105_O_2_1_1; // @[Top.scala 775:22]
  wire [31:0] n105_O_2_1_2; // @[Top.scala 775:22]
  wire [31:0] n105_O_2_2_0; // @[Top.scala 775:22]
  wire [31:0] n105_O_2_2_1; // @[Top.scala 775:22]
  wire [31:0] n105_O_2_2_2; // @[Top.scala 775:22]
  wire [31:0] n105_O_3_0_0; // @[Top.scala 775:22]
  wire [31:0] n105_O_3_0_1; // @[Top.scala 775:22]
  wire [31:0] n105_O_3_0_2; // @[Top.scala 775:22]
  wire [31:0] n105_O_3_1_0; // @[Top.scala 775:22]
  wire [31:0] n105_O_3_1_1; // @[Top.scala 775:22]
  wire [31:0] n105_O_3_1_2; // @[Top.scala 775:22]
  wire [31:0] n105_O_3_2_0; // @[Top.scala 775:22]
  wire [31:0] n105_O_3_2_1; // @[Top.scala 775:22]
  wire [31:0] n105_O_3_2_2; // @[Top.scala 775:22]
  wire [31:0] n105_O_4_0_0; // @[Top.scala 775:22]
  wire [31:0] n105_O_4_0_1; // @[Top.scala 775:22]
  wire [31:0] n105_O_4_0_2; // @[Top.scala 775:22]
  wire [31:0] n105_O_4_1_0; // @[Top.scala 775:22]
  wire [31:0] n105_O_4_1_1; // @[Top.scala 775:22]
  wire [31:0] n105_O_4_1_2; // @[Top.scala 775:22]
  wire [31:0] n105_O_4_2_0; // @[Top.scala 775:22]
  wire [31:0] n105_O_4_2_1; // @[Top.scala 775:22]
  wire [31:0] n105_O_4_2_2; // @[Top.scala 775:22]
  wire [31:0] n105_O_5_0_0; // @[Top.scala 775:22]
  wire [31:0] n105_O_5_0_1; // @[Top.scala 775:22]
  wire [31:0] n105_O_5_0_2; // @[Top.scala 775:22]
  wire [31:0] n105_O_5_1_0; // @[Top.scala 775:22]
  wire [31:0] n105_O_5_1_1; // @[Top.scala 775:22]
  wire [31:0] n105_O_5_1_2; // @[Top.scala 775:22]
  wire [31:0] n105_O_5_2_0; // @[Top.scala 775:22]
  wire [31:0] n105_O_5_2_1; // @[Top.scala 775:22]
  wire [31:0] n105_O_5_2_2; // @[Top.scala 775:22]
  wire [31:0] n105_O_6_0_0; // @[Top.scala 775:22]
  wire [31:0] n105_O_6_0_1; // @[Top.scala 775:22]
  wire [31:0] n105_O_6_0_2; // @[Top.scala 775:22]
  wire [31:0] n105_O_6_1_0; // @[Top.scala 775:22]
  wire [31:0] n105_O_6_1_1; // @[Top.scala 775:22]
  wire [31:0] n105_O_6_1_2; // @[Top.scala 775:22]
  wire [31:0] n105_O_6_2_0; // @[Top.scala 775:22]
  wire [31:0] n105_O_6_2_1; // @[Top.scala 775:22]
  wire [31:0] n105_O_6_2_2; // @[Top.scala 775:22]
  wire [31:0] n105_O_7_0_0; // @[Top.scala 775:22]
  wire [31:0] n105_O_7_0_1; // @[Top.scala 775:22]
  wire [31:0] n105_O_7_0_2; // @[Top.scala 775:22]
  wire [31:0] n105_O_7_1_0; // @[Top.scala 775:22]
  wire [31:0] n105_O_7_1_1; // @[Top.scala 775:22]
  wire [31:0] n105_O_7_1_2; // @[Top.scala 775:22]
  wire [31:0] n105_O_7_2_0; // @[Top.scala 775:22]
  wire [31:0] n105_O_7_2_1; // @[Top.scala 775:22]
  wire [31:0] n105_O_7_2_2; // @[Top.scala 775:22]
  wire  n106_valid_up; // @[Top.scala 778:22]
  wire  n106_valid_down; // @[Top.scala 778:22]
  wire [31:0] n106_I_0_0_0; // @[Top.scala 778:22]
  wire [31:0] n106_I_0_0_1; // @[Top.scala 778:22]
  wire [31:0] n106_I_0_0_2; // @[Top.scala 778:22]
  wire [31:0] n106_I_0_1_0; // @[Top.scala 778:22]
  wire [31:0] n106_I_0_1_1; // @[Top.scala 778:22]
  wire [31:0] n106_I_0_1_2; // @[Top.scala 778:22]
  wire [31:0] n106_I_0_2_0; // @[Top.scala 778:22]
  wire [31:0] n106_I_0_2_1; // @[Top.scala 778:22]
  wire [31:0] n106_I_0_2_2; // @[Top.scala 778:22]
  wire [31:0] n106_I_1_0_0; // @[Top.scala 778:22]
  wire [31:0] n106_I_1_0_1; // @[Top.scala 778:22]
  wire [31:0] n106_I_1_0_2; // @[Top.scala 778:22]
  wire [31:0] n106_I_1_1_0; // @[Top.scala 778:22]
  wire [31:0] n106_I_1_1_1; // @[Top.scala 778:22]
  wire [31:0] n106_I_1_1_2; // @[Top.scala 778:22]
  wire [31:0] n106_I_1_2_0; // @[Top.scala 778:22]
  wire [31:0] n106_I_1_2_1; // @[Top.scala 778:22]
  wire [31:0] n106_I_1_2_2; // @[Top.scala 778:22]
  wire [31:0] n106_I_2_0_0; // @[Top.scala 778:22]
  wire [31:0] n106_I_2_0_1; // @[Top.scala 778:22]
  wire [31:0] n106_I_2_0_2; // @[Top.scala 778:22]
  wire [31:0] n106_I_2_1_0; // @[Top.scala 778:22]
  wire [31:0] n106_I_2_1_1; // @[Top.scala 778:22]
  wire [31:0] n106_I_2_1_2; // @[Top.scala 778:22]
  wire [31:0] n106_I_2_2_0; // @[Top.scala 778:22]
  wire [31:0] n106_I_2_2_1; // @[Top.scala 778:22]
  wire [31:0] n106_I_2_2_2; // @[Top.scala 778:22]
  wire [31:0] n106_I_3_0_0; // @[Top.scala 778:22]
  wire [31:0] n106_I_3_0_1; // @[Top.scala 778:22]
  wire [31:0] n106_I_3_0_2; // @[Top.scala 778:22]
  wire [31:0] n106_I_3_1_0; // @[Top.scala 778:22]
  wire [31:0] n106_I_3_1_1; // @[Top.scala 778:22]
  wire [31:0] n106_I_3_1_2; // @[Top.scala 778:22]
  wire [31:0] n106_I_3_2_0; // @[Top.scala 778:22]
  wire [31:0] n106_I_3_2_1; // @[Top.scala 778:22]
  wire [31:0] n106_I_3_2_2; // @[Top.scala 778:22]
  wire [31:0] n106_I_4_0_0; // @[Top.scala 778:22]
  wire [31:0] n106_I_4_0_1; // @[Top.scala 778:22]
  wire [31:0] n106_I_4_0_2; // @[Top.scala 778:22]
  wire [31:0] n106_I_4_1_0; // @[Top.scala 778:22]
  wire [31:0] n106_I_4_1_1; // @[Top.scala 778:22]
  wire [31:0] n106_I_4_1_2; // @[Top.scala 778:22]
  wire [31:0] n106_I_4_2_0; // @[Top.scala 778:22]
  wire [31:0] n106_I_4_2_1; // @[Top.scala 778:22]
  wire [31:0] n106_I_4_2_2; // @[Top.scala 778:22]
  wire [31:0] n106_I_5_0_0; // @[Top.scala 778:22]
  wire [31:0] n106_I_5_0_1; // @[Top.scala 778:22]
  wire [31:0] n106_I_5_0_2; // @[Top.scala 778:22]
  wire [31:0] n106_I_5_1_0; // @[Top.scala 778:22]
  wire [31:0] n106_I_5_1_1; // @[Top.scala 778:22]
  wire [31:0] n106_I_5_1_2; // @[Top.scala 778:22]
  wire [31:0] n106_I_5_2_0; // @[Top.scala 778:22]
  wire [31:0] n106_I_5_2_1; // @[Top.scala 778:22]
  wire [31:0] n106_I_5_2_2; // @[Top.scala 778:22]
  wire [31:0] n106_I_6_0_0; // @[Top.scala 778:22]
  wire [31:0] n106_I_6_0_1; // @[Top.scala 778:22]
  wire [31:0] n106_I_6_0_2; // @[Top.scala 778:22]
  wire [31:0] n106_I_6_1_0; // @[Top.scala 778:22]
  wire [31:0] n106_I_6_1_1; // @[Top.scala 778:22]
  wire [31:0] n106_I_6_1_2; // @[Top.scala 778:22]
  wire [31:0] n106_I_6_2_0; // @[Top.scala 778:22]
  wire [31:0] n106_I_6_2_1; // @[Top.scala 778:22]
  wire [31:0] n106_I_6_2_2; // @[Top.scala 778:22]
  wire [31:0] n106_I_7_0_0; // @[Top.scala 778:22]
  wire [31:0] n106_I_7_0_1; // @[Top.scala 778:22]
  wire [31:0] n106_I_7_0_2; // @[Top.scala 778:22]
  wire [31:0] n106_I_7_1_0; // @[Top.scala 778:22]
  wire [31:0] n106_I_7_1_1; // @[Top.scala 778:22]
  wire [31:0] n106_I_7_1_2; // @[Top.scala 778:22]
  wire [31:0] n106_I_7_2_0; // @[Top.scala 778:22]
  wire [31:0] n106_I_7_2_1; // @[Top.scala 778:22]
  wire [31:0] n106_I_7_2_2; // @[Top.scala 778:22]
  wire [31:0] n106_O_0_0_0; // @[Top.scala 778:22]
  wire [31:0] n106_O_0_0_1; // @[Top.scala 778:22]
  wire [31:0] n106_O_0_0_2; // @[Top.scala 778:22]
  wire [31:0] n106_O_0_1_0; // @[Top.scala 778:22]
  wire [31:0] n106_O_0_1_1; // @[Top.scala 778:22]
  wire [31:0] n106_O_0_1_2; // @[Top.scala 778:22]
  wire [31:0] n106_O_0_2_0; // @[Top.scala 778:22]
  wire [31:0] n106_O_0_2_1; // @[Top.scala 778:22]
  wire [31:0] n106_O_0_2_2; // @[Top.scala 778:22]
  wire [31:0] n106_O_1_0_0; // @[Top.scala 778:22]
  wire [31:0] n106_O_1_0_1; // @[Top.scala 778:22]
  wire [31:0] n106_O_1_0_2; // @[Top.scala 778:22]
  wire [31:0] n106_O_1_1_0; // @[Top.scala 778:22]
  wire [31:0] n106_O_1_1_1; // @[Top.scala 778:22]
  wire [31:0] n106_O_1_1_2; // @[Top.scala 778:22]
  wire [31:0] n106_O_1_2_0; // @[Top.scala 778:22]
  wire [31:0] n106_O_1_2_1; // @[Top.scala 778:22]
  wire [31:0] n106_O_1_2_2; // @[Top.scala 778:22]
  wire [31:0] n106_O_2_0_0; // @[Top.scala 778:22]
  wire [31:0] n106_O_2_0_1; // @[Top.scala 778:22]
  wire [31:0] n106_O_2_0_2; // @[Top.scala 778:22]
  wire [31:0] n106_O_2_1_0; // @[Top.scala 778:22]
  wire [31:0] n106_O_2_1_1; // @[Top.scala 778:22]
  wire [31:0] n106_O_2_1_2; // @[Top.scala 778:22]
  wire [31:0] n106_O_2_2_0; // @[Top.scala 778:22]
  wire [31:0] n106_O_2_2_1; // @[Top.scala 778:22]
  wire [31:0] n106_O_2_2_2; // @[Top.scala 778:22]
  wire [31:0] n106_O_3_0_0; // @[Top.scala 778:22]
  wire [31:0] n106_O_3_0_1; // @[Top.scala 778:22]
  wire [31:0] n106_O_3_0_2; // @[Top.scala 778:22]
  wire [31:0] n106_O_3_1_0; // @[Top.scala 778:22]
  wire [31:0] n106_O_3_1_1; // @[Top.scala 778:22]
  wire [31:0] n106_O_3_1_2; // @[Top.scala 778:22]
  wire [31:0] n106_O_3_2_0; // @[Top.scala 778:22]
  wire [31:0] n106_O_3_2_1; // @[Top.scala 778:22]
  wire [31:0] n106_O_3_2_2; // @[Top.scala 778:22]
  wire [31:0] n106_O_4_0_0; // @[Top.scala 778:22]
  wire [31:0] n106_O_4_0_1; // @[Top.scala 778:22]
  wire [31:0] n106_O_4_0_2; // @[Top.scala 778:22]
  wire [31:0] n106_O_4_1_0; // @[Top.scala 778:22]
  wire [31:0] n106_O_4_1_1; // @[Top.scala 778:22]
  wire [31:0] n106_O_4_1_2; // @[Top.scala 778:22]
  wire [31:0] n106_O_4_2_0; // @[Top.scala 778:22]
  wire [31:0] n106_O_4_2_1; // @[Top.scala 778:22]
  wire [31:0] n106_O_4_2_2; // @[Top.scala 778:22]
  wire [31:0] n106_O_5_0_0; // @[Top.scala 778:22]
  wire [31:0] n106_O_5_0_1; // @[Top.scala 778:22]
  wire [31:0] n106_O_5_0_2; // @[Top.scala 778:22]
  wire [31:0] n106_O_5_1_0; // @[Top.scala 778:22]
  wire [31:0] n106_O_5_1_1; // @[Top.scala 778:22]
  wire [31:0] n106_O_5_1_2; // @[Top.scala 778:22]
  wire [31:0] n106_O_5_2_0; // @[Top.scala 778:22]
  wire [31:0] n106_O_5_2_1; // @[Top.scala 778:22]
  wire [31:0] n106_O_5_2_2; // @[Top.scala 778:22]
  wire [31:0] n106_O_6_0_0; // @[Top.scala 778:22]
  wire [31:0] n106_O_6_0_1; // @[Top.scala 778:22]
  wire [31:0] n106_O_6_0_2; // @[Top.scala 778:22]
  wire [31:0] n106_O_6_1_0; // @[Top.scala 778:22]
  wire [31:0] n106_O_6_1_1; // @[Top.scala 778:22]
  wire [31:0] n106_O_6_1_2; // @[Top.scala 778:22]
  wire [31:0] n106_O_6_2_0; // @[Top.scala 778:22]
  wire [31:0] n106_O_6_2_1; // @[Top.scala 778:22]
  wire [31:0] n106_O_6_2_2; // @[Top.scala 778:22]
  wire [31:0] n106_O_7_0_0; // @[Top.scala 778:22]
  wire [31:0] n106_O_7_0_1; // @[Top.scala 778:22]
  wire [31:0] n106_O_7_0_2; // @[Top.scala 778:22]
  wire [31:0] n106_O_7_1_0; // @[Top.scala 778:22]
  wire [31:0] n106_O_7_1_1; // @[Top.scala 778:22]
  wire [31:0] n106_O_7_1_2; // @[Top.scala 778:22]
  wire [31:0] n106_O_7_2_0; // @[Top.scala 778:22]
  wire [31:0] n106_O_7_2_1; // @[Top.scala 778:22]
  wire [31:0] n106_O_7_2_2; // @[Top.scala 778:22]
  wire  n443_clock; // @[Top.scala 781:22]
  wire  n443_reset; // @[Top.scala 781:22]
  wire  n443_valid_up; // @[Top.scala 781:22]
  wire  n443_valid_down; // @[Top.scala 781:22]
  wire [31:0] n443_I_0_0_0; // @[Top.scala 781:22]
  wire [31:0] n443_I_0_0_1; // @[Top.scala 781:22]
  wire [31:0] n443_I_0_0_2; // @[Top.scala 781:22]
  wire [31:0] n443_I_0_1_0; // @[Top.scala 781:22]
  wire [31:0] n443_I_0_1_1; // @[Top.scala 781:22]
  wire [31:0] n443_I_0_1_2; // @[Top.scala 781:22]
  wire [31:0] n443_I_0_2_0; // @[Top.scala 781:22]
  wire [31:0] n443_I_0_2_1; // @[Top.scala 781:22]
  wire [31:0] n443_I_0_2_2; // @[Top.scala 781:22]
  wire [31:0] n443_I_1_0_0; // @[Top.scala 781:22]
  wire [31:0] n443_I_1_0_1; // @[Top.scala 781:22]
  wire [31:0] n443_I_1_0_2; // @[Top.scala 781:22]
  wire [31:0] n443_I_1_1_0; // @[Top.scala 781:22]
  wire [31:0] n443_I_1_1_1; // @[Top.scala 781:22]
  wire [31:0] n443_I_1_1_2; // @[Top.scala 781:22]
  wire [31:0] n443_I_1_2_0; // @[Top.scala 781:22]
  wire [31:0] n443_I_1_2_1; // @[Top.scala 781:22]
  wire [31:0] n443_I_1_2_2; // @[Top.scala 781:22]
  wire [31:0] n443_I_2_0_0; // @[Top.scala 781:22]
  wire [31:0] n443_I_2_0_1; // @[Top.scala 781:22]
  wire [31:0] n443_I_2_0_2; // @[Top.scala 781:22]
  wire [31:0] n443_I_2_1_0; // @[Top.scala 781:22]
  wire [31:0] n443_I_2_1_1; // @[Top.scala 781:22]
  wire [31:0] n443_I_2_1_2; // @[Top.scala 781:22]
  wire [31:0] n443_I_2_2_0; // @[Top.scala 781:22]
  wire [31:0] n443_I_2_2_1; // @[Top.scala 781:22]
  wire [31:0] n443_I_2_2_2; // @[Top.scala 781:22]
  wire [31:0] n443_I_3_0_0; // @[Top.scala 781:22]
  wire [31:0] n443_I_3_0_1; // @[Top.scala 781:22]
  wire [31:0] n443_I_3_0_2; // @[Top.scala 781:22]
  wire [31:0] n443_I_3_1_0; // @[Top.scala 781:22]
  wire [31:0] n443_I_3_1_1; // @[Top.scala 781:22]
  wire [31:0] n443_I_3_1_2; // @[Top.scala 781:22]
  wire [31:0] n443_I_3_2_0; // @[Top.scala 781:22]
  wire [31:0] n443_I_3_2_1; // @[Top.scala 781:22]
  wire [31:0] n443_I_3_2_2; // @[Top.scala 781:22]
  wire [31:0] n443_I_4_0_0; // @[Top.scala 781:22]
  wire [31:0] n443_I_4_0_1; // @[Top.scala 781:22]
  wire [31:0] n443_I_4_0_2; // @[Top.scala 781:22]
  wire [31:0] n443_I_4_1_0; // @[Top.scala 781:22]
  wire [31:0] n443_I_4_1_1; // @[Top.scala 781:22]
  wire [31:0] n443_I_4_1_2; // @[Top.scala 781:22]
  wire [31:0] n443_I_4_2_0; // @[Top.scala 781:22]
  wire [31:0] n443_I_4_2_1; // @[Top.scala 781:22]
  wire [31:0] n443_I_4_2_2; // @[Top.scala 781:22]
  wire [31:0] n443_I_5_0_0; // @[Top.scala 781:22]
  wire [31:0] n443_I_5_0_1; // @[Top.scala 781:22]
  wire [31:0] n443_I_5_0_2; // @[Top.scala 781:22]
  wire [31:0] n443_I_5_1_0; // @[Top.scala 781:22]
  wire [31:0] n443_I_5_1_1; // @[Top.scala 781:22]
  wire [31:0] n443_I_5_1_2; // @[Top.scala 781:22]
  wire [31:0] n443_I_5_2_0; // @[Top.scala 781:22]
  wire [31:0] n443_I_5_2_1; // @[Top.scala 781:22]
  wire [31:0] n443_I_5_2_2; // @[Top.scala 781:22]
  wire [31:0] n443_I_6_0_0; // @[Top.scala 781:22]
  wire [31:0] n443_I_6_0_1; // @[Top.scala 781:22]
  wire [31:0] n443_I_6_0_2; // @[Top.scala 781:22]
  wire [31:0] n443_I_6_1_0; // @[Top.scala 781:22]
  wire [31:0] n443_I_6_1_1; // @[Top.scala 781:22]
  wire [31:0] n443_I_6_1_2; // @[Top.scala 781:22]
  wire [31:0] n443_I_6_2_0; // @[Top.scala 781:22]
  wire [31:0] n443_I_6_2_1; // @[Top.scala 781:22]
  wire [31:0] n443_I_6_2_2; // @[Top.scala 781:22]
  wire [31:0] n443_I_7_0_0; // @[Top.scala 781:22]
  wire [31:0] n443_I_7_0_1; // @[Top.scala 781:22]
  wire [31:0] n443_I_7_0_2; // @[Top.scala 781:22]
  wire [31:0] n443_I_7_1_0; // @[Top.scala 781:22]
  wire [31:0] n443_I_7_1_1; // @[Top.scala 781:22]
  wire [31:0] n443_I_7_1_2; // @[Top.scala 781:22]
  wire [31:0] n443_I_7_2_0; // @[Top.scala 781:22]
  wire [31:0] n443_I_7_2_1; // @[Top.scala 781:22]
  wire [31:0] n443_I_7_2_2; // @[Top.scala 781:22]
  wire [31:0] n443_O_0_0_0_t0b; // @[Top.scala 781:22]
  wire [31:0] n443_O_0_0_0_t1b_t0b; // @[Top.scala 781:22]
  wire [31:0] n443_O_0_0_0_t1b_t1b; // @[Top.scala 781:22]
  wire [31:0] n443_O_1_0_0_t0b; // @[Top.scala 781:22]
  wire [31:0] n443_O_1_0_0_t1b_t0b; // @[Top.scala 781:22]
  wire [31:0] n443_O_1_0_0_t1b_t1b; // @[Top.scala 781:22]
  wire [31:0] n443_O_2_0_0_t0b; // @[Top.scala 781:22]
  wire [31:0] n443_O_2_0_0_t1b_t0b; // @[Top.scala 781:22]
  wire [31:0] n443_O_2_0_0_t1b_t1b; // @[Top.scala 781:22]
  wire [31:0] n443_O_3_0_0_t0b; // @[Top.scala 781:22]
  wire [31:0] n443_O_3_0_0_t1b_t0b; // @[Top.scala 781:22]
  wire [31:0] n443_O_3_0_0_t1b_t1b; // @[Top.scala 781:22]
  wire [31:0] n443_O_4_0_0_t0b; // @[Top.scala 781:22]
  wire [31:0] n443_O_4_0_0_t1b_t0b; // @[Top.scala 781:22]
  wire [31:0] n443_O_4_0_0_t1b_t1b; // @[Top.scala 781:22]
  wire [31:0] n443_O_5_0_0_t0b; // @[Top.scala 781:22]
  wire [31:0] n443_O_5_0_0_t1b_t0b; // @[Top.scala 781:22]
  wire [31:0] n443_O_5_0_0_t1b_t1b; // @[Top.scala 781:22]
  wire [31:0] n443_O_6_0_0_t0b; // @[Top.scala 781:22]
  wire [31:0] n443_O_6_0_0_t1b_t0b; // @[Top.scala 781:22]
  wire [31:0] n443_O_6_0_0_t1b_t1b; // @[Top.scala 781:22]
  wire [31:0] n443_O_7_0_0_t0b; // @[Top.scala 781:22]
  wire [31:0] n443_O_7_0_0_t1b_t0b; // @[Top.scala 781:22]
  wire [31:0] n443_O_7_0_0_t1b_t1b; // @[Top.scala 781:22]
  wire  n444_valid_up; // @[Top.scala 784:22]
  wire  n444_valid_down; // @[Top.scala 784:22]
  wire [31:0] n444_I_0_0_0_t0b; // @[Top.scala 784:22]
  wire [31:0] n444_I_0_0_0_t1b_t0b; // @[Top.scala 784:22]
  wire [31:0] n444_I_0_0_0_t1b_t1b; // @[Top.scala 784:22]
  wire [31:0] n444_I_1_0_0_t0b; // @[Top.scala 784:22]
  wire [31:0] n444_I_1_0_0_t1b_t0b; // @[Top.scala 784:22]
  wire [31:0] n444_I_1_0_0_t1b_t1b; // @[Top.scala 784:22]
  wire [31:0] n444_I_2_0_0_t0b; // @[Top.scala 784:22]
  wire [31:0] n444_I_2_0_0_t1b_t0b; // @[Top.scala 784:22]
  wire [31:0] n444_I_2_0_0_t1b_t1b; // @[Top.scala 784:22]
  wire [31:0] n444_I_3_0_0_t0b; // @[Top.scala 784:22]
  wire [31:0] n444_I_3_0_0_t1b_t0b; // @[Top.scala 784:22]
  wire [31:0] n444_I_3_0_0_t1b_t1b; // @[Top.scala 784:22]
  wire [31:0] n444_I_4_0_0_t0b; // @[Top.scala 784:22]
  wire [31:0] n444_I_4_0_0_t1b_t0b; // @[Top.scala 784:22]
  wire [31:0] n444_I_4_0_0_t1b_t1b; // @[Top.scala 784:22]
  wire [31:0] n444_I_5_0_0_t0b; // @[Top.scala 784:22]
  wire [31:0] n444_I_5_0_0_t1b_t0b; // @[Top.scala 784:22]
  wire [31:0] n444_I_5_0_0_t1b_t1b; // @[Top.scala 784:22]
  wire [31:0] n444_I_6_0_0_t0b; // @[Top.scala 784:22]
  wire [31:0] n444_I_6_0_0_t1b_t0b; // @[Top.scala 784:22]
  wire [31:0] n444_I_6_0_0_t1b_t1b; // @[Top.scala 784:22]
  wire [31:0] n444_I_7_0_0_t0b; // @[Top.scala 784:22]
  wire [31:0] n444_I_7_0_0_t1b_t0b; // @[Top.scala 784:22]
  wire [31:0] n444_I_7_0_0_t1b_t1b; // @[Top.scala 784:22]
  wire [31:0] n444_O_0_0_0_t0b; // @[Top.scala 784:22]
  wire [31:0] n444_O_0_0_0_t1b_t0b; // @[Top.scala 784:22]
  wire [31:0] n444_O_0_0_0_t1b_t1b; // @[Top.scala 784:22]
  wire [31:0] n444_O_1_0_0_t0b; // @[Top.scala 784:22]
  wire [31:0] n444_O_1_0_0_t1b_t0b; // @[Top.scala 784:22]
  wire [31:0] n444_O_1_0_0_t1b_t1b; // @[Top.scala 784:22]
  wire [31:0] n444_O_2_0_0_t0b; // @[Top.scala 784:22]
  wire [31:0] n444_O_2_0_0_t1b_t0b; // @[Top.scala 784:22]
  wire [31:0] n444_O_2_0_0_t1b_t1b; // @[Top.scala 784:22]
  wire [31:0] n444_O_3_0_0_t0b; // @[Top.scala 784:22]
  wire [31:0] n444_O_3_0_0_t1b_t0b; // @[Top.scala 784:22]
  wire [31:0] n444_O_3_0_0_t1b_t1b; // @[Top.scala 784:22]
  wire [31:0] n444_O_4_0_0_t0b; // @[Top.scala 784:22]
  wire [31:0] n444_O_4_0_0_t1b_t0b; // @[Top.scala 784:22]
  wire [31:0] n444_O_4_0_0_t1b_t1b; // @[Top.scala 784:22]
  wire [31:0] n444_O_5_0_0_t0b; // @[Top.scala 784:22]
  wire [31:0] n444_O_5_0_0_t1b_t0b; // @[Top.scala 784:22]
  wire [31:0] n444_O_5_0_0_t1b_t1b; // @[Top.scala 784:22]
  wire [31:0] n444_O_6_0_0_t0b; // @[Top.scala 784:22]
  wire [31:0] n444_O_6_0_0_t1b_t0b; // @[Top.scala 784:22]
  wire [31:0] n444_O_6_0_0_t1b_t1b; // @[Top.scala 784:22]
  wire [31:0] n444_O_7_0_0_t0b; // @[Top.scala 784:22]
  wire [31:0] n444_O_7_0_0_t1b_t0b; // @[Top.scala 784:22]
  wire [31:0] n444_O_7_0_0_t1b_t1b; // @[Top.scala 784:22]
  wire  n445_valid_up; // @[Top.scala 787:22]
  wire  n445_valid_down; // @[Top.scala 787:22]
  wire [31:0] n445_I_0_0_0_t0b; // @[Top.scala 787:22]
  wire [31:0] n445_I_0_0_0_t1b_t0b; // @[Top.scala 787:22]
  wire [31:0] n445_I_0_0_0_t1b_t1b; // @[Top.scala 787:22]
  wire [31:0] n445_I_1_0_0_t0b; // @[Top.scala 787:22]
  wire [31:0] n445_I_1_0_0_t1b_t0b; // @[Top.scala 787:22]
  wire [31:0] n445_I_1_0_0_t1b_t1b; // @[Top.scala 787:22]
  wire [31:0] n445_I_2_0_0_t0b; // @[Top.scala 787:22]
  wire [31:0] n445_I_2_0_0_t1b_t0b; // @[Top.scala 787:22]
  wire [31:0] n445_I_2_0_0_t1b_t1b; // @[Top.scala 787:22]
  wire [31:0] n445_I_3_0_0_t0b; // @[Top.scala 787:22]
  wire [31:0] n445_I_3_0_0_t1b_t0b; // @[Top.scala 787:22]
  wire [31:0] n445_I_3_0_0_t1b_t1b; // @[Top.scala 787:22]
  wire [31:0] n445_I_4_0_0_t0b; // @[Top.scala 787:22]
  wire [31:0] n445_I_4_0_0_t1b_t0b; // @[Top.scala 787:22]
  wire [31:0] n445_I_4_0_0_t1b_t1b; // @[Top.scala 787:22]
  wire [31:0] n445_I_5_0_0_t0b; // @[Top.scala 787:22]
  wire [31:0] n445_I_5_0_0_t1b_t0b; // @[Top.scala 787:22]
  wire [31:0] n445_I_5_0_0_t1b_t1b; // @[Top.scala 787:22]
  wire [31:0] n445_I_6_0_0_t0b; // @[Top.scala 787:22]
  wire [31:0] n445_I_6_0_0_t1b_t0b; // @[Top.scala 787:22]
  wire [31:0] n445_I_6_0_0_t1b_t1b; // @[Top.scala 787:22]
  wire [31:0] n445_I_7_0_0_t0b; // @[Top.scala 787:22]
  wire [31:0] n445_I_7_0_0_t1b_t0b; // @[Top.scala 787:22]
  wire [31:0] n445_I_7_0_0_t1b_t1b; // @[Top.scala 787:22]
  wire [31:0] n445_O_0_0_t0b; // @[Top.scala 787:22]
  wire [31:0] n445_O_0_0_t1b_t0b; // @[Top.scala 787:22]
  wire [31:0] n445_O_0_0_t1b_t1b; // @[Top.scala 787:22]
  wire [31:0] n445_O_1_0_t0b; // @[Top.scala 787:22]
  wire [31:0] n445_O_1_0_t1b_t0b; // @[Top.scala 787:22]
  wire [31:0] n445_O_1_0_t1b_t1b; // @[Top.scala 787:22]
  wire [31:0] n445_O_2_0_t0b; // @[Top.scala 787:22]
  wire [31:0] n445_O_2_0_t1b_t0b; // @[Top.scala 787:22]
  wire [31:0] n445_O_2_0_t1b_t1b; // @[Top.scala 787:22]
  wire [31:0] n445_O_3_0_t0b; // @[Top.scala 787:22]
  wire [31:0] n445_O_3_0_t1b_t0b; // @[Top.scala 787:22]
  wire [31:0] n445_O_3_0_t1b_t1b; // @[Top.scala 787:22]
  wire [31:0] n445_O_4_0_t0b; // @[Top.scala 787:22]
  wire [31:0] n445_O_4_0_t1b_t0b; // @[Top.scala 787:22]
  wire [31:0] n445_O_4_0_t1b_t1b; // @[Top.scala 787:22]
  wire [31:0] n445_O_5_0_t0b; // @[Top.scala 787:22]
  wire [31:0] n445_O_5_0_t1b_t0b; // @[Top.scala 787:22]
  wire [31:0] n445_O_5_0_t1b_t1b; // @[Top.scala 787:22]
  wire [31:0] n445_O_6_0_t0b; // @[Top.scala 787:22]
  wire [31:0] n445_O_6_0_t1b_t0b; // @[Top.scala 787:22]
  wire [31:0] n445_O_6_0_t1b_t1b; // @[Top.scala 787:22]
  wire [31:0] n445_O_7_0_t0b; // @[Top.scala 787:22]
  wire [31:0] n445_O_7_0_t1b_t0b; // @[Top.scala 787:22]
  wire [31:0] n445_O_7_0_t1b_t1b; // @[Top.scala 787:22]
  wire  n446_valid_up; // @[Top.scala 790:22]
  wire  n446_valid_down; // @[Top.scala 790:22]
  wire [31:0] n446_I_0_0_t0b; // @[Top.scala 790:22]
  wire [31:0] n446_I_0_0_t1b_t0b; // @[Top.scala 790:22]
  wire [31:0] n446_I_0_0_t1b_t1b; // @[Top.scala 790:22]
  wire [31:0] n446_I_1_0_t0b; // @[Top.scala 790:22]
  wire [31:0] n446_I_1_0_t1b_t0b; // @[Top.scala 790:22]
  wire [31:0] n446_I_1_0_t1b_t1b; // @[Top.scala 790:22]
  wire [31:0] n446_I_2_0_t0b; // @[Top.scala 790:22]
  wire [31:0] n446_I_2_0_t1b_t0b; // @[Top.scala 790:22]
  wire [31:0] n446_I_2_0_t1b_t1b; // @[Top.scala 790:22]
  wire [31:0] n446_I_3_0_t0b; // @[Top.scala 790:22]
  wire [31:0] n446_I_3_0_t1b_t0b; // @[Top.scala 790:22]
  wire [31:0] n446_I_3_0_t1b_t1b; // @[Top.scala 790:22]
  wire [31:0] n446_I_4_0_t0b; // @[Top.scala 790:22]
  wire [31:0] n446_I_4_0_t1b_t0b; // @[Top.scala 790:22]
  wire [31:0] n446_I_4_0_t1b_t1b; // @[Top.scala 790:22]
  wire [31:0] n446_I_5_0_t0b; // @[Top.scala 790:22]
  wire [31:0] n446_I_5_0_t1b_t0b; // @[Top.scala 790:22]
  wire [31:0] n446_I_5_0_t1b_t1b; // @[Top.scala 790:22]
  wire [31:0] n446_I_6_0_t0b; // @[Top.scala 790:22]
  wire [31:0] n446_I_6_0_t1b_t0b; // @[Top.scala 790:22]
  wire [31:0] n446_I_6_0_t1b_t1b; // @[Top.scala 790:22]
  wire [31:0] n446_I_7_0_t0b; // @[Top.scala 790:22]
  wire [31:0] n446_I_7_0_t1b_t0b; // @[Top.scala 790:22]
  wire [31:0] n446_I_7_0_t1b_t1b; // @[Top.scala 790:22]
  wire [31:0] n446_O_0_t0b; // @[Top.scala 790:22]
  wire [31:0] n446_O_0_t1b_t0b; // @[Top.scala 790:22]
  wire [31:0] n446_O_0_t1b_t1b; // @[Top.scala 790:22]
  wire [31:0] n446_O_1_t0b; // @[Top.scala 790:22]
  wire [31:0] n446_O_1_t1b_t0b; // @[Top.scala 790:22]
  wire [31:0] n446_O_1_t1b_t1b; // @[Top.scala 790:22]
  wire [31:0] n446_O_2_t0b; // @[Top.scala 790:22]
  wire [31:0] n446_O_2_t1b_t0b; // @[Top.scala 790:22]
  wire [31:0] n446_O_2_t1b_t1b; // @[Top.scala 790:22]
  wire [31:0] n446_O_3_t0b; // @[Top.scala 790:22]
  wire [31:0] n446_O_3_t1b_t0b; // @[Top.scala 790:22]
  wire [31:0] n446_O_3_t1b_t1b; // @[Top.scala 790:22]
  wire [31:0] n446_O_4_t0b; // @[Top.scala 790:22]
  wire [31:0] n446_O_4_t1b_t0b; // @[Top.scala 790:22]
  wire [31:0] n446_O_4_t1b_t1b; // @[Top.scala 790:22]
  wire [31:0] n446_O_5_t0b; // @[Top.scala 790:22]
  wire [31:0] n446_O_5_t1b_t0b; // @[Top.scala 790:22]
  wire [31:0] n446_O_5_t1b_t1b; // @[Top.scala 790:22]
  wire [31:0] n446_O_6_t0b; // @[Top.scala 790:22]
  wire [31:0] n446_O_6_t1b_t0b; // @[Top.scala 790:22]
  wire [31:0] n446_O_6_t1b_t1b; // @[Top.scala 790:22]
  wire [31:0] n446_O_7_t0b; // @[Top.scala 790:22]
  wire [31:0] n446_O_7_t1b_t0b; // @[Top.scala 790:22]
  wire [31:0] n446_O_7_t1b_t1b; // @[Top.scala 790:22]
  wire  n451_valid_up; // @[Top.scala 793:22]
  wire  n451_valid_down; // @[Top.scala 793:22]
  wire [31:0] n451_I_0_t0b; // @[Top.scala 793:22]
  wire [31:0] n451_I_1_t0b; // @[Top.scala 793:22]
  wire [31:0] n451_I_2_t0b; // @[Top.scala 793:22]
  wire [31:0] n451_I_3_t0b; // @[Top.scala 793:22]
  wire [31:0] n451_I_4_t0b; // @[Top.scala 793:22]
  wire [31:0] n451_I_5_t0b; // @[Top.scala 793:22]
  wire [31:0] n451_I_6_t0b; // @[Top.scala 793:22]
  wire [31:0] n451_I_7_t0b; // @[Top.scala 793:22]
  wire [31:0] n451_O_0; // @[Top.scala 793:22]
  wire [31:0] n451_O_1; // @[Top.scala 793:22]
  wire [31:0] n451_O_2; // @[Top.scala 793:22]
  wire [31:0] n451_O_3; // @[Top.scala 793:22]
  wire [31:0] n451_O_4; // @[Top.scala 793:22]
  wire [31:0] n451_O_5; // @[Top.scala 793:22]
  wire [31:0] n451_O_6; // @[Top.scala 793:22]
  wire [31:0] n451_O_7; // @[Top.scala 793:22]
  wire  n452_clock; // @[Top.scala 796:22]
  wire  n452_reset; // @[Top.scala 796:22]
  wire  n452_valid_up; // @[Top.scala 796:22]
  wire  n452_valid_down; // @[Top.scala 796:22]
  wire [31:0] n452_I_0; // @[Top.scala 796:22]
  wire [31:0] n452_I_1; // @[Top.scala 796:22]
  wire [31:0] n452_I_2; // @[Top.scala 796:22]
  wire [31:0] n452_I_3; // @[Top.scala 796:22]
  wire [31:0] n452_I_4; // @[Top.scala 796:22]
  wire [31:0] n452_I_5; // @[Top.scala 796:22]
  wire [31:0] n452_I_6; // @[Top.scala 796:22]
  wire [31:0] n452_I_7; // @[Top.scala 796:22]
  wire [31:0] n452_O_0; // @[Top.scala 796:22]
  wire [31:0] n452_O_1; // @[Top.scala 796:22]
  wire [31:0] n452_O_2; // @[Top.scala 796:22]
  wire [31:0] n452_O_3; // @[Top.scala 796:22]
  wire [31:0] n452_O_4; // @[Top.scala 796:22]
  wire [31:0] n452_O_5; // @[Top.scala 796:22]
  wire [31:0] n452_O_6; // @[Top.scala 796:22]
  wire [31:0] n452_O_7; // @[Top.scala 796:22]
  wire  n453_clock; // @[Top.scala 799:22]
  wire  n453_reset; // @[Top.scala 799:22]
  wire  n453_valid_up; // @[Top.scala 799:22]
  wire  n453_valid_down; // @[Top.scala 799:22]
  wire [31:0] n453_I_0; // @[Top.scala 799:22]
  wire [31:0] n453_I_1; // @[Top.scala 799:22]
  wire [31:0] n453_I_2; // @[Top.scala 799:22]
  wire [31:0] n453_I_3; // @[Top.scala 799:22]
  wire [31:0] n453_I_4; // @[Top.scala 799:22]
  wire [31:0] n453_I_5; // @[Top.scala 799:22]
  wire [31:0] n453_I_6; // @[Top.scala 799:22]
  wire [31:0] n453_I_7; // @[Top.scala 799:22]
  wire [31:0] n453_O_0; // @[Top.scala 799:22]
  wire [31:0] n453_O_1; // @[Top.scala 799:22]
  wire [31:0] n453_O_2; // @[Top.scala 799:22]
  wire [31:0] n453_O_3; // @[Top.scala 799:22]
  wire [31:0] n453_O_4; // @[Top.scala 799:22]
  wire [31:0] n453_O_5; // @[Top.scala 799:22]
  wire [31:0] n453_O_6; // @[Top.scala 799:22]
  wire [31:0] n453_O_7; // @[Top.scala 799:22]
  wire  n454_clock; // @[Top.scala 802:22]
  wire  n454_valid_up; // @[Top.scala 802:22]
  wire  n454_valid_down; // @[Top.scala 802:22]
  wire [31:0] n454_I_0; // @[Top.scala 802:22]
  wire [31:0] n454_I_1; // @[Top.scala 802:22]
  wire [31:0] n454_I_2; // @[Top.scala 802:22]
  wire [31:0] n454_I_3; // @[Top.scala 802:22]
  wire [31:0] n454_I_4; // @[Top.scala 802:22]
  wire [31:0] n454_I_5; // @[Top.scala 802:22]
  wire [31:0] n454_I_6; // @[Top.scala 802:22]
  wire [31:0] n454_I_7; // @[Top.scala 802:22]
  wire [31:0] n454_O_0; // @[Top.scala 802:22]
  wire [31:0] n454_O_1; // @[Top.scala 802:22]
  wire [31:0] n454_O_2; // @[Top.scala 802:22]
  wire [31:0] n454_O_3; // @[Top.scala 802:22]
  wire [31:0] n454_O_4; // @[Top.scala 802:22]
  wire [31:0] n454_O_5; // @[Top.scala 802:22]
  wire [31:0] n454_O_6; // @[Top.scala 802:22]
  wire [31:0] n454_O_7; // @[Top.scala 802:22]
  wire  n455_clock; // @[Top.scala 805:22]
  wire  n455_valid_up; // @[Top.scala 805:22]
  wire  n455_valid_down; // @[Top.scala 805:22]
  wire [31:0] n455_I_0; // @[Top.scala 805:22]
  wire [31:0] n455_I_1; // @[Top.scala 805:22]
  wire [31:0] n455_I_2; // @[Top.scala 805:22]
  wire [31:0] n455_I_3; // @[Top.scala 805:22]
  wire [31:0] n455_I_4; // @[Top.scala 805:22]
  wire [31:0] n455_I_5; // @[Top.scala 805:22]
  wire [31:0] n455_I_6; // @[Top.scala 805:22]
  wire [31:0] n455_I_7; // @[Top.scala 805:22]
  wire [31:0] n455_O_0; // @[Top.scala 805:22]
  wire [31:0] n455_O_1; // @[Top.scala 805:22]
  wire [31:0] n455_O_2; // @[Top.scala 805:22]
  wire [31:0] n455_O_3; // @[Top.scala 805:22]
  wire [31:0] n455_O_4; // @[Top.scala 805:22]
  wire [31:0] n455_O_5; // @[Top.scala 805:22]
  wire [31:0] n455_O_6; // @[Top.scala 805:22]
  wire [31:0] n455_O_7; // @[Top.scala 805:22]
  wire  n456_valid_up; // @[Top.scala 808:22]
  wire  n456_valid_down; // @[Top.scala 808:22]
  wire [31:0] n456_I0_0; // @[Top.scala 808:22]
  wire [31:0] n456_I0_1; // @[Top.scala 808:22]
  wire [31:0] n456_I0_2; // @[Top.scala 808:22]
  wire [31:0] n456_I0_3; // @[Top.scala 808:22]
  wire [31:0] n456_I0_4; // @[Top.scala 808:22]
  wire [31:0] n456_I0_5; // @[Top.scala 808:22]
  wire [31:0] n456_I0_6; // @[Top.scala 808:22]
  wire [31:0] n456_I0_7; // @[Top.scala 808:22]
  wire [31:0] n456_I1_0; // @[Top.scala 808:22]
  wire [31:0] n456_I1_1; // @[Top.scala 808:22]
  wire [31:0] n456_I1_2; // @[Top.scala 808:22]
  wire [31:0] n456_I1_3; // @[Top.scala 808:22]
  wire [31:0] n456_I1_4; // @[Top.scala 808:22]
  wire [31:0] n456_I1_5; // @[Top.scala 808:22]
  wire [31:0] n456_I1_6; // @[Top.scala 808:22]
  wire [31:0] n456_I1_7; // @[Top.scala 808:22]
  wire [31:0] n456_O_0_0; // @[Top.scala 808:22]
  wire [31:0] n456_O_0_1; // @[Top.scala 808:22]
  wire [31:0] n456_O_1_0; // @[Top.scala 808:22]
  wire [31:0] n456_O_1_1; // @[Top.scala 808:22]
  wire [31:0] n456_O_2_0; // @[Top.scala 808:22]
  wire [31:0] n456_O_2_1; // @[Top.scala 808:22]
  wire [31:0] n456_O_3_0; // @[Top.scala 808:22]
  wire [31:0] n456_O_3_1; // @[Top.scala 808:22]
  wire [31:0] n456_O_4_0; // @[Top.scala 808:22]
  wire [31:0] n456_O_4_1; // @[Top.scala 808:22]
  wire [31:0] n456_O_5_0; // @[Top.scala 808:22]
  wire [31:0] n456_O_5_1; // @[Top.scala 808:22]
  wire [31:0] n456_O_6_0; // @[Top.scala 808:22]
  wire [31:0] n456_O_6_1; // @[Top.scala 808:22]
  wire [31:0] n456_O_7_0; // @[Top.scala 808:22]
  wire [31:0] n456_O_7_1; // @[Top.scala 808:22]
  wire  n463_valid_up; // @[Top.scala 812:22]
  wire  n463_valid_down; // @[Top.scala 812:22]
  wire [31:0] n463_I0_0_0; // @[Top.scala 812:22]
  wire [31:0] n463_I0_0_1; // @[Top.scala 812:22]
  wire [31:0] n463_I0_1_0; // @[Top.scala 812:22]
  wire [31:0] n463_I0_1_1; // @[Top.scala 812:22]
  wire [31:0] n463_I0_2_0; // @[Top.scala 812:22]
  wire [31:0] n463_I0_2_1; // @[Top.scala 812:22]
  wire [31:0] n463_I0_3_0; // @[Top.scala 812:22]
  wire [31:0] n463_I0_3_1; // @[Top.scala 812:22]
  wire [31:0] n463_I0_4_0; // @[Top.scala 812:22]
  wire [31:0] n463_I0_4_1; // @[Top.scala 812:22]
  wire [31:0] n463_I0_5_0; // @[Top.scala 812:22]
  wire [31:0] n463_I0_5_1; // @[Top.scala 812:22]
  wire [31:0] n463_I0_6_0; // @[Top.scala 812:22]
  wire [31:0] n463_I0_6_1; // @[Top.scala 812:22]
  wire [31:0] n463_I0_7_0; // @[Top.scala 812:22]
  wire [31:0] n463_I0_7_1; // @[Top.scala 812:22]
  wire [31:0] n463_I1_0; // @[Top.scala 812:22]
  wire [31:0] n463_I1_1; // @[Top.scala 812:22]
  wire [31:0] n463_I1_2; // @[Top.scala 812:22]
  wire [31:0] n463_I1_3; // @[Top.scala 812:22]
  wire [31:0] n463_I1_4; // @[Top.scala 812:22]
  wire [31:0] n463_I1_5; // @[Top.scala 812:22]
  wire [31:0] n463_I1_6; // @[Top.scala 812:22]
  wire [31:0] n463_I1_7; // @[Top.scala 812:22]
  wire [31:0] n463_O_0_0; // @[Top.scala 812:22]
  wire [31:0] n463_O_0_1; // @[Top.scala 812:22]
  wire [31:0] n463_O_0_2; // @[Top.scala 812:22]
  wire [31:0] n463_O_1_0; // @[Top.scala 812:22]
  wire [31:0] n463_O_1_1; // @[Top.scala 812:22]
  wire [31:0] n463_O_1_2; // @[Top.scala 812:22]
  wire [31:0] n463_O_2_0; // @[Top.scala 812:22]
  wire [31:0] n463_O_2_1; // @[Top.scala 812:22]
  wire [31:0] n463_O_2_2; // @[Top.scala 812:22]
  wire [31:0] n463_O_3_0; // @[Top.scala 812:22]
  wire [31:0] n463_O_3_1; // @[Top.scala 812:22]
  wire [31:0] n463_O_3_2; // @[Top.scala 812:22]
  wire [31:0] n463_O_4_0; // @[Top.scala 812:22]
  wire [31:0] n463_O_4_1; // @[Top.scala 812:22]
  wire [31:0] n463_O_4_2; // @[Top.scala 812:22]
  wire [31:0] n463_O_5_0; // @[Top.scala 812:22]
  wire [31:0] n463_O_5_1; // @[Top.scala 812:22]
  wire [31:0] n463_O_5_2; // @[Top.scala 812:22]
  wire [31:0] n463_O_6_0; // @[Top.scala 812:22]
  wire [31:0] n463_O_6_1; // @[Top.scala 812:22]
  wire [31:0] n463_O_6_2; // @[Top.scala 812:22]
  wire [31:0] n463_O_7_0; // @[Top.scala 812:22]
  wire [31:0] n463_O_7_1; // @[Top.scala 812:22]
  wire [31:0] n463_O_7_2; // @[Top.scala 812:22]
  wire  n472_valid_up; // @[Top.scala 816:22]
  wire  n472_valid_down; // @[Top.scala 816:22]
  wire [31:0] n472_I_0_0; // @[Top.scala 816:22]
  wire [31:0] n472_I_0_1; // @[Top.scala 816:22]
  wire [31:0] n472_I_0_2; // @[Top.scala 816:22]
  wire [31:0] n472_I_1_0; // @[Top.scala 816:22]
  wire [31:0] n472_I_1_1; // @[Top.scala 816:22]
  wire [31:0] n472_I_1_2; // @[Top.scala 816:22]
  wire [31:0] n472_I_2_0; // @[Top.scala 816:22]
  wire [31:0] n472_I_2_1; // @[Top.scala 816:22]
  wire [31:0] n472_I_2_2; // @[Top.scala 816:22]
  wire [31:0] n472_I_3_0; // @[Top.scala 816:22]
  wire [31:0] n472_I_3_1; // @[Top.scala 816:22]
  wire [31:0] n472_I_3_2; // @[Top.scala 816:22]
  wire [31:0] n472_I_4_0; // @[Top.scala 816:22]
  wire [31:0] n472_I_4_1; // @[Top.scala 816:22]
  wire [31:0] n472_I_4_2; // @[Top.scala 816:22]
  wire [31:0] n472_I_5_0; // @[Top.scala 816:22]
  wire [31:0] n472_I_5_1; // @[Top.scala 816:22]
  wire [31:0] n472_I_5_2; // @[Top.scala 816:22]
  wire [31:0] n472_I_6_0; // @[Top.scala 816:22]
  wire [31:0] n472_I_6_1; // @[Top.scala 816:22]
  wire [31:0] n472_I_6_2; // @[Top.scala 816:22]
  wire [31:0] n472_I_7_0; // @[Top.scala 816:22]
  wire [31:0] n472_I_7_1; // @[Top.scala 816:22]
  wire [31:0] n472_I_7_2; // @[Top.scala 816:22]
  wire [31:0] n472_O_0_0_0; // @[Top.scala 816:22]
  wire [31:0] n472_O_0_0_1; // @[Top.scala 816:22]
  wire [31:0] n472_O_0_0_2; // @[Top.scala 816:22]
  wire [31:0] n472_O_1_0_0; // @[Top.scala 816:22]
  wire [31:0] n472_O_1_0_1; // @[Top.scala 816:22]
  wire [31:0] n472_O_1_0_2; // @[Top.scala 816:22]
  wire [31:0] n472_O_2_0_0; // @[Top.scala 816:22]
  wire [31:0] n472_O_2_0_1; // @[Top.scala 816:22]
  wire [31:0] n472_O_2_0_2; // @[Top.scala 816:22]
  wire [31:0] n472_O_3_0_0; // @[Top.scala 816:22]
  wire [31:0] n472_O_3_0_1; // @[Top.scala 816:22]
  wire [31:0] n472_O_3_0_2; // @[Top.scala 816:22]
  wire [31:0] n472_O_4_0_0; // @[Top.scala 816:22]
  wire [31:0] n472_O_4_0_1; // @[Top.scala 816:22]
  wire [31:0] n472_O_4_0_2; // @[Top.scala 816:22]
  wire [31:0] n472_O_5_0_0; // @[Top.scala 816:22]
  wire [31:0] n472_O_5_0_1; // @[Top.scala 816:22]
  wire [31:0] n472_O_5_0_2; // @[Top.scala 816:22]
  wire [31:0] n472_O_6_0_0; // @[Top.scala 816:22]
  wire [31:0] n472_O_6_0_1; // @[Top.scala 816:22]
  wire [31:0] n472_O_6_0_2; // @[Top.scala 816:22]
  wire [31:0] n472_O_7_0_0; // @[Top.scala 816:22]
  wire [31:0] n472_O_7_0_1; // @[Top.scala 816:22]
  wire [31:0] n472_O_7_0_2; // @[Top.scala 816:22]
  wire  n479_valid_up; // @[Top.scala 819:22]
  wire  n479_valid_down; // @[Top.scala 819:22]
  wire [31:0] n479_I_0_0_0; // @[Top.scala 819:22]
  wire [31:0] n479_I_0_0_1; // @[Top.scala 819:22]
  wire [31:0] n479_I_0_0_2; // @[Top.scala 819:22]
  wire [31:0] n479_I_1_0_0; // @[Top.scala 819:22]
  wire [31:0] n479_I_1_0_1; // @[Top.scala 819:22]
  wire [31:0] n479_I_1_0_2; // @[Top.scala 819:22]
  wire [31:0] n479_I_2_0_0; // @[Top.scala 819:22]
  wire [31:0] n479_I_2_0_1; // @[Top.scala 819:22]
  wire [31:0] n479_I_2_0_2; // @[Top.scala 819:22]
  wire [31:0] n479_I_3_0_0; // @[Top.scala 819:22]
  wire [31:0] n479_I_3_0_1; // @[Top.scala 819:22]
  wire [31:0] n479_I_3_0_2; // @[Top.scala 819:22]
  wire [31:0] n479_I_4_0_0; // @[Top.scala 819:22]
  wire [31:0] n479_I_4_0_1; // @[Top.scala 819:22]
  wire [31:0] n479_I_4_0_2; // @[Top.scala 819:22]
  wire [31:0] n479_I_5_0_0; // @[Top.scala 819:22]
  wire [31:0] n479_I_5_0_1; // @[Top.scala 819:22]
  wire [31:0] n479_I_5_0_2; // @[Top.scala 819:22]
  wire [31:0] n479_I_6_0_0; // @[Top.scala 819:22]
  wire [31:0] n479_I_6_0_1; // @[Top.scala 819:22]
  wire [31:0] n479_I_6_0_2; // @[Top.scala 819:22]
  wire [31:0] n479_I_7_0_0; // @[Top.scala 819:22]
  wire [31:0] n479_I_7_0_1; // @[Top.scala 819:22]
  wire [31:0] n479_I_7_0_2; // @[Top.scala 819:22]
  wire [31:0] n479_O_0_0; // @[Top.scala 819:22]
  wire [31:0] n479_O_0_1; // @[Top.scala 819:22]
  wire [31:0] n479_O_0_2; // @[Top.scala 819:22]
  wire [31:0] n479_O_1_0; // @[Top.scala 819:22]
  wire [31:0] n479_O_1_1; // @[Top.scala 819:22]
  wire [31:0] n479_O_1_2; // @[Top.scala 819:22]
  wire [31:0] n479_O_2_0; // @[Top.scala 819:22]
  wire [31:0] n479_O_2_1; // @[Top.scala 819:22]
  wire [31:0] n479_O_2_2; // @[Top.scala 819:22]
  wire [31:0] n479_O_3_0; // @[Top.scala 819:22]
  wire [31:0] n479_O_3_1; // @[Top.scala 819:22]
  wire [31:0] n479_O_3_2; // @[Top.scala 819:22]
  wire [31:0] n479_O_4_0; // @[Top.scala 819:22]
  wire [31:0] n479_O_4_1; // @[Top.scala 819:22]
  wire [31:0] n479_O_4_2; // @[Top.scala 819:22]
  wire [31:0] n479_O_5_0; // @[Top.scala 819:22]
  wire [31:0] n479_O_5_1; // @[Top.scala 819:22]
  wire [31:0] n479_O_5_2; // @[Top.scala 819:22]
  wire [31:0] n479_O_6_0; // @[Top.scala 819:22]
  wire [31:0] n479_O_6_1; // @[Top.scala 819:22]
  wire [31:0] n479_O_6_2; // @[Top.scala 819:22]
  wire [31:0] n479_O_7_0; // @[Top.scala 819:22]
  wire [31:0] n479_O_7_1; // @[Top.scala 819:22]
  wire [31:0] n479_O_7_2; // @[Top.scala 819:22]
  wire  n480_clock; // @[Top.scala 822:22]
  wire  n480_valid_up; // @[Top.scala 822:22]
  wire  n480_valid_down; // @[Top.scala 822:22]
  wire [31:0] n480_I_0; // @[Top.scala 822:22]
  wire [31:0] n480_I_1; // @[Top.scala 822:22]
  wire [31:0] n480_I_2; // @[Top.scala 822:22]
  wire [31:0] n480_I_3; // @[Top.scala 822:22]
  wire [31:0] n480_I_4; // @[Top.scala 822:22]
  wire [31:0] n480_I_5; // @[Top.scala 822:22]
  wire [31:0] n480_I_6; // @[Top.scala 822:22]
  wire [31:0] n480_I_7; // @[Top.scala 822:22]
  wire [31:0] n480_O_0; // @[Top.scala 822:22]
  wire [31:0] n480_O_1; // @[Top.scala 822:22]
  wire [31:0] n480_O_2; // @[Top.scala 822:22]
  wire [31:0] n480_O_3; // @[Top.scala 822:22]
  wire [31:0] n480_O_4; // @[Top.scala 822:22]
  wire [31:0] n480_O_5; // @[Top.scala 822:22]
  wire [31:0] n480_O_6; // @[Top.scala 822:22]
  wire [31:0] n480_O_7; // @[Top.scala 822:22]
  wire  n481_clock; // @[Top.scala 825:22]
  wire  n481_valid_up; // @[Top.scala 825:22]
  wire  n481_valid_down; // @[Top.scala 825:22]
  wire [31:0] n481_I_0; // @[Top.scala 825:22]
  wire [31:0] n481_I_1; // @[Top.scala 825:22]
  wire [31:0] n481_I_2; // @[Top.scala 825:22]
  wire [31:0] n481_I_3; // @[Top.scala 825:22]
  wire [31:0] n481_I_4; // @[Top.scala 825:22]
  wire [31:0] n481_I_5; // @[Top.scala 825:22]
  wire [31:0] n481_I_6; // @[Top.scala 825:22]
  wire [31:0] n481_I_7; // @[Top.scala 825:22]
  wire [31:0] n481_O_0; // @[Top.scala 825:22]
  wire [31:0] n481_O_1; // @[Top.scala 825:22]
  wire [31:0] n481_O_2; // @[Top.scala 825:22]
  wire [31:0] n481_O_3; // @[Top.scala 825:22]
  wire [31:0] n481_O_4; // @[Top.scala 825:22]
  wire [31:0] n481_O_5; // @[Top.scala 825:22]
  wire [31:0] n481_O_6; // @[Top.scala 825:22]
  wire [31:0] n481_O_7; // @[Top.scala 825:22]
  wire  n482_valid_up; // @[Top.scala 828:22]
  wire  n482_valid_down; // @[Top.scala 828:22]
  wire [31:0] n482_I0_0; // @[Top.scala 828:22]
  wire [31:0] n482_I0_1; // @[Top.scala 828:22]
  wire [31:0] n482_I0_2; // @[Top.scala 828:22]
  wire [31:0] n482_I0_3; // @[Top.scala 828:22]
  wire [31:0] n482_I0_4; // @[Top.scala 828:22]
  wire [31:0] n482_I0_5; // @[Top.scala 828:22]
  wire [31:0] n482_I0_6; // @[Top.scala 828:22]
  wire [31:0] n482_I0_7; // @[Top.scala 828:22]
  wire [31:0] n482_I1_0; // @[Top.scala 828:22]
  wire [31:0] n482_I1_1; // @[Top.scala 828:22]
  wire [31:0] n482_I1_2; // @[Top.scala 828:22]
  wire [31:0] n482_I1_3; // @[Top.scala 828:22]
  wire [31:0] n482_I1_4; // @[Top.scala 828:22]
  wire [31:0] n482_I1_5; // @[Top.scala 828:22]
  wire [31:0] n482_I1_6; // @[Top.scala 828:22]
  wire [31:0] n482_I1_7; // @[Top.scala 828:22]
  wire [31:0] n482_O_0_0; // @[Top.scala 828:22]
  wire [31:0] n482_O_0_1; // @[Top.scala 828:22]
  wire [31:0] n482_O_1_0; // @[Top.scala 828:22]
  wire [31:0] n482_O_1_1; // @[Top.scala 828:22]
  wire [31:0] n482_O_2_0; // @[Top.scala 828:22]
  wire [31:0] n482_O_2_1; // @[Top.scala 828:22]
  wire [31:0] n482_O_3_0; // @[Top.scala 828:22]
  wire [31:0] n482_O_3_1; // @[Top.scala 828:22]
  wire [31:0] n482_O_4_0; // @[Top.scala 828:22]
  wire [31:0] n482_O_4_1; // @[Top.scala 828:22]
  wire [31:0] n482_O_5_0; // @[Top.scala 828:22]
  wire [31:0] n482_O_5_1; // @[Top.scala 828:22]
  wire [31:0] n482_O_6_0; // @[Top.scala 828:22]
  wire [31:0] n482_O_6_1; // @[Top.scala 828:22]
  wire [31:0] n482_O_7_0; // @[Top.scala 828:22]
  wire [31:0] n482_O_7_1; // @[Top.scala 828:22]
  wire  n489_valid_up; // @[Top.scala 832:22]
  wire  n489_valid_down; // @[Top.scala 832:22]
  wire [31:0] n489_I0_0_0; // @[Top.scala 832:22]
  wire [31:0] n489_I0_0_1; // @[Top.scala 832:22]
  wire [31:0] n489_I0_1_0; // @[Top.scala 832:22]
  wire [31:0] n489_I0_1_1; // @[Top.scala 832:22]
  wire [31:0] n489_I0_2_0; // @[Top.scala 832:22]
  wire [31:0] n489_I0_2_1; // @[Top.scala 832:22]
  wire [31:0] n489_I0_3_0; // @[Top.scala 832:22]
  wire [31:0] n489_I0_3_1; // @[Top.scala 832:22]
  wire [31:0] n489_I0_4_0; // @[Top.scala 832:22]
  wire [31:0] n489_I0_4_1; // @[Top.scala 832:22]
  wire [31:0] n489_I0_5_0; // @[Top.scala 832:22]
  wire [31:0] n489_I0_5_1; // @[Top.scala 832:22]
  wire [31:0] n489_I0_6_0; // @[Top.scala 832:22]
  wire [31:0] n489_I0_6_1; // @[Top.scala 832:22]
  wire [31:0] n489_I0_7_0; // @[Top.scala 832:22]
  wire [31:0] n489_I0_7_1; // @[Top.scala 832:22]
  wire [31:0] n489_I1_0; // @[Top.scala 832:22]
  wire [31:0] n489_I1_1; // @[Top.scala 832:22]
  wire [31:0] n489_I1_2; // @[Top.scala 832:22]
  wire [31:0] n489_I1_3; // @[Top.scala 832:22]
  wire [31:0] n489_I1_4; // @[Top.scala 832:22]
  wire [31:0] n489_I1_5; // @[Top.scala 832:22]
  wire [31:0] n489_I1_6; // @[Top.scala 832:22]
  wire [31:0] n489_I1_7; // @[Top.scala 832:22]
  wire [31:0] n489_O_0_0; // @[Top.scala 832:22]
  wire [31:0] n489_O_0_1; // @[Top.scala 832:22]
  wire [31:0] n489_O_0_2; // @[Top.scala 832:22]
  wire [31:0] n489_O_1_0; // @[Top.scala 832:22]
  wire [31:0] n489_O_1_1; // @[Top.scala 832:22]
  wire [31:0] n489_O_1_2; // @[Top.scala 832:22]
  wire [31:0] n489_O_2_0; // @[Top.scala 832:22]
  wire [31:0] n489_O_2_1; // @[Top.scala 832:22]
  wire [31:0] n489_O_2_2; // @[Top.scala 832:22]
  wire [31:0] n489_O_3_0; // @[Top.scala 832:22]
  wire [31:0] n489_O_3_1; // @[Top.scala 832:22]
  wire [31:0] n489_O_3_2; // @[Top.scala 832:22]
  wire [31:0] n489_O_4_0; // @[Top.scala 832:22]
  wire [31:0] n489_O_4_1; // @[Top.scala 832:22]
  wire [31:0] n489_O_4_2; // @[Top.scala 832:22]
  wire [31:0] n489_O_5_0; // @[Top.scala 832:22]
  wire [31:0] n489_O_5_1; // @[Top.scala 832:22]
  wire [31:0] n489_O_5_2; // @[Top.scala 832:22]
  wire [31:0] n489_O_6_0; // @[Top.scala 832:22]
  wire [31:0] n489_O_6_1; // @[Top.scala 832:22]
  wire [31:0] n489_O_6_2; // @[Top.scala 832:22]
  wire [31:0] n489_O_7_0; // @[Top.scala 832:22]
  wire [31:0] n489_O_7_1; // @[Top.scala 832:22]
  wire [31:0] n489_O_7_2; // @[Top.scala 832:22]
  wire  n498_valid_up; // @[Top.scala 836:22]
  wire  n498_valid_down; // @[Top.scala 836:22]
  wire [31:0] n498_I_0_0; // @[Top.scala 836:22]
  wire [31:0] n498_I_0_1; // @[Top.scala 836:22]
  wire [31:0] n498_I_0_2; // @[Top.scala 836:22]
  wire [31:0] n498_I_1_0; // @[Top.scala 836:22]
  wire [31:0] n498_I_1_1; // @[Top.scala 836:22]
  wire [31:0] n498_I_1_2; // @[Top.scala 836:22]
  wire [31:0] n498_I_2_0; // @[Top.scala 836:22]
  wire [31:0] n498_I_2_1; // @[Top.scala 836:22]
  wire [31:0] n498_I_2_2; // @[Top.scala 836:22]
  wire [31:0] n498_I_3_0; // @[Top.scala 836:22]
  wire [31:0] n498_I_3_1; // @[Top.scala 836:22]
  wire [31:0] n498_I_3_2; // @[Top.scala 836:22]
  wire [31:0] n498_I_4_0; // @[Top.scala 836:22]
  wire [31:0] n498_I_4_1; // @[Top.scala 836:22]
  wire [31:0] n498_I_4_2; // @[Top.scala 836:22]
  wire [31:0] n498_I_5_0; // @[Top.scala 836:22]
  wire [31:0] n498_I_5_1; // @[Top.scala 836:22]
  wire [31:0] n498_I_5_2; // @[Top.scala 836:22]
  wire [31:0] n498_I_6_0; // @[Top.scala 836:22]
  wire [31:0] n498_I_6_1; // @[Top.scala 836:22]
  wire [31:0] n498_I_6_2; // @[Top.scala 836:22]
  wire [31:0] n498_I_7_0; // @[Top.scala 836:22]
  wire [31:0] n498_I_7_1; // @[Top.scala 836:22]
  wire [31:0] n498_I_7_2; // @[Top.scala 836:22]
  wire [31:0] n498_O_0_0_0; // @[Top.scala 836:22]
  wire [31:0] n498_O_0_0_1; // @[Top.scala 836:22]
  wire [31:0] n498_O_0_0_2; // @[Top.scala 836:22]
  wire [31:0] n498_O_1_0_0; // @[Top.scala 836:22]
  wire [31:0] n498_O_1_0_1; // @[Top.scala 836:22]
  wire [31:0] n498_O_1_0_2; // @[Top.scala 836:22]
  wire [31:0] n498_O_2_0_0; // @[Top.scala 836:22]
  wire [31:0] n498_O_2_0_1; // @[Top.scala 836:22]
  wire [31:0] n498_O_2_0_2; // @[Top.scala 836:22]
  wire [31:0] n498_O_3_0_0; // @[Top.scala 836:22]
  wire [31:0] n498_O_3_0_1; // @[Top.scala 836:22]
  wire [31:0] n498_O_3_0_2; // @[Top.scala 836:22]
  wire [31:0] n498_O_4_0_0; // @[Top.scala 836:22]
  wire [31:0] n498_O_4_0_1; // @[Top.scala 836:22]
  wire [31:0] n498_O_4_0_2; // @[Top.scala 836:22]
  wire [31:0] n498_O_5_0_0; // @[Top.scala 836:22]
  wire [31:0] n498_O_5_0_1; // @[Top.scala 836:22]
  wire [31:0] n498_O_5_0_2; // @[Top.scala 836:22]
  wire [31:0] n498_O_6_0_0; // @[Top.scala 836:22]
  wire [31:0] n498_O_6_0_1; // @[Top.scala 836:22]
  wire [31:0] n498_O_6_0_2; // @[Top.scala 836:22]
  wire [31:0] n498_O_7_0_0; // @[Top.scala 836:22]
  wire [31:0] n498_O_7_0_1; // @[Top.scala 836:22]
  wire [31:0] n498_O_7_0_2; // @[Top.scala 836:22]
  wire  n505_valid_up; // @[Top.scala 839:22]
  wire  n505_valid_down; // @[Top.scala 839:22]
  wire [31:0] n505_I_0_0_0; // @[Top.scala 839:22]
  wire [31:0] n505_I_0_0_1; // @[Top.scala 839:22]
  wire [31:0] n505_I_0_0_2; // @[Top.scala 839:22]
  wire [31:0] n505_I_1_0_0; // @[Top.scala 839:22]
  wire [31:0] n505_I_1_0_1; // @[Top.scala 839:22]
  wire [31:0] n505_I_1_0_2; // @[Top.scala 839:22]
  wire [31:0] n505_I_2_0_0; // @[Top.scala 839:22]
  wire [31:0] n505_I_2_0_1; // @[Top.scala 839:22]
  wire [31:0] n505_I_2_0_2; // @[Top.scala 839:22]
  wire [31:0] n505_I_3_0_0; // @[Top.scala 839:22]
  wire [31:0] n505_I_3_0_1; // @[Top.scala 839:22]
  wire [31:0] n505_I_3_0_2; // @[Top.scala 839:22]
  wire [31:0] n505_I_4_0_0; // @[Top.scala 839:22]
  wire [31:0] n505_I_4_0_1; // @[Top.scala 839:22]
  wire [31:0] n505_I_4_0_2; // @[Top.scala 839:22]
  wire [31:0] n505_I_5_0_0; // @[Top.scala 839:22]
  wire [31:0] n505_I_5_0_1; // @[Top.scala 839:22]
  wire [31:0] n505_I_5_0_2; // @[Top.scala 839:22]
  wire [31:0] n505_I_6_0_0; // @[Top.scala 839:22]
  wire [31:0] n505_I_6_0_1; // @[Top.scala 839:22]
  wire [31:0] n505_I_6_0_2; // @[Top.scala 839:22]
  wire [31:0] n505_I_7_0_0; // @[Top.scala 839:22]
  wire [31:0] n505_I_7_0_1; // @[Top.scala 839:22]
  wire [31:0] n505_I_7_0_2; // @[Top.scala 839:22]
  wire [31:0] n505_O_0_0; // @[Top.scala 839:22]
  wire [31:0] n505_O_0_1; // @[Top.scala 839:22]
  wire [31:0] n505_O_0_2; // @[Top.scala 839:22]
  wire [31:0] n505_O_1_0; // @[Top.scala 839:22]
  wire [31:0] n505_O_1_1; // @[Top.scala 839:22]
  wire [31:0] n505_O_1_2; // @[Top.scala 839:22]
  wire [31:0] n505_O_2_0; // @[Top.scala 839:22]
  wire [31:0] n505_O_2_1; // @[Top.scala 839:22]
  wire [31:0] n505_O_2_2; // @[Top.scala 839:22]
  wire [31:0] n505_O_3_0; // @[Top.scala 839:22]
  wire [31:0] n505_O_3_1; // @[Top.scala 839:22]
  wire [31:0] n505_O_3_2; // @[Top.scala 839:22]
  wire [31:0] n505_O_4_0; // @[Top.scala 839:22]
  wire [31:0] n505_O_4_1; // @[Top.scala 839:22]
  wire [31:0] n505_O_4_2; // @[Top.scala 839:22]
  wire [31:0] n505_O_5_0; // @[Top.scala 839:22]
  wire [31:0] n505_O_5_1; // @[Top.scala 839:22]
  wire [31:0] n505_O_5_2; // @[Top.scala 839:22]
  wire [31:0] n505_O_6_0; // @[Top.scala 839:22]
  wire [31:0] n505_O_6_1; // @[Top.scala 839:22]
  wire [31:0] n505_O_6_2; // @[Top.scala 839:22]
  wire [31:0] n505_O_7_0; // @[Top.scala 839:22]
  wire [31:0] n505_O_7_1; // @[Top.scala 839:22]
  wire [31:0] n505_O_7_2; // @[Top.scala 839:22]
  wire  n506_valid_up; // @[Top.scala 842:22]
  wire  n506_valid_down; // @[Top.scala 842:22]
  wire [31:0] n506_I0_0_0; // @[Top.scala 842:22]
  wire [31:0] n506_I0_0_1; // @[Top.scala 842:22]
  wire [31:0] n506_I0_0_2; // @[Top.scala 842:22]
  wire [31:0] n506_I0_1_0; // @[Top.scala 842:22]
  wire [31:0] n506_I0_1_1; // @[Top.scala 842:22]
  wire [31:0] n506_I0_1_2; // @[Top.scala 842:22]
  wire [31:0] n506_I0_2_0; // @[Top.scala 842:22]
  wire [31:0] n506_I0_2_1; // @[Top.scala 842:22]
  wire [31:0] n506_I0_2_2; // @[Top.scala 842:22]
  wire [31:0] n506_I0_3_0; // @[Top.scala 842:22]
  wire [31:0] n506_I0_3_1; // @[Top.scala 842:22]
  wire [31:0] n506_I0_3_2; // @[Top.scala 842:22]
  wire [31:0] n506_I0_4_0; // @[Top.scala 842:22]
  wire [31:0] n506_I0_4_1; // @[Top.scala 842:22]
  wire [31:0] n506_I0_4_2; // @[Top.scala 842:22]
  wire [31:0] n506_I0_5_0; // @[Top.scala 842:22]
  wire [31:0] n506_I0_5_1; // @[Top.scala 842:22]
  wire [31:0] n506_I0_5_2; // @[Top.scala 842:22]
  wire [31:0] n506_I0_6_0; // @[Top.scala 842:22]
  wire [31:0] n506_I0_6_1; // @[Top.scala 842:22]
  wire [31:0] n506_I0_6_2; // @[Top.scala 842:22]
  wire [31:0] n506_I0_7_0; // @[Top.scala 842:22]
  wire [31:0] n506_I0_7_1; // @[Top.scala 842:22]
  wire [31:0] n506_I0_7_2; // @[Top.scala 842:22]
  wire [31:0] n506_I1_0_0; // @[Top.scala 842:22]
  wire [31:0] n506_I1_0_1; // @[Top.scala 842:22]
  wire [31:0] n506_I1_0_2; // @[Top.scala 842:22]
  wire [31:0] n506_I1_1_0; // @[Top.scala 842:22]
  wire [31:0] n506_I1_1_1; // @[Top.scala 842:22]
  wire [31:0] n506_I1_1_2; // @[Top.scala 842:22]
  wire [31:0] n506_I1_2_0; // @[Top.scala 842:22]
  wire [31:0] n506_I1_2_1; // @[Top.scala 842:22]
  wire [31:0] n506_I1_2_2; // @[Top.scala 842:22]
  wire [31:0] n506_I1_3_0; // @[Top.scala 842:22]
  wire [31:0] n506_I1_3_1; // @[Top.scala 842:22]
  wire [31:0] n506_I1_3_2; // @[Top.scala 842:22]
  wire [31:0] n506_I1_4_0; // @[Top.scala 842:22]
  wire [31:0] n506_I1_4_1; // @[Top.scala 842:22]
  wire [31:0] n506_I1_4_2; // @[Top.scala 842:22]
  wire [31:0] n506_I1_5_0; // @[Top.scala 842:22]
  wire [31:0] n506_I1_5_1; // @[Top.scala 842:22]
  wire [31:0] n506_I1_5_2; // @[Top.scala 842:22]
  wire [31:0] n506_I1_6_0; // @[Top.scala 842:22]
  wire [31:0] n506_I1_6_1; // @[Top.scala 842:22]
  wire [31:0] n506_I1_6_2; // @[Top.scala 842:22]
  wire [31:0] n506_I1_7_0; // @[Top.scala 842:22]
  wire [31:0] n506_I1_7_1; // @[Top.scala 842:22]
  wire [31:0] n506_I1_7_2; // @[Top.scala 842:22]
  wire [31:0] n506_O_0_0_0; // @[Top.scala 842:22]
  wire [31:0] n506_O_0_0_1; // @[Top.scala 842:22]
  wire [31:0] n506_O_0_0_2; // @[Top.scala 842:22]
  wire [31:0] n506_O_0_1_0; // @[Top.scala 842:22]
  wire [31:0] n506_O_0_1_1; // @[Top.scala 842:22]
  wire [31:0] n506_O_0_1_2; // @[Top.scala 842:22]
  wire [31:0] n506_O_1_0_0; // @[Top.scala 842:22]
  wire [31:0] n506_O_1_0_1; // @[Top.scala 842:22]
  wire [31:0] n506_O_1_0_2; // @[Top.scala 842:22]
  wire [31:0] n506_O_1_1_0; // @[Top.scala 842:22]
  wire [31:0] n506_O_1_1_1; // @[Top.scala 842:22]
  wire [31:0] n506_O_1_1_2; // @[Top.scala 842:22]
  wire [31:0] n506_O_2_0_0; // @[Top.scala 842:22]
  wire [31:0] n506_O_2_0_1; // @[Top.scala 842:22]
  wire [31:0] n506_O_2_0_2; // @[Top.scala 842:22]
  wire [31:0] n506_O_2_1_0; // @[Top.scala 842:22]
  wire [31:0] n506_O_2_1_1; // @[Top.scala 842:22]
  wire [31:0] n506_O_2_1_2; // @[Top.scala 842:22]
  wire [31:0] n506_O_3_0_0; // @[Top.scala 842:22]
  wire [31:0] n506_O_3_0_1; // @[Top.scala 842:22]
  wire [31:0] n506_O_3_0_2; // @[Top.scala 842:22]
  wire [31:0] n506_O_3_1_0; // @[Top.scala 842:22]
  wire [31:0] n506_O_3_1_1; // @[Top.scala 842:22]
  wire [31:0] n506_O_3_1_2; // @[Top.scala 842:22]
  wire [31:0] n506_O_4_0_0; // @[Top.scala 842:22]
  wire [31:0] n506_O_4_0_1; // @[Top.scala 842:22]
  wire [31:0] n506_O_4_0_2; // @[Top.scala 842:22]
  wire [31:0] n506_O_4_1_0; // @[Top.scala 842:22]
  wire [31:0] n506_O_4_1_1; // @[Top.scala 842:22]
  wire [31:0] n506_O_4_1_2; // @[Top.scala 842:22]
  wire [31:0] n506_O_5_0_0; // @[Top.scala 842:22]
  wire [31:0] n506_O_5_0_1; // @[Top.scala 842:22]
  wire [31:0] n506_O_5_0_2; // @[Top.scala 842:22]
  wire [31:0] n506_O_5_1_0; // @[Top.scala 842:22]
  wire [31:0] n506_O_5_1_1; // @[Top.scala 842:22]
  wire [31:0] n506_O_5_1_2; // @[Top.scala 842:22]
  wire [31:0] n506_O_6_0_0; // @[Top.scala 842:22]
  wire [31:0] n506_O_6_0_1; // @[Top.scala 842:22]
  wire [31:0] n506_O_6_0_2; // @[Top.scala 842:22]
  wire [31:0] n506_O_6_1_0; // @[Top.scala 842:22]
  wire [31:0] n506_O_6_1_1; // @[Top.scala 842:22]
  wire [31:0] n506_O_6_1_2; // @[Top.scala 842:22]
  wire [31:0] n506_O_7_0_0; // @[Top.scala 842:22]
  wire [31:0] n506_O_7_0_1; // @[Top.scala 842:22]
  wire [31:0] n506_O_7_0_2; // @[Top.scala 842:22]
  wire [31:0] n506_O_7_1_0; // @[Top.scala 842:22]
  wire [31:0] n506_O_7_1_1; // @[Top.scala 842:22]
  wire [31:0] n506_O_7_1_2; // @[Top.scala 842:22]
  wire  n513_clock; // @[Top.scala 846:22]
  wire  n513_valid_up; // @[Top.scala 846:22]
  wire  n513_valid_down; // @[Top.scala 846:22]
  wire [31:0] n513_I_0; // @[Top.scala 846:22]
  wire [31:0] n513_I_1; // @[Top.scala 846:22]
  wire [31:0] n513_I_2; // @[Top.scala 846:22]
  wire [31:0] n513_I_3; // @[Top.scala 846:22]
  wire [31:0] n513_I_4; // @[Top.scala 846:22]
  wire [31:0] n513_I_5; // @[Top.scala 846:22]
  wire [31:0] n513_I_6; // @[Top.scala 846:22]
  wire [31:0] n513_I_7; // @[Top.scala 846:22]
  wire [31:0] n513_O_0; // @[Top.scala 846:22]
  wire [31:0] n513_O_1; // @[Top.scala 846:22]
  wire [31:0] n513_O_2; // @[Top.scala 846:22]
  wire [31:0] n513_O_3; // @[Top.scala 846:22]
  wire [31:0] n513_O_4; // @[Top.scala 846:22]
  wire [31:0] n513_O_5; // @[Top.scala 846:22]
  wire [31:0] n513_O_6; // @[Top.scala 846:22]
  wire [31:0] n513_O_7; // @[Top.scala 846:22]
  wire  n514_clock; // @[Top.scala 849:22]
  wire  n514_valid_up; // @[Top.scala 849:22]
  wire  n514_valid_down; // @[Top.scala 849:22]
  wire [31:0] n514_I_0; // @[Top.scala 849:22]
  wire [31:0] n514_I_1; // @[Top.scala 849:22]
  wire [31:0] n514_I_2; // @[Top.scala 849:22]
  wire [31:0] n514_I_3; // @[Top.scala 849:22]
  wire [31:0] n514_I_4; // @[Top.scala 849:22]
  wire [31:0] n514_I_5; // @[Top.scala 849:22]
  wire [31:0] n514_I_6; // @[Top.scala 849:22]
  wire [31:0] n514_I_7; // @[Top.scala 849:22]
  wire [31:0] n514_O_0; // @[Top.scala 849:22]
  wire [31:0] n514_O_1; // @[Top.scala 849:22]
  wire [31:0] n514_O_2; // @[Top.scala 849:22]
  wire [31:0] n514_O_3; // @[Top.scala 849:22]
  wire [31:0] n514_O_4; // @[Top.scala 849:22]
  wire [31:0] n514_O_5; // @[Top.scala 849:22]
  wire [31:0] n514_O_6; // @[Top.scala 849:22]
  wire [31:0] n514_O_7; // @[Top.scala 849:22]
  wire  n515_valid_up; // @[Top.scala 852:22]
  wire  n515_valid_down; // @[Top.scala 852:22]
  wire [31:0] n515_I0_0; // @[Top.scala 852:22]
  wire [31:0] n515_I0_1; // @[Top.scala 852:22]
  wire [31:0] n515_I0_2; // @[Top.scala 852:22]
  wire [31:0] n515_I0_3; // @[Top.scala 852:22]
  wire [31:0] n515_I0_4; // @[Top.scala 852:22]
  wire [31:0] n515_I0_5; // @[Top.scala 852:22]
  wire [31:0] n515_I0_6; // @[Top.scala 852:22]
  wire [31:0] n515_I0_7; // @[Top.scala 852:22]
  wire [31:0] n515_I1_0; // @[Top.scala 852:22]
  wire [31:0] n515_I1_1; // @[Top.scala 852:22]
  wire [31:0] n515_I1_2; // @[Top.scala 852:22]
  wire [31:0] n515_I1_3; // @[Top.scala 852:22]
  wire [31:0] n515_I1_4; // @[Top.scala 852:22]
  wire [31:0] n515_I1_5; // @[Top.scala 852:22]
  wire [31:0] n515_I1_6; // @[Top.scala 852:22]
  wire [31:0] n515_I1_7; // @[Top.scala 852:22]
  wire [31:0] n515_O_0_0; // @[Top.scala 852:22]
  wire [31:0] n515_O_0_1; // @[Top.scala 852:22]
  wire [31:0] n515_O_1_0; // @[Top.scala 852:22]
  wire [31:0] n515_O_1_1; // @[Top.scala 852:22]
  wire [31:0] n515_O_2_0; // @[Top.scala 852:22]
  wire [31:0] n515_O_2_1; // @[Top.scala 852:22]
  wire [31:0] n515_O_3_0; // @[Top.scala 852:22]
  wire [31:0] n515_O_3_1; // @[Top.scala 852:22]
  wire [31:0] n515_O_4_0; // @[Top.scala 852:22]
  wire [31:0] n515_O_4_1; // @[Top.scala 852:22]
  wire [31:0] n515_O_5_0; // @[Top.scala 852:22]
  wire [31:0] n515_O_5_1; // @[Top.scala 852:22]
  wire [31:0] n515_O_6_0; // @[Top.scala 852:22]
  wire [31:0] n515_O_6_1; // @[Top.scala 852:22]
  wire [31:0] n515_O_7_0; // @[Top.scala 852:22]
  wire [31:0] n515_O_7_1; // @[Top.scala 852:22]
  wire  n522_valid_up; // @[Top.scala 856:22]
  wire  n522_valid_down; // @[Top.scala 856:22]
  wire [31:0] n522_I0_0_0; // @[Top.scala 856:22]
  wire [31:0] n522_I0_0_1; // @[Top.scala 856:22]
  wire [31:0] n522_I0_1_0; // @[Top.scala 856:22]
  wire [31:0] n522_I0_1_1; // @[Top.scala 856:22]
  wire [31:0] n522_I0_2_0; // @[Top.scala 856:22]
  wire [31:0] n522_I0_2_1; // @[Top.scala 856:22]
  wire [31:0] n522_I0_3_0; // @[Top.scala 856:22]
  wire [31:0] n522_I0_3_1; // @[Top.scala 856:22]
  wire [31:0] n522_I0_4_0; // @[Top.scala 856:22]
  wire [31:0] n522_I0_4_1; // @[Top.scala 856:22]
  wire [31:0] n522_I0_5_0; // @[Top.scala 856:22]
  wire [31:0] n522_I0_5_1; // @[Top.scala 856:22]
  wire [31:0] n522_I0_6_0; // @[Top.scala 856:22]
  wire [31:0] n522_I0_6_1; // @[Top.scala 856:22]
  wire [31:0] n522_I0_7_0; // @[Top.scala 856:22]
  wire [31:0] n522_I0_7_1; // @[Top.scala 856:22]
  wire [31:0] n522_I1_0; // @[Top.scala 856:22]
  wire [31:0] n522_I1_1; // @[Top.scala 856:22]
  wire [31:0] n522_I1_2; // @[Top.scala 856:22]
  wire [31:0] n522_I1_3; // @[Top.scala 856:22]
  wire [31:0] n522_I1_4; // @[Top.scala 856:22]
  wire [31:0] n522_I1_5; // @[Top.scala 856:22]
  wire [31:0] n522_I1_6; // @[Top.scala 856:22]
  wire [31:0] n522_I1_7; // @[Top.scala 856:22]
  wire [31:0] n522_O_0_0; // @[Top.scala 856:22]
  wire [31:0] n522_O_0_1; // @[Top.scala 856:22]
  wire [31:0] n522_O_0_2; // @[Top.scala 856:22]
  wire [31:0] n522_O_1_0; // @[Top.scala 856:22]
  wire [31:0] n522_O_1_1; // @[Top.scala 856:22]
  wire [31:0] n522_O_1_2; // @[Top.scala 856:22]
  wire [31:0] n522_O_2_0; // @[Top.scala 856:22]
  wire [31:0] n522_O_2_1; // @[Top.scala 856:22]
  wire [31:0] n522_O_2_2; // @[Top.scala 856:22]
  wire [31:0] n522_O_3_0; // @[Top.scala 856:22]
  wire [31:0] n522_O_3_1; // @[Top.scala 856:22]
  wire [31:0] n522_O_3_2; // @[Top.scala 856:22]
  wire [31:0] n522_O_4_0; // @[Top.scala 856:22]
  wire [31:0] n522_O_4_1; // @[Top.scala 856:22]
  wire [31:0] n522_O_4_2; // @[Top.scala 856:22]
  wire [31:0] n522_O_5_0; // @[Top.scala 856:22]
  wire [31:0] n522_O_5_1; // @[Top.scala 856:22]
  wire [31:0] n522_O_5_2; // @[Top.scala 856:22]
  wire [31:0] n522_O_6_0; // @[Top.scala 856:22]
  wire [31:0] n522_O_6_1; // @[Top.scala 856:22]
  wire [31:0] n522_O_6_2; // @[Top.scala 856:22]
  wire [31:0] n522_O_7_0; // @[Top.scala 856:22]
  wire [31:0] n522_O_7_1; // @[Top.scala 856:22]
  wire [31:0] n522_O_7_2; // @[Top.scala 856:22]
  wire  n531_valid_up; // @[Top.scala 860:22]
  wire  n531_valid_down; // @[Top.scala 860:22]
  wire [31:0] n531_I_0_0; // @[Top.scala 860:22]
  wire [31:0] n531_I_0_1; // @[Top.scala 860:22]
  wire [31:0] n531_I_0_2; // @[Top.scala 860:22]
  wire [31:0] n531_I_1_0; // @[Top.scala 860:22]
  wire [31:0] n531_I_1_1; // @[Top.scala 860:22]
  wire [31:0] n531_I_1_2; // @[Top.scala 860:22]
  wire [31:0] n531_I_2_0; // @[Top.scala 860:22]
  wire [31:0] n531_I_2_1; // @[Top.scala 860:22]
  wire [31:0] n531_I_2_2; // @[Top.scala 860:22]
  wire [31:0] n531_I_3_0; // @[Top.scala 860:22]
  wire [31:0] n531_I_3_1; // @[Top.scala 860:22]
  wire [31:0] n531_I_3_2; // @[Top.scala 860:22]
  wire [31:0] n531_I_4_0; // @[Top.scala 860:22]
  wire [31:0] n531_I_4_1; // @[Top.scala 860:22]
  wire [31:0] n531_I_4_2; // @[Top.scala 860:22]
  wire [31:0] n531_I_5_0; // @[Top.scala 860:22]
  wire [31:0] n531_I_5_1; // @[Top.scala 860:22]
  wire [31:0] n531_I_5_2; // @[Top.scala 860:22]
  wire [31:0] n531_I_6_0; // @[Top.scala 860:22]
  wire [31:0] n531_I_6_1; // @[Top.scala 860:22]
  wire [31:0] n531_I_6_2; // @[Top.scala 860:22]
  wire [31:0] n531_I_7_0; // @[Top.scala 860:22]
  wire [31:0] n531_I_7_1; // @[Top.scala 860:22]
  wire [31:0] n531_I_7_2; // @[Top.scala 860:22]
  wire [31:0] n531_O_0_0_0; // @[Top.scala 860:22]
  wire [31:0] n531_O_0_0_1; // @[Top.scala 860:22]
  wire [31:0] n531_O_0_0_2; // @[Top.scala 860:22]
  wire [31:0] n531_O_1_0_0; // @[Top.scala 860:22]
  wire [31:0] n531_O_1_0_1; // @[Top.scala 860:22]
  wire [31:0] n531_O_1_0_2; // @[Top.scala 860:22]
  wire [31:0] n531_O_2_0_0; // @[Top.scala 860:22]
  wire [31:0] n531_O_2_0_1; // @[Top.scala 860:22]
  wire [31:0] n531_O_2_0_2; // @[Top.scala 860:22]
  wire [31:0] n531_O_3_0_0; // @[Top.scala 860:22]
  wire [31:0] n531_O_3_0_1; // @[Top.scala 860:22]
  wire [31:0] n531_O_3_0_2; // @[Top.scala 860:22]
  wire [31:0] n531_O_4_0_0; // @[Top.scala 860:22]
  wire [31:0] n531_O_4_0_1; // @[Top.scala 860:22]
  wire [31:0] n531_O_4_0_2; // @[Top.scala 860:22]
  wire [31:0] n531_O_5_0_0; // @[Top.scala 860:22]
  wire [31:0] n531_O_5_0_1; // @[Top.scala 860:22]
  wire [31:0] n531_O_5_0_2; // @[Top.scala 860:22]
  wire [31:0] n531_O_6_0_0; // @[Top.scala 860:22]
  wire [31:0] n531_O_6_0_1; // @[Top.scala 860:22]
  wire [31:0] n531_O_6_0_2; // @[Top.scala 860:22]
  wire [31:0] n531_O_7_0_0; // @[Top.scala 860:22]
  wire [31:0] n531_O_7_0_1; // @[Top.scala 860:22]
  wire [31:0] n531_O_7_0_2; // @[Top.scala 860:22]
  wire  n538_valid_up; // @[Top.scala 863:22]
  wire  n538_valid_down; // @[Top.scala 863:22]
  wire [31:0] n538_I_0_0_0; // @[Top.scala 863:22]
  wire [31:0] n538_I_0_0_1; // @[Top.scala 863:22]
  wire [31:0] n538_I_0_0_2; // @[Top.scala 863:22]
  wire [31:0] n538_I_1_0_0; // @[Top.scala 863:22]
  wire [31:0] n538_I_1_0_1; // @[Top.scala 863:22]
  wire [31:0] n538_I_1_0_2; // @[Top.scala 863:22]
  wire [31:0] n538_I_2_0_0; // @[Top.scala 863:22]
  wire [31:0] n538_I_2_0_1; // @[Top.scala 863:22]
  wire [31:0] n538_I_2_0_2; // @[Top.scala 863:22]
  wire [31:0] n538_I_3_0_0; // @[Top.scala 863:22]
  wire [31:0] n538_I_3_0_1; // @[Top.scala 863:22]
  wire [31:0] n538_I_3_0_2; // @[Top.scala 863:22]
  wire [31:0] n538_I_4_0_0; // @[Top.scala 863:22]
  wire [31:0] n538_I_4_0_1; // @[Top.scala 863:22]
  wire [31:0] n538_I_4_0_2; // @[Top.scala 863:22]
  wire [31:0] n538_I_5_0_0; // @[Top.scala 863:22]
  wire [31:0] n538_I_5_0_1; // @[Top.scala 863:22]
  wire [31:0] n538_I_5_0_2; // @[Top.scala 863:22]
  wire [31:0] n538_I_6_0_0; // @[Top.scala 863:22]
  wire [31:0] n538_I_6_0_1; // @[Top.scala 863:22]
  wire [31:0] n538_I_6_0_2; // @[Top.scala 863:22]
  wire [31:0] n538_I_7_0_0; // @[Top.scala 863:22]
  wire [31:0] n538_I_7_0_1; // @[Top.scala 863:22]
  wire [31:0] n538_I_7_0_2; // @[Top.scala 863:22]
  wire [31:0] n538_O_0_0; // @[Top.scala 863:22]
  wire [31:0] n538_O_0_1; // @[Top.scala 863:22]
  wire [31:0] n538_O_0_2; // @[Top.scala 863:22]
  wire [31:0] n538_O_1_0; // @[Top.scala 863:22]
  wire [31:0] n538_O_1_1; // @[Top.scala 863:22]
  wire [31:0] n538_O_1_2; // @[Top.scala 863:22]
  wire [31:0] n538_O_2_0; // @[Top.scala 863:22]
  wire [31:0] n538_O_2_1; // @[Top.scala 863:22]
  wire [31:0] n538_O_2_2; // @[Top.scala 863:22]
  wire [31:0] n538_O_3_0; // @[Top.scala 863:22]
  wire [31:0] n538_O_3_1; // @[Top.scala 863:22]
  wire [31:0] n538_O_3_2; // @[Top.scala 863:22]
  wire [31:0] n538_O_4_0; // @[Top.scala 863:22]
  wire [31:0] n538_O_4_1; // @[Top.scala 863:22]
  wire [31:0] n538_O_4_2; // @[Top.scala 863:22]
  wire [31:0] n538_O_5_0; // @[Top.scala 863:22]
  wire [31:0] n538_O_5_1; // @[Top.scala 863:22]
  wire [31:0] n538_O_5_2; // @[Top.scala 863:22]
  wire [31:0] n538_O_6_0; // @[Top.scala 863:22]
  wire [31:0] n538_O_6_1; // @[Top.scala 863:22]
  wire [31:0] n538_O_6_2; // @[Top.scala 863:22]
  wire [31:0] n538_O_7_0; // @[Top.scala 863:22]
  wire [31:0] n538_O_7_1; // @[Top.scala 863:22]
  wire [31:0] n538_O_7_2; // @[Top.scala 863:22]
  wire  n539_valid_up; // @[Top.scala 866:22]
  wire  n539_valid_down; // @[Top.scala 866:22]
  wire [31:0] n539_I0_0_0_0; // @[Top.scala 866:22]
  wire [31:0] n539_I0_0_0_1; // @[Top.scala 866:22]
  wire [31:0] n539_I0_0_0_2; // @[Top.scala 866:22]
  wire [31:0] n539_I0_0_1_0; // @[Top.scala 866:22]
  wire [31:0] n539_I0_0_1_1; // @[Top.scala 866:22]
  wire [31:0] n539_I0_0_1_2; // @[Top.scala 866:22]
  wire [31:0] n539_I0_1_0_0; // @[Top.scala 866:22]
  wire [31:0] n539_I0_1_0_1; // @[Top.scala 866:22]
  wire [31:0] n539_I0_1_0_2; // @[Top.scala 866:22]
  wire [31:0] n539_I0_1_1_0; // @[Top.scala 866:22]
  wire [31:0] n539_I0_1_1_1; // @[Top.scala 866:22]
  wire [31:0] n539_I0_1_1_2; // @[Top.scala 866:22]
  wire [31:0] n539_I0_2_0_0; // @[Top.scala 866:22]
  wire [31:0] n539_I0_2_0_1; // @[Top.scala 866:22]
  wire [31:0] n539_I0_2_0_2; // @[Top.scala 866:22]
  wire [31:0] n539_I0_2_1_0; // @[Top.scala 866:22]
  wire [31:0] n539_I0_2_1_1; // @[Top.scala 866:22]
  wire [31:0] n539_I0_2_1_2; // @[Top.scala 866:22]
  wire [31:0] n539_I0_3_0_0; // @[Top.scala 866:22]
  wire [31:0] n539_I0_3_0_1; // @[Top.scala 866:22]
  wire [31:0] n539_I0_3_0_2; // @[Top.scala 866:22]
  wire [31:0] n539_I0_3_1_0; // @[Top.scala 866:22]
  wire [31:0] n539_I0_3_1_1; // @[Top.scala 866:22]
  wire [31:0] n539_I0_3_1_2; // @[Top.scala 866:22]
  wire [31:0] n539_I0_4_0_0; // @[Top.scala 866:22]
  wire [31:0] n539_I0_4_0_1; // @[Top.scala 866:22]
  wire [31:0] n539_I0_4_0_2; // @[Top.scala 866:22]
  wire [31:0] n539_I0_4_1_0; // @[Top.scala 866:22]
  wire [31:0] n539_I0_4_1_1; // @[Top.scala 866:22]
  wire [31:0] n539_I0_4_1_2; // @[Top.scala 866:22]
  wire [31:0] n539_I0_5_0_0; // @[Top.scala 866:22]
  wire [31:0] n539_I0_5_0_1; // @[Top.scala 866:22]
  wire [31:0] n539_I0_5_0_2; // @[Top.scala 866:22]
  wire [31:0] n539_I0_5_1_0; // @[Top.scala 866:22]
  wire [31:0] n539_I0_5_1_1; // @[Top.scala 866:22]
  wire [31:0] n539_I0_5_1_2; // @[Top.scala 866:22]
  wire [31:0] n539_I0_6_0_0; // @[Top.scala 866:22]
  wire [31:0] n539_I0_6_0_1; // @[Top.scala 866:22]
  wire [31:0] n539_I0_6_0_2; // @[Top.scala 866:22]
  wire [31:0] n539_I0_6_1_0; // @[Top.scala 866:22]
  wire [31:0] n539_I0_6_1_1; // @[Top.scala 866:22]
  wire [31:0] n539_I0_6_1_2; // @[Top.scala 866:22]
  wire [31:0] n539_I0_7_0_0; // @[Top.scala 866:22]
  wire [31:0] n539_I0_7_0_1; // @[Top.scala 866:22]
  wire [31:0] n539_I0_7_0_2; // @[Top.scala 866:22]
  wire [31:0] n539_I0_7_1_0; // @[Top.scala 866:22]
  wire [31:0] n539_I0_7_1_1; // @[Top.scala 866:22]
  wire [31:0] n539_I0_7_1_2; // @[Top.scala 866:22]
  wire [31:0] n539_I1_0_0; // @[Top.scala 866:22]
  wire [31:0] n539_I1_0_1; // @[Top.scala 866:22]
  wire [31:0] n539_I1_0_2; // @[Top.scala 866:22]
  wire [31:0] n539_I1_1_0; // @[Top.scala 866:22]
  wire [31:0] n539_I1_1_1; // @[Top.scala 866:22]
  wire [31:0] n539_I1_1_2; // @[Top.scala 866:22]
  wire [31:0] n539_I1_2_0; // @[Top.scala 866:22]
  wire [31:0] n539_I1_2_1; // @[Top.scala 866:22]
  wire [31:0] n539_I1_2_2; // @[Top.scala 866:22]
  wire [31:0] n539_I1_3_0; // @[Top.scala 866:22]
  wire [31:0] n539_I1_3_1; // @[Top.scala 866:22]
  wire [31:0] n539_I1_3_2; // @[Top.scala 866:22]
  wire [31:0] n539_I1_4_0; // @[Top.scala 866:22]
  wire [31:0] n539_I1_4_1; // @[Top.scala 866:22]
  wire [31:0] n539_I1_4_2; // @[Top.scala 866:22]
  wire [31:0] n539_I1_5_0; // @[Top.scala 866:22]
  wire [31:0] n539_I1_5_1; // @[Top.scala 866:22]
  wire [31:0] n539_I1_5_2; // @[Top.scala 866:22]
  wire [31:0] n539_I1_6_0; // @[Top.scala 866:22]
  wire [31:0] n539_I1_6_1; // @[Top.scala 866:22]
  wire [31:0] n539_I1_6_2; // @[Top.scala 866:22]
  wire [31:0] n539_I1_7_0; // @[Top.scala 866:22]
  wire [31:0] n539_I1_7_1; // @[Top.scala 866:22]
  wire [31:0] n539_I1_7_2; // @[Top.scala 866:22]
  wire [31:0] n539_O_0_0_0; // @[Top.scala 866:22]
  wire [31:0] n539_O_0_0_1; // @[Top.scala 866:22]
  wire [31:0] n539_O_0_0_2; // @[Top.scala 866:22]
  wire [31:0] n539_O_0_1_0; // @[Top.scala 866:22]
  wire [31:0] n539_O_0_1_1; // @[Top.scala 866:22]
  wire [31:0] n539_O_0_1_2; // @[Top.scala 866:22]
  wire [31:0] n539_O_0_2_0; // @[Top.scala 866:22]
  wire [31:0] n539_O_0_2_1; // @[Top.scala 866:22]
  wire [31:0] n539_O_0_2_2; // @[Top.scala 866:22]
  wire [31:0] n539_O_1_0_0; // @[Top.scala 866:22]
  wire [31:0] n539_O_1_0_1; // @[Top.scala 866:22]
  wire [31:0] n539_O_1_0_2; // @[Top.scala 866:22]
  wire [31:0] n539_O_1_1_0; // @[Top.scala 866:22]
  wire [31:0] n539_O_1_1_1; // @[Top.scala 866:22]
  wire [31:0] n539_O_1_1_2; // @[Top.scala 866:22]
  wire [31:0] n539_O_1_2_0; // @[Top.scala 866:22]
  wire [31:0] n539_O_1_2_1; // @[Top.scala 866:22]
  wire [31:0] n539_O_1_2_2; // @[Top.scala 866:22]
  wire [31:0] n539_O_2_0_0; // @[Top.scala 866:22]
  wire [31:0] n539_O_2_0_1; // @[Top.scala 866:22]
  wire [31:0] n539_O_2_0_2; // @[Top.scala 866:22]
  wire [31:0] n539_O_2_1_0; // @[Top.scala 866:22]
  wire [31:0] n539_O_2_1_1; // @[Top.scala 866:22]
  wire [31:0] n539_O_2_1_2; // @[Top.scala 866:22]
  wire [31:0] n539_O_2_2_0; // @[Top.scala 866:22]
  wire [31:0] n539_O_2_2_1; // @[Top.scala 866:22]
  wire [31:0] n539_O_2_2_2; // @[Top.scala 866:22]
  wire [31:0] n539_O_3_0_0; // @[Top.scala 866:22]
  wire [31:0] n539_O_3_0_1; // @[Top.scala 866:22]
  wire [31:0] n539_O_3_0_2; // @[Top.scala 866:22]
  wire [31:0] n539_O_3_1_0; // @[Top.scala 866:22]
  wire [31:0] n539_O_3_1_1; // @[Top.scala 866:22]
  wire [31:0] n539_O_3_1_2; // @[Top.scala 866:22]
  wire [31:0] n539_O_3_2_0; // @[Top.scala 866:22]
  wire [31:0] n539_O_3_2_1; // @[Top.scala 866:22]
  wire [31:0] n539_O_3_2_2; // @[Top.scala 866:22]
  wire [31:0] n539_O_4_0_0; // @[Top.scala 866:22]
  wire [31:0] n539_O_4_0_1; // @[Top.scala 866:22]
  wire [31:0] n539_O_4_0_2; // @[Top.scala 866:22]
  wire [31:0] n539_O_4_1_0; // @[Top.scala 866:22]
  wire [31:0] n539_O_4_1_1; // @[Top.scala 866:22]
  wire [31:0] n539_O_4_1_2; // @[Top.scala 866:22]
  wire [31:0] n539_O_4_2_0; // @[Top.scala 866:22]
  wire [31:0] n539_O_4_2_1; // @[Top.scala 866:22]
  wire [31:0] n539_O_4_2_2; // @[Top.scala 866:22]
  wire [31:0] n539_O_5_0_0; // @[Top.scala 866:22]
  wire [31:0] n539_O_5_0_1; // @[Top.scala 866:22]
  wire [31:0] n539_O_5_0_2; // @[Top.scala 866:22]
  wire [31:0] n539_O_5_1_0; // @[Top.scala 866:22]
  wire [31:0] n539_O_5_1_1; // @[Top.scala 866:22]
  wire [31:0] n539_O_5_1_2; // @[Top.scala 866:22]
  wire [31:0] n539_O_5_2_0; // @[Top.scala 866:22]
  wire [31:0] n539_O_5_2_1; // @[Top.scala 866:22]
  wire [31:0] n539_O_5_2_2; // @[Top.scala 866:22]
  wire [31:0] n539_O_6_0_0; // @[Top.scala 866:22]
  wire [31:0] n539_O_6_0_1; // @[Top.scala 866:22]
  wire [31:0] n539_O_6_0_2; // @[Top.scala 866:22]
  wire [31:0] n539_O_6_1_0; // @[Top.scala 866:22]
  wire [31:0] n539_O_6_1_1; // @[Top.scala 866:22]
  wire [31:0] n539_O_6_1_2; // @[Top.scala 866:22]
  wire [31:0] n539_O_6_2_0; // @[Top.scala 866:22]
  wire [31:0] n539_O_6_2_1; // @[Top.scala 866:22]
  wire [31:0] n539_O_6_2_2; // @[Top.scala 866:22]
  wire [31:0] n539_O_7_0_0; // @[Top.scala 866:22]
  wire [31:0] n539_O_7_0_1; // @[Top.scala 866:22]
  wire [31:0] n539_O_7_0_2; // @[Top.scala 866:22]
  wire [31:0] n539_O_7_1_0; // @[Top.scala 866:22]
  wire [31:0] n539_O_7_1_1; // @[Top.scala 866:22]
  wire [31:0] n539_O_7_1_2; // @[Top.scala 866:22]
  wire [31:0] n539_O_7_2_0; // @[Top.scala 866:22]
  wire [31:0] n539_O_7_2_1; // @[Top.scala 866:22]
  wire [31:0] n539_O_7_2_2; // @[Top.scala 866:22]
  wire  n548_valid_up; // @[Top.scala 870:22]
  wire  n548_valid_down; // @[Top.scala 870:22]
  wire [31:0] n548_I_0_0_0; // @[Top.scala 870:22]
  wire [31:0] n548_I_0_0_1; // @[Top.scala 870:22]
  wire [31:0] n548_I_0_0_2; // @[Top.scala 870:22]
  wire [31:0] n548_I_0_1_0; // @[Top.scala 870:22]
  wire [31:0] n548_I_0_1_1; // @[Top.scala 870:22]
  wire [31:0] n548_I_0_1_2; // @[Top.scala 870:22]
  wire [31:0] n548_I_0_2_0; // @[Top.scala 870:22]
  wire [31:0] n548_I_0_2_1; // @[Top.scala 870:22]
  wire [31:0] n548_I_0_2_2; // @[Top.scala 870:22]
  wire [31:0] n548_I_1_0_0; // @[Top.scala 870:22]
  wire [31:0] n548_I_1_0_1; // @[Top.scala 870:22]
  wire [31:0] n548_I_1_0_2; // @[Top.scala 870:22]
  wire [31:0] n548_I_1_1_0; // @[Top.scala 870:22]
  wire [31:0] n548_I_1_1_1; // @[Top.scala 870:22]
  wire [31:0] n548_I_1_1_2; // @[Top.scala 870:22]
  wire [31:0] n548_I_1_2_0; // @[Top.scala 870:22]
  wire [31:0] n548_I_1_2_1; // @[Top.scala 870:22]
  wire [31:0] n548_I_1_2_2; // @[Top.scala 870:22]
  wire [31:0] n548_I_2_0_0; // @[Top.scala 870:22]
  wire [31:0] n548_I_2_0_1; // @[Top.scala 870:22]
  wire [31:0] n548_I_2_0_2; // @[Top.scala 870:22]
  wire [31:0] n548_I_2_1_0; // @[Top.scala 870:22]
  wire [31:0] n548_I_2_1_1; // @[Top.scala 870:22]
  wire [31:0] n548_I_2_1_2; // @[Top.scala 870:22]
  wire [31:0] n548_I_2_2_0; // @[Top.scala 870:22]
  wire [31:0] n548_I_2_2_1; // @[Top.scala 870:22]
  wire [31:0] n548_I_2_2_2; // @[Top.scala 870:22]
  wire [31:0] n548_I_3_0_0; // @[Top.scala 870:22]
  wire [31:0] n548_I_3_0_1; // @[Top.scala 870:22]
  wire [31:0] n548_I_3_0_2; // @[Top.scala 870:22]
  wire [31:0] n548_I_3_1_0; // @[Top.scala 870:22]
  wire [31:0] n548_I_3_1_1; // @[Top.scala 870:22]
  wire [31:0] n548_I_3_1_2; // @[Top.scala 870:22]
  wire [31:0] n548_I_3_2_0; // @[Top.scala 870:22]
  wire [31:0] n548_I_3_2_1; // @[Top.scala 870:22]
  wire [31:0] n548_I_3_2_2; // @[Top.scala 870:22]
  wire [31:0] n548_I_4_0_0; // @[Top.scala 870:22]
  wire [31:0] n548_I_4_0_1; // @[Top.scala 870:22]
  wire [31:0] n548_I_4_0_2; // @[Top.scala 870:22]
  wire [31:0] n548_I_4_1_0; // @[Top.scala 870:22]
  wire [31:0] n548_I_4_1_1; // @[Top.scala 870:22]
  wire [31:0] n548_I_4_1_2; // @[Top.scala 870:22]
  wire [31:0] n548_I_4_2_0; // @[Top.scala 870:22]
  wire [31:0] n548_I_4_2_1; // @[Top.scala 870:22]
  wire [31:0] n548_I_4_2_2; // @[Top.scala 870:22]
  wire [31:0] n548_I_5_0_0; // @[Top.scala 870:22]
  wire [31:0] n548_I_5_0_1; // @[Top.scala 870:22]
  wire [31:0] n548_I_5_0_2; // @[Top.scala 870:22]
  wire [31:0] n548_I_5_1_0; // @[Top.scala 870:22]
  wire [31:0] n548_I_5_1_1; // @[Top.scala 870:22]
  wire [31:0] n548_I_5_1_2; // @[Top.scala 870:22]
  wire [31:0] n548_I_5_2_0; // @[Top.scala 870:22]
  wire [31:0] n548_I_5_2_1; // @[Top.scala 870:22]
  wire [31:0] n548_I_5_2_2; // @[Top.scala 870:22]
  wire [31:0] n548_I_6_0_0; // @[Top.scala 870:22]
  wire [31:0] n548_I_6_0_1; // @[Top.scala 870:22]
  wire [31:0] n548_I_6_0_2; // @[Top.scala 870:22]
  wire [31:0] n548_I_6_1_0; // @[Top.scala 870:22]
  wire [31:0] n548_I_6_1_1; // @[Top.scala 870:22]
  wire [31:0] n548_I_6_1_2; // @[Top.scala 870:22]
  wire [31:0] n548_I_6_2_0; // @[Top.scala 870:22]
  wire [31:0] n548_I_6_2_1; // @[Top.scala 870:22]
  wire [31:0] n548_I_6_2_2; // @[Top.scala 870:22]
  wire [31:0] n548_I_7_0_0; // @[Top.scala 870:22]
  wire [31:0] n548_I_7_0_1; // @[Top.scala 870:22]
  wire [31:0] n548_I_7_0_2; // @[Top.scala 870:22]
  wire [31:0] n548_I_7_1_0; // @[Top.scala 870:22]
  wire [31:0] n548_I_7_1_1; // @[Top.scala 870:22]
  wire [31:0] n548_I_7_1_2; // @[Top.scala 870:22]
  wire [31:0] n548_I_7_2_0; // @[Top.scala 870:22]
  wire [31:0] n548_I_7_2_1; // @[Top.scala 870:22]
  wire [31:0] n548_I_7_2_2; // @[Top.scala 870:22]
  wire [31:0] n548_O_0_0_0_0; // @[Top.scala 870:22]
  wire [31:0] n548_O_0_0_0_1; // @[Top.scala 870:22]
  wire [31:0] n548_O_0_0_0_2; // @[Top.scala 870:22]
  wire [31:0] n548_O_0_0_1_0; // @[Top.scala 870:22]
  wire [31:0] n548_O_0_0_1_1; // @[Top.scala 870:22]
  wire [31:0] n548_O_0_0_1_2; // @[Top.scala 870:22]
  wire [31:0] n548_O_0_0_2_0; // @[Top.scala 870:22]
  wire [31:0] n548_O_0_0_2_1; // @[Top.scala 870:22]
  wire [31:0] n548_O_0_0_2_2; // @[Top.scala 870:22]
  wire [31:0] n548_O_1_0_0_0; // @[Top.scala 870:22]
  wire [31:0] n548_O_1_0_0_1; // @[Top.scala 870:22]
  wire [31:0] n548_O_1_0_0_2; // @[Top.scala 870:22]
  wire [31:0] n548_O_1_0_1_0; // @[Top.scala 870:22]
  wire [31:0] n548_O_1_0_1_1; // @[Top.scala 870:22]
  wire [31:0] n548_O_1_0_1_2; // @[Top.scala 870:22]
  wire [31:0] n548_O_1_0_2_0; // @[Top.scala 870:22]
  wire [31:0] n548_O_1_0_2_1; // @[Top.scala 870:22]
  wire [31:0] n548_O_1_0_2_2; // @[Top.scala 870:22]
  wire [31:0] n548_O_2_0_0_0; // @[Top.scala 870:22]
  wire [31:0] n548_O_2_0_0_1; // @[Top.scala 870:22]
  wire [31:0] n548_O_2_0_0_2; // @[Top.scala 870:22]
  wire [31:0] n548_O_2_0_1_0; // @[Top.scala 870:22]
  wire [31:0] n548_O_2_0_1_1; // @[Top.scala 870:22]
  wire [31:0] n548_O_2_0_1_2; // @[Top.scala 870:22]
  wire [31:0] n548_O_2_0_2_0; // @[Top.scala 870:22]
  wire [31:0] n548_O_2_0_2_1; // @[Top.scala 870:22]
  wire [31:0] n548_O_2_0_2_2; // @[Top.scala 870:22]
  wire [31:0] n548_O_3_0_0_0; // @[Top.scala 870:22]
  wire [31:0] n548_O_3_0_0_1; // @[Top.scala 870:22]
  wire [31:0] n548_O_3_0_0_2; // @[Top.scala 870:22]
  wire [31:0] n548_O_3_0_1_0; // @[Top.scala 870:22]
  wire [31:0] n548_O_3_0_1_1; // @[Top.scala 870:22]
  wire [31:0] n548_O_3_0_1_2; // @[Top.scala 870:22]
  wire [31:0] n548_O_3_0_2_0; // @[Top.scala 870:22]
  wire [31:0] n548_O_3_0_2_1; // @[Top.scala 870:22]
  wire [31:0] n548_O_3_0_2_2; // @[Top.scala 870:22]
  wire [31:0] n548_O_4_0_0_0; // @[Top.scala 870:22]
  wire [31:0] n548_O_4_0_0_1; // @[Top.scala 870:22]
  wire [31:0] n548_O_4_0_0_2; // @[Top.scala 870:22]
  wire [31:0] n548_O_4_0_1_0; // @[Top.scala 870:22]
  wire [31:0] n548_O_4_0_1_1; // @[Top.scala 870:22]
  wire [31:0] n548_O_4_0_1_2; // @[Top.scala 870:22]
  wire [31:0] n548_O_4_0_2_0; // @[Top.scala 870:22]
  wire [31:0] n548_O_4_0_2_1; // @[Top.scala 870:22]
  wire [31:0] n548_O_4_0_2_2; // @[Top.scala 870:22]
  wire [31:0] n548_O_5_0_0_0; // @[Top.scala 870:22]
  wire [31:0] n548_O_5_0_0_1; // @[Top.scala 870:22]
  wire [31:0] n548_O_5_0_0_2; // @[Top.scala 870:22]
  wire [31:0] n548_O_5_0_1_0; // @[Top.scala 870:22]
  wire [31:0] n548_O_5_0_1_1; // @[Top.scala 870:22]
  wire [31:0] n548_O_5_0_1_2; // @[Top.scala 870:22]
  wire [31:0] n548_O_5_0_2_0; // @[Top.scala 870:22]
  wire [31:0] n548_O_5_0_2_1; // @[Top.scala 870:22]
  wire [31:0] n548_O_5_0_2_2; // @[Top.scala 870:22]
  wire [31:0] n548_O_6_0_0_0; // @[Top.scala 870:22]
  wire [31:0] n548_O_6_0_0_1; // @[Top.scala 870:22]
  wire [31:0] n548_O_6_0_0_2; // @[Top.scala 870:22]
  wire [31:0] n548_O_6_0_1_0; // @[Top.scala 870:22]
  wire [31:0] n548_O_6_0_1_1; // @[Top.scala 870:22]
  wire [31:0] n548_O_6_0_1_2; // @[Top.scala 870:22]
  wire [31:0] n548_O_6_0_2_0; // @[Top.scala 870:22]
  wire [31:0] n548_O_6_0_2_1; // @[Top.scala 870:22]
  wire [31:0] n548_O_6_0_2_2; // @[Top.scala 870:22]
  wire [31:0] n548_O_7_0_0_0; // @[Top.scala 870:22]
  wire [31:0] n548_O_7_0_0_1; // @[Top.scala 870:22]
  wire [31:0] n548_O_7_0_0_2; // @[Top.scala 870:22]
  wire [31:0] n548_O_7_0_1_0; // @[Top.scala 870:22]
  wire [31:0] n548_O_7_0_1_1; // @[Top.scala 870:22]
  wire [31:0] n548_O_7_0_1_2; // @[Top.scala 870:22]
  wire [31:0] n548_O_7_0_2_0; // @[Top.scala 870:22]
  wire [31:0] n548_O_7_0_2_1; // @[Top.scala 870:22]
  wire [31:0] n548_O_7_0_2_2; // @[Top.scala 870:22]
  wire  n555_valid_up; // @[Top.scala 873:22]
  wire  n555_valid_down; // @[Top.scala 873:22]
  wire [31:0] n555_I_0_0_0_0; // @[Top.scala 873:22]
  wire [31:0] n555_I_0_0_0_1; // @[Top.scala 873:22]
  wire [31:0] n555_I_0_0_0_2; // @[Top.scala 873:22]
  wire [31:0] n555_I_0_0_1_0; // @[Top.scala 873:22]
  wire [31:0] n555_I_0_0_1_1; // @[Top.scala 873:22]
  wire [31:0] n555_I_0_0_1_2; // @[Top.scala 873:22]
  wire [31:0] n555_I_0_0_2_0; // @[Top.scala 873:22]
  wire [31:0] n555_I_0_0_2_1; // @[Top.scala 873:22]
  wire [31:0] n555_I_0_0_2_2; // @[Top.scala 873:22]
  wire [31:0] n555_I_1_0_0_0; // @[Top.scala 873:22]
  wire [31:0] n555_I_1_0_0_1; // @[Top.scala 873:22]
  wire [31:0] n555_I_1_0_0_2; // @[Top.scala 873:22]
  wire [31:0] n555_I_1_0_1_0; // @[Top.scala 873:22]
  wire [31:0] n555_I_1_0_1_1; // @[Top.scala 873:22]
  wire [31:0] n555_I_1_0_1_2; // @[Top.scala 873:22]
  wire [31:0] n555_I_1_0_2_0; // @[Top.scala 873:22]
  wire [31:0] n555_I_1_0_2_1; // @[Top.scala 873:22]
  wire [31:0] n555_I_1_0_2_2; // @[Top.scala 873:22]
  wire [31:0] n555_I_2_0_0_0; // @[Top.scala 873:22]
  wire [31:0] n555_I_2_0_0_1; // @[Top.scala 873:22]
  wire [31:0] n555_I_2_0_0_2; // @[Top.scala 873:22]
  wire [31:0] n555_I_2_0_1_0; // @[Top.scala 873:22]
  wire [31:0] n555_I_2_0_1_1; // @[Top.scala 873:22]
  wire [31:0] n555_I_2_0_1_2; // @[Top.scala 873:22]
  wire [31:0] n555_I_2_0_2_0; // @[Top.scala 873:22]
  wire [31:0] n555_I_2_0_2_1; // @[Top.scala 873:22]
  wire [31:0] n555_I_2_0_2_2; // @[Top.scala 873:22]
  wire [31:0] n555_I_3_0_0_0; // @[Top.scala 873:22]
  wire [31:0] n555_I_3_0_0_1; // @[Top.scala 873:22]
  wire [31:0] n555_I_3_0_0_2; // @[Top.scala 873:22]
  wire [31:0] n555_I_3_0_1_0; // @[Top.scala 873:22]
  wire [31:0] n555_I_3_0_1_1; // @[Top.scala 873:22]
  wire [31:0] n555_I_3_0_1_2; // @[Top.scala 873:22]
  wire [31:0] n555_I_3_0_2_0; // @[Top.scala 873:22]
  wire [31:0] n555_I_3_0_2_1; // @[Top.scala 873:22]
  wire [31:0] n555_I_3_0_2_2; // @[Top.scala 873:22]
  wire [31:0] n555_I_4_0_0_0; // @[Top.scala 873:22]
  wire [31:0] n555_I_4_0_0_1; // @[Top.scala 873:22]
  wire [31:0] n555_I_4_0_0_2; // @[Top.scala 873:22]
  wire [31:0] n555_I_4_0_1_0; // @[Top.scala 873:22]
  wire [31:0] n555_I_4_0_1_1; // @[Top.scala 873:22]
  wire [31:0] n555_I_4_0_1_2; // @[Top.scala 873:22]
  wire [31:0] n555_I_4_0_2_0; // @[Top.scala 873:22]
  wire [31:0] n555_I_4_0_2_1; // @[Top.scala 873:22]
  wire [31:0] n555_I_4_0_2_2; // @[Top.scala 873:22]
  wire [31:0] n555_I_5_0_0_0; // @[Top.scala 873:22]
  wire [31:0] n555_I_5_0_0_1; // @[Top.scala 873:22]
  wire [31:0] n555_I_5_0_0_2; // @[Top.scala 873:22]
  wire [31:0] n555_I_5_0_1_0; // @[Top.scala 873:22]
  wire [31:0] n555_I_5_0_1_1; // @[Top.scala 873:22]
  wire [31:0] n555_I_5_0_1_2; // @[Top.scala 873:22]
  wire [31:0] n555_I_5_0_2_0; // @[Top.scala 873:22]
  wire [31:0] n555_I_5_0_2_1; // @[Top.scala 873:22]
  wire [31:0] n555_I_5_0_2_2; // @[Top.scala 873:22]
  wire [31:0] n555_I_6_0_0_0; // @[Top.scala 873:22]
  wire [31:0] n555_I_6_0_0_1; // @[Top.scala 873:22]
  wire [31:0] n555_I_6_0_0_2; // @[Top.scala 873:22]
  wire [31:0] n555_I_6_0_1_0; // @[Top.scala 873:22]
  wire [31:0] n555_I_6_0_1_1; // @[Top.scala 873:22]
  wire [31:0] n555_I_6_0_1_2; // @[Top.scala 873:22]
  wire [31:0] n555_I_6_0_2_0; // @[Top.scala 873:22]
  wire [31:0] n555_I_6_0_2_1; // @[Top.scala 873:22]
  wire [31:0] n555_I_6_0_2_2; // @[Top.scala 873:22]
  wire [31:0] n555_I_7_0_0_0; // @[Top.scala 873:22]
  wire [31:0] n555_I_7_0_0_1; // @[Top.scala 873:22]
  wire [31:0] n555_I_7_0_0_2; // @[Top.scala 873:22]
  wire [31:0] n555_I_7_0_1_0; // @[Top.scala 873:22]
  wire [31:0] n555_I_7_0_1_1; // @[Top.scala 873:22]
  wire [31:0] n555_I_7_0_1_2; // @[Top.scala 873:22]
  wire [31:0] n555_I_7_0_2_0; // @[Top.scala 873:22]
  wire [31:0] n555_I_7_0_2_1; // @[Top.scala 873:22]
  wire [31:0] n555_I_7_0_2_2; // @[Top.scala 873:22]
  wire [31:0] n555_O_0_0_0; // @[Top.scala 873:22]
  wire [31:0] n555_O_0_0_1; // @[Top.scala 873:22]
  wire [31:0] n555_O_0_0_2; // @[Top.scala 873:22]
  wire [31:0] n555_O_0_1_0; // @[Top.scala 873:22]
  wire [31:0] n555_O_0_1_1; // @[Top.scala 873:22]
  wire [31:0] n555_O_0_1_2; // @[Top.scala 873:22]
  wire [31:0] n555_O_0_2_0; // @[Top.scala 873:22]
  wire [31:0] n555_O_0_2_1; // @[Top.scala 873:22]
  wire [31:0] n555_O_0_2_2; // @[Top.scala 873:22]
  wire [31:0] n555_O_1_0_0; // @[Top.scala 873:22]
  wire [31:0] n555_O_1_0_1; // @[Top.scala 873:22]
  wire [31:0] n555_O_1_0_2; // @[Top.scala 873:22]
  wire [31:0] n555_O_1_1_0; // @[Top.scala 873:22]
  wire [31:0] n555_O_1_1_1; // @[Top.scala 873:22]
  wire [31:0] n555_O_1_1_2; // @[Top.scala 873:22]
  wire [31:0] n555_O_1_2_0; // @[Top.scala 873:22]
  wire [31:0] n555_O_1_2_1; // @[Top.scala 873:22]
  wire [31:0] n555_O_1_2_2; // @[Top.scala 873:22]
  wire [31:0] n555_O_2_0_0; // @[Top.scala 873:22]
  wire [31:0] n555_O_2_0_1; // @[Top.scala 873:22]
  wire [31:0] n555_O_2_0_2; // @[Top.scala 873:22]
  wire [31:0] n555_O_2_1_0; // @[Top.scala 873:22]
  wire [31:0] n555_O_2_1_1; // @[Top.scala 873:22]
  wire [31:0] n555_O_2_1_2; // @[Top.scala 873:22]
  wire [31:0] n555_O_2_2_0; // @[Top.scala 873:22]
  wire [31:0] n555_O_2_2_1; // @[Top.scala 873:22]
  wire [31:0] n555_O_2_2_2; // @[Top.scala 873:22]
  wire [31:0] n555_O_3_0_0; // @[Top.scala 873:22]
  wire [31:0] n555_O_3_0_1; // @[Top.scala 873:22]
  wire [31:0] n555_O_3_0_2; // @[Top.scala 873:22]
  wire [31:0] n555_O_3_1_0; // @[Top.scala 873:22]
  wire [31:0] n555_O_3_1_1; // @[Top.scala 873:22]
  wire [31:0] n555_O_3_1_2; // @[Top.scala 873:22]
  wire [31:0] n555_O_3_2_0; // @[Top.scala 873:22]
  wire [31:0] n555_O_3_2_1; // @[Top.scala 873:22]
  wire [31:0] n555_O_3_2_2; // @[Top.scala 873:22]
  wire [31:0] n555_O_4_0_0; // @[Top.scala 873:22]
  wire [31:0] n555_O_4_0_1; // @[Top.scala 873:22]
  wire [31:0] n555_O_4_0_2; // @[Top.scala 873:22]
  wire [31:0] n555_O_4_1_0; // @[Top.scala 873:22]
  wire [31:0] n555_O_4_1_1; // @[Top.scala 873:22]
  wire [31:0] n555_O_4_1_2; // @[Top.scala 873:22]
  wire [31:0] n555_O_4_2_0; // @[Top.scala 873:22]
  wire [31:0] n555_O_4_2_1; // @[Top.scala 873:22]
  wire [31:0] n555_O_4_2_2; // @[Top.scala 873:22]
  wire [31:0] n555_O_5_0_0; // @[Top.scala 873:22]
  wire [31:0] n555_O_5_0_1; // @[Top.scala 873:22]
  wire [31:0] n555_O_5_0_2; // @[Top.scala 873:22]
  wire [31:0] n555_O_5_1_0; // @[Top.scala 873:22]
  wire [31:0] n555_O_5_1_1; // @[Top.scala 873:22]
  wire [31:0] n555_O_5_1_2; // @[Top.scala 873:22]
  wire [31:0] n555_O_5_2_0; // @[Top.scala 873:22]
  wire [31:0] n555_O_5_2_1; // @[Top.scala 873:22]
  wire [31:0] n555_O_5_2_2; // @[Top.scala 873:22]
  wire [31:0] n555_O_6_0_0; // @[Top.scala 873:22]
  wire [31:0] n555_O_6_0_1; // @[Top.scala 873:22]
  wire [31:0] n555_O_6_0_2; // @[Top.scala 873:22]
  wire [31:0] n555_O_6_1_0; // @[Top.scala 873:22]
  wire [31:0] n555_O_6_1_1; // @[Top.scala 873:22]
  wire [31:0] n555_O_6_1_2; // @[Top.scala 873:22]
  wire [31:0] n555_O_6_2_0; // @[Top.scala 873:22]
  wire [31:0] n555_O_6_2_1; // @[Top.scala 873:22]
  wire [31:0] n555_O_6_2_2; // @[Top.scala 873:22]
  wire [31:0] n555_O_7_0_0; // @[Top.scala 873:22]
  wire [31:0] n555_O_7_0_1; // @[Top.scala 873:22]
  wire [31:0] n555_O_7_0_2; // @[Top.scala 873:22]
  wire [31:0] n555_O_7_1_0; // @[Top.scala 873:22]
  wire [31:0] n555_O_7_1_1; // @[Top.scala 873:22]
  wire [31:0] n555_O_7_1_2; // @[Top.scala 873:22]
  wire [31:0] n555_O_7_2_0; // @[Top.scala 873:22]
  wire [31:0] n555_O_7_2_1; // @[Top.scala 873:22]
  wire [31:0] n555_O_7_2_2; // @[Top.scala 873:22]
  wire  n597_clock; // @[Top.scala 876:22]
  wire  n597_reset; // @[Top.scala 876:22]
  wire  n597_valid_up; // @[Top.scala 876:22]
  wire  n597_valid_down; // @[Top.scala 876:22]
  wire [31:0] n597_I_0_0_0; // @[Top.scala 876:22]
  wire [31:0] n597_I_0_0_1; // @[Top.scala 876:22]
  wire [31:0] n597_I_0_0_2; // @[Top.scala 876:22]
  wire [31:0] n597_I_0_1_0; // @[Top.scala 876:22]
  wire [31:0] n597_I_0_1_1; // @[Top.scala 876:22]
  wire [31:0] n597_I_0_1_2; // @[Top.scala 876:22]
  wire [31:0] n597_I_0_2_0; // @[Top.scala 876:22]
  wire [31:0] n597_I_0_2_1; // @[Top.scala 876:22]
  wire [31:0] n597_I_0_2_2; // @[Top.scala 876:22]
  wire [31:0] n597_I_1_0_0; // @[Top.scala 876:22]
  wire [31:0] n597_I_1_0_1; // @[Top.scala 876:22]
  wire [31:0] n597_I_1_0_2; // @[Top.scala 876:22]
  wire [31:0] n597_I_1_1_0; // @[Top.scala 876:22]
  wire [31:0] n597_I_1_1_1; // @[Top.scala 876:22]
  wire [31:0] n597_I_1_1_2; // @[Top.scala 876:22]
  wire [31:0] n597_I_1_2_0; // @[Top.scala 876:22]
  wire [31:0] n597_I_1_2_1; // @[Top.scala 876:22]
  wire [31:0] n597_I_1_2_2; // @[Top.scala 876:22]
  wire [31:0] n597_I_2_0_0; // @[Top.scala 876:22]
  wire [31:0] n597_I_2_0_1; // @[Top.scala 876:22]
  wire [31:0] n597_I_2_0_2; // @[Top.scala 876:22]
  wire [31:0] n597_I_2_1_0; // @[Top.scala 876:22]
  wire [31:0] n597_I_2_1_1; // @[Top.scala 876:22]
  wire [31:0] n597_I_2_1_2; // @[Top.scala 876:22]
  wire [31:0] n597_I_2_2_0; // @[Top.scala 876:22]
  wire [31:0] n597_I_2_2_1; // @[Top.scala 876:22]
  wire [31:0] n597_I_2_2_2; // @[Top.scala 876:22]
  wire [31:0] n597_I_3_0_0; // @[Top.scala 876:22]
  wire [31:0] n597_I_3_0_1; // @[Top.scala 876:22]
  wire [31:0] n597_I_3_0_2; // @[Top.scala 876:22]
  wire [31:0] n597_I_3_1_0; // @[Top.scala 876:22]
  wire [31:0] n597_I_3_1_1; // @[Top.scala 876:22]
  wire [31:0] n597_I_3_1_2; // @[Top.scala 876:22]
  wire [31:0] n597_I_3_2_0; // @[Top.scala 876:22]
  wire [31:0] n597_I_3_2_1; // @[Top.scala 876:22]
  wire [31:0] n597_I_3_2_2; // @[Top.scala 876:22]
  wire [31:0] n597_I_4_0_0; // @[Top.scala 876:22]
  wire [31:0] n597_I_4_0_1; // @[Top.scala 876:22]
  wire [31:0] n597_I_4_0_2; // @[Top.scala 876:22]
  wire [31:0] n597_I_4_1_0; // @[Top.scala 876:22]
  wire [31:0] n597_I_4_1_1; // @[Top.scala 876:22]
  wire [31:0] n597_I_4_1_2; // @[Top.scala 876:22]
  wire [31:0] n597_I_4_2_0; // @[Top.scala 876:22]
  wire [31:0] n597_I_4_2_1; // @[Top.scala 876:22]
  wire [31:0] n597_I_4_2_2; // @[Top.scala 876:22]
  wire [31:0] n597_I_5_0_0; // @[Top.scala 876:22]
  wire [31:0] n597_I_5_0_1; // @[Top.scala 876:22]
  wire [31:0] n597_I_5_0_2; // @[Top.scala 876:22]
  wire [31:0] n597_I_5_1_0; // @[Top.scala 876:22]
  wire [31:0] n597_I_5_1_1; // @[Top.scala 876:22]
  wire [31:0] n597_I_5_1_2; // @[Top.scala 876:22]
  wire [31:0] n597_I_5_2_0; // @[Top.scala 876:22]
  wire [31:0] n597_I_5_2_1; // @[Top.scala 876:22]
  wire [31:0] n597_I_5_2_2; // @[Top.scala 876:22]
  wire [31:0] n597_I_6_0_0; // @[Top.scala 876:22]
  wire [31:0] n597_I_6_0_1; // @[Top.scala 876:22]
  wire [31:0] n597_I_6_0_2; // @[Top.scala 876:22]
  wire [31:0] n597_I_6_1_0; // @[Top.scala 876:22]
  wire [31:0] n597_I_6_1_1; // @[Top.scala 876:22]
  wire [31:0] n597_I_6_1_2; // @[Top.scala 876:22]
  wire [31:0] n597_I_6_2_0; // @[Top.scala 876:22]
  wire [31:0] n597_I_6_2_1; // @[Top.scala 876:22]
  wire [31:0] n597_I_6_2_2; // @[Top.scala 876:22]
  wire [31:0] n597_I_7_0_0; // @[Top.scala 876:22]
  wire [31:0] n597_I_7_0_1; // @[Top.scala 876:22]
  wire [31:0] n597_I_7_0_2; // @[Top.scala 876:22]
  wire [31:0] n597_I_7_1_0; // @[Top.scala 876:22]
  wire [31:0] n597_I_7_1_1; // @[Top.scala 876:22]
  wire [31:0] n597_I_7_1_2; // @[Top.scala 876:22]
  wire [31:0] n597_I_7_2_0; // @[Top.scala 876:22]
  wire [31:0] n597_I_7_2_1; // @[Top.scala 876:22]
  wire [31:0] n597_I_7_2_2; // @[Top.scala 876:22]
  wire [31:0] n597_O_0_0_0; // @[Top.scala 876:22]
  wire [31:0] n597_O_1_0_0; // @[Top.scala 876:22]
  wire [31:0] n597_O_2_0_0; // @[Top.scala 876:22]
  wire [31:0] n597_O_3_0_0; // @[Top.scala 876:22]
  wire [31:0] n597_O_4_0_0; // @[Top.scala 876:22]
  wire [31:0] n597_O_5_0_0; // @[Top.scala 876:22]
  wire [31:0] n597_O_6_0_0; // @[Top.scala 876:22]
  wire [31:0] n597_O_7_0_0; // @[Top.scala 876:22]
  wire  n598_valid_up; // @[Top.scala 879:22]
  wire  n598_valid_down; // @[Top.scala 879:22]
  wire [31:0] n598_I_0_0_0; // @[Top.scala 879:22]
  wire [31:0] n598_I_1_0_0; // @[Top.scala 879:22]
  wire [31:0] n598_I_2_0_0; // @[Top.scala 879:22]
  wire [31:0] n598_I_3_0_0; // @[Top.scala 879:22]
  wire [31:0] n598_I_4_0_0; // @[Top.scala 879:22]
  wire [31:0] n598_I_5_0_0; // @[Top.scala 879:22]
  wire [31:0] n598_I_6_0_0; // @[Top.scala 879:22]
  wire [31:0] n598_I_7_0_0; // @[Top.scala 879:22]
  wire [31:0] n598_O_0_0; // @[Top.scala 879:22]
  wire [31:0] n598_O_1_0; // @[Top.scala 879:22]
  wire [31:0] n598_O_2_0; // @[Top.scala 879:22]
  wire [31:0] n598_O_3_0; // @[Top.scala 879:22]
  wire [31:0] n598_O_4_0; // @[Top.scala 879:22]
  wire [31:0] n598_O_5_0; // @[Top.scala 879:22]
  wire [31:0] n598_O_6_0; // @[Top.scala 879:22]
  wire [31:0] n598_O_7_0; // @[Top.scala 879:22]
  wire  n599_valid_up; // @[Top.scala 882:22]
  wire  n599_valid_down; // @[Top.scala 882:22]
  wire [31:0] n599_I_0_0; // @[Top.scala 882:22]
  wire [31:0] n599_I_1_0; // @[Top.scala 882:22]
  wire [31:0] n599_I_2_0; // @[Top.scala 882:22]
  wire [31:0] n599_I_3_0; // @[Top.scala 882:22]
  wire [31:0] n599_I_4_0; // @[Top.scala 882:22]
  wire [31:0] n599_I_5_0; // @[Top.scala 882:22]
  wire [31:0] n599_I_6_0; // @[Top.scala 882:22]
  wire [31:0] n599_I_7_0; // @[Top.scala 882:22]
  wire [31:0] n599_O_0; // @[Top.scala 882:22]
  wire [31:0] n599_O_1; // @[Top.scala 882:22]
  wire [31:0] n599_O_2; // @[Top.scala 882:22]
  wire [31:0] n599_O_3; // @[Top.scala 882:22]
  wire [31:0] n599_O_4; // @[Top.scala 882:22]
  wire [31:0] n599_O_5; // @[Top.scala 882:22]
  wire [31:0] n599_O_6; // @[Top.scala 882:22]
  wire [31:0] n599_O_7; // @[Top.scala 882:22]
  wire  n600_clock; // @[Top.scala 885:22]
  wire  n600_reset; // @[Top.scala 885:22]
  wire  n600_valid_up; // @[Top.scala 885:22]
  wire  n600_valid_down; // @[Top.scala 885:22]
  wire [31:0] n600_I_0; // @[Top.scala 885:22]
  wire [31:0] n600_I_1; // @[Top.scala 885:22]
  wire [31:0] n600_I_2; // @[Top.scala 885:22]
  wire [31:0] n600_I_3; // @[Top.scala 885:22]
  wire [31:0] n600_I_4; // @[Top.scala 885:22]
  wire [31:0] n600_I_5; // @[Top.scala 885:22]
  wire [31:0] n600_I_6; // @[Top.scala 885:22]
  wire [31:0] n600_I_7; // @[Top.scala 885:22]
  wire [31:0] n600_O_0; // @[Top.scala 885:22]
  wire [31:0] n600_O_1; // @[Top.scala 885:22]
  wire [31:0] n600_O_2; // @[Top.scala 885:22]
  wire [31:0] n600_O_3; // @[Top.scala 885:22]
  wire [31:0] n600_O_4; // @[Top.scala 885:22]
  wire [31:0] n600_O_5; // @[Top.scala 885:22]
  wire [31:0] n600_O_6; // @[Top.scala 885:22]
  wire [31:0] n600_O_7; // @[Top.scala 885:22]
  wire  n601_clock; // @[Top.scala 888:22]
  wire  n601_reset; // @[Top.scala 888:22]
  wire  n601_valid_up; // @[Top.scala 888:22]
  wire  n601_valid_down; // @[Top.scala 888:22]
  wire [31:0] n601_I0_0; // @[Top.scala 888:22]
  wire [31:0] n601_I0_1; // @[Top.scala 888:22]
  wire [31:0] n601_I0_2; // @[Top.scala 888:22]
  wire [31:0] n601_I0_3; // @[Top.scala 888:22]
  wire [31:0] n601_I0_4; // @[Top.scala 888:22]
  wire [31:0] n601_I0_5; // @[Top.scala 888:22]
  wire [31:0] n601_I0_6; // @[Top.scala 888:22]
  wire [31:0] n601_I0_7; // @[Top.scala 888:22]
  wire [31:0] n601_I1_0; // @[Top.scala 888:22]
  wire [31:0] n601_I1_1; // @[Top.scala 888:22]
  wire [31:0] n601_I1_2; // @[Top.scala 888:22]
  wire [31:0] n601_I1_3; // @[Top.scala 888:22]
  wire [31:0] n601_I1_4; // @[Top.scala 888:22]
  wire [31:0] n601_I1_5; // @[Top.scala 888:22]
  wire [31:0] n601_I1_6; // @[Top.scala 888:22]
  wire [31:0] n601_I1_7; // @[Top.scala 888:22]
  wire [31:0] n601_O_0; // @[Top.scala 888:22]
  wire [31:0] n601_O_1; // @[Top.scala 888:22]
  wire [31:0] n601_O_2; // @[Top.scala 888:22]
  wire [31:0] n601_O_3; // @[Top.scala 888:22]
  wire [31:0] n601_O_4; // @[Top.scala 888:22]
  wire [31:0] n601_O_5; // @[Top.scala 888:22]
  wire [31:0] n601_O_6; // @[Top.scala 888:22]
  wire [31:0] n601_O_7; // @[Top.scala 888:22]
  wire  n637_valid_up; // @[Top.scala 892:22]
  wire  n637_valid_down; // @[Top.scala 892:22]
  wire [31:0] n637_I_0_t1b_t0b; // @[Top.scala 892:22]
  wire [31:0] n637_I_0_t1b_t1b; // @[Top.scala 892:22]
  wire [31:0] n637_I_1_t1b_t0b; // @[Top.scala 892:22]
  wire [31:0] n637_I_1_t1b_t1b; // @[Top.scala 892:22]
  wire [31:0] n637_I_2_t1b_t0b; // @[Top.scala 892:22]
  wire [31:0] n637_I_2_t1b_t1b; // @[Top.scala 892:22]
  wire [31:0] n637_I_3_t1b_t0b; // @[Top.scala 892:22]
  wire [31:0] n637_I_3_t1b_t1b; // @[Top.scala 892:22]
  wire [31:0] n637_I_4_t1b_t0b; // @[Top.scala 892:22]
  wire [31:0] n637_I_4_t1b_t1b; // @[Top.scala 892:22]
  wire [31:0] n637_I_5_t1b_t0b; // @[Top.scala 892:22]
  wire [31:0] n637_I_5_t1b_t1b; // @[Top.scala 892:22]
  wire [31:0] n637_I_6_t1b_t0b; // @[Top.scala 892:22]
  wire [31:0] n637_I_6_t1b_t1b; // @[Top.scala 892:22]
  wire [31:0] n637_I_7_t1b_t0b; // @[Top.scala 892:22]
  wire [31:0] n637_I_7_t1b_t1b; // @[Top.scala 892:22]
  wire [31:0] n637_O_0; // @[Top.scala 892:22]
  wire [31:0] n637_O_1; // @[Top.scala 892:22]
  wire [31:0] n637_O_2; // @[Top.scala 892:22]
  wire [31:0] n637_O_3; // @[Top.scala 892:22]
  wire [31:0] n637_O_4; // @[Top.scala 892:22]
  wire [31:0] n637_O_5; // @[Top.scala 892:22]
  wire [31:0] n637_O_6; // @[Top.scala 892:22]
  wire [31:0] n637_O_7; // @[Top.scala 892:22]
  wire  n638_clock; // @[Top.scala 895:22]
  wire  n638_reset; // @[Top.scala 895:22]
  wire  n638_valid_up; // @[Top.scala 895:22]
  wire  n638_valid_down; // @[Top.scala 895:22]
  wire [31:0] n638_I_0; // @[Top.scala 895:22]
  wire [31:0] n638_I_1; // @[Top.scala 895:22]
  wire [31:0] n638_I_2; // @[Top.scala 895:22]
  wire [31:0] n638_I_3; // @[Top.scala 895:22]
  wire [31:0] n638_I_4; // @[Top.scala 895:22]
  wire [31:0] n638_I_5; // @[Top.scala 895:22]
  wire [31:0] n638_I_6; // @[Top.scala 895:22]
  wire [31:0] n638_I_7; // @[Top.scala 895:22]
  wire [31:0] n638_O_0; // @[Top.scala 895:22]
  wire [31:0] n638_O_1; // @[Top.scala 895:22]
  wire [31:0] n638_O_2; // @[Top.scala 895:22]
  wire [31:0] n638_O_3; // @[Top.scala 895:22]
  wire [31:0] n638_O_4; // @[Top.scala 895:22]
  wire [31:0] n638_O_5; // @[Top.scala 895:22]
  wire [31:0] n638_O_6; // @[Top.scala 895:22]
  wire [31:0] n638_O_7; // @[Top.scala 895:22]
  wire  n639_clock; // @[Top.scala 898:22]
  wire  n639_reset; // @[Top.scala 898:22]
  wire  n639_valid_up; // @[Top.scala 898:22]
  wire  n639_valid_down; // @[Top.scala 898:22]
  wire [31:0] n639_I_0; // @[Top.scala 898:22]
  wire [31:0] n639_I_1; // @[Top.scala 898:22]
  wire [31:0] n639_I_2; // @[Top.scala 898:22]
  wire [31:0] n639_I_3; // @[Top.scala 898:22]
  wire [31:0] n639_I_4; // @[Top.scala 898:22]
  wire [31:0] n639_I_5; // @[Top.scala 898:22]
  wire [31:0] n639_I_6; // @[Top.scala 898:22]
  wire [31:0] n639_I_7; // @[Top.scala 898:22]
  wire [31:0] n639_O_0; // @[Top.scala 898:22]
  wire [31:0] n639_O_1; // @[Top.scala 898:22]
  wire [31:0] n639_O_2; // @[Top.scala 898:22]
  wire [31:0] n639_O_3; // @[Top.scala 898:22]
  wire [31:0] n639_O_4; // @[Top.scala 898:22]
  wire [31:0] n639_O_5; // @[Top.scala 898:22]
  wire [31:0] n639_O_6; // @[Top.scala 898:22]
  wire [31:0] n639_O_7; // @[Top.scala 898:22]
  wire  n640_clock; // @[Top.scala 901:22]
  wire  n640_valid_up; // @[Top.scala 901:22]
  wire  n640_valid_down; // @[Top.scala 901:22]
  wire [31:0] n640_I_0; // @[Top.scala 901:22]
  wire [31:0] n640_I_1; // @[Top.scala 901:22]
  wire [31:0] n640_I_2; // @[Top.scala 901:22]
  wire [31:0] n640_I_3; // @[Top.scala 901:22]
  wire [31:0] n640_I_4; // @[Top.scala 901:22]
  wire [31:0] n640_I_5; // @[Top.scala 901:22]
  wire [31:0] n640_I_6; // @[Top.scala 901:22]
  wire [31:0] n640_I_7; // @[Top.scala 901:22]
  wire [31:0] n640_O_0; // @[Top.scala 901:22]
  wire [31:0] n640_O_1; // @[Top.scala 901:22]
  wire [31:0] n640_O_2; // @[Top.scala 901:22]
  wire [31:0] n640_O_3; // @[Top.scala 901:22]
  wire [31:0] n640_O_4; // @[Top.scala 901:22]
  wire [31:0] n640_O_5; // @[Top.scala 901:22]
  wire [31:0] n640_O_6; // @[Top.scala 901:22]
  wire [31:0] n640_O_7; // @[Top.scala 901:22]
  wire  n641_clock; // @[Top.scala 904:22]
  wire  n641_valid_up; // @[Top.scala 904:22]
  wire  n641_valid_down; // @[Top.scala 904:22]
  wire [31:0] n641_I_0; // @[Top.scala 904:22]
  wire [31:0] n641_I_1; // @[Top.scala 904:22]
  wire [31:0] n641_I_2; // @[Top.scala 904:22]
  wire [31:0] n641_I_3; // @[Top.scala 904:22]
  wire [31:0] n641_I_4; // @[Top.scala 904:22]
  wire [31:0] n641_I_5; // @[Top.scala 904:22]
  wire [31:0] n641_I_6; // @[Top.scala 904:22]
  wire [31:0] n641_I_7; // @[Top.scala 904:22]
  wire [31:0] n641_O_0; // @[Top.scala 904:22]
  wire [31:0] n641_O_1; // @[Top.scala 904:22]
  wire [31:0] n641_O_2; // @[Top.scala 904:22]
  wire [31:0] n641_O_3; // @[Top.scala 904:22]
  wire [31:0] n641_O_4; // @[Top.scala 904:22]
  wire [31:0] n641_O_5; // @[Top.scala 904:22]
  wire [31:0] n641_O_6; // @[Top.scala 904:22]
  wire [31:0] n641_O_7; // @[Top.scala 904:22]
  wire  n642_valid_up; // @[Top.scala 907:22]
  wire  n642_valid_down; // @[Top.scala 907:22]
  wire [31:0] n642_I0_0; // @[Top.scala 907:22]
  wire [31:0] n642_I0_1; // @[Top.scala 907:22]
  wire [31:0] n642_I0_2; // @[Top.scala 907:22]
  wire [31:0] n642_I0_3; // @[Top.scala 907:22]
  wire [31:0] n642_I0_4; // @[Top.scala 907:22]
  wire [31:0] n642_I0_5; // @[Top.scala 907:22]
  wire [31:0] n642_I0_6; // @[Top.scala 907:22]
  wire [31:0] n642_I0_7; // @[Top.scala 907:22]
  wire [31:0] n642_I1_0; // @[Top.scala 907:22]
  wire [31:0] n642_I1_1; // @[Top.scala 907:22]
  wire [31:0] n642_I1_2; // @[Top.scala 907:22]
  wire [31:0] n642_I1_3; // @[Top.scala 907:22]
  wire [31:0] n642_I1_4; // @[Top.scala 907:22]
  wire [31:0] n642_I1_5; // @[Top.scala 907:22]
  wire [31:0] n642_I1_6; // @[Top.scala 907:22]
  wire [31:0] n642_I1_7; // @[Top.scala 907:22]
  wire [31:0] n642_O_0_0; // @[Top.scala 907:22]
  wire [31:0] n642_O_0_1; // @[Top.scala 907:22]
  wire [31:0] n642_O_1_0; // @[Top.scala 907:22]
  wire [31:0] n642_O_1_1; // @[Top.scala 907:22]
  wire [31:0] n642_O_2_0; // @[Top.scala 907:22]
  wire [31:0] n642_O_2_1; // @[Top.scala 907:22]
  wire [31:0] n642_O_3_0; // @[Top.scala 907:22]
  wire [31:0] n642_O_3_1; // @[Top.scala 907:22]
  wire [31:0] n642_O_4_0; // @[Top.scala 907:22]
  wire [31:0] n642_O_4_1; // @[Top.scala 907:22]
  wire [31:0] n642_O_5_0; // @[Top.scala 907:22]
  wire [31:0] n642_O_5_1; // @[Top.scala 907:22]
  wire [31:0] n642_O_6_0; // @[Top.scala 907:22]
  wire [31:0] n642_O_6_1; // @[Top.scala 907:22]
  wire [31:0] n642_O_7_0; // @[Top.scala 907:22]
  wire [31:0] n642_O_7_1; // @[Top.scala 907:22]
  wire  n649_valid_up; // @[Top.scala 911:22]
  wire  n649_valid_down; // @[Top.scala 911:22]
  wire [31:0] n649_I0_0_0; // @[Top.scala 911:22]
  wire [31:0] n649_I0_0_1; // @[Top.scala 911:22]
  wire [31:0] n649_I0_1_0; // @[Top.scala 911:22]
  wire [31:0] n649_I0_1_1; // @[Top.scala 911:22]
  wire [31:0] n649_I0_2_0; // @[Top.scala 911:22]
  wire [31:0] n649_I0_2_1; // @[Top.scala 911:22]
  wire [31:0] n649_I0_3_0; // @[Top.scala 911:22]
  wire [31:0] n649_I0_3_1; // @[Top.scala 911:22]
  wire [31:0] n649_I0_4_0; // @[Top.scala 911:22]
  wire [31:0] n649_I0_4_1; // @[Top.scala 911:22]
  wire [31:0] n649_I0_5_0; // @[Top.scala 911:22]
  wire [31:0] n649_I0_5_1; // @[Top.scala 911:22]
  wire [31:0] n649_I0_6_0; // @[Top.scala 911:22]
  wire [31:0] n649_I0_6_1; // @[Top.scala 911:22]
  wire [31:0] n649_I0_7_0; // @[Top.scala 911:22]
  wire [31:0] n649_I0_7_1; // @[Top.scala 911:22]
  wire [31:0] n649_I1_0; // @[Top.scala 911:22]
  wire [31:0] n649_I1_1; // @[Top.scala 911:22]
  wire [31:0] n649_I1_2; // @[Top.scala 911:22]
  wire [31:0] n649_I1_3; // @[Top.scala 911:22]
  wire [31:0] n649_I1_4; // @[Top.scala 911:22]
  wire [31:0] n649_I1_5; // @[Top.scala 911:22]
  wire [31:0] n649_I1_6; // @[Top.scala 911:22]
  wire [31:0] n649_I1_7; // @[Top.scala 911:22]
  wire [31:0] n649_O_0_0; // @[Top.scala 911:22]
  wire [31:0] n649_O_0_1; // @[Top.scala 911:22]
  wire [31:0] n649_O_0_2; // @[Top.scala 911:22]
  wire [31:0] n649_O_1_0; // @[Top.scala 911:22]
  wire [31:0] n649_O_1_1; // @[Top.scala 911:22]
  wire [31:0] n649_O_1_2; // @[Top.scala 911:22]
  wire [31:0] n649_O_2_0; // @[Top.scala 911:22]
  wire [31:0] n649_O_2_1; // @[Top.scala 911:22]
  wire [31:0] n649_O_2_2; // @[Top.scala 911:22]
  wire [31:0] n649_O_3_0; // @[Top.scala 911:22]
  wire [31:0] n649_O_3_1; // @[Top.scala 911:22]
  wire [31:0] n649_O_3_2; // @[Top.scala 911:22]
  wire [31:0] n649_O_4_0; // @[Top.scala 911:22]
  wire [31:0] n649_O_4_1; // @[Top.scala 911:22]
  wire [31:0] n649_O_4_2; // @[Top.scala 911:22]
  wire [31:0] n649_O_5_0; // @[Top.scala 911:22]
  wire [31:0] n649_O_5_1; // @[Top.scala 911:22]
  wire [31:0] n649_O_5_2; // @[Top.scala 911:22]
  wire [31:0] n649_O_6_0; // @[Top.scala 911:22]
  wire [31:0] n649_O_6_1; // @[Top.scala 911:22]
  wire [31:0] n649_O_6_2; // @[Top.scala 911:22]
  wire [31:0] n649_O_7_0; // @[Top.scala 911:22]
  wire [31:0] n649_O_7_1; // @[Top.scala 911:22]
  wire [31:0] n649_O_7_2; // @[Top.scala 911:22]
  wire  n658_valid_up; // @[Top.scala 915:22]
  wire  n658_valid_down; // @[Top.scala 915:22]
  wire [31:0] n658_I_0_0; // @[Top.scala 915:22]
  wire [31:0] n658_I_0_1; // @[Top.scala 915:22]
  wire [31:0] n658_I_0_2; // @[Top.scala 915:22]
  wire [31:0] n658_I_1_0; // @[Top.scala 915:22]
  wire [31:0] n658_I_1_1; // @[Top.scala 915:22]
  wire [31:0] n658_I_1_2; // @[Top.scala 915:22]
  wire [31:0] n658_I_2_0; // @[Top.scala 915:22]
  wire [31:0] n658_I_2_1; // @[Top.scala 915:22]
  wire [31:0] n658_I_2_2; // @[Top.scala 915:22]
  wire [31:0] n658_I_3_0; // @[Top.scala 915:22]
  wire [31:0] n658_I_3_1; // @[Top.scala 915:22]
  wire [31:0] n658_I_3_2; // @[Top.scala 915:22]
  wire [31:0] n658_I_4_0; // @[Top.scala 915:22]
  wire [31:0] n658_I_4_1; // @[Top.scala 915:22]
  wire [31:0] n658_I_4_2; // @[Top.scala 915:22]
  wire [31:0] n658_I_5_0; // @[Top.scala 915:22]
  wire [31:0] n658_I_5_1; // @[Top.scala 915:22]
  wire [31:0] n658_I_5_2; // @[Top.scala 915:22]
  wire [31:0] n658_I_6_0; // @[Top.scala 915:22]
  wire [31:0] n658_I_6_1; // @[Top.scala 915:22]
  wire [31:0] n658_I_6_2; // @[Top.scala 915:22]
  wire [31:0] n658_I_7_0; // @[Top.scala 915:22]
  wire [31:0] n658_I_7_1; // @[Top.scala 915:22]
  wire [31:0] n658_I_7_2; // @[Top.scala 915:22]
  wire [31:0] n658_O_0_0_0; // @[Top.scala 915:22]
  wire [31:0] n658_O_0_0_1; // @[Top.scala 915:22]
  wire [31:0] n658_O_0_0_2; // @[Top.scala 915:22]
  wire [31:0] n658_O_1_0_0; // @[Top.scala 915:22]
  wire [31:0] n658_O_1_0_1; // @[Top.scala 915:22]
  wire [31:0] n658_O_1_0_2; // @[Top.scala 915:22]
  wire [31:0] n658_O_2_0_0; // @[Top.scala 915:22]
  wire [31:0] n658_O_2_0_1; // @[Top.scala 915:22]
  wire [31:0] n658_O_2_0_2; // @[Top.scala 915:22]
  wire [31:0] n658_O_3_0_0; // @[Top.scala 915:22]
  wire [31:0] n658_O_3_0_1; // @[Top.scala 915:22]
  wire [31:0] n658_O_3_0_2; // @[Top.scala 915:22]
  wire [31:0] n658_O_4_0_0; // @[Top.scala 915:22]
  wire [31:0] n658_O_4_0_1; // @[Top.scala 915:22]
  wire [31:0] n658_O_4_0_2; // @[Top.scala 915:22]
  wire [31:0] n658_O_5_0_0; // @[Top.scala 915:22]
  wire [31:0] n658_O_5_0_1; // @[Top.scala 915:22]
  wire [31:0] n658_O_5_0_2; // @[Top.scala 915:22]
  wire [31:0] n658_O_6_0_0; // @[Top.scala 915:22]
  wire [31:0] n658_O_6_0_1; // @[Top.scala 915:22]
  wire [31:0] n658_O_6_0_2; // @[Top.scala 915:22]
  wire [31:0] n658_O_7_0_0; // @[Top.scala 915:22]
  wire [31:0] n658_O_7_0_1; // @[Top.scala 915:22]
  wire [31:0] n658_O_7_0_2; // @[Top.scala 915:22]
  wire  n665_valid_up; // @[Top.scala 918:22]
  wire  n665_valid_down; // @[Top.scala 918:22]
  wire [31:0] n665_I_0_0_0; // @[Top.scala 918:22]
  wire [31:0] n665_I_0_0_1; // @[Top.scala 918:22]
  wire [31:0] n665_I_0_0_2; // @[Top.scala 918:22]
  wire [31:0] n665_I_1_0_0; // @[Top.scala 918:22]
  wire [31:0] n665_I_1_0_1; // @[Top.scala 918:22]
  wire [31:0] n665_I_1_0_2; // @[Top.scala 918:22]
  wire [31:0] n665_I_2_0_0; // @[Top.scala 918:22]
  wire [31:0] n665_I_2_0_1; // @[Top.scala 918:22]
  wire [31:0] n665_I_2_0_2; // @[Top.scala 918:22]
  wire [31:0] n665_I_3_0_0; // @[Top.scala 918:22]
  wire [31:0] n665_I_3_0_1; // @[Top.scala 918:22]
  wire [31:0] n665_I_3_0_2; // @[Top.scala 918:22]
  wire [31:0] n665_I_4_0_0; // @[Top.scala 918:22]
  wire [31:0] n665_I_4_0_1; // @[Top.scala 918:22]
  wire [31:0] n665_I_4_0_2; // @[Top.scala 918:22]
  wire [31:0] n665_I_5_0_0; // @[Top.scala 918:22]
  wire [31:0] n665_I_5_0_1; // @[Top.scala 918:22]
  wire [31:0] n665_I_5_0_2; // @[Top.scala 918:22]
  wire [31:0] n665_I_6_0_0; // @[Top.scala 918:22]
  wire [31:0] n665_I_6_0_1; // @[Top.scala 918:22]
  wire [31:0] n665_I_6_0_2; // @[Top.scala 918:22]
  wire [31:0] n665_I_7_0_0; // @[Top.scala 918:22]
  wire [31:0] n665_I_7_0_1; // @[Top.scala 918:22]
  wire [31:0] n665_I_7_0_2; // @[Top.scala 918:22]
  wire [31:0] n665_O_0_0; // @[Top.scala 918:22]
  wire [31:0] n665_O_0_1; // @[Top.scala 918:22]
  wire [31:0] n665_O_0_2; // @[Top.scala 918:22]
  wire [31:0] n665_O_1_0; // @[Top.scala 918:22]
  wire [31:0] n665_O_1_1; // @[Top.scala 918:22]
  wire [31:0] n665_O_1_2; // @[Top.scala 918:22]
  wire [31:0] n665_O_2_0; // @[Top.scala 918:22]
  wire [31:0] n665_O_2_1; // @[Top.scala 918:22]
  wire [31:0] n665_O_2_2; // @[Top.scala 918:22]
  wire [31:0] n665_O_3_0; // @[Top.scala 918:22]
  wire [31:0] n665_O_3_1; // @[Top.scala 918:22]
  wire [31:0] n665_O_3_2; // @[Top.scala 918:22]
  wire [31:0] n665_O_4_0; // @[Top.scala 918:22]
  wire [31:0] n665_O_4_1; // @[Top.scala 918:22]
  wire [31:0] n665_O_4_2; // @[Top.scala 918:22]
  wire [31:0] n665_O_5_0; // @[Top.scala 918:22]
  wire [31:0] n665_O_5_1; // @[Top.scala 918:22]
  wire [31:0] n665_O_5_2; // @[Top.scala 918:22]
  wire [31:0] n665_O_6_0; // @[Top.scala 918:22]
  wire [31:0] n665_O_6_1; // @[Top.scala 918:22]
  wire [31:0] n665_O_6_2; // @[Top.scala 918:22]
  wire [31:0] n665_O_7_0; // @[Top.scala 918:22]
  wire [31:0] n665_O_7_1; // @[Top.scala 918:22]
  wire [31:0] n665_O_7_2; // @[Top.scala 918:22]
  wire  n666_clock; // @[Top.scala 921:22]
  wire  n666_valid_up; // @[Top.scala 921:22]
  wire  n666_valid_down; // @[Top.scala 921:22]
  wire [31:0] n666_I_0; // @[Top.scala 921:22]
  wire [31:0] n666_I_1; // @[Top.scala 921:22]
  wire [31:0] n666_I_2; // @[Top.scala 921:22]
  wire [31:0] n666_I_3; // @[Top.scala 921:22]
  wire [31:0] n666_I_4; // @[Top.scala 921:22]
  wire [31:0] n666_I_5; // @[Top.scala 921:22]
  wire [31:0] n666_I_6; // @[Top.scala 921:22]
  wire [31:0] n666_I_7; // @[Top.scala 921:22]
  wire [31:0] n666_O_0; // @[Top.scala 921:22]
  wire [31:0] n666_O_1; // @[Top.scala 921:22]
  wire [31:0] n666_O_2; // @[Top.scala 921:22]
  wire [31:0] n666_O_3; // @[Top.scala 921:22]
  wire [31:0] n666_O_4; // @[Top.scala 921:22]
  wire [31:0] n666_O_5; // @[Top.scala 921:22]
  wire [31:0] n666_O_6; // @[Top.scala 921:22]
  wire [31:0] n666_O_7; // @[Top.scala 921:22]
  wire  n667_clock; // @[Top.scala 924:22]
  wire  n667_valid_up; // @[Top.scala 924:22]
  wire  n667_valid_down; // @[Top.scala 924:22]
  wire [31:0] n667_I_0; // @[Top.scala 924:22]
  wire [31:0] n667_I_1; // @[Top.scala 924:22]
  wire [31:0] n667_I_2; // @[Top.scala 924:22]
  wire [31:0] n667_I_3; // @[Top.scala 924:22]
  wire [31:0] n667_I_4; // @[Top.scala 924:22]
  wire [31:0] n667_I_5; // @[Top.scala 924:22]
  wire [31:0] n667_I_6; // @[Top.scala 924:22]
  wire [31:0] n667_I_7; // @[Top.scala 924:22]
  wire [31:0] n667_O_0; // @[Top.scala 924:22]
  wire [31:0] n667_O_1; // @[Top.scala 924:22]
  wire [31:0] n667_O_2; // @[Top.scala 924:22]
  wire [31:0] n667_O_3; // @[Top.scala 924:22]
  wire [31:0] n667_O_4; // @[Top.scala 924:22]
  wire [31:0] n667_O_5; // @[Top.scala 924:22]
  wire [31:0] n667_O_6; // @[Top.scala 924:22]
  wire [31:0] n667_O_7; // @[Top.scala 924:22]
  wire  n668_valid_up; // @[Top.scala 927:22]
  wire  n668_valid_down; // @[Top.scala 927:22]
  wire [31:0] n668_I0_0; // @[Top.scala 927:22]
  wire [31:0] n668_I0_1; // @[Top.scala 927:22]
  wire [31:0] n668_I0_2; // @[Top.scala 927:22]
  wire [31:0] n668_I0_3; // @[Top.scala 927:22]
  wire [31:0] n668_I0_4; // @[Top.scala 927:22]
  wire [31:0] n668_I0_5; // @[Top.scala 927:22]
  wire [31:0] n668_I0_6; // @[Top.scala 927:22]
  wire [31:0] n668_I0_7; // @[Top.scala 927:22]
  wire [31:0] n668_I1_0; // @[Top.scala 927:22]
  wire [31:0] n668_I1_1; // @[Top.scala 927:22]
  wire [31:0] n668_I1_2; // @[Top.scala 927:22]
  wire [31:0] n668_I1_3; // @[Top.scala 927:22]
  wire [31:0] n668_I1_4; // @[Top.scala 927:22]
  wire [31:0] n668_I1_5; // @[Top.scala 927:22]
  wire [31:0] n668_I1_6; // @[Top.scala 927:22]
  wire [31:0] n668_I1_7; // @[Top.scala 927:22]
  wire [31:0] n668_O_0_0; // @[Top.scala 927:22]
  wire [31:0] n668_O_0_1; // @[Top.scala 927:22]
  wire [31:0] n668_O_1_0; // @[Top.scala 927:22]
  wire [31:0] n668_O_1_1; // @[Top.scala 927:22]
  wire [31:0] n668_O_2_0; // @[Top.scala 927:22]
  wire [31:0] n668_O_2_1; // @[Top.scala 927:22]
  wire [31:0] n668_O_3_0; // @[Top.scala 927:22]
  wire [31:0] n668_O_3_1; // @[Top.scala 927:22]
  wire [31:0] n668_O_4_0; // @[Top.scala 927:22]
  wire [31:0] n668_O_4_1; // @[Top.scala 927:22]
  wire [31:0] n668_O_5_0; // @[Top.scala 927:22]
  wire [31:0] n668_O_5_1; // @[Top.scala 927:22]
  wire [31:0] n668_O_6_0; // @[Top.scala 927:22]
  wire [31:0] n668_O_6_1; // @[Top.scala 927:22]
  wire [31:0] n668_O_7_0; // @[Top.scala 927:22]
  wire [31:0] n668_O_7_1; // @[Top.scala 927:22]
  wire  n675_valid_up; // @[Top.scala 931:22]
  wire  n675_valid_down; // @[Top.scala 931:22]
  wire [31:0] n675_I0_0_0; // @[Top.scala 931:22]
  wire [31:0] n675_I0_0_1; // @[Top.scala 931:22]
  wire [31:0] n675_I0_1_0; // @[Top.scala 931:22]
  wire [31:0] n675_I0_1_1; // @[Top.scala 931:22]
  wire [31:0] n675_I0_2_0; // @[Top.scala 931:22]
  wire [31:0] n675_I0_2_1; // @[Top.scala 931:22]
  wire [31:0] n675_I0_3_0; // @[Top.scala 931:22]
  wire [31:0] n675_I0_3_1; // @[Top.scala 931:22]
  wire [31:0] n675_I0_4_0; // @[Top.scala 931:22]
  wire [31:0] n675_I0_4_1; // @[Top.scala 931:22]
  wire [31:0] n675_I0_5_0; // @[Top.scala 931:22]
  wire [31:0] n675_I0_5_1; // @[Top.scala 931:22]
  wire [31:0] n675_I0_6_0; // @[Top.scala 931:22]
  wire [31:0] n675_I0_6_1; // @[Top.scala 931:22]
  wire [31:0] n675_I0_7_0; // @[Top.scala 931:22]
  wire [31:0] n675_I0_7_1; // @[Top.scala 931:22]
  wire [31:0] n675_I1_0; // @[Top.scala 931:22]
  wire [31:0] n675_I1_1; // @[Top.scala 931:22]
  wire [31:0] n675_I1_2; // @[Top.scala 931:22]
  wire [31:0] n675_I1_3; // @[Top.scala 931:22]
  wire [31:0] n675_I1_4; // @[Top.scala 931:22]
  wire [31:0] n675_I1_5; // @[Top.scala 931:22]
  wire [31:0] n675_I1_6; // @[Top.scala 931:22]
  wire [31:0] n675_I1_7; // @[Top.scala 931:22]
  wire [31:0] n675_O_0_0; // @[Top.scala 931:22]
  wire [31:0] n675_O_0_1; // @[Top.scala 931:22]
  wire [31:0] n675_O_0_2; // @[Top.scala 931:22]
  wire [31:0] n675_O_1_0; // @[Top.scala 931:22]
  wire [31:0] n675_O_1_1; // @[Top.scala 931:22]
  wire [31:0] n675_O_1_2; // @[Top.scala 931:22]
  wire [31:0] n675_O_2_0; // @[Top.scala 931:22]
  wire [31:0] n675_O_2_1; // @[Top.scala 931:22]
  wire [31:0] n675_O_2_2; // @[Top.scala 931:22]
  wire [31:0] n675_O_3_0; // @[Top.scala 931:22]
  wire [31:0] n675_O_3_1; // @[Top.scala 931:22]
  wire [31:0] n675_O_3_2; // @[Top.scala 931:22]
  wire [31:0] n675_O_4_0; // @[Top.scala 931:22]
  wire [31:0] n675_O_4_1; // @[Top.scala 931:22]
  wire [31:0] n675_O_4_2; // @[Top.scala 931:22]
  wire [31:0] n675_O_5_0; // @[Top.scala 931:22]
  wire [31:0] n675_O_5_1; // @[Top.scala 931:22]
  wire [31:0] n675_O_5_2; // @[Top.scala 931:22]
  wire [31:0] n675_O_6_0; // @[Top.scala 931:22]
  wire [31:0] n675_O_6_1; // @[Top.scala 931:22]
  wire [31:0] n675_O_6_2; // @[Top.scala 931:22]
  wire [31:0] n675_O_7_0; // @[Top.scala 931:22]
  wire [31:0] n675_O_7_1; // @[Top.scala 931:22]
  wire [31:0] n675_O_7_2; // @[Top.scala 931:22]
  wire  n684_valid_up; // @[Top.scala 935:22]
  wire  n684_valid_down; // @[Top.scala 935:22]
  wire [31:0] n684_I_0_0; // @[Top.scala 935:22]
  wire [31:0] n684_I_0_1; // @[Top.scala 935:22]
  wire [31:0] n684_I_0_2; // @[Top.scala 935:22]
  wire [31:0] n684_I_1_0; // @[Top.scala 935:22]
  wire [31:0] n684_I_1_1; // @[Top.scala 935:22]
  wire [31:0] n684_I_1_2; // @[Top.scala 935:22]
  wire [31:0] n684_I_2_0; // @[Top.scala 935:22]
  wire [31:0] n684_I_2_1; // @[Top.scala 935:22]
  wire [31:0] n684_I_2_2; // @[Top.scala 935:22]
  wire [31:0] n684_I_3_0; // @[Top.scala 935:22]
  wire [31:0] n684_I_3_1; // @[Top.scala 935:22]
  wire [31:0] n684_I_3_2; // @[Top.scala 935:22]
  wire [31:0] n684_I_4_0; // @[Top.scala 935:22]
  wire [31:0] n684_I_4_1; // @[Top.scala 935:22]
  wire [31:0] n684_I_4_2; // @[Top.scala 935:22]
  wire [31:0] n684_I_5_0; // @[Top.scala 935:22]
  wire [31:0] n684_I_5_1; // @[Top.scala 935:22]
  wire [31:0] n684_I_5_2; // @[Top.scala 935:22]
  wire [31:0] n684_I_6_0; // @[Top.scala 935:22]
  wire [31:0] n684_I_6_1; // @[Top.scala 935:22]
  wire [31:0] n684_I_6_2; // @[Top.scala 935:22]
  wire [31:0] n684_I_7_0; // @[Top.scala 935:22]
  wire [31:0] n684_I_7_1; // @[Top.scala 935:22]
  wire [31:0] n684_I_7_2; // @[Top.scala 935:22]
  wire [31:0] n684_O_0_0_0; // @[Top.scala 935:22]
  wire [31:0] n684_O_0_0_1; // @[Top.scala 935:22]
  wire [31:0] n684_O_0_0_2; // @[Top.scala 935:22]
  wire [31:0] n684_O_1_0_0; // @[Top.scala 935:22]
  wire [31:0] n684_O_1_0_1; // @[Top.scala 935:22]
  wire [31:0] n684_O_1_0_2; // @[Top.scala 935:22]
  wire [31:0] n684_O_2_0_0; // @[Top.scala 935:22]
  wire [31:0] n684_O_2_0_1; // @[Top.scala 935:22]
  wire [31:0] n684_O_2_0_2; // @[Top.scala 935:22]
  wire [31:0] n684_O_3_0_0; // @[Top.scala 935:22]
  wire [31:0] n684_O_3_0_1; // @[Top.scala 935:22]
  wire [31:0] n684_O_3_0_2; // @[Top.scala 935:22]
  wire [31:0] n684_O_4_0_0; // @[Top.scala 935:22]
  wire [31:0] n684_O_4_0_1; // @[Top.scala 935:22]
  wire [31:0] n684_O_4_0_2; // @[Top.scala 935:22]
  wire [31:0] n684_O_5_0_0; // @[Top.scala 935:22]
  wire [31:0] n684_O_5_0_1; // @[Top.scala 935:22]
  wire [31:0] n684_O_5_0_2; // @[Top.scala 935:22]
  wire [31:0] n684_O_6_0_0; // @[Top.scala 935:22]
  wire [31:0] n684_O_6_0_1; // @[Top.scala 935:22]
  wire [31:0] n684_O_6_0_2; // @[Top.scala 935:22]
  wire [31:0] n684_O_7_0_0; // @[Top.scala 935:22]
  wire [31:0] n684_O_7_0_1; // @[Top.scala 935:22]
  wire [31:0] n684_O_7_0_2; // @[Top.scala 935:22]
  wire  n691_valid_up; // @[Top.scala 938:22]
  wire  n691_valid_down; // @[Top.scala 938:22]
  wire [31:0] n691_I_0_0_0; // @[Top.scala 938:22]
  wire [31:0] n691_I_0_0_1; // @[Top.scala 938:22]
  wire [31:0] n691_I_0_0_2; // @[Top.scala 938:22]
  wire [31:0] n691_I_1_0_0; // @[Top.scala 938:22]
  wire [31:0] n691_I_1_0_1; // @[Top.scala 938:22]
  wire [31:0] n691_I_1_0_2; // @[Top.scala 938:22]
  wire [31:0] n691_I_2_0_0; // @[Top.scala 938:22]
  wire [31:0] n691_I_2_0_1; // @[Top.scala 938:22]
  wire [31:0] n691_I_2_0_2; // @[Top.scala 938:22]
  wire [31:0] n691_I_3_0_0; // @[Top.scala 938:22]
  wire [31:0] n691_I_3_0_1; // @[Top.scala 938:22]
  wire [31:0] n691_I_3_0_2; // @[Top.scala 938:22]
  wire [31:0] n691_I_4_0_0; // @[Top.scala 938:22]
  wire [31:0] n691_I_4_0_1; // @[Top.scala 938:22]
  wire [31:0] n691_I_4_0_2; // @[Top.scala 938:22]
  wire [31:0] n691_I_5_0_0; // @[Top.scala 938:22]
  wire [31:0] n691_I_5_0_1; // @[Top.scala 938:22]
  wire [31:0] n691_I_5_0_2; // @[Top.scala 938:22]
  wire [31:0] n691_I_6_0_0; // @[Top.scala 938:22]
  wire [31:0] n691_I_6_0_1; // @[Top.scala 938:22]
  wire [31:0] n691_I_6_0_2; // @[Top.scala 938:22]
  wire [31:0] n691_I_7_0_0; // @[Top.scala 938:22]
  wire [31:0] n691_I_7_0_1; // @[Top.scala 938:22]
  wire [31:0] n691_I_7_0_2; // @[Top.scala 938:22]
  wire [31:0] n691_O_0_0; // @[Top.scala 938:22]
  wire [31:0] n691_O_0_1; // @[Top.scala 938:22]
  wire [31:0] n691_O_0_2; // @[Top.scala 938:22]
  wire [31:0] n691_O_1_0; // @[Top.scala 938:22]
  wire [31:0] n691_O_1_1; // @[Top.scala 938:22]
  wire [31:0] n691_O_1_2; // @[Top.scala 938:22]
  wire [31:0] n691_O_2_0; // @[Top.scala 938:22]
  wire [31:0] n691_O_2_1; // @[Top.scala 938:22]
  wire [31:0] n691_O_2_2; // @[Top.scala 938:22]
  wire [31:0] n691_O_3_0; // @[Top.scala 938:22]
  wire [31:0] n691_O_3_1; // @[Top.scala 938:22]
  wire [31:0] n691_O_3_2; // @[Top.scala 938:22]
  wire [31:0] n691_O_4_0; // @[Top.scala 938:22]
  wire [31:0] n691_O_4_1; // @[Top.scala 938:22]
  wire [31:0] n691_O_4_2; // @[Top.scala 938:22]
  wire [31:0] n691_O_5_0; // @[Top.scala 938:22]
  wire [31:0] n691_O_5_1; // @[Top.scala 938:22]
  wire [31:0] n691_O_5_2; // @[Top.scala 938:22]
  wire [31:0] n691_O_6_0; // @[Top.scala 938:22]
  wire [31:0] n691_O_6_1; // @[Top.scala 938:22]
  wire [31:0] n691_O_6_2; // @[Top.scala 938:22]
  wire [31:0] n691_O_7_0; // @[Top.scala 938:22]
  wire [31:0] n691_O_7_1; // @[Top.scala 938:22]
  wire [31:0] n691_O_7_2; // @[Top.scala 938:22]
  wire  n692_valid_up; // @[Top.scala 941:22]
  wire  n692_valid_down; // @[Top.scala 941:22]
  wire [31:0] n692_I0_0_0; // @[Top.scala 941:22]
  wire [31:0] n692_I0_0_1; // @[Top.scala 941:22]
  wire [31:0] n692_I0_0_2; // @[Top.scala 941:22]
  wire [31:0] n692_I0_1_0; // @[Top.scala 941:22]
  wire [31:0] n692_I0_1_1; // @[Top.scala 941:22]
  wire [31:0] n692_I0_1_2; // @[Top.scala 941:22]
  wire [31:0] n692_I0_2_0; // @[Top.scala 941:22]
  wire [31:0] n692_I0_2_1; // @[Top.scala 941:22]
  wire [31:0] n692_I0_2_2; // @[Top.scala 941:22]
  wire [31:0] n692_I0_3_0; // @[Top.scala 941:22]
  wire [31:0] n692_I0_3_1; // @[Top.scala 941:22]
  wire [31:0] n692_I0_3_2; // @[Top.scala 941:22]
  wire [31:0] n692_I0_4_0; // @[Top.scala 941:22]
  wire [31:0] n692_I0_4_1; // @[Top.scala 941:22]
  wire [31:0] n692_I0_4_2; // @[Top.scala 941:22]
  wire [31:0] n692_I0_5_0; // @[Top.scala 941:22]
  wire [31:0] n692_I0_5_1; // @[Top.scala 941:22]
  wire [31:0] n692_I0_5_2; // @[Top.scala 941:22]
  wire [31:0] n692_I0_6_0; // @[Top.scala 941:22]
  wire [31:0] n692_I0_6_1; // @[Top.scala 941:22]
  wire [31:0] n692_I0_6_2; // @[Top.scala 941:22]
  wire [31:0] n692_I0_7_0; // @[Top.scala 941:22]
  wire [31:0] n692_I0_7_1; // @[Top.scala 941:22]
  wire [31:0] n692_I0_7_2; // @[Top.scala 941:22]
  wire [31:0] n692_I1_0_0; // @[Top.scala 941:22]
  wire [31:0] n692_I1_0_1; // @[Top.scala 941:22]
  wire [31:0] n692_I1_0_2; // @[Top.scala 941:22]
  wire [31:0] n692_I1_1_0; // @[Top.scala 941:22]
  wire [31:0] n692_I1_1_1; // @[Top.scala 941:22]
  wire [31:0] n692_I1_1_2; // @[Top.scala 941:22]
  wire [31:0] n692_I1_2_0; // @[Top.scala 941:22]
  wire [31:0] n692_I1_2_1; // @[Top.scala 941:22]
  wire [31:0] n692_I1_2_2; // @[Top.scala 941:22]
  wire [31:0] n692_I1_3_0; // @[Top.scala 941:22]
  wire [31:0] n692_I1_3_1; // @[Top.scala 941:22]
  wire [31:0] n692_I1_3_2; // @[Top.scala 941:22]
  wire [31:0] n692_I1_4_0; // @[Top.scala 941:22]
  wire [31:0] n692_I1_4_1; // @[Top.scala 941:22]
  wire [31:0] n692_I1_4_2; // @[Top.scala 941:22]
  wire [31:0] n692_I1_5_0; // @[Top.scala 941:22]
  wire [31:0] n692_I1_5_1; // @[Top.scala 941:22]
  wire [31:0] n692_I1_5_2; // @[Top.scala 941:22]
  wire [31:0] n692_I1_6_0; // @[Top.scala 941:22]
  wire [31:0] n692_I1_6_1; // @[Top.scala 941:22]
  wire [31:0] n692_I1_6_2; // @[Top.scala 941:22]
  wire [31:0] n692_I1_7_0; // @[Top.scala 941:22]
  wire [31:0] n692_I1_7_1; // @[Top.scala 941:22]
  wire [31:0] n692_I1_7_2; // @[Top.scala 941:22]
  wire [31:0] n692_O_0_0_0; // @[Top.scala 941:22]
  wire [31:0] n692_O_0_0_1; // @[Top.scala 941:22]
  wire [31:0] n692_O_0_0_2; // @[Top.scala 941:22]
  wire [31:0] n692_O_0_1_0; // @[Top.scala 941:22]
  wire [31:0] n692_O_0_1_1; // @[Top.scala 941:22]
  wire [31:0] n692_O_0_1_2; // @[Top.scala 941:22]
  wire [31:0] n692_O_1_0_0; // @[Top.scala 941:22]
  wire [31:0] n692_O_1_0_1; // @[Top.scala 941:22]
  wire [31:0] n692_O_1_0_2; // @[Top.scala 941:22]
  wire [31:0] n692_O_1_1_0; // @[Top.scala 941:22]
  wire [31:0] n692_O_1_1_1; // @[Top.scala 941:22]
  wire [31:0] n692_O_1_1_2; // @[Top.scala 941:22]
  wire [31:0] n692_O_2_0_0; // @[Top.scala 941:22]
  wire [31:0] n692_O_2_0_1; // @[Top.scala 941:22]
  wire [31:0] n692_O_2_0_2; // @[Top.scala 941:22]
  wire [31:0] n692_O_2_1_0; // @[Top.scala 941:22]
  wire [31:0] n692_O_2_1_1; // @[Top.scala 941:22]
  wire [31:0] n692_O_2_1_2; // @[Top.scala 941:22]
  wire [31:0] n692_O_3_0_0; // @[Top.scala 941:22]
  wire [31:0] n692_O_3_0_1; // @[Top.scala 941:22]
  wire [31:0] n692_O_3_0_2; // @[Top.scala 941:22]
  wire [31:0] n692_O_3_1_0; // @[Top.scala 941:22]
  wire [31:0] n692_O_3_1_1; // @[Top.scala 941:22]
  wire [31:0] n692_O_3_1_2; // @[Top.scala 941:22]
  wire [31:0] n692_O_4_0_0; // @[Top.scala 941:22]
  wire [31:0] n692_O_4_0_1; // @[Top.scala 941:22]
  wire [31:0] n692_O_4_0_2; // @[Top.scala 941:22]
  wire [31:0] n692_O_4_1_0; // @[Top.scala 941:22]
  wire [31:0] n692_O_4_1_1; // @[Top.scala 941:22]
  wire [31:0] n692_O_4_1_2; // @[Top.scala 941:22]
  wire [31:0] n692_O_5_0_0; // @[Top.scala 941:22]
  wire [31:0] n692_O_5_0_1; // @[Top.scala 941:22]
  wire [31:0] n692_O_5_0_2; // @[Top.scala 941:22]
  wire [31:0] n692_O_5_1_0; // @[Top.scala 941:22]
  wire [31:0] n692_O_5_1_1; // @[Top.scala 941:22]
  wire [31:0] n692_O_5_1_2; // @[Top.scala 941:22]
  wire [31:0] n692_O_6_0_0; // @[Top.scala 941:22]
  wire [31:0] n692_O_6_0_1; // @[Top.scala 941:22]
  wire [31:0] n692_O_6_0_2; // @[Top.scala 941:22]
  wire [31:0] n692_O_6_1_0; // @[Top.scala 941:22]
  wire [31:0] n692_O_6_1_1; // @[Top.scala 941:22]
  wire [31:0] n692_O_6_1_2; // @[Top.scala 941:22]
  wire [31:0] n692_O_7_0_0; // @[Top.scala 941:22]
  wire [31:0] n692_O_7_0_1; // @[Top.scala 941:22]
  wire [31:0] n692_O_7_0_2; // @[Top.scala 941:22]
  wire [31:0] n692_O_7_1_0; // @[Top.scala 941:22]
  wire [31:0] n692_O_7_1_1; // @[Top.scala 941:22]
  wire [31:0] n692_O_7_1_2; // @[Top.scala 941:22]
  wire  n699_clock; // @[Top.scala 945:22]
  wire  n699_valid_up; // @[Top.scala 945:22]
  wire  n699_valid_down; // @[Top.scala 945:22]
  wire [31:0] n699_I_0; // @[Top.scala 945:22]
  wire [31:0] n699_I_1; // @[Top.scala 945:22]
  wire [31:0] n699_I_2; // @[Top.scala 945:22]
  wire [31:0] n699_I_3; // @[Top.scala 945:22]
  wire [31:0] n699_I_4; // @[Top.scala 945:22]
  wire [31:0] n699_I_5; // @[Top.scala 945:22]
  wire [31:0] n699_I_6; // @[Top.scala 945:22]
  wire [31:0] n699_I_7; // @[Top.scala 945:22]
  wire [31:0] n699_O_0; // @[Top.scala 945:22]
  wire [31:0] n699_O_1; // @[Top.scala 945:22]
  wire [31:0] n699_O_2; // @[Top.scala 945:22]
  wire [31:0] n699_O_3; // @[Top.scala 945:22]
  wire [31:0] n699_O_4; // @[Top.scala 945:22]
  wire [31:0] n699_O_5; // @[Top.scala 945:22]
  wire [31:0] n699_O_6; // @[Top.scala 945:22]
  wire [31:0] n699_O_7; // @[Top.scala 945:22]
  wire  n700_clock; // @[Top.scala 948:22]
  wire  n700_valid_up; // @[Top.scala 948:22]
  wire  n700_valid_down; // @[Top.scala 948:22]
  wire [31:0] n700_I_0; // @[Top.scala 948:22]
  wire [31:0] n700_I_1; // @[Top.scala 948:22]
  wire [31:0] n700_I_2; // @[Top.scala 948:22]
  wire [31:0] n700_I_3; // @[Top.scala 948:22]
  wire [31:0] n700_I_4; // @[Top.scala 948:22]
  wire [31:0] n700_I_5; // @[Top.scala 948:22]
  wire [31:0] n700_I_6; // @[Top.scala 948:22]
  wire [31:0] n700_I_7; // @[Top.scala 948:22]
  wire [31:0] n700_O_0; // @[Top.scala 948:22]
  wire [31:0] n700_O_1; // @[Top.scala 948:22]
  wire [31:0] n700_O_2; // @[Top.scala 948:22]
  wire [31:0] n700_O_3; // @[Top.scala 948:22]
  wire [31:0] n700_O_4; // @[Top.scala 948:22]
  wire [31:0] n700_O_5; // @[Top.scala 948:22]
  wire [31:0] n700_O_6; // @[Top.scala 948:22]
  wire [31:0] n700_O_7; // @[Top.scala 948:22]
  wire  n701_valid_up; // @[Top.scala 951:22]
  wire  n701_valid_down; // @[Top.scala 951:22]
  wire [31:0] n701_I0_0; // @[Top.scala 951:22]
  wire [31:0] n701_I0_1; // @[Top.scala 951:22]
  wire [31:0] n701_I0_2; // @[Top.scala 951:22]
  wire [31:0] n701_I0_3; // @[Top.scala 951:22]
  wire [31:0] n701_I0_4; // @[Top.scala 951:22]
  wire [31:0] n701_I0_5; // @[Top.scala 951:22]
  wire [31:0] n701_I0_6; // @[Top.scala 951:22]
  wire [31:0] n701_I0_7; // @[Top.scala 951:22]
  wire [31:0] n701_I1_0; // @[Top.scala 951:22]
  wire [31:0] n701_I1_1; // @[Top.scala 951:22]
  wire [31:0] n701_I1_2; // @[Top.scala 951:22]
  wire [31:0] n701_I1_3; // @[Top.scala 951:22]
  wire [31:0] n701_I1_4; // @[Top.scala 951:22]
  wire [31:0] n701_I1_5; // @[Top.scala 951:22]
  wire [31:0] n701_I1_6; // @[Top.scala 951:22]
  wire [31:0] n701_I1_7; // @[Top.scala 951:22]
  wire [31:0] n701_O_0_0; // @[Top.scala 951:22]
  wire [31:0] n701_O_0_1; // @[Top.scala 951:22]
  wire [31:0] n701_O_1_0; // @[Top.scala 951:22]
  wire [31:0] n701_O_1_1; // @[Top.scala 951:22]
  wire [31:0] n701_O_2_0; // @[Top.scala 951:22]
  wire [31:0] n701_O_2_1; // @[Top.scala 951:22]
  wire [31:0] n701_O_3_0; // @[Top.scala 951:22]
  wire [31:0] n701_O_3_1; // @[Top.scala 951:22]
  wire [31:0] n701_O_4_0; // @[Top.scala 951:22]
  wire [31:0] n701_O_4_1; // @[Top.scala 951:22]
  wire [31:0] n701_O_5_0; // @[Top.scala 951:22]
  wire [31:0] n701_O_5_1; // @[Top.scala 951:22]
  wire [31:0] n701_O_6_0; // @[Top.scala 951:22]
  wire [31:0] n701_O_6_1; // @[Top.scala 951:22]
  wire [31:0] n701_O_7_0; // @[Top.scala 951:22]
  wire [31:0] n701_O_7_1; // @[Top.scala 951:22]
  wire  n708_valid_up; // @[Top.scala 955:22]
  wire  n708_valid_down; // @[Top.scala 955:22]
  wire [31:0] n708_I0_0_0; // @[Top.scala 955:22]
  wire [31:0] n708_I0_0_1; // @[Top.scala 955:22]
  wire [31:0] n708_I0_1_0; // @[Top.scala 955:22]
  wire [31:0] n708_I0_1_1; // @[Top.scala 955:22]
  wire [31:0] n708_I0_2_0; // @[Top.scala 955:22]
  wire [31:0] n708_I0_2_1; // @[Top.scala 955:22]
  wire [31:0] n708_I0_3_0; // @[Top.scala 955:22]
  wire [31:0] n708_I0_3_1; // @[Top.scala 955:22]
  wire [31:0] n708_I0_4_0; // @[Top.scala 955:22]
  wire [31:0] n708_I0_4_1; // @[Top.scala 955:22]
  wire [31:0] n708_I0_5_0; // @[Top.scala 955:22]
  wire [31:0] n708_I0_5_1; // @[Top.scala 955:22]
  wire [31:0] n708_I0_6_0; // @[Top.scala 955:22]
  wire [31:0] n708_I0_6_1; // @[Top.scala 955:22]
  wire [31:0] n708_I0_7_0; // @[Top.scala 955:22]
  wire [31:0] n708_I0_7_1; // @[Top.scala 955:22]
  wire [31:0] n708_I1_0; // @[Top.scala 955:22]
  wire [31:0] n708_I1_1; // @[Top.scala 955:22]
  wire [31:0] n708_I1_2; // @[Top.scala 955:22]
  wire [31:0] n708_I1_3; // @[Top.scala 955:22]
  wire [31:0] n708_I1_4; // @[Top.scala 955:22]
  wire [31:0] n708_I1_5; // @[Top.scala 955:22]
  wire [31:0] n708_I1_6; // @[Top.scala 955:22]
  wire [31:0] n708_I1_7; // @[Top.scala 955:22]
  wire [31:0] n708_O_0_0; // @[Top.scala 955:22]
  wire [31:0] n708_O_0_1; // @[Top.scala 955:22]
  wire [31:0] n708_O_0_2; // @[Top.scala 955:22]
  wire [31:0] n708_O_1_0; // @[Top.scala 955:22]
  wire [31:0] n708_O_1_1; // @[Top.scala 955:22]
  wire [31:0] n708_O_1_2; // @[Top.scala 955:22]
  wire [31:0] n708_O_2_0; // @[Top.scala 955:22]
  wire [31:0] n708_O_2_1; // @[Top.scala 955:22]
  wire [31:0] n708_O_2_2; // @[Top.scala 955:22]
  wire [31:0] n708_O_3_0; // @[Top.scala 955:22]
  wire [31:0] n708_O_3_1; // @[Top.scala 955:22]
  wire [31:0] n708_O_3_2; // @[Top.scala 955:22]
  wire [31:0] n708_O_4_0; // @[Top.scala 955:22]
  wire [31:0] n708_O_4_1; // @[Top.scala 955:22]
  wire [31:0] n708_O_4_2; // @[Top.scala 955:22]
  wire [31:0] n708_O_5_0; // @[Top.scala 955:22]
  wire [31:0] n708_O_5_1; // @[Top.scala 955:22]
  wire [31:0] n708_O_5_2; // @[Top.scala 955:22]
  wire [31:0] n708_O_6_0; // @[Top.scala 955:22]
  wire [31:0] n708_O_6_1; // @[Top.scala 955:22]
  wire [31:0] n708_O_6_2; // @[Top.scala 955:22]
  wire [31:0] n708_O_7_0; // @[Top.scala 955:22]
  wire [31:0] n708_O_7_1; // @[Top.scala 955:22]
  wire [31:0] n708_O_7_2; // @[Top.scala 955:22]
  wire  n717_valid_up; // @[Top.scala 959:22]
  wire  n717_valid_down; // @[Top.scala 959:22]
  wire [31:0] n717_I_0_0; // @[Top.scala 959:22]
  wire [31:0] n717_I_0_1; // @[Top.scala 959:22]
  wire [31:0] n717_I_0_2; // @[Top.scala 959:22]
  wire [31:0] n717_I_1_0; // @[Top.scala 959:22]
  wire [31:0] n717_I_1_1; // @[Top.scala 959:22]
  wire [31:0] n717_I_1_2; // @[Top.scala 959:22]
  wire [31:0] n717_I_2_0; // @[Top.scala 959:22]
  wire [31:0] n717_I_2_1; // @[Top.scala 959:22]
  wire [31:0] n717_I_2_2; // @[Top.scala 959:22]
  wire [31:0] n717_I_3_0; // @[Top.scala 959:22]
  wire [31:0] n717_I_3_1; // @[Top.scala 959:22]
  wire [31:0] n717_I_3_2; // @[Top.scala 959:22]
  wire [31:0] n717_I_4_0; // @[Top.scala 959:22]
  wire [31:0] n717_I_4_1; // @[Top.scala 959:22]
  wire [31:0] n717_I_4_2; // @[Top.scala 959:22]
  wire [31:0] n717_I_5_0; // @[Top.scala 959:22]
  wire [31:0] n717_I_5_1; // @[Top.scala 959:22]
  wire [31:0] n717_I_5_2; // @[Top.scala 959:22]
  wire [31:0] n717_I_6_0; // @[Top.scala 959:22]
  wire [31:0] n717_I_6_1; // @[Top.scala 959:22]
  wire [31:0] n717_I_6_2; // @[Top.scala 959:22]
  wire [31:0] n717_I_7_0; // @[Top.scala 959:22]
  wire [31:0] n717_I_7_1; // @[Top.scala 959:22]
  wire [31:0] n717_I_7_2; // @[Top.scala 959:22]
  wire [31:0] n717_O_0_0_0; // @[Top.scala 959:22]
  wire [31:0] n717_O_0_0_1; // @[Top.scala 959:22]
  wire [31:0] n717_O_0_0_2; // @[Top.scala 959:22]
  wire [31:0] n717_O_1_0_0; // @[Top.scala 959:22]
  wire [31:0] n717_O_1_0_1; // @[Top.scala 959:22]
  wire [31:0] n717_O_1_0_2; // @[Top.scala 959:22]
  wire [31:0] n717_O_2_0_0; // @[Top.scala 959:22]
  wire [31:0] n717_O_2_0_1; // @[Top.scala 959:22]
  wire [31:0] n717_O_2_0_2; // @[Top.scala 959:22]
  wire [31:0] n717_O_3_0_0; // @[Top.scala 959:22]
  wire [31:0] n717_O_3_0_1; // @[Top.scala 959:22]
  wire [31:0] n717_O_3_0_2; // @[Top.scala 959:22]
  wire [31:0] n717_O_4_0_0; // @[Top.scala 959:22]
  wire [31:0] n717_O_4_0_1; // @[Top.scala 959:22]
  wire [31:0] n717_O_4_0_2; // @[Top.scala 959:22]
  wire [31:0] n717_O_5_0_0; // @[Top.scala 959:22]
  wire [31:0] n717_O_5_0_1; // @[Top.scala 959:22]
  wire [31:0] n717_O_5_0_2; // @[Top.scala 959:22]
  wire [31:0] n717_O_6_0_0; // @[Top.scala 959:22]
  wire [31:0] n717_O_6_0_1; // @[Top.scala 959:22]
  wire [31:0] n717_O_6_0_2; // @[Top.scala 959:22]
  wire [31:0] n717_O_7_0_0; // @[Top.scala 959:22]
  wire [31:0] n717_O_7_0_1; // @[Top.scala 959:22]
  wire [31:0] n717_O_7_0_2; // @[Top.scala 959:22]
  wire  n724_valid_up; // @[Top.scala 962:22]
  wire  n724_valid_down; // @[Top.scala 962:22]
  wire [31:0] n724_I_0_0_0; // @[Top.scala 962:22]
  wire [31:0] n724_I_0_0_1; // @[Top.scala 962:22]
  wire [31:0] n724_I_0_0_2; // @[Top.scala 962:22]
  wire [31:0] n724_I_1_0_0; // @[Top.scala 962:22]
  wire [31:0] n724_I_1_0_1; // @[Top.scala 962:22]
  wire [31:0] n724_I_1_0_2; // @[Top.scala 962:22]
  wire [31:0] n724_I_2_0_0; // @[Top.scala 962:22]
  wire [31:0] n724_I_2_0_1; // @[Top.scala 962:22]
  wire [31:0] n724_I_2_0_2; // @[Top.scala 962:22]
  wire [31:0] n724_I_3_0_0; // @[Top.scala 962:22]
  wire [31:0] n724_I_3_0_1; // @[Top.scala 962:22]
  wire [31:0] n724_I_3_0_2; // @[Top.scala 962:22]
  wire [31:0] n724_I_4_0_0; // @[Top.scala 962:22]
  wire [31:0] n724_I_4_0_1; // @[Top.scala 962:22]
  wire [31:0] n724_I_4_0_2; // @[Top.scala 962:22]
  wire [31:0] n724_I_5_0_0; // @[Top.scala 962:22]
  wire [31:0] n724_I_5_0_1; // @[Top.scala 962:22]
  wire [31:0] n724_I_5_0_2; // @[Top.scala 962:22]
  wire [31:0] n724_I_6_0_0; // @[Top.scala 962:22]
  wire [31:0] n724_I_6_0_1; // @[Top.scala 962:22]
  wire [31:0] n724_I_6_0_2; // @[Top.scala 962:22]
  wire [31:0] n724_I_7_0_0; // @[Top.scala 962:22]
  wire [31:0] n724_I_7_0_1; // @[Top.scala 962:22]
  wire [31:0] n724_I_7_0_2; // @[Top.scala 962:22]
  wire [31:0] n724_O_0_0; // @[Top.scala 962:22]
  wire [31:0] n724_O_0_1; // @[Top.scala 962:22]
  wire [31:0] n724_O_0_2; // @[Top.scala 962:22]
  wire [31:0] n724_O_1_0; // @[Top.scala 962:22]
  wire [31:0] n724_O_1_1; // @[Top.scala 962:22]
  wire [31:0] n724_O_1_2; // @[Top.scala 962:22]
  wire [31:0] n724_O_2_0; // @[Top.scala 962:22]
  wire [31:0] n724_O_2_1; // @[Top.scala 962:22]
  wire [31:0] n724_O_2_2; // @[Top.scala 962:22]
  wire [31:0] n724_O_3_0; // @[Top.scala 962:22]
  wire [31:0] n724_O_3_1; // @[Top.scala 962:22]
  wire [31:0] n724_O_3_2; // @[Top.scala 962:22]
  wire [31:0] n724_O_4_0; // @[Top.scala 962:22]
  wire [31:0] n724_O_4_1; // @[Top.scala 962:22]
  wire [31:0] n724_O_4_2; // @[Top.scala 962:22]
  wire [31:0] n724_O_5_0; // @[Top.scala 962:22]
  wire [31:0] n724_O_5_1; // @[Top.scala 962:22]
  wire [31:0] n724_O_5_2; // @[Top.scala 962:22]
  wire [31:0] n724_O_6_0; // @[Top.scala 962:22]
  wire [31:0] n724_O_6_1; // @[Top.scala 962:22]
  wire [31:0] n724_O_6_2; // @[Top.scala 962:22]
  wire [31:0] n724_O_7_0; // @[Top.scala 962:22]
  wire [31:0] n724_O_7_1; // @[Top.scala 962:22]
  wire [31:0] n724_O_7_2; // @[Top.scala 962:22]
  wire  n725_valid_up; // @[Top.scala 965:22]
  wire  n725_valid_down; // @[Top.scala 965:22]
  wire [31:0] n725_I0_0_0_0; // @[Top.scala 965:22]
  wire [31:0] n725_I0_0_0_1; // @[Top.scala 965:22]
  wire [31:0] n725_I0_0_0_2; // @[Top.scala 965:22]
  wire [31:0] n725_I0_0_1_0; // @[Top.scala 965:22]
  wire [31:0] n725_I0_0_1_1; // @[Top.scala 965:22]
  wire [31:0] n725_I0_0_1_2; // @[Top.scala 965:22]
  wire [31:0] n725_I0_1_0_0; // @[Top.scala 965:22]
  wire [31:0] n725_I0_1_0_1; // @[Top.scala 965:22]
  wire [31:0] n725_I0_1_0_2; // @[Top.scala 965:22]
  wire [31:0] n725_I0_1_1_0; // @[Top.scala 965:22]
  wire [31:0] n725_I0_1_1_1; // @[Top.scala 965:22]
  wire [31:0] n725_I0_1_1_2; // @[Top.scala 965:22]
  wire [31:0] n725_I0_2_0_0; // @[Top.scala 965:22]
  wire [31:0] n725_I0_2_0_1; // @[Top.scala 965:22]
  wire [31:0] n725_I0_2_0_2; // @[Top.scala 965:22]
  wire [31:0] n725_I0_2_1_0; // @[Top.scala 965:22]
  wire [31:0] n725_I0_2_1_1; // @[Top.scala 965:22]
  wire [31:0] n725_I0_2_1_2; // @[Top.scala 965:22]
  wire [31:0] n725_I0_3_0_0; // @[Top.scala 965:22]
  wire [31:0] n725_I0_3_0_1; // @[Top.scala 965:22]
  wire [31:0] n725_I0_3_0_2; // @[Top.scala 965:22]
  wire [31:0] n725_I0_3_1_0; // @[Top.scala 965:22]
  wire [31:0] n725_I0_3_1_1; // @[Top.scala 965:22]
  wire [31:0] n725_I0_3_1_2; // @[Top.scala 965:22]
  wire [31:0] n725_I0_4_0_0; // @[Top.scala 965:22]
  wire [31:0] n725_I0_4_0_1; // @[Top.scala 965:22]
  wire [31:0] n725_I0_4_0_2; // @[Top.scala 965:22]
  wire [31:0] n725_I0_4_1_0; // @[Top.scala 965:22]
  wire [31:0] n725_I0_4_1_1; // @[Top.scala 965:22]
  wire [31:0] n725_I0_4_1_2; // @[Top.scala 965:22]
  wire [31:0] n725_I0_5_0_0; // @[Top.scala 965:22]
  wire [31:0] n725_I0_5_0_1; // @[Top.scala 965:22]
  wire [31:0] n725_I0_5_0_2; // @[Top.scala 965:22]
  wire [31:0] n725_I0_5_1_0; // @[Top.scala 965:22]
  wire [31:0] n725_I0_5_1_1; // @[Top.scala 965:22]
  wire [31:0] n725_I0_5_1_2; // @[Top.scala 965:22]
  wire [31:0] n725_I0_6_0_0; // @[Top.scala 965:22]
  wire [31:0] n725_I0_6_0_1; // @[Top.scala 965:22]
  wire [31:0] n725_I0_6_0_2; // @[Top.scala 965:22]
  wire [31:0] n725_I0_6_1_0; // @[Top.scala 965:22]
  wire [31:0] n725_I0_6_1_1; // @[Top.scala 965:22]
  wire [31:0] n725_I0_6_1_2; // @[Top.scala 965:22]
  wire [31:0] n725_I0_7_0_0; // @[Top.scala 965:22]
  wire [31:0] n725_I0_7_0_1; // @[Top.scala 965:22]
  wire [31:0] n725_I0_7_0_2; // @[Top.scala 965:22]
  wire [31:0] n725_I0_7_1_0; // @[Top.scala 965:22]
  wire [31:0] n725_I0_7_1_1; // @[Top.scala 965:22]
  wire [31:0] n725_I0_7_1_2; // @[Top.scala 965:22]
  wire [31:0] n725_I1_0_0; // @[Top.scala 965:22]
  wire [31:0] n725_I1_0_1; // @[Top.scala 965:22]
  wire [31:0] n725_I1_0_2; // @[Top.scala 965:22]
  wire [31:0] n725_I1_1_0; // @[Top.scala 965:22]
  wire [31:0] n725_I1_1_1; // @[Top.scala 965:22]
  wire [31:0] n725_I1_1_2; // @[Top.scala 965:22]
  wire [31:0] n725_I1_2_0; // @[Top.scala 965:22]
  wire [31:0] n725_I1_2_1; // @[Top.scala 965:22]
  wire [31:0] n725_I1_2_2; // @[Top.scala 965:22]
  wire [31:0] n725_I1_3_0; // @[Top.scala 965:22]
  wire [31:0] n725_I1_3_1; // @[Top.scala 965:22]
  wire [31:0] n725_I1_3_2; // @[Top.scala 965:22]
  wire [31:0] n725_I1_4_0; // @[Top.scala 965:22]
  wire [31:0] n725_I1_4_1; // @[Top.scala 965:22]
  wire [31:0] n725_I1_4_2; // @[Top.scala 965:22]
  wire [31:0] n725_I1_5_0; // @[Top.scala 965:22]
  wire [31:0] n725_I1_5_1; // @[Top.scala 965:22]
  wire [31:0] n725_I1_5_2; // @[Top.scala 965:22]
  wire [31:0] n725_I1_6_0; // @[Top.scala 965:22]
  wire [31:0] n725_I1_6_1; // @[Top.scala 965:22]
  wire [31:0] n725_I1_6_2; // @[Top.scala 965:22]
  wire [31:0] n725_I1_7_0; // @[Top.scala 965:22]
  wire [31:0] n725_I1_7_1; // @[Top.scala 965:22]
  wire [31:0] n725_I1_7_2; // @[Top.scala 965:22]
  wire [31:0] n725_O_0_0_0; // @[Top.scala 965:22]
  wire [31:0] n725_O_0_0_1; // @[Top.scala 965:22]
  wire [31:0] n725_O_0_0_2; // @[Top.scala 965:22]
  wire [31:0] n725_O_0_1_0; // @[Top.scala 965:22]
  wire [31:0] n725_O_0_1_1; // @[Top.scala 965:22]
  wire [31:0] n725_O_0_1_2; // @[Top.scala 965:22]
  wire [31:0] n725_O_0_2_0; // @[Top.scala 965:22]
  wire [31:0] n725_O_0_2_1; // @[Top.scala 965:22]
  wire [31:0] n725_O_0_2_2; // @[Top.scala 965:22]
  wire [31:0] n725_O_1_0_0; // @[Top.scala 965:22]
  wire [31:0] n725_O_1_0_1; // @[Top.scala 965:22]
  wire [31:0] n725_O_1_0_2; // @[Top.scala 965:22]
  wire [31:0] n725_O_1_1_0; // @[Top.scala 965:22]
  wire [31:0] n725_O_1_1_1; // @[Top.scala 965:22]
  wire [31:0] n725_O_1_1_2; // @[Top.scala 965:22]
  wire [31:0] n725_O_1_2_0; // @[Top.scala 965:22]
  wire [31:0] n725_O_1_2_1; // @[Top.scala 965:22]
  wire [31:0] n725_O_1_2_2; // @[Top.scala 965:22]
  wire [31:0] n725_O_2_0_0; // @[Top.scala 965:22]
  wire [31:0] n725_O_2_0_1; // @[Top.scala 965:22]
  wire [31:0] n725_O_2_0_2; // @[Top.scala 965:22]
  wire [31:0] n725_O_2_1_0; // @[Top.scala 965:22]
  wire [31:0] n725_O_2_1_1; // @[Top.scala 965:22]
  wire [31:0] n725_O_2_1_2; // @[Top.scala 965:22]
  wire [31:0] n725_O_2_2_0; // @[Top.scala 965:22]
  wire [31:0] n725_O_2_2_1; // @[Top.scala 965:22]
  wire [31:0] n725_O_2_2_2; // @[Top.scala 965:22]
  wire [31:0] n725_O_3_0_0; // @[Top.scala 965:22]
  wire [31:0] n725_O_3_0_1; // @[Top.scala 965:22]
  wire [31:0] n725_O_3_0_2; // @[Top.scala 965:22]
  wire [31:0] n725_O_3_1_0; // @[Top.scala 965:22]
  wire [31:0] n725_O_3_1_1; // @[Top.scala 965:22]
  wire [31:0] n725_O_3_1_2; // @[Top.scala 965:22]
  wire [31:0] n725_O_3_2_0; // @[Top.scala 965:22]
  wire [31:0] n725_O_3_2_1; // @[Top.scala 965:22]
  wire [31:0] n725_O_3_2_2; // @[Top.scala 965:22]
  wire [31:0] n725_O_4_0_0; // @[Top.scala 965:22]
  wire [31:0] n725_O_4_0_1; // @[Top.scala 965:22]
  wire [31:0] n725_O_4_0_2; // @[Top.scala 965:22]
  wire [31:0] n725_O_4_1_0; // @[Top.scala 965:22]
  wire [31:0] n725_O_4_1_1; // @[Top.scala 965:22]
  wire [31:0] n725_O_4_1_2; // @[Top.scala 965:22]
  wire [31:0] n725_O_4_2_0; // @[Top.scala 965:22]
  wire [31:0] n725_O_4_2_1; // @[Top.scala 965:22]
  wire [31:0] n725_O_4_2_2; // @[Top.scala 965:22]
  wire [31:0] n725_O_5_0_0; // @[Top.scala 965:22]
  wire [31:0] n725_O_5_0_1; // @[Top.scala 965:22]
  wire [31:0] n725_O_5_0_2; // @[Top.scala 965:22]
  wire [31:0] n725_O_5_1_0; // @[Top.scala 965:22]
  wire [31:0] n725_O_5_1_1; // @[Top.scala 965:22]
  wire [31:0] n725_O_5_1_2; // @[Top.scala 965:22]
  wire [31:0] n725_O_5_2_0; // @[Top.scala 965:22]
  wire [31:0] n725_O_5_2_1; // @[Top.scala 965:22]
  wire [31:0] n725_O_5_2_2; // @[Top.scala 965:22]
  wire [31:0] n725_O_6_0_0; // @[Top.scala 965:22]
  wire [31:0] n725_O_6_0_1; // @[Top.scala 965:22]
  wire [31:0] n725_O_6_0_2; // @[Top.scala 965:22]
  wire [31:0] n725_O_6_1_0; // @[Top.scala 965:22]
  wire [31:0] n725_O_6_1_1; // @[Top.scala 965:22]
  wire [31:0] n725_O_6_1_2; // @[Top.scala 965:22]
  wire [31:0] n725_O_6_2_0; // @[Top.scala 965:22]
  wire [31:0] n725_O_6_2_1; // @[Top.scala 965:22]
  wire [31:0] n725_O_6_2_2; // @[Top.scala 965:22]
  wire [31:0] n725_O_7_0_0; // @[Top.scala 965:22]
  wire [31:0] n725_O_7_0_1; // @[Top.scala 965:22]
  wire [31:0] n725_O_7_0_2; // @[Top.scala 965:22]
  wire [31:0] n725_O_7_1_0; // @[Top.scala 965:22]
  wire [31:0] n725_O_7_1_1; // @[Top.scala 965:22]
  wire [31:0] n725_O_7_1_2; // @[Top.scala 965:22]
  wire [31:0] n725_O_7_2_0; // @[Top.scala 965:22]
  wire [31:0] n725_O_7_2_1; // @[Top.scala 965:22]
  wire [31:0] n725_O_7_2_2; // @[Top.scala 965:22]
  wire  n734_valid_up; // @[Top.scala 969:22]
  wire  n734_valid_down; // @[Top.scala 969:22]
  wire [31:0] n734_I_0_0_0; // @[Top.scala 969:22]
  wire [31:0] n734_I_0_0_1; // @[Top.scala 969:22]
  wire [31:0] n734_I_0_0_2; // @[Top.scala 969:22]
  wire [31:0] n734_I_0_1_0; // @[Top.scala 969:22]
  wire [31:0] n734_I_0_1_1; // @[Top.scala 969:22]
  wire [31:0] n734_I_0_1_2; // @[Top.scala 969:22]
  wire [31:0] n734_I_0_2_0; // @[Top.scala 969:22]
  wire [31:0] n734_I_0_2_1; // @[Top.scala 969:22]
  wire [31:0] n734_I_0_2_2; // @[Top.scala 969:22]
  wire [31:0] n734_I_1_0_0; // @[Top.scala 969:22]
  wire [31:0] n734_I_1_0_1; // @[Top.scala 969:22]
  wire [31:0] n734_I_1_0_2; // @[Top.scala 969:22]
  wire [31:0] n734_I_1_1_0; // @[Top.scala 969:22]
  wire [31:0] n734_I_1_1_1; // @[Top.scala 969:22]
  wire [31:0] n734_I_1_1_2; // @[Top.scala 969:22]
  wire [31:0] n734_I_1_2_0; // @[Top.scala 969:22]
  wire [31:0] n734_I_1_2_1; // @[Top.scala 969:22]
  wire [31:0] n734_I_1_2_2; // @[Top.scala 969:22]
  wire [31:0] n734_I_2_0_0; // @[Top.scala 969:22]
  wire [31:0] n734_I_2_0_1; // @[Top.scala 969:22]
  wire [31:0] n734_I_2_0_2; // @[Top.scala 969:22]
  wire [31:0] n734_I_2_1_0; // @[Top.scala 969:22]
  wire [31:0] n734_I_2_1_1; // @[Top.scala 969:22]
  wire [31:0] n734_I_2_1_2; // @[Top.scala 969:22]
  wire [31:0] n734_I_2_2_0; // @[Top.scala 969:22]
  wire [31:0] n734_I_2_2_1; // @[Top.scala 969:22]
  wire [31:0] n734_I_2_2_2; // @[Top.scala 969:22]
  wire [31:0] n734_I_3_0_0; // @[Top.scala 969:22]
  wire [31:0] n734_I_3_0_1; // @[Top.scala 969:22]
  wire [31:0] n734_I_3_0_2; // @[Top.scala 969:22]
  wire [31:0] n734_I_3_1_0; // @[Top.scala 969:22]
  wire [31:0] n734_I_3_1_1; // @[Top.scala 969:22]
  wire [31:0] n734_I_3_1_2; // @[Top.scala 969:22]
  wire [31:0] n734_I_3_2_0; // @[Top.scala 969:22]
  wire [31:0] n734_I_3_2_1; // @[Top.scala 969:22]
  wire [31:0] n734_I_3_2_2; // @[Top.scala 969:22]
  wire [31:0] n734_I_4_0_0; // @[Top.scala 969:22]
  wire [31:0] n734_I_4_0_1; // @[Top.scala 969:22]
  wire [31:0] n734_I_4_0_2; // @[Top.scala 969:22]
  wire [31:0] n734_I_4_1_0; // @[Top.scala 969:22]
  wire [31:0] n734_I_4_1_1; // @[Top.scala 969:22]
  wire [31:0] n734_I_4_1_2; // @[Top.scala 969:22]
  wire [31:0] n734_I_4_2_0; // @[Top.scala 969:22]
  wire [31:0] n734_I_4_2_1; // @[Top.scala 969:22]
  wire [31:0] n734_I_4_2_2; // @[Top.scala 969:22]
  wire [31:0] n734_I_5_0_0; // @[Top.scala 969:22]
  wire [31:0] n734_I_5_0_1; // @[Top.scala 969:22]
  wire [31:0] n734_I_5_0_2; // @[Top.scala 969:22]
  wire [31:0] n734_I_5_1_0; // @[Top.scala 969:22]
  wire [31:0] n734_I_5_1_1; // @[Top.scala 969:22]
  wire [31:0] n734_I_5_1_2; // @[Top.scala 969:22]
  wire [31:0] n734_I_5_2_0; // @[Top.scala 969:22]
  wire [31:0] n734_I_5_2_1; // @[Top.scala 969:22]
  wire [31:0] n734_I_5_2_2; // @[Top.scala 969:22]
  wire [31:0] n734_I_6_0_0; // @[Top.scala 969:22]
  wire [31:0] n734_I_6_0_1; // @[Top.scala 969:22]
  wire [31:0] n734_I_6_0_2; // @[Top.scala 969:22]
  wire [31:0] n734_I_6_1_0; // @[Top.scala 969:22]
  wire [31:0] n734_I_6_1_1; // @[Top.scala 969:22]
  wire [31:0] n734_I_6_1_2; // @[Top.scala 969:22]
  wire [31:0] n734_I_6_2_0; // @[Top.scala 969:22]
  wire [31:0] n734_I_6_2_1; // @[Top.scala 969:22]
  wire [31:0] n734_I_6_2_2; // @[Top.scala 969:22]
  wire [31:0] n734_I_7_0_0; // @[Top.scala 969:22]
  wire [31:0] n734_I_7_0_1; // @[Top.scala 969:22]
  wire [31:0] n734_I_7_0_2; // @[Top.scala 969:22]
  wire [31:0] n734_I_7_1_0; // @[Top.scala 969:22]
  wire [31:0] n734_I_7_1_1; // @[Top.scala 969:22]
  wire [31:0] n734_I_7_1_2; // @[Top.scala 969:22]
  wire [31:0] n734_I_7_2_0; // @[Top.scala 969:22]
  wire [31:0] n734_I_7_2_1; // @[Top.scala 969:22]
  wire [31:0] n734_I_7_2_2; // @[Top.scala 969:22]
  wire [31:0] n734_O_0_0_0_0; // @[Top.scala 969:22]
  wire [31:0] n734_O_0_0_0_1; // @[Top.scala 969:22]
  wire [31:0] n734_O_0_0_0_2; // @[Top.scala 969:22]
  wire [31:0] n734_O_0_0_1_0; // @[Top.scala 969:22]
  wire [31:0] n734_O_0_0_1_1; // @[Top.scala 969:22]
  wire [31:0] n734_O_0_0_1_2; // @[Top.scala 969:22]
  wire [31:0] n734_O_0_0_2_0; // @[Top.scala 969:22]
  wire [31:0] n734_O_0_0_2_1; // @[Top.scala 969:22]
  wire [31:0] n734_O_0_0_2_2; // @[Top.scala 969:22]
  wire [31:0] n734_O_1_0_0_0; // @[Top.scala 969:22]
  wire [31:0] n734_O_1_0_0_1; // @[Top.scala 969:22]
  wire [31:0] n734_O_1_0_0_2; // @[Top.scala 969:22]
  wire [31:0] n734_O_1_0_1_0; // @[Top.scala 969:22]
  wire [31:0] n734_O_1_0_1_1; // @[Top.scala 969:22]
  wire [31:0] n734_O_1_0_1_2; // @[Top.scala 969:22]
  wire [31:0] n734_O_1_0_2_0; // @[Top.scala 969:22]
  wire [31:0] n734_O_1_0_2_1; // @[Top.scala 969:22]
  wire [31:0] n734_O_1_0_2_2; // @[Top.scala 969:22]
  wire [31:0] n734_O_2_0_0_0; // @[Top.scala 969:22]
  wire [31:0] n734_O_2_0_0_1; // @[Top.scala 969:22]
  wire [31:0] n734_O_2_0_0_2; // @[Top.scala 969:22]
  wire [31:0] n734_O_2_0_1_0; // @[Top.scala 969:22]
  wire [31:0] n734_O_2_0_1_1; // @[Top.scala 969:22]
  wire [31:0] n734_O_2_0_1_2; // @[Top.scala 969:22]
  wire [31:0] n734_O_2_0_2_0; // @[Top.scala 969:22]
  wire [31:0] n734_O_2_0_2_1; // @[Top.scala 969:22]
  wire [31:0] n734_O_2_0_2_2; // @[Top.scala 969:22]
  wire [31:0] n734_O_3_0_0_0; // @[Top.scala 969:22]
  wire [31:0] n734_O_3_0_0_1; // @[Top.scala 969:22]
  wire [31:0] n734_O_3_0_0_2; // @[Top.scala 969:22]
  wire [31:0] n734_O_3_0_1_0; // @[Top.scala 969:22]
  wire [31:0] n734_O_3_0_1_1; // @[Top.scala 969:22]
  wire [31:0] n734_O_3_0_1_2; // @[Top.scala 969:22]
  wire [31:0] n734_O_3_0_2_0; // @[Top.scala 969:22]
  wire [31:0] n734_O_3_0_2_1; // @[Top.scala 969:22]
  wire [31:0] n734_O_3_0_2_2; // @[Top.scala 969:22]
  wire [31:0] n734_O_4_0_0_0; // @[Top.scala 969:22]
  wire [31:0] n734_O_4_0_0_1; // @[Top.scala 969:22]
  wire [31:0] n734_O_4_0_0_2; // @[Top.scala 969:22]
  wire [31:0] n734_O_4_0_1_0; // @[Top.scala 969:22]
  wire [31:0] n734_O_4_0_1_1; // @[Top.scala 969:22]
  wire [31:0] n734_O_4_0_1_2; // @[Top.scala 969:22]
  wire [31:0] n734_O_4_0_2_0; // @[Top.scala 969:22]
  wire [31:0] n734_O_4_0_2_1; // @[Top.scala 969:22]
  wire [31:0] n734_O_4_0_2_2; // @[Top.scala 969:22]
  wire [31:0] n734_O_5_0_0_0; // @[Top.scala 969:22]
  wire [31:0] n734_O_5_0_0_1; // @[Top.scala 969:22]
  wire [31:0] n734_O_5_0_0_2; // @[Top.scala 969:22]
  wire [31:0] n734_O_5_0_1_0; // @[Top.scala 969:22]
  wire [31:0] n734_O_5_0_1_1; // @[Top.scala 969:22]
  wire [31:0] n734_O_5_0_1_2; // @[Top.scala 969:22]
  wire [31:0] n734_O_5_0_2_0; // @[Top.scala 969:22]
  wire [31:0] n734_O_5_0_2_1; // @[Top.scala 969:22]
  wire [31:0] n734_O_5_0_2_2; // @[Top.scala 969:22]
  wire [31:0] n734_O_6_0_0_0; // @[Top.scala 969:22]
  wire [31:0] n734_O_6_0_0_1; // @[Top.scala 969:22]
  wire [31:0] n734_O_6_0_0_2; // @[Top.scala 969:22]
  wire [31:0] n734_O_6_0_1_0; // @[Top.scala 969:22]
  wire [31:0] n734_O_6_0_1_1; // @[Top.scala 969:22]
  wire [31:0] n734_O_6_0_1_2; // @[Top.scala 969:22]
  wire [31:0] n734_O_6_0_2_0; // @[Top.scala 969:22]
  wire [31:0] n734_O_6_0_2_1; // @[Top.scala 969:22]
  wire [31:0] n734_O_6_0_2_2; // @[Top.scala 969:22]
  wire [31:0] n734_O_7_0_0_0; // @[Top.scala 969:22]
  wire [31:0] n734_O_7_0_0_1; // @[Top.scala 969:22]
  wire [31:0] n734_O_7_0_0_2; // @[Top.scala 969:22]
  wire [31:0] n734_O_7_0_1_0; // @[Top.scala 969:22]
  wire [31:0] n734_O_7_0_1_1; // @[Top.scala 969:22]
  wire [31:0] n734_O_7_0_1_2; // @[Top.scala 969:22]
  wire [31:0] n734_O_7_0_2_0; // @[Top.scala 969:22]
  wire [31:0] n734_O_7_0_2_1; // @[Top.scala 969:22]
  wire [31:0] n734_O_7_0_2_2; // @[Top.scala 969:22]
  wire  n741_valid_up; // @[Top.scala 972:22]
  wire  n741_valid_down; // @[Top.scala 972:22]
  wire [31:0] n741_I_0_0_0_0; // @[Top.scala 972:22]
  wire [31:0] n741_I_0_0_0_1; // @[Top.scala 972:22]
  wire [31:0] n741_I_0_0_0_2; // @[Top.scala 972:22]
  wire [31:0] n741_I_0_0_1_0; // @[Top.scala 972:22]
  wire [31:0] n741_I_0_0_1_1; // @[Top.scala 972:22]
  wire [31:0] n741_I_0_0_1_2; // @[Top.scala 972:22]
  wire [31:0] n741_I_0_0_2_0; // @[Top.scala 972:22]
  wire [31:0] n741_I_0_0_2_1; // @[Top.scala 972:22]
  wire [31:0] n741_I_0_0_2_2; // @[Top.scala 972:22]
  wire [31:0] n741_I_1_0_0_0; // @[Top.scala 972:22]
  wire [31:0] n741_I_1_0_0_1; // @[Top.scala 972:22]
  wire [31:0] n741_I_1_0_0_2; // @[Top.scala 972:22]
  wire [31:0] n741_I_1_0_1_0; // @[Top.scala 972:22]
  wire [31:0] n741_I_1_0_1_1; // @[Top.scala 972:22]
  wire [31:0] n741_I_1_0_1_2; // @[Top.scala 972:22]
  wire [31:0] n741_I_1_0_2_0; // @[Top.scala 972:22]
  wire [31:0] n741_I_1_0_2_1; // @[Top.scala 972:22]
  wire [31:0] n741_I_1_0_2_2; // @[Top.scala 972:22]
  wire [31:0] n741_I_2_0_0_0; // @[Top.scala 972:22]
  wire [31:0] n741_I_2_0_0_1; // @[Top.scala 972:22]
  wire [31:0] n741_I_2_0_0_2; // @[Top.scala 972:22]
  wire [31:0] n741_I_2_0_1_0; // @[Top.scala 972:22]
  wire [31:0] n741_I_2_0_1_1; // @[Top.scala 972:22]
  wire [31:0] n741_I_2_0_1_2; // @[Top.scala 972:22]
  wire [31:0] n741_I_2_0_2_0; // @[Top.scala 972:22]
  wire [31:0] n741_I_2_0_2_1; // @[Top.scala 972:22]
  wire [31:0] n741_I_2_0_2_2; // @[Top.scala 972:22]
  wire [31:0] n741_I_3_0_0_0; // @[Top.scala 972:22]
  wire [31:0] n741_I_3_0_0_1; // @[Top.scala 972:22]
  wire [31:0] n741_I_3_0_0_2; // @[Top.scala 972:22]
  wire [31:0] n741_I_3_0_1_0; // @[Top.scala 972:22]
  wire [31:0] n741_I_3_0_1_1; // @[Top.scala 972:22]
  wire [31:0] n741_I_3_0_1_2; // @[Top.scala 972:22]
  wire [31:0] n741_I_3_0_2_0; // @[Top.scala 972:22]
  wire [31:0] n741_I_3_0_2_1; // @[Top.scala 972:22]
  wire [31:0] n741_I_3_0_2_2; // @[Top.scala 972:22]
  wire [31:0] n741_I_4_0_0_0; // @[Top.scala 972:22]
  wire [31:0] n741_I_4_0_0_1; // @[Top.scala 972:22]
  wire [31:0] n741_I_4_0_0_2; // @[Top.scala 972:22]
  wire [31:0] n741_I_4_0_1_0; // @[Top.scala 972:22]
  wire [31:0] n741_I_4_0_1_1; // @[Top.scala 972:22]
  wire [31:0] n741_I_4_0_1_2; // @[Top.scala 972:22]
  wire [31:0] n741_I_4_0_2_0; // @[Top.scala 972:22]
  wire [31:0] n741_I_4_0_2_1; // @[Top.scala 972:22]
  wire [31:0] n741_I_4_0_2_2; // @[Top.scala 972:22]
  wire [31:0] n741_I_5_0_0_0; // @[Top.scala 972:22]
  wire [31:0] n741_I_5_0_0_1; // @[Top.scala 972:22]
  wire [31:0] n741_I_5_0_0_2; // @[Top.scala 972:22]
  wire [31:0] n741_I_5_0_1_0; // @[Top.scala 972:22]
  wire [31:0] n741_I_5_0_1_1; // @[Top.scala 972:22]
  wire [31:0] n741_I_5_0_1_2; // @[Top.scala 972:22]
  wire [31:0] n741_I_5_0_2_0; // @[Top.scala 972:22]
  wire [31:0] n741_I_5_0_2_1; // @[Top.scala 972:22]
  wire [31:0] n741_I_5_0_2_2; // @[Top.scala 972:22]
  wire [31:0] n741_I_6_0_0_0; // @[Top.scala 972:22]
  wire [31:0] n741_I_6_0_0_1; // @[Top.scala 972:22]
  wire [31:0] n741_I_6_0_0_2; // @[Top.scala 972:22]
  wire [31:0] n741_I_6_0_1_0; // @[Top.scala 972:22]
  wire [31:0] n741_I_6_0_1_1; // @[Top.scala 972:22]
  wire [31:0] n741_I_6_0_1_2; // @[Top.scala 972:22]
  wire [31:0] n741_I_6_0_2_0; // @[Top.scala 972:22]
  wire [31:0] n741_I_6_0_2_1; // @[Top.scala 972:22]
  wire [31:0] n741_I_6_0_2_2; // @[Top.scala 972:22]
  wire [31:0] n741_I_7_0_0_0; // @[Top.scala 972:22]
  wire [31:0] n741_I_7_0_0_1; // @[Top.scala 972:22]
  wire [31:0] n741_I_7_0_0_2; // @[Top.scala 972:22]
  wire [31:0] n741_I_7_0_1_0; // @[Top.scala 972:22]
  wire [31:0] n741_I_7_0_1_1; // @[Top.scala 972:22]
  wire [31:0] n741_I_7_0_1_2; // @[Top.scala 972:22]
  wire [31:0] n741_I_7_0_2_0; // @[Top.scala 972:22]
  wire [31:0] n741_I_7_0_2_1; // @[Top.scala 972:22]
  wire [31:0] n741_I_7_0_2_2; // @[Top.scala 972:22]
  wire [31:0] n741_O_0_0_0; // @[Top.scala 972:22]
  wire [31:0] n741_O_0_0_1; // @[Top.scala 972:22]
  wire [31:0] n741_O_0_0_2; // @[Top.scala 972:22]
  wire [31:0] n741_O_0_1_0; // @[Top.scala 972:22]
  wire [31:0] n741_O_0_1_1; // @[Top.scala 972:22]
  wire [31:0] n741_O_0_1_2; // @[Top.scala 972:22]
  wire [31:0] n741_O_0_2_0; // @[Top.scala 972:22]
  wire [31:0] n741_O_0_2_1; // @[Top.scala 972:22]
  wire [31:0] n741_O_0_2_2; // @[Top.scala 972:22]
  wire [31:0] n741_O_1_0_0; // @[Top.scala 972:22]
  wire [31:0] n741_O_1_0_1; // @[Top.scala 972:22]
  wire [31:0] n741_O_1_0_2; // @[Top.scala 972:22]
  wire [31:0] n741_O_1_1_0; // @[Top.scala 972:22]
  wire [31:0] n741_O_1_1_1; // @[Top.scala 972:22]
  wire [31:0] n741_O_1_1_2; // @[Top.scala 972:22]
  wire [31:0] n741_O_1_2_0; // @[Top.scala 972:22]
  wire [31:0] n741_O_1_2_1; // @[Top.scala 972:22]
  wire [31:0] n741_O_1_2_2; // @[Top.scala 972:22]
  wire [31:0] n741_O_2_0_0; // @[Top.scala 972:22]
  wire [31:0] n741_O_2_0_1; // @[Top.scala 972:22]
  wire [31:0] n741_O_2_0_2; // @[Top.scala 972:22]
  wire [31:0] n741_O_2_1_0; // @[Top.scala 972:22]
  wire [31:0] n741_O_2_1_1; // @[Top.scala 972:22]
  wire [31:0] n741_O_2_1_2; // @[Top.scala 972:22]
  wire [31:0] n741_O_2_2_0; // @[Top.scala 972:22]
  wire [31:0] n741_O_2_2_1; // @[Top.scala 972:22]
  wire [31:0] n741_O_2_2_2; // @[Top.scala 972:22]
  wire [31:0] n741_O_3_0_0; // @[Top.scala 972:22]
  wire [31:0] n741_O_3_0_1; // @[Top.scala 972:22]
  wire [31:0] n741_O_3_0_2; // @[Top.scala 972:22]
  wire [31:0] n741_O_3_1_0; // @[Top.scala 972:22]
  wire [31:0] n741_O_3_1_1; // @[Top.scala 972:22]
  wire [31:0] n741_O_3_1_2; // @[Top.scala 972:22]
  wire [31:0] n741_O_3_2_0; // @[Top.scala 972:22]
  wire [31:0] n741_O_3_2_1; // @[Top.scala 972:22]
  wire [31:0] n741_O_3_2_2; // @[Top.scala 972:22]
  wire [31:0] n741_O_4_0_0; // @[Top.scala 972:22]
  wire [31:0] n741_O_4_0_1; // @[Top.scala 972:22]
  wire [31:0] n741_O_4_0_2; // @[Top.scala 972:22]
  wire [31:0] n741_O_4_1_0; // @[Top.scala 972:22]
  wire [31:0] n741_O_4_1_1; // @[Top.scala 972:22]
  wire [31:0] n741_O_4_1_2; // @[Top.scala 972:22]
  wire [31:0] n741_O_4_2_0; // @[Top.scala 972:22]
  wire [31:0] n741_O_4_2_1; // @[Top.scala 972:22]
  wire [31:0] n741_O_4_2_2; // @[Top.scala 972:22]
  wire [31:0] n741_O_5_0_0; // @[Top.scala 972:22]
  wire [31:0] n741_O_5_0_1; // @[Top.scala 972:22]
  wire [31:0] n741_O_5_0_2; // @[Top.scala 972:22]
  wire [31:0] n741_O_5_1_0; // @[Top.scala 972:22]
  wire [31:0] n741_O_5_1_1; // @[Top.scala 972:22]
  wire [31:0] n741_O_5_1_2; // @[Top.scala 972:22]
  wire [31:0] n741_O_5_2_0; // @[Top.scala 972:22]
  wire [31:0] n741_O_5_2_1; // @[Top.scala 972:22]
  wire [31:0] n741_O_5_2_2; // @[Top.scala 972:22]
  wire [31:0] n741_O_6_0_0; // @[Top.scala 972:22]
  wire [31:0] n741_O_6_0_1; // @[Top.scala 972:22]
  wire [31:0] n741_O_6_0_2; // @[Top.scala 972:22]
  wire [31:0] n741_O_6_1_0; // @[Top.scala 972:22]
  wire [31:0] n741_O_6_1_1; // @[Top.scala 972:22]
  wire [31:0] n741_O_6_1_2; // @[Top.scala 972:22]
  wire [31:0] n741_O_6_2_0; // @[Top.scala 972:22]
  wire [31:0] n741_O_6_2_1; // @[Top.scala 972:22]
  wire [31:0] n741_O_6_2_2; // @[Top.scala 972:22]
  wire [31:0] n741_O_7_0_0; // @[Top.scala 972:22]
  wire [31:0] n741_O_7_0_1; // @[Top.scala 972:22]
  wire [31:0] n741_O_7_0_2; // @[Top.scala 972:22]
  wire [31:0] n741_O_7_1_0; // @[Top.scala 972:22]
  wire [31:0] n741_O_7_1_1; // @[Top.scala 972:22]
  wire [31:0] n741_O_7_1_2; // @[Top.scala 972:22]
  wire [31:0] n741_O_7_2_0; // @[Top.scala 972:22]
  wire [31:0] n741_O_7_2_1; // @[Top.scala 972:22]
  wire [31:0] n741_O_7_2_2; // @[Top.scala 972:22]
  wire  n783_clock; // @[Top.scala 975:22]
  wire  n783_reset; // @[Top.scala 975:22]
  wire  n783_valid_up; // @[Top.scala 975:22]
  wire  n783_valid_down; // @[Top.scala 975:22]
  wire [31:0] n783_I_0_0_0; // @[Top.scala 975:22]
  wire [31:0] n783_I_0_0_1; // @[Top.scala 975:22]
  wire [31:0] n783_I_0_0_2; // @[Top.scala 975:22]
  wire [31:0] n783_I_0_1_0; // @[Top.scala 975:22]
  wire [31:0] n783_I_0_1_1; // @[Top.scala 975:22]
  wire [31:0] n783_I_0_1_2; // @[Top.scala 975:22]
  wire [31:0] n783_I_0_2_0; // @[Top.scala 975:22]
  wire [31:0] n783_I_0_2_1; // @[Top.scala 975:22]
  wire [31:0] n783_I_0_2_2; // @[Top.scala 975:22]
  wire [31:0] n783_I_1_0_0; // @[Top.scala 975:22]
  wire [31:0] n783_I_1_0_1; // @[Top.scala 975:22]
  wire [31:0] n783_I_1_0_2; // @[Top.scala 975:22]
  wire [31:0] n783_I_1_1_0; // @[Top.scala 975:22]
  wire [31:0] n783_I_1_1_1; // @[Top.scala 975:22]
  wire [31:0] n783_I_1_1_2; // @[Top.scala 975:22]
  wire [31:0] n783_I_1_2_0; // @[Top.scala 975:22]
  wire [31:0] n783_I_1_2_1; // @[Top.scala 975:22]
  wire [31:0] n783_I_1_2_2; // @[Top.scala 975:22]
  wire [31:0] n783_I_2_0_0; // @[Top.scala 975:22]
  wire [31:0] n783_I_2_0_1; // @[Top.scala 975:22]
  wire [31:0] n783_I_2_0_2; // @[Top.scala 975:22]
  wire [31:0] n783_I_2_1_0; // @[Top.scala 975:22]
  wire [31:0] n783_I_2_1_1; // @[Top.scala 975:22]
  wire [31:0] n783_I_2_1_2; // @[Top.scala 975:22]
  wire [31:0] n783_I_2_2_0; // @[Top.scala 975:22]
  wire [31:0] n783_I_2_2_1; // @[Top.scala 975:22]
  wire [31:0] n783_I_2_2_2; // @[Top.scala 975:22]
  wire [31:0] n783_I_3_0_0; // @[Top.scala 975:22]
  wire [31:0] n783_I_3_0_1; // @[Top.scala 975:22]
  wire [31:0] n783_I_3_0_2; // @[Top.scala 975:22]
  wire [31:0] n783_I_3_1_0; // @[Top.scala 975:22]
  wire [31:0] n783_I_3_1_1; // @[Top.scala 975:22]
  wire [31:0] n783_I_3_1_2; // @[Top.scala 975:22]
  wire [31:0] n783_I_3_2_0; // @[Top.scala 975:22]
  wire [31:0] n783_I_3_2_1; // @[Top.scala 975:22]
  wire [31:0] n783_I_3_2_2; // @[Top.scala 975:22]
  wire [31:0] n783_I_4_0_0; // @[Top.scala 975:22]
  wire [31:0] n783_I_4_0_1; // @[Top.scala 975:22]
  wire [31:0] n783_I_4_0_2; // @[Top.scala 975:22]
  wire [31:0] n783_I_4_1_0; // @[Top.scala 975:22]
  wire [31:0] n783_I_4_1_1; // @[Top.scala 975:22]
  wire [31:0] n783_I_4_1_2; // @[Top.scala 975:22]
  wire [31:0] n783_I_4_2_0; // @[Top.scala 975:22]
  wire [31:0] n783_I_4_2_1; // @[Top.scala 975:22]
  wire [31:0] n783_I_4_2_2; // @[Top.scala 975:22]
  wire [31:0] n783_I_5_0_0; // @[Top.scala 975:22]
  wire [31:0] n783_I_5_0_1; // @[Top.scala 975:22]
  wire [31:0] n783_I_5_0_2; // @[Top.scala 975:22]
  wire [31:0] n783_I_5_1_0; // @[Top.scala 975:22]
  wire [31:0] n783_I_5_1_1; // @[Top.scala 975:22]
  wire [31:0] n783_I_5_1_2; // @[Top.scala 975:22]
  wire [31:0] n783_I_5_2_0; // @[Top.scala 975:22]
  wire [31:0] n783_I_5_2_1; // @[Top.scala 975:22]
  wire [31:0] n783_I_5_2_2; // @[Top.scala 975:22]
  wire [31:0] n783_I_6_0_0; // @[Top.scala 975:22]
  wire [31:0] n783_I_6_0_1; // @[Top.scala 975:22]
  wire [31:0] n783_I_6_0_2; // @[Top.scala 975:22]
  wire [31:0] n783_I_6_1_0; // @[Top.scala 975:22]
  wire [31:0] n783_I_6_1_1; // @[Top.scala 975:22]
  wire [31:0] n783_I_6_1_2; // @[Top.scala 975:22]
  wire [31:0] n783_I_6_2_0; // @[Top.scala 975:22]
  wire [31:0] n783_I_6_2_1; // @[Top.scala 975:22]
  wire [31:0] n783_I_6_2_2; // @[Top.scala 975:22]
  wire [31:0] n783_I_7_0_0; // @[Top.scala 975:22]
  wire [31:0] n783_I_7_0_1; // @[Top.scala 975:22]
  wire [31:0] n783_I_7_0_2; // @[Top.scala 975:22]
  wire [31:0] n783_I_7_1_0; // @[Top.scala 975:22]
  wire [31:0] n783_I_7_1_1; // @[Top.scala 975:22]
  wire [31:0] n783_I_7_1_2; // @[Top.scala 975:22]
  wire [31:0] n783_I_7_2_0; // @[Top.scala 975:22]
  wire [31:0] n783_I_7_2_1; // @[Top.scala 975:22]
  wire [31:0] n783_I_7_2_2; // @[Top.scala 975:22]
  wire [31:0] n783_O_0_0_0; // @[Top.scala 975:22]
  wire [31:0] n783_O_1_0_0; // @[Top.scala 975:22]
  wire [31:0] n783_O_2_0_0; // @[Top.scala 975:22]
  wire [31:0] n783_O_3_0_0; // @[Top.scala 975:22]
  wire [31:0] n783_O_4_0_0; // @[Top.scala 975:22]
  wire [31:0] n783_O_5_0_0; // @[Top.scala 975:22]
  wire [31:0] n783_O_6_0_0; // @[Top.scala 975:22]
  wire [31:0] n783_O_7_0_0; // @[Top.scala 975:22]
  wire  n784_valid_up; // @[Top.scala 978:22]
  wire  n784_valid_down; // @[Top.scala 978:22]
  wire [31:0] n784_I_0_0_0; // @[Top.scala 978:22]
  wire [31:0] n784_I_1_0_0; // @[Top.scala 978:22]
  wire [31:0] n784_I_2_0_0; // @[Top.scala 978:22]
  wire [31:0] n784_I_3_0_0; // @[Top.scala 978:22]
  wire [31:0] n784_I_4_0_0; // @[Top.scala 978:22]
  wire [31:0] n784_I_5_0_0; // @[Top.scala 978:22]
  wire [31:0] n784_I_6_0_0; // @[Top.scala 978:22]
  wire [31:0] n784_I_7_0_0; // @[Top.scala 978:22]
  wire [31:0] n784_O_0_0; // @[Top.scala 978:22]
  wire [31:0] n784_O_1_0; // @[Top.scala 978:22]
  wire [31:0] n784_O_2_0; // @[Top.scala 978:22]
  wire [31:0] n784_O_3_0; // @[Top.scala 978:22]
  wire [31:0] n784_O_4_0; // @[Top.scala 978:22]
  wire [31:0] n784_O_5_0; // @[Top.scala 978:22]
  wire [31:0] n784_O_6_0; // @[Top.scala 978:22]
  wire [31:0] n784_O_7_0; // @[Top.scala 978:22]
  wire  n785_valid_up; // @[Top.scala 981:22]
  wire  n785_valid_down; // @[Top.scala 981:22]
  wire [31:0] n785_I_0_0; // @[Top.scala 981:22]
  wire [31:0] n785_I_1_0; // @[Top.scala 981:22]
  wire [31:0] n785_I_2_0; // @[Top.scala 981:22]
  wire [31:0] n785_I_3_0; // @[Top.scala 981:22]
  wire [31:0] n785_I_4_0; // @[Top.scala 981:22]
  wire [31:0] n785_I_5_0; // @[Top.scala 981:22]
  wire [31:0] n785_I_6_0; // @[Top.scala 981:22]
  wire [31:0] n785_I_7_0; // @[Top.scala 981:22]
  wire [31:0] n785_O_0; // @[Top.scala 981:22]
  wire [31:0] n785_O_1; // @[Top.scala 981:22]
  wire [31:0] n785_O_2; // @[Top.scala 981:22]
  wire [31:0] n785_O_3; // @[Top.scala 981:22]
  wire [31:0] n785_O_4; // @[Top.scala 981:22]
  wire [31:0] n785_O_5; // @[Top.scala 981:22]
  wire [31:0] n785_O_6; // @[Top.scala 981:22]
  wire [31:0] n785_O_7; // @[Top.scala 981:22]
  wire  n786_clock; // @[Top.scala 984:22]
  wire  n786_reset; // @[Top.scala 984:22]
  wire  n786_valid_up; // @[Top.scala 984:22]
  wire  n786_valid_down; // @[Top.scala 984:22]
  wire [31:0] n786_I_0; // @[Top.scala 984:22]
  wire [31:0] n786_I_1; // @[Top.scala 984:22]
  wire [31:0] n786_I_2; // @[Top.scala 984:22]
  wire [31:0] n786_I_3; // @[Top.scala 984:22]
  wire [31:0] n786_I_4; // @[Top.scala 984:22]
  wire [31:0] n786_I_5; // @[Top.scala 984:22]
  wire [31:0] n786_I_6; // @[Top.scala 984:22]
  wire [31:0] n786_I_7; // @[Top.scala 984:22]
  wire [31:0] n786_O_0; // @[Top.scala 984:22]
  wire [31:0] n786_O_1; // @[Top.scala 984:22]
  wire [31:0] n786_O_2; // @[Top.scala 984:22]
  wire [31:0] n786_O_3; // @[Top.scala 984:22]
  wire [31:0] n786_O_4; // @[Top.scala 984:22]
  wire [31:0] n786_O_5; // @[Top.scala 984:22]
  wire [31:0] n786_O_6; // @[Top.scala 984:22]
  wire [31:0] n786_O_7; // @[Top.scala 984:22]
  wire  n787_clock; // @[Top.scala 987:22]
  wire  n787_reset; // @[Top.scala 987:22]
  wire  n787_valid_up; // @[Top.scala 987:22]
  wire  n787_valid_down; // @[Top.scala 987:22]
  wire [31:0] n787_I0_0; // @[Top.scala 987:22]
  wire [31:0] n787_I0_1; // @[Top.scala 987:22]
  wire [31:0] n787_I0_2; // @[Top.scala 987:22]
  wire [31:0] n787_I0_3; // @[Top.scala 987:22]
  wire [31:0] n787_I0_4; // @[Top.scala 987:22]
  wire [31:0] n787_I0_5; // @[Top.scala 987:22]
  wire [31:0] n787_I0_6; // @[Top.scala 987:22]
  wire [31:0] n787_I0_7; // @[Top.scala 987:22]
  wire [31:0] n787_I1_0; // @[Top.scala 987:22]
  wire [31:0] n787_I1_1; // @[Top.scala 987:22]
  wire [31:0] n787_I1_2; // @[Top.scala 987:22]
  wire [31:0] n787_I1_3; // @[Top.scala 987:22]
  wire [31:0] n787_I1_4; // @[Top.scala 987:22]
  wire [31:0] n787_I1_5; // @[Top.scala 987:22]
  wire [31:0] n787_I1_6; // @[Top.scala 987:22]
  wire [31:0] n787_I1_7; // @[Top.scala 987:22]
  wire [31:0] n787_O_0; // @[Top.scala 987:22]
  wire [31:0] n787_O_1; // @[Top.scala 987:22]
  wire [31:0] n787_O_2; // @[Top.scala 987:22]
  wire [31:0] n787_O_3; // @[Top.scala 987:22]
  wire [31:0] n787_O_4; // @[Top.scala 987:22]
  wire [31:0] n787_O_5; // @[Top.scala 987:22]
  wire [31:0] n787_O_6; // @[Top.scala 987:22]
  wire [31:0] n787_O_7; // @[Top.scala 987:22]
  wire  n823_valid_up; // @[Top.scala 991:22]
  wire  n823_valid_down; // @[Top.scala 991:22]
  wire [31:0] n823_I_0_t1b_t0b; // @[Top.scala 991:22]
  wire [31:0] n823_I_0_t1b_t1b; // @[Top.scala 991:22]
  wire [31:0] n823_I_1_t1b_t0b; // @[Top.scala 991:22]
  wire [31:0] n823_I_1_t1b_t1b; // @[Top.scala 991:22]
  wire [31:0] n823_I_2_t1b_t0b; // @[Top.scala 991:22]
  wire [31:0] n823_I_2_t1b_t1b; // @[Top.scala 991:22]
  wire [31:0] n823_I_3_t1b_t0b; // @[Top.scala 991:22]
  wire [31:0] n823_I_3_t1b_t1b; // @[Top.scala 991:22]
  wire [31:0] n823_I_4_t1b_t0b; // @[Top.scala 991:22]
  wire [31:0] n823_I_4_t1b_t1b; // @[Top.scala 991:22]
  wire [31:0] n823_I_5_t1b_t0b; // @[Top.scala 991:22]
  wire [31:0] n823_I_5_t1b_t1b; // @[Top.scala 991:22]
  wire [31:0] n823_I_6_t1b_t0b; // @[Top.scala 991:22]
  wire [31:0] n823_I_6_t1b_t1b; // @[Top.scala 991:22]
  wire [31:0] n823_I_7_t1b_t0b; // @[Top.scala 991:22]
  wire [31:0] n823_I_7_t1b_t1b; // @[Top.scala 991:22]
  wire [31:0] n823_O_0; // @[Top.scala 991:22]
  wire [31:0] n823_O_1; // @[Top.scala 991:22]
  wire [31:0] n823_O_2; // @[Top.scala 991:22]
  wire [31:0] n823_O_3; // @[Top.scala 991:22]
  wire [31:0] n823_O_4; // @[Top.scala 991:22]
  wire [31:0] n823_O_5; // @[Top.scala 991:22]
  wire [31:0] n823_O_6; // @[Top.scala 991:22]
  wire [31:0] n823_O_7; // @[Top.scala 991:22]
  wire  n824_clock; // @[Top.scala 994:22]
  wire  n824_reset; // @[Top.scala 994:22]
  wire  n824_valid_up; // @[Top.scala 994:22]
  wire  n824_valid_down; // @[Top.scala 994:22]
  wire [31:0] n824_I_0; // @[Top.scala 994:22]
  wire [31:0] n824_I_1; // @[Top.scala 994:22]
  wire [31:0] n824_I_2; // @[Top.scala 994:22]
  wire [31:0] n824_I_3; // @[Top.scala 994:22]
  wire [31:0] n824_I_4; // @[Top.scala 994:22]
  wire [31:0] n824_I_5; // @[Top.scala 994:22]
  wire [31:0] n824_I_6; // @[Top.scala 994:22]
  wire [31:0] n824_I_7; // @[Top.scala 994:22]
  wire [31:0] n824_O_0; // @[Top.scala 994:22]
  wire [31:0] n824_O_1; // @[Top.scala 994:22]
  wire [31:0] n824_O_2; // @[Top.scala 994:22]
  wire [31:0] n824_O_3; // @[Top.scala 994:22]
  wire [31:0] n824_O_4; // @[Top.scala 994:22]
  wire [31:0] n824_O_5; // @[Top.scala 994:22]
  wire [31:0] n824_O_6; // @[Top.scala 994:22]
  wire [31:0] n824_O_7; // @[Top.scala 994:22]
  wire  n825_clock; // @[Top.scala 997:22]
  wire  n825_reset; // @[Top.scala 997:22]
  wire  n825_valid_up; // @[Top.scala 997:22]
  wire  n825_valid_down; // @[Top.scala 997:22]
  wire [31:0] n825_I_0; // @[Top.scala 997:22]
  wire [31:0] n825_I_1; // @[Top.scala 997:22]
  wire [31:0] n825_I_2; // @[Top.scala 997:22]
  wire [31:0] n825_I_3; // @[Top.scala 997:22]
  wire [31:0] n825_I_4; // @[Top.scala 997:22]
  wire [31:0] n825_I_5; // @[Top.scala 997:22]
  wire [31:0] n825_I_6; // @[Top.scala 997:22]
  wire [31:0] n825_I_7; // @[Top.scala 997:22]
  wire [31:0] n825_O_0; // @[Top.scala 997:22]
  wire [31:0] n825_O_1; // @[Top.scala 997:22]
  wire [31:0] n825_O_2; // @[Top.scala 997:22]
  wire [31:0] n825_O_3; // @[Top.scala 997:22]
  wire [31:0] n825_O_4; // @[Top.scala 997:22]
  wire [31:0] n825_O_5; // @[Top.scala 997:22]
  wire [31:0] n825_O_6; // @[Top.scala 997:22]
  wire [31:0] n825_O_7; // @[Top.scala 997:22]
  wire  n826_clock; // @[Top.scala 1000:22]
  wire  n826_valid_up; // @[Top.scala 1000:22]
  wire  n826_valid_down; // @[Top.scala 1000:22]
  wire [31:0] n826_I_0; // @[Top.scala 1000:22]
  wire [31:0] n826_I_1; // @[Top.scala 1000:22]
  wire [31:0] n826_I_2; // @[Top.scala 1000:22]
  wire [31:0] n826_I_3; // @[Top.scala 1000:22]
  wire [31:0] n826_I_4; // @[Top.scala 1000:22]
  wire [31:0] n826_I_5; // @[Top.scala 1000:22]
  wire [31:0] n826_I_6; // @[Top.scala 1000:22]
  wire [31:0] n826_I_7; // @[Top.scala 1000:22]
  wire [31:0] n826_O_0; // @[Top.scala 1000:22]
  wire [31:0] n826_O_1; // @[Top.scala 1000:22]
  wire [31:0] n826_O_2; // @[Top.scala 1000:22]
  wire [31:0] n826_O_3; // @[Top.scala 1000:22]
  wire [31:0] n826_O_4; // @[Top.scala 1000:22]
  wire [31:0] n826_O_5; // @[Top.scala 1000:22]
  wire [31:0] n826_O_6; // @[Top.scala 1000:22]
  wire [31:0] n826_O_7; // @[Top.scala 1000:22]
  wire  n827_clock; // @[Top.scala 1003:22]
  wire  n827_valid_up; // @[Top.scala 1003:22]
  wire  n827_valid_down; // @[Top.scala 1003:22]
  wire [31:0] n827_I_0; // @[Top.scala 1003:22]
  wire [31:0] n827_I_1; // @[Top.scala 1003:22]
  wire [31:0] n827_I_2; // @[Top.scala 1003:22]
  wire [31:0] n827_I_3; // @[Top.scala 1003:22]
  wire [31:0] n827_I_4; // @[Top.scala 1003:22]
  wire [31:0] n827_I_5; // @[Top.scala 1003:22]
  wire [31:0] n827_I_6; // @[Top.scala 1003:22]
  wire [31:0] n827_I_7; // @[Top.scala 1003:22]
  wire [31:0] n827_O_0; // @[Top.scala 1003:22]
  wire [31:0] n827_O_1; // @[Top.scala 1003:22]
  wire [31:0] n827_O_2; // @[Top.scala 1003:22]
  wire [31:0] n827_O_3; // @[Top.scala 1003:22]
  wire [31:0] n827_O_4; // @[Top.scala 1003:22]
  wire [31:0] n827_O_5; // @[Top.scala 1003:22]
  wire [31:0] n827_O_6; // @[Top.scala 1003:22]
  wire [31:0] n827_O_7; // @[Top.scala 1003:22]
  wire  n828_valid_up; // @[Top.scala 1006:22]
  wire  n828_valid_down; // @[Top.scala 1006:22]
  wire [31:0] n828_I0_0; // @[Top.scala 1006:22]
  wire [31:0] n828_I0_1; // @[Top.scala 1006:22]
  wire [31:0] n828_I0_2; // @[Top.scala 1006:22]
  wire [31:0] n828_I0_3; // @[Top.scala 1006:22]
  wire [31:0] n828_I0_4; // @[Top.scala 1006:22]
  wire [31:0] n828_I0_5; // @[Top.scala 1006:22]
  wire [31:0] n828_I0_6; // @[Top.scala 1006:22]
  wire [31:0] n828_I0_7; // @[Top.scala 1006:22]
  wire [31:0] n828_I1_0; // @[Top.scala 1006:22]
  wire [31:0] n828_I1_1; // @[Top.scala 1006:22]
  wire [31:0] n828_I1_2; // @[Top.scala 1006:22]
  wire [31:0] n828_I1_3; // @[Top.scala 1006:22]
  wire [31:0] n828_I1_4; // @[Top.scala 1006:22]
  wire [31:0] n828_I1_5; // @[Top.scala 1006:22]
  wire [31:0] n828_I1_6; // @[Top.scala 1006:22]
  wire [31:0] n828_I1_7; // @[Top.scala 1006:22]
  wire [31:0] n828_O_0_0; // @[Top.scala 1006:22]
  wire [31:0] n828_O_0_1; // @[Top.scala 1006:22]
  wire [31:0] n828_O_1_0; // @[Top.scala 1006:22]
  wire [31:0] n828_O_1_1; // @[Top.scala 1006:22]
  wire [31:0] n828_O_2_0; // @[Top.scala 1006:22]
  wire [31:0] n828_O_2_1; // @[Top.scala 1006:22]
  wire [31:0] n828_O_3_0; // @[Top.scala 1006:22]
  wire [31:0] n828_O_3_1; // @[Top.scala 1006:22]
  wire [31:0] n828_O_4_0; // @[Top.scala 1006:22]
  wire [31:0] n828_O_4_1; // @[Top.scala 1006:22]
  wire [31:0] n828_O_5_0; // @[Top.scala 1006:22]
  wire [31:0] n828_O_5_1; // @[Top.scala 1006:22]
  wire [31:0] n828_O_6_0; // @[Top.scala 1006:22]
  wire [31:0] n828_O_6_1; // @[Top.scala 1006:22]
  wire [31:0] n828_O_7_0; // @[Top.scala 1006:22]
  wire [31:0] n828_O_7_1; // @[Top.scala 1006:22]
  wire  n835_valid_up; // @[Top.scala 1010:22]
  wire  n835_valid_down; // @[Top.scala 1010:22]
  wire [31:0] n835_I0_0_0; // @[Top.scala 1010:22]
  wire [31:0] n835_I0_0_1; // @[Top.scala 1010:22]
  wire [31:0] n835_I0_1_0; // @[Top.scala 1010:22]
  wire [31:0] n835_I0_1_1; // @[Top.scala 1010:22]
  wire [31:0] n835_I0_2_0; // @[Top.scala 1010:22]
  wire [31:0] n835_I0_2_1; // @[Top.scala 1010:22]
  wire [31:0] n835_I0_3_0; // @[Top.scala 1010:22]
  wire [31:0] n835_I0_3_1; // @[Top.scala 1010:22]
  wire [31:0] n835_I0_4_0; // @[Top.scala 1010:22]
  wire [31:0] n835_I0_4_1; // @[Top.scala 1010:22]
  wire [31:0] n835_I0_5_0; // @[Top.scala 1010:22]
  wire [31:0] n835_I0_5_1; // @[Top.scala 1010:22]
  wire [31:0] n835_I0_6_0; // @[Top.scala 1010:22]
  wire [31:0] n835_I0_6_1; // @[Top.scala 1010:22]
  wire [31:0] n835_I0_7_0; // @[Top.scala 1010:22]
  wire [31:0] n835_I0_7_1; // @[Top.scala 1010:22]
  wire [31:0] n835_I1_0; // @[Top.scala 1010:22]
  wire [31:0] n835_I1_1; // @[Top.scala 1010:22]
  wire [31:0] n835_I1_2; // @[Top.scala 1010:22]
  wire [31:0] n835_I1_3; // @[Top.scala 1010:22]
  wire [31:0] n835_I1_4; // @[Top.scala 1010:22]
  wire [31:0] n835_I1_5; // @[Top.scala 1010:22]
  wire [31:0] n835_I1_6; // @[Top.scala 1010:22]
  wire [31:0] n835_I1_7; // @[Top.scala 1010:22]
  wire [31:0] n835_O_0_0; // @[Top.scala 1010:22]
  wire [31:0] n835_O_0_1; // @[Top.scala 1010:22]
  wire [31:0] n835_O_0_2; // @[Top.scala 1010:22]
  wire [31:0] n835_O_1_0; // @[Top.scala 1010:22]
  wire [31:0] n835_O_1_1; // @[Top.scala 1010:22]
  wire [31:0] n835_O_1_2; // @[Top.scala 1010:22]
  wire [31:0] n835_O_2_0; // @[Top.scala 1010:22]
  wire [31:0] n835_O_2_1; // @[Top.scala 1010:22]
  wire [31:0] n835_O_2_2; // @[Top.scala 1010:22]
  wire [31:0] n835_O_3_0; // @[Top.scala 1010:22]
  wire [31:0] n835_O_3_1; // @[Top.scala 1010:22]
  wire [31:0] n835_O_3_2; // @[Top.scala 1010:22]
  wire [31:0] n835_O_4_0; // @[Top.scala 1010:22]
  wire [31:0] n835_O_4_1; // @[Top.scala 1010:22]
  wire [31:0] n835_O_4_2; // @[Top.scala 1010:22]
  wire [31:0] n835_O_5_0; // @[Top.scala 1010:22]
  wire [31:0] n835_O_5_1; // @[Top.scala 1010:22]
  wire [31:0] n835_O_5_2; // @[Top.scala 1010:22]
  wire [31:0] n835_O_6_0; // @[Top.scala 1010:22]
  wire [31:0] n835_O_6_1; // @[Top.scala 1010:22]
  wire [31:0] n835_O_6_2; // @[Top.scala 1010:22]
  wire [31:0] n835_O_7_0; // @[Top.scala 1010:22]
  wire [31:0] n835_O_7_1; // @[Top.scala 1010:22]
  wire [31:0] n835_O_7_2; // @[Top.scala 1010:22]
  wire  n844_valid_up; // @[Top.scala 1014:22]
  wire  n844_valid_down; // @[Top.scala 1014:22]
  wire [31:0] n844_I_0_0; // @[Top.scala 1014:22]
  wire [31:0] n844_I_0_1; // @[Top.scala 1014:22]
  wire [31:0] n844_I_0_2; // @[Top.scala 1014:22]
  wire [31:0] n844_I_1_0; // @[Top.scala 1014:22]
  wire [31:0] n844_I_1_1; // @[Top.scala 1014:22]
  wire [31:0] n844_I_1_2; // @[Top.scala 1014:22]
  wire [31:0] n844_I_2_0; // @[Top.scala 1014:22]
  wire [31:0] n844_I_2_1; // @[Top.scala 1014:22]
  wire [31:0] n844_I_2_2; // @[Top.scala 1014:22]
  wire [31:0] n844_I_3_0; // @[Top.scala 1014:22]
  wire [31:0] n844_I_3_1; // @[Top.scala 1014:22]
  wire [31:0] n844_I_3_2; // @[Top.scala 1014:22]
  wire [31:0] n844_I_4_0; // @[Top.scala 1014:22]
  wire [31:0] n844_I_4_1; // @[Top.scala 1014:22]
  wire [31:0] n844_I_4_2; // @[Top.scala 1014:22]
  wire [31:0] n844_I_5_0; // @[Top.scala 1014:22]
  wire [31:0] n844_I_5_1; // @[Top.scala 1014:22]
  wire [31:0] n844_I_5_2; // @[Top.scala 1014:22]
  wire [31:0] n844_I_6_0; // @[Top.scala 1014:22]
  wire [31:0] n844_I_6_1; // @[Top.scala 1014:22]
  wire [31:0] n844_I_6_2; // @[Top.scala 1014:22]
  wire [31:0] n844_I_7_0; // @[Top.scala 1014:22]
  wire [31:0] n844_I_7_1; // @[Top.scala 1014:22]
  wire [31:0] n844_I_7_2; // @[Top.scala 1014:22]
  wire [31:0] n844_O_0_0_0; // @[Top.scala 1014:22]
  wire [31:0] n844_O_0_0_1; // @[Top.scala 1014:22]
  wire [31:0] n844_O_0_0_2; // @[Top.scala 1014:22]
  wire [31:0] n844_O_1_0_0; // @[Top.scala 1014:22]
  wire [31:0] n844_O_1_0_1; // @[Top.scala 1014:22]
  wire [31:0] n844_O_1_0_2; // @[Top.scala 1014:22]
  wire [31:0] n844_O_2_0_0; // @[Top.scala 1014:22]
  wire [31:0] n844_O_2_0_1; // @[Top.scala 1014:22]
  wire [31:0] n844_O_2_0_2; // @[Top.scala 1014:22]
  wire [31:0] n844_O_3_0_0; // @[Top.scala 1014:22]
  wire [31:0] n844_O_3_0_1; // @[Top.scala 1014:22]
  wire [31:0] n844_O_3_0_2; // @[Top.scala 1014:22]
  wire [31:0] n844_O_4_0_0; // @[Top.scala 1014:22]
  wire [31:0] n844_O_4_0_1; // @[Top.scala 1014:22]
  wire [31:0] n844_O_4_0_2; // @[Top.scala 1014:22]
  wire [31:0] n844_O_5_0_0; // @[Top.scala 1014:22]
  wire [31:0] n844_O_5_0_1; // @[Top.scala 1014:22]
  wire [31:0] n844_O_5_0_2; // @[Top.scala 1014:22]
  wire [31:0] n844_O_6_0_0; // @[Top.scala 1014:22]
  wire [31:0] n844_O_6_0_1; // @[Top.scala 1014:22]
  wire [31:0] n844_O_6_0_2; // @[Top.scala 1014:22]
  wire [31:0] n844_O_7_0_0; // @[Top.scala 1014:22]
  wire [31:0] n844_O_7_0_1; // @[Top.scala 1014:22]
  wire [31:0] n844_O_7_0_2; // @[Top.scala 1014:22]
  wire  n851_valid_up; // @[Top.scala 1017:22]
  wire  n851_valid_down; // @[Top.scala 1017:22]
  wire [31:0] n851_I_0_0_0; // @[Top.scala 1017:22]
  wire [31:0] n851_I_0_0_1; // @[Top.scala 1017:22]
  wire [31:0] n851_I_0_0_2; // @[Top.scala 1017:22]
  wire [31:0] n851_I_1_0_0; // @[Top.scala 1017:22]
  wire [31:0] n851_I_1_0_1; // @[Top.scala 1017:22]
  wire [31:0] n851_I_1_0_2; // @[Top.scala 1017:22]
  wire [31:0] n851_I_2_0_0; // @[Top.scala 1017:22]
  wire [31:0] n851_I_2_0_1; // @[Top.scala 1017:22]
  wire [31:0] n851_I_2_0_2; // @[Top.scala 1017:22]
  wire [31:0] n851_I_3_0_0; // @[Top.scala 1017:22]
  wire [31:0] n851_I_3_0_1; // @[Top.scala 1017:22]
  wire [31:0] n851_I_3_0_2; // @[Top.scala 1017:22]
  wire [31:0] n851_I_4_0_0; // @[Top.scala 1017:22]
  wire [31:0] n851_I_4_0_1; // @[Top.scala 1017:22]
  wire [31:0] n851_I_4_0_2; // @[Top.scala 1017:22]
  wire [31:0] n851_I_5_0_0; // @[Top.scala 1017:22]
  wire [31:0] n851_I_5_0_1; // @[Top.scala 1017:22]
  wire [31:0] n851_I_5_0_2; // @[Top.scala 1017:22]
  wire [31:0] n851_I_6_0_0; // @[Top.scala 1017:22]
  wire [31:0] n851_I_6_0_1; // @[Top.scala 1017:22]
  wire [31:0] n851_I_6_0_2; // @[Top.scala 1017:22]
  wire [31:0] n851_I_7_0_0; // @[Top.scala 1017:22]
  wire [31:0] n851_I_7_0_1; // @[Top.scala 1017:22]
  wire [31:0] n851_I_7_0_2; // @[Top.scala 1017:22]
  wire [31:0] n851_O_0_0; // @[Top.scala 1017:22]
  wire [31:0] n851_O_0_1; // @[Top.scala 1017:22]
  wire [31:0] n851_O_0_2; // @[Top.scala 1017:22]
  wire [31:0] n851_O_1_0; // @[Top.scala 1017:22]
  wire [31:0] n851_O_1_1; // @[Top.scala 1017:22]
  wire [31:0] n851_O_1_2; // @[Top.scala 1017:22]
  wire [31:0] n851_O_2_0; // @[Top.scala 1017:22]
  wire [31:0] n851_O_2_1; // @[Top.scala 1017:22]
  wire [31:0] n851_O_2_2; // @[Top.scala 1017:22]
  wire [31:0] n851_O_3_0; // @[Top.scala 1017:22]
  wire [31:0] n851_O_3_1; // @[Top.scala 1017:22]
  wire [31:0] n851_O_3_2; // @[Top.scala 1017:22]
  wire [31:0] n851_O_4_0; // @[Top.scala 1017:22]
  wire [31:0] n851_O_4_1; // @[Top.scala 1017:22]
  wire [31:0] n851_O_4_2; // @[Top.scala 1017:22]
  wire [31:0] n851_O_5_0; // @[Top.scala 1017:22]
  wire [31:0] n851_O_5_1; // @[Top.scala 1017:22]
  wire [31:0] n851_O_5_2; // @[Top.scala 1017:22]
  wire [31:0] n851_O_6_0; // @[Top.scala 1017:22]
  wire [31:0] n851_O_6_1; // @[Top.scala 1017:22]
  wire [31:0] n851_O_6_2; // @[Top.scala 1017:22]
  wire [31:0] n851_O_7_0; // @[Top.scala 1017:22]
  wire [31:0] n851_O_7_1; // @[Top.scala 1017:22]
  wire [31:0] n851_O_7_2; // @[Top.scala 1017:22]
  wire  n852_clock; // @[Top.scala 1020:22]
  wire  n852_valid_up; // @[Top.scala 1020:22]
  wire  n852_valid_down; // @[Top.scala 1020:22]
  wire [31:0] n852_I_0; // @[Top.scala 1020:22]
  wire [31:0] n852_I_1; // @[Top.scala 1020:22]
  wire [31:0] n852_I_2; // @[Top.scala 1020:22]
  wire [31:0] n852_I_3; // @[Top.scala 1020:22]
  wire [31:0] n852_I_4; // @[Top.scala 1020:22]
  wire [31:0] n852_I_5; // @[Top.scala 1020:22]
  wire [31:0] n852_I_6; // @[Top.scala 1020:22]
  wire [31:0] n852_I_7; // @[Top.scala 1020:22]
  wire [31:0] n852_O_0; // @[Top.scala 1020:22]
  wire [31:0] n852_O_1; // @[Top.scala 1020:22]
  wire [31:0] n852_O_2; // @[Top.scala 1020:22]
  wire [31:0] n852_O_3; // @[Top.scala 1020:22]
  wire [31:0] n852_O_4; // @[Top.scala 1020:22]
  wire [31:0] n852_O_5; // @[Top.scala 1020:22]
  wire [31:0] n852_O_6; // @[Top.scala 1020:22]
  wire [31:0] n852_O_7; // @[Top.scala 1020:22]
  wire  n853_clock; // @[Top.scala 1023:22]
  wire  n853_valid_up; // @[Top.scala 1023:22]
  wire  n853_valid_down; // @[Top.scala 1023:22]
  wire [31:0] n853_I_0; // @[Top.scala 1023:22]
  wire [31:0] n853_I_1; // @[Top.scala 1023:22]
  wire [31:0] n853_I_2; // @[Top.scala 1023:22]
  wire [31:0] n853_I_3; // @[Top.scala 1023:22]
  wire [31:0] n853_I_4; // @[Top.scala 1023:22]
  wire [31:0] n853_I_5; // @[Top.scala 1023:22]
  wire [31:0] n853_I_6; // @[Top.scala 1023:22]
  wire [31:0] n853_I_7; // @[Top.scala 1023:22]
  wire [31:0] n853_O_0; // @[Top.scala 1023:22]
  wire [31:0] n853_O_1; // @[Top.scala 1023:22]
  wire [31:0] n853_O_2; // @[Top.scala 1023:22]
  wire [31:0] n853_O_3; // @[Top.scala 1023:22]
  wire [31:0] n853_O_4; // @[Top.scala 1023:22]
  wire [31:0] n853_O_5; // @[Top.scala 1023:22]
  wire [31:0] n853_O_6; // @[Top.scala 1023:22]
  wire [31:0] n853_O_7; // @[Top.scala 1023:22]
  wire  n854_valid_up; // @[Top.scala 1026:22]
  wire  n854_valid_down; // @[Top.scala 1026:22]
  wire [31:0] n854_I0_0; // @[Top.scala 1026:22]
  wire [31:0] n854_I0_1; // @[Top.scala 1026:22]
  wire [31:0] n854_I0_2; // @[Top.scala 1026:22]
  wire [31:0] n854_I0_3; // @[Top.scala 1026:22]
  wire [31:0] n854_I0_4; // @[Top.scala 1026:22]
  wire [31:0] n854_I0_5; // @[Top.scala 1026:22]
  wire [31:0] n854_I0_6; // @[Top.scala 1026:22]
  wire [31:0] n854_I0_7; // @[Top.scala 1026:22]
  wire [31:0] n854_I1_0; // @[Top.scala 1026:22]
  wire [31:0] n854_I1_1; // @[Top.scala 1026:22]
  wire [31:0] n854_I1_2; // @[Top.scala 1026:22]
  wire [31:0] n854_I1_3; // @[Top.scala 1026:22]
  wire [31:0] n854_I1_4; // @[Top.scala 1026:22]
  wire [31:0] n854_I1_5; // @[Top.scala 1026:22]
  wire [31:0] n854_I1_6; // @[Top.scala 1026:22]
  wire [31:0] n854_I1_7; // @[Top.scala 1026:22]
  wire [31:0] n854_O_0_0; // @[Top.scala 1026:22]
  wire [31:0] n854_O_0_1; // @[Top.scala 1026:22]
  wire [31:0] n854_O_1_0; // @[Top.scala 1026:22]
  wire [31:0] n854_O_1_1; // @[Top.scala 1026:22]
  wire [31:0] n854_O_2_0; // @[Top.scala 1026:22]
  wire [31:0] n854_O_2_1; // @[Top.scala 1026:22]
  wire [31:0] n854_O_3_0; // @[Top.scala 1026:22]
  wire [31:0] n854_O_3_1; // @[Top.scala 1026:22]
  wire [31:0] n854_O_4_0; // @[Top.scala 1026:22]
  wire [31:0] n854_O_4_1; // @[Top.scala 1026:22]
  wire [31:0] n854_O_5_0; // @[Top.scala 1026:22]
  wire [31:0] n854_O_5_1; // @[Top.scala 1026:22]
  wire [31:0] n854_O_6_0; // @[Top.scala 1026:22]
  wire [31:0] n854_O_6_1; // @[Top.scala 1026:22]
  wire [31:0] n854_O_7_0; // @[Top.scala 1026:22]
  wire [31:0] n854_O_7_1; // @[Top.scala 1026:22]
  wire  n861_valid_up; // @[Top.scala 1030:22]
  wire  n861_valid_down; // @[Top.scala 1030:22]
  wire [31:0] n861_I0_0_0; // @[Top.scala 1030:22]
  wire [31:0] n861_I0_0_1; // @[Top.scala 1030:22]
  wire [31:0] n861_I0_1_0; // @[Top.scala 1030:22]
  wire [31:0] n861_I0_1_1; // @[Top.scala 1030:22]
  wire [31:0] n861_I0_2_0; // @[Top.scala 1030:22]
  wire [31:0] n861_I0_2_1; // @[Top.scala 1030:22]
  wire [31:0] n861_I0_3_0; // @[Top.scala 1030:22]
  wire [31:0] n861_I0_3_1; // @[Top.scala 1030:22]
  wire [31:0] n861_I0_4_0; // @[Top.scala 1030:22]
  wire [31:0] n861_I0_4_1; // @[Top.scala 1030:22]
  wire [31:0] n861_I0_5_0; // @[Top.scala 1030:22]
  wire [31:0] n861_I0_5_1; // @[Top.scala 1030:22]
  wire [31:0] n861_I0_6_0; // @[Top.scala 1030:22]
  wire [31:0] n861_I0_6_1; // @[Top.scala 1030:22]
  wire [31:0] n861_I0_7_0; // @[Top.scala 1030:22]
  wire [31:0] n861_I0_7_1; // @[Top.scala 1030:22]
  wire [31:0] n861_I1_0; // @[Top.scala 1030:22]
  wire [31:0] n861_I1_1; // @[Top.scala 1030:22]
  wire [31:0] n861_I1_2; // @[Top.scala 1030:22]
  wire [31:0] n861_I1_3; // @[Top.scala 1030:22]
  wire [31:0] n861_I1_4; // @[Top.scala 1030:22]
  wire [31:0] n861_I1_5; // @[Top.scala 1030:22]
  wire [31:0] n861_I1_6; // @[Top.scala 1030:22]
  wire [31:0] n861_I1_7; // @[Top.scala 1030:22]
  wire [31:0] n861_O_0_0; // @[Top.scala 1030:22]
  wire [31:0] n861_O_0_1; // @[Top.scala 1030:22]
  wire [31:0] n861_O_0_2; // @[Top.scala 1030:22]
  wire [31:0] n861_O_1_0; // @[Top.scala 1030:22]
  wire [31:0] n861_O_1_1; // @[Top.scala 1030:22]
  wire [31:0] n861_O_1_2; // @[Top.scala 1030:22]
  wire [31:0] n861_O_2_0; // @[Top.scala 1030:22]
  wire [31:0] n861_O_2_1; // @[Top.scala 1030:22]
  wire [31:0] n861_O_2_2; // @[Top.scala 1030:22]
  wire [31:0] n861_O_3_0; // @[Top.scala 1030:22]
  wire [31:0] n861_O_3_1; // @[Top.scala 1030:22]
  wire [31:0] n861_O_3_2; // @[Top.scala 1030:22]
  wire [31:0] n861_O_4_0; // @[Top.scala 1030:22]
  wire [31:0] n861_O_4_1; // @[Top.scala 1030:22]
  wire [31:0] n861_O_4_2; // @[Top.scala 1030:22]
  wire [31:0] n861_O_5_0; // @[Top.scala 1030:22]
  wire [31:0] n861_O_5_1; // @[Top.scala 1030:22]
  wire [31:0] n861_O_5_2; // @[Top.scala 1030:22]
  wire [31:0] n861_O_6_0; // @[Top.scala 1030:22]
  wire [31:0] n861_O_6_1; // @[Top.scala 1030:22]
  wire [31:0] n861_O_6_2; // @[Top.scala 1030:22]
  wire [31:0] n861_O_7_0; // @[Top.scala 1030:22]
  wire [31:0] n861_O_7_1; // @[Top.scala 1030:22]
  wire [31:0] n861_O_7_2; // @[Top.scala 1030:22]
  wire  n870_valid_up; // @[Top.scala 1034:22]
  wire  n870_valid_down; // @[Top.scala 1034:22]
  wire [31:0] n870_I_0_0; // @[Top.scala 1034:22]
  wire [31:0] n870_I_0_1; // @[Top.scala 1034:22]
  wire [31:0] n870_I_0_2; // @[Top.scala 1034:22]
  wire [31:0] n870_I_1_0; // @[Top.scala 1034:22]
  wire [31:0] n870_I_1_1; // @[Top.scala 1034:22]
  wire [31:0] n870_I_1_2; // @[Top.scala 1034:22]
  wire [31:0] n870_I_2_0; // @[Top.scala 1034:22]
  wire [31:0] n870_I_2_1; // @[Top.scala 1034:22]
  wire [31:0] n870_I_2_2; // @[Top.scala 1034:22]
  wire [31:0] n870_I_3_0; // @[Top.scala 1034:22]
  wire [31:0] n870_I_3_1; // @[Top.scala 1034:22]
  wire [31:0] n870_I_3_2; // @[Top.scala 1034:22]
  wire [31:0] n870_I_4_0; // @[Top.scala 1034:22]
  wire [31:0] n870_I_4_1; // @[Top.scala 1034:22]
  wire [31:0] n870_I_4_2; // @[Top.scala 1034:22]
  wire [31:0] n870_I_5_0; // @[Top.scala 1034:22]
  wire [31:0] n870_I_5_1; // @[Top.scala 1034:22]
  wire [31:0] n870_I_5_2; // @[Top.scala 1034:22]
  wire [31:0] n870_I_6_0; // @[Top.scala 1034:22]
  wire [31:0] n870_I_6_1; // @[Top.scala 1034:22]
  wire [31:0] n870_I_6_2; // @[Top.scala 1034:22]
  wire [31:0] n870_I_7_0; // @[Top.scala 1034:22]
  wire [31:0] n870_I_7_1; // @[Top.scala 1034:22]
  wire [31:0] n870_I_7_2; // @[Top.scala 1034:22]
  wire [31:0] n870_O_0_0_0; // @[Top.scala 1034:22]
  wire [31:0] n870_O_0_0_1; // @[Top.scala 1034:22]
  wire [31:0] n870_O_0_0_2; // @[Top.scala 1034:22]
  wire [31:0] n870_O_1_0_0; // @[Top.scala 1034:22]
  wire [31:0] n870_O_1_0_1; // @[Top.scala 1034:22]
  wire [31:0] n870_O_1_0_2; // @[Top.scala 1034:22]
  wire [31:0] n870_O_2_0_0; // @[Top.scala 1034:22]
  wire [31:0] n870_O_2_0_1; // @[Top.scala 1034:22]
  wire [31:0] n870_O_2_0_2; // @[Top.scala 1034:22]
  wire [31:0] n870_O_3_0_0; // @[Top.scala 1034:22]
  wire [31:0] n870_O_3_0_1; // @[Top.scala 1034:22]
  wire [31:0] n870_O_3_0_2; // @[Top.scala 1034:22]
  wire [31:0] n870_O_4_0_0; // @[Top.scala 1034:22]
  wire [31:0] n870_O_4_0_1; // @[Top.scala 1034:22]
  wire [31:0] n870_O_4_0_2; // @[Top.scala 1034:22]
  wire [31:0] n870_O_5_0_0; // @[Top.scala 1034:22]
  wire [31:0] n870_O_5_0_1; // @[Top.scala 1034:22]
  wire [31:0] n870_O_5_0_2; // @[Top.scala 1034:22]
  wire [31:0] n870_O_6_0_0; // @[Top.scala 1034:22]
  wire [31:0] n870_O_6_0_1; // @[Top.scala 1034:22]
  wire [31:0] n870_O_6_0_2; // @[Top.scala 1034:22]
  wire [31:0] n870_O_7_0_0; // @[Top.scala 1034:22]
  wire [31:0] n870_O_7_0_1; // @[Top.scala 1034:22]
  wire [31:0] n870_O_7_0_2; // @[Top.scala 1034:22]
  wire  n877_valid_up; // @[Top.scala 1037:22]
  wire  n877_valid_down; // @[Top.scala 1037:22]
  wire [31:0] n877_I_0_0_0; // @[Top.scala 1037:22]
  wire [31:0] n877_I_0_0_1; // @[Top.scala 1037:22]
  wire [31:0] n877_I_0_0_2; // @[Top.scala 1037:22]
  wire [31:0] n877_I_1_0_0; // @[Top.scala 1037:22]
  wire [31:0] n877_I_1_0_1; // @[Top.scala 1037:22]
  wire [31:0] n877_I_1_0_2; // @[Top.scala 1037:22]
  wire [31:0] n877_I_2_0_0; // @[Top.scala 1037:22]
  wire [31:0] n877_I_2_0_1; // @[Top.scala 1037:22]
  wire [31:0] n877_I_2_0_2; // @[Top.scala 1037:22]
  wire [31:0] n877_I_3_0_0; // @[Top.scala 1037:22]
  wire [31:0] n877_I_3_0_1; // @[Top.scala 1037:22]
  wire [31:0] n877_I_3_0_2; // @[Top.scala 1037:22]
  wire [31:0] n877_I_4_0_0; // @[Top.scala 1037:22]
  wire [31:0] n877_I_4_0_1; // @[Top.scala 1037:22]
  wire [31:0] n877_I_4_0_2; // @[Top.scala 1037:22]
  wire [31:0] n877_I_5_0_0; // @[Top.scala 1037:22]
  wire [31:0] n877_I_5_0_1; // @[Top.scala 1037:22]
  wire [31:0] n877_I_5_0_2; // @[Top.scala 1037:22]
  wire [31:0] n877_I_6_0_0; // @[Top.scala 1037:22]
  wire [31:0] n877_I_6_0_1; // @[Top.scala 1037:22]
  wire [31:0] n877_I_6_0_2; // @[Top.scala 1037:22]
  wire [31:0] n877_I_7_0_0; // @[Top.scala 1037:22]
  wire [31:0] n877_I_7_0_1; // @[Top.scala 1037:22]
  wire [31:0] n877_I_7_0_2; // @[Top.scala 1037:22]
  wire [31:0] n877_O_0_0; // @[Top.scala 1037:22]
  wire [31:0] n877_O_0_1; // @[Top.scala 1037:22]
  wire [31:0] n877_O_0_2; // @[Top.scala 1037:22]
  wire [31:0] n877_O_1_0; // @[Top.scala 1037:22]
  wire [31:0] n877_O_1_1; // @[Top.scala 1037:22]
  wire [31:0] n877_O_1_2; // @[Top.scala 1037:22]
  wire [31:0] n877_O_2_0; // @[Top.scala 1037:22]
  wire [31:0] n877_O_2_1; // @[Top.scala 1037:22]
  wire [31:0] n877_O_2_2; // @[Top.scala 1037:22]
  wire [31:0] n877_O_3_0; // @[Top.scala 1037:22]
  wire [31:0] n877_O_3_1; // @[Top.scala 1037:22]
  wire [31:0] n877_O_3_2; // @[Top.scala 1037:22]
  wire [31:0] n877_O_4_0; // @[Top.scala 1037:22]
  wire [31:0] n877_O_4_1; // @[Top.scala 1037:22]
  wire [31:0] n877_O_4_2; // @[Top.scala 1037:22]
  wire [31:0] n877_O_5_0; // @[Top.scala 1037:22]
  wire [31:0] n877_O_5_1; // @[Top.scala 1037:22]
  wire [31:0] n877_O_5_2; // @[Top.scala 1037:22]
  wire [31:0] n877_O_6_0; // @[Top.scala 1037:22]
  wire [31:0] n877_O_6_1; // @[Top.scala 1037:22]
  wire [31:0] n877_O_6_2; // @[Top.scala 1037:22]
  wire [31:0] n877_O_7_0; // @[Top.scala 1037:22]
  wire [31:0] n877_O_7_1; // @[Top.scala 1037:22]
  wire [31:0] n877_O_7_2; // @[Top.scala 1037:22]
  wire  n878_valid_up; // @[Top.scala 1040:22]
  wire  n878_valid_down; // @[Top.scala 1040:22]
  wire [31:0] n878_I0_0_0; // @[Top.scala 1040:22]
  wire [31:0] n878_I0_0_1; // @[Top.scala 1040:22]
  wire [31:0] n878_I0_0_2; // @[Top.scala 1040:22]
  wire [31:0] n878_I0_1_0; // @[Top.scala 1040:22]
  wire [31:0] n878_I0_1_1; // @[Top.scala 1040:22]
  wire [31:0] n878_I0_1_2; // @[Top.scala 1040:22]
  wire [31:0] n878_I0_2_0; // @[Top.scala 1040:22]
  wire [31:0] n878_I0_2_1; // @[Top.scala 1040:22]
  wire [31:0] n878_I0_2_2; // @[Top.scala 1040:22]
  wire [31:0] n878_I0_3_0; // @[Top.scala 1040:22]
  wire [31:0] n878_I0_3_1; // @[Top.scala 1040:22]
  wire [31:0] n878_I0_3_2; // @[Top.scala 1040:22]
  wire [31:0] n878_I0_4_0; // @[Top.scala 1040:22]
  wire [31:0] n878_I0_4_1; // @[Top.scala 1040:22]
  wire [31:0] n878_I0_4_2; // @[Top.scala 1040:22]
  wire [31:0] n878_I0_5_0; // @[Top.scala 1040:22]
  wire [31:0] n878_I0_5_1; // @[Top.scala 1040:22]
  wire [31:0] n878_I0_5_2; // @[Top.scala 1040:22]
  wire [31:0] n878_I0_6_0; // @[Top.scala 1040:22]
  wire [31:0] n878_I0_6_1; // @[Top.scala 1040:22]
  wire [31:0] n878_I0_6_2; // @[Top.scala 1040:22]
  wire [31:0] n878_I0_7_0; // @[Top.scala 1040:22]
  wire [31:0] n878_I0_7_1; // @[Top.scala 1040:22]
  wire [31:0] n878_I0_7_2; // @[Top.scala 1040:22]
  wire [31:0] n878_I1_0_0; // @[Top.scala 1040:22]
  wire [31:0] n878_I1_0_1; // @[Top.scala 1040:22]
  wire [31:0] n878_I1_0_2; // @[Top.scala 1040:22]
  wire [31:0] n878_I1_1_0; // @[Top.scala 1040:22]
  wire [31:0] n878_I1_1_1; // @[Top.scala 1040:22]
  wire [31:0] n878_I1_1_2; // @[Top.scala 1040:22]
  wire [31:0] n878_I1_2_0; // @[Top.scala 1040:22]
  wire [31:0] n878_I1_2_1; // @[Top.scala 1040:22]
  wire [31:0] n878_I1_2_2; // @[Top.scala 1040:22]
  wire [31:0] n878_I1_3_0; // @[Top.scala 1040:22]
  wire [31:0] n878_I1_3_1; // @[Top.scala 1040:22]
  wire [31:0] n878_I1_3_2; // @[Top.scala 1040:22]
  wire [31:0] n878_I1_4_0; // @[Top.scala 1040:22]
  wire [31:0] n878_I1_4_1; // @[Top.scala 1040:22]
  wire [31:0] n878_I1_4_2; // @[Top.scala 1040:22]
  wire [31:0] n878_I1_5_0; // @[Top.scala 1040:22]
  wire [31:0] n878_I1_5_1; // @[Top.scala 1040:22]
  wire [31:0] n878_I1_5_2; // @[Top.scala 1040:22]
  wire [31:0] n878_I1_6_0; // @[Top.scala 1040:22]
  wire [31:0] n878_I1_6_1; // @[Top.scala 1040:22]
  wire [31:0] n878_I1_6_2; // @[Top.scala 1040:22]
  wire [31:0] n878_I1_7_0; // @[Top.scala 1040:22]
  wire [31:0] n878_I1_7_1; // @[Top.scala 1040:22]
  wire [31:0] n878_I1_7_2; // @[Top.scala 1040:22]
  wire [31:0] n878_O_0_0_0; // @[Top.scala 1040:22]
  wire [31:0] n878_O_0_0_1; // @[Top.scala 1040:22]
  wire [31:0] n878_O_0_0_2; // @[Top.scala 1040:22]
  wire [31:0] n878_O_0_1_0; // @[Top.scala 1040:22]
  wire [31:0] n878_O_0_1_1; // @[Top.scala 1040:22]
  wire [31:0] n878_O_0_1_2; // @[Top.scala 1040:22]
  wire [31:0] n878_O_1_0_0; // @[Top.scala 1040:22]
  wire [31:0] n878_O_1_0_1; // @[Top.scala 1040:22]
  wire [31:0] n878_O_1_0_2; // @[Top.scala 1040:22]
  wire [31:0] n878_O_1_1_0; // @[Top.scala 1040:22]
  wire [31:0] n878_O_1_1_1; // @[Top.scala 1040:22]
  wire [31:0] n878_O_1_1_2; // @[Top.scala 1040:22]
  wire [31:0] n878_O_2_0_0; // @[Top.scala 1040:22]
  wire [31:0] n878_O_2_0_1; // @[Top.scala 1040:22]
  wire [31:0] n878_O_2_0_2; // @[Top.scala 1040:22]
  wire [31:0] n878_O_2_1_0; // @[Top.scala 1040:22]
  wire [31:0] n878_O_2_1_1; // @[Top.scala 1040:22]
  wire [31:0] n878_O_2_1_2; // @[Top.scala 1040:22]
  wire [31:0] n878_O_3_0_0; // @[Top.scala 1040:22]
  wire [31:0] n878_O_3_0_1; // @[Top.scala 1040:22]
  wire [31:0] n878_O_3_0_2; // @[Top.scala 1040:22]
  wire [31:0] n878_O_3_1_0; // @[Top.scala 1040:22]
  wire [31:0] n878_O_3_1_1; // @[Top.scala 1040:22]
  wire [31:0] n878_O_3_1_2; // @[Top.scala 1040:22]
  wire [31:0] n878_O_4_0_0; // @[Top.scala 1040:22]
  wire [31:0] n878_O_4_0_1; // @[Top.scala 1040:22]
  wire [31:0] n878_O_4_0_2; // @[Top.scala 1040:22]
  wire [31:0] n878_O_4_1_0; // @[Top.scala 1040:22]
  wire [31:0] n878_O_4_1_1; // @[Top.scala 1040:22]
  wire [31:0] n878_O_4_1_2; // @[Top.scala 1040:22]
  wire [31:0] n878_O_5_0_0; // @[Top.scala 1040:22]
  wire [31:0] n878_O_5_0_1; // @[Top.scala 1040:22]
  wire [31:0] n878_O_5_0_2; // @[Top.scala 1040:22]
  wire [31:0] n878_O_5_1_0; // @[Top.scala 1040:22]
  wire [31:0] n878_O_5_1_1; // @[Top.scala 1040:22]
  wire [31:0] n878_O_5_1_2; // @[Top.scala 1040:22]
  wire [31:0] n878_O_6_0_0; // @[Top.scala 1040:22]
  wire [31:0] n878_O_6_0_1; // @[Top.scala 1040:22]
  wire [31:0] n878_O_6_0_2; // @[Top.scala 1040:22]
  wire [31:0] n878_O_6_1_0; // @[Top.scala 1040:22]
  wire [31:0] n878_O_6_1_1; // @[Top.scala 1040:22]
  wire [31:0] n878_O_6_1_2; // @[Top.scala 1040:22]
  wire [31:0] n878_O_7_0_0; // @[Top.scala 1040:22]
  wire [31:0] n878_O_7_0_1; // @[Top.scala 1040:22]
  wire [31:0] n878_O_7_0_2; // @[Top.scala 1040:22]
  wire [31:0] n878_O_7_1_0; // @[Top.scala 1040:22]
  wire [31:0] n878_O_7_1_1; // @[Top.scala 1040:22]
  wire [31:0] n878_O_7_1_2; // @[Top.scala 1040:22]
  wire  n885_clock; // @[Top.scala 1044:22]
  wire  n885_valid_up; // @[Top.scala 1044:22]
  wire  n885_valid_down; // @[Top.scala 1044:22]
  wire [31:0] n885_I_0; // @[Top.scala 1044:22]
  wire [31:0] n885_I_1; // @[Top.scala 1044:22]
  wire [31:0] n885_I_2; // @[Top.scala 1044:22]
  wire [31:0] n885_I_3; // @[Top.scala 1044:22]
  wire [31:0] n885_I_4; // @[Top.scala 1044:22]
  wire [31:0] n885_I_5; // @[Top.scala 1044:22]
  wire [31:0] n885_I_6; // @[Top.scala 1044:22]
  wire [31:0] n885_I_7; // @[Top.scala 1044:22]
  wire [31:0] n885_O_0; // @[Top.scala 1044:22]
  wire [31:0] n885_O_1; // @[Top.scala 1044:22]
  wire [31:0] n885_O_2; // @[Top.scala 1044:22]
  wire [31:0] n885_O_3; // @[Top.scala 1044:22]
  wire [31:0] n885_O_4; // @[Top.scala 1044:22]
  wire [31:0] n885_O_5; // @[Top.scala 1044:22]
  wire [31:0] n885_O_6; // @[Top.scala 1044:22]
  wire [31:0] n885_O_7; // @[Top.scala 1044:22]
  wire  n886_clock; // @[Top.scala 1047:22]
  wire  n886_valid_up; // @[Top.scala 1047:22]
  wire  n886_valid_down; // @[Top.scala 1047:22]
  wire [31:0] n886_I_0; // @[Top.scala 1047:22]
  wire [31:0] n886_I_1; // @[Top.scala 1047:22]
  wire [31:0] n886_I_2; // @[Top.scala 1047:22]
  wire [31:0] n886_I_3; // @[Top.scala 1047:22]
  wire [31:0] n886_I_4; // @[Top.scala 1047:22]
  wire [31:0] n886_I_5; // @[Top.scala 1047:22]
  wire [31:0] n886_I_6; // @[Top.scala 1047:22]
  wire [31:0] n886_I_7; // @[Top.scala 1047:22]
  wire [31:0] n886_O_0; // @[Top.scala 1047:22]
  wire [31:0] n886_O_1; // @[Top.scala 1047:22]
  wire [31:0] n886_O_2; // @[Top.scala 1047:22]
  wire [31:0] n886_O_3; // @[Top.scala 1047:22]
  wire [31:0] n886_O_4; // @[Top.scala 1047:22]
  wire [31:0] n886_O_5; // @[Top.scala 1047:22]
  wire [31:0] n886_O_6; // @[Top.scala 1047:22]
  wire [31:0] n886_O_7; // @[Top.scala 1047:22]
  wire  n887_valid_up; // @[Top.scala 1050:22]
  wire  n887_valid_down; // @[Top.scala 1050:22]
  wire [31:0] n887_I0_0; // @[Top.scala 1050:22]
  wire [31:0] n887_I0_1; // @[Top.scala 1050:22]
  wire [31:0] n887_I0_2; // @[Top.scala 1050:22]
  wire [31:0] n887_I0_3; // @[Top.scala 1050:22]
  wire [31:0] n887_I0_4; // @[Top.scala 1050:22]
  wire [31:0] n887_I0_5; // @[Top.scala 1050:22]
  wire [31:0] n887_I0_6; // @[Top.scala 1050:22]
  wire [31:0] n887_I0_7; // @[Top.scala 1050:22]
  wire [31:0] n887_I1_0; // @[Top.scala 1050:22]
  wire [31:0] n887_I1_1; // @[Top.scala 1050:22]
  wire [31:0] n887_I1_2; // @[Top.scala 1050:22]
  wire [31:0] n887_I1_3; // @[Top.scala 1050:22]
  wire [31:0] n887_I1_4; // @[Top.scala 1050:22]
  wire [31:0] n887_I1_5; // @[Top.scala 1050:22]
  wire [31:0] n887_I1_6; // @[Top.scala 1050:22]
  wire [31:0] n887_I1_7; // @[Top.scala 1050:22]
  wire [31:0] n887_O_0_0; // @[Top.scala 1050:22]
  wire [31:0] n887_O_0_1; // @[Top.scala 1050:22]
  wire [31:0] n887_O_1_0; // @[Top.scala 1050:22]
  wire [31:0] n887_O_1_1; // @[Top.scala 1050:22]
  wire [31:0] n887_O_2_0; // @[Top.scala 1050:22]
  wire [31:0] n887_O_2_1; // @[Top.scala 1050:22]
  wire [31:0] n887_O_3_0; // @[Top.scala 1050:22]
  wire [31:0] n887_O_3_1; // @[Top.scala 1050:22]
  wire [31:0] n887_O_4_0; // @[Top.scala 1050:22]
  wire [31:0] n887_O_4_1; // @[Top.scala 1050:22]
  wire [31:0] n887_O_5_0; // @[Top.scala 1050:22]
  wire [31:0] n887_O_5_1; // @[Top.scala 1050:22]
  wire [31:0] n887_O_6_0; // @[Top.scala 1050:22]
  wire [31:0] n887_O_6_1; // @[Top.scala 1050:22]
  wire [31:0] n887_O_7_0; // @[Top.scala 1050:22]
  wire [31:0] n887_O_7_1; // @[Top.scala 1050:22]
  wire  n894_valid_up; // @[Top.scala 1054:22]
  wire  n894_valid_down; // @[Top.scala 1054:22]
  wire [31:0] n894_I0_0_0; // @[Top.scala 1054:22]
  wire [31:0] n894_I0_0_1; // @[Top.scala 1054:22]
  wire [31:0] n894_I0_1_0; // @[Top.scala 1054:22]
  wire [31:0] n894_I0_1_1; // @[Top.scala 1054:22]
  wire [31:0] n894_I0_2_0; // @[Top.scala 1054:22]
  wire [31:0] n894_I0_2_1; // @[Top.scala 1054:22]
  wire [31:0] n894_I0_3_0; // @[Top.scala 1054:22]
  wire [31:0] n894_I0_3_1; // @[Top.scala 1054:22]
  wire [31:0] n894_I0_4_0; // @[Top.scala 1054:22]
  wire [31:0] n894_I0_4_1; // @[Top.scala 1054:22]
  wire [31:0] n894_I0_5_0; // @[Top.scala 1054:22]
  wire [31:0] n894_I0_5_1; // @[Top.scala 1054:22]
  wire [31:0] n894_I0_6_0; // @[Top.scala 1054:22]
  wire [31:0] n894_I0_6_1; // @[Top.scala 1054:22]
  wire [31:0] n894_I0_7_0; // @[Top.scala 1054:22]
  wire [31:0] n894_I0_7_1; // @[Top.scala 1054:22]
  wire [31:0] n894_I1_0; // @[Top.scala 1054:22]
  wire [31:0] n894_I1_1; // @[Top.scala 1054:22]
  wire [31:0] n894_I1_2; // @[Top.scala 1054:22]
  wire [31:0] n894_I1_3; // @[Top.scala 1054:22]
  wire [31:0] n894_I1_4; // @[Top.scala 1054:22]
  wire [31:0] n894_I1_5; // @[Top.scala 1054:22]
  wire [31:0] n894_I1_6; // @[Top.scala 1054:22]
  wire [31:0] n894_I1_7; // @[Top.scala 1054:22]
  wire [31:0] n894_O_0_0; // @[Top.scala 1054:22]
  wire [31:0] n894_O_0_1; // @[Top.scala 1054:22]
  wire [31:0] n894_O_0_2; // @[Top.scala 1054:22]
  wire [31:0] n894_O_1_0; // @[Top.scala 1054:22]
  wire [31:0] n894_O_1_1; // @[Top.scala 1054:22]
  wire [31:0] n894_O_1_2; // @[Top.scala 1054:22]
  wire [31:0] n894_O_2_0; // @[Top.scala 1054:22]
  wire [31:0] n894_O_2_1; // @[Top.scala 1054:22]
  wire [31:0] n894_O_2_2; // @[Top.scala 1054:22]
  wire [31:0] n894_O_3_0; // @[Top.scala 1054:22]
  wire [31:0] n894_O_3_1; // @[Top.scala 1054:22]
  wire [31:0] n894_O_3_2; // @[Top.scala 1054:22]
  wire [31:0] n894_O_4_0; // @[Top.scala 1054:22]
  wire [31:0] n894_O_4_1; // @[Top.scala 1054:22]
  wire [31:0] n894_O_4_2; // @[Top.scala 1054:22]
  wire [31:0] n894_O_5_0; // @[Top.scala 1054:22]
  wire [31:0] n894_O_5_1; // @[Top.scala 1054:22]
  wire [31:0] n894_O_5_2; // @[Top.scala 1054:22]
  wire [31:0] n894_O_6_0; // @[Top.scala 1054:22]
  wire [31:0] n894_O_6_1; // @[Top.scala 1054:22]
  wire [31:0] n894_O_6_2; // @[Top.scala 1054:22]
  wire [31:0] n894_O_7_0; // @[Top.scala 1054:22]
  wire [31:0] n894_O_7_1; // @[Top.scala 1054:22]
  wire [31:0] n894_O_7_2; // @[Top.scala 1054:22]
  wire  n903_valid_up; // @[Top.scala 1058:22]
  wire  n903_valid_down; // @[Top.scala 1058:22]
  wire [31:0] n903_I_0_0; // @[Top.scala 1058:22]
  wire [31:0] n903_I_0_1; // @[Top.scala 1058:22]
  wire [31:0] n903_I_0_2; // @[Top.scala 1058:22]
  wire [31:0] n903_I_1_0; // @[Top.scala 1058:22]
  wire [31:0] n903_I_1_1; // @[Top.scala 1058:22]
  wire [31:0] n903_I_1_2; // @[Top.scala 1058:22]
  wire [31:0] n903_I_2_0; // @[Top.scala 1058:22]
  wire [31:0] n903_I_2_1; // @[Top.scala 1058:22]
  wire [31:0] n903_I_2_2; // @[Top.scala 1058:22]
  wire [31:0] n903_I_3_0; // @[Top.scala 1058:22]
  wire [31:0] n903_I_3_1; // @[Top.scala 1058:22]
  wire [31:0] n903_I_3_2; // @[Top.scala 1058:22]
  wire [31:0] n903_I_4_0; // @[Top.scala 1058:22]
  wire [31:0] n903_I_4_1; // @[Top.scala 1058:22]
  wire [31:0] n903_I_4_2; // @[Top.scala 1058:22]
  wire [31:0] n903_I_5_0; // @[Top.scala 1058:22]
  wire [31:0] n903_I_5_1; // @[Top.scala 1058:22]
  wire [31:0] n903_I_5_2; // @[Top.scala 1058:22]
  wire [31:0] n903_I_6_0; // @[Top.scala 1058:22]
  wire [31:0] n903_I_6_1; // @[Top.scala 1058:22]
  wire [31:0] n903_I_6_2; // @[Top.scala 1058:22]
  wire [31:0] n903_I_7_0; // @[Top.scala 1058:22]
  wire [31:0] n903_I_7_1; // @[Top.scala 1058:22]
  wire [31:0] n903_I_7_2; // @[Top.scala 1058:22]
  wire [31:0] n903_O_0_0_0; // @[Top.scala 1058:22]
  wire [31:0] n903_O_0_0_1; // @[Top.scala 1058:22]
  wire [31:0] n903_O_0_0_2; // @[Top.scala 1058:22]
  wire [31:0] n903_O_1_0_0; // @[Top.scala 1058:22]
  wire [31:0] n903_O_1_0_1; // @[Top.scala 1058:22]
  wire [31:0] n903_O_1_0_2; // @[Top.scala 1058:22]
  wire [31:0] n903_O_2_0_0; // @[Top.scala 1058:22]
  wire [31:0] n903_O_2_0_1; // @[Top.scala 1058:22]
  wire [31:0] n903_O_2_0_2; // @[Top.scala 1058:22]
  wire [31:0] n903_O_3_0_0; // @[Top.scala 1058:22]
  wire [31:0] n903_O_3_0_1; // @[Top.scala 1058:22]
  wire [31:0] n903_O_3_0_2; // @[Top.scala 1058:22]
  wire [31:0] n903_O_4_0_0; // @[Top.scala 1058:22]
  wire [31:0] n903_O_4_0_1; // @[Top.scala 1058:22]
  wire [31:0] n903_O_4_0_2; // @[Top.scala 1058:22]
  wire [31:0] n903_O_5_0_0; // @[Top.scala 1058:22]
  wire [31:0] n903_O_5_0_1; // @[Top.scala 1058:22]
  wire [31:0] n903_O_5_0_2; // @[Top.scala 1058:22]
  wire [31:0] n903_O_6_0_0; // @[Top.scala 1058:22]
  wire [31:0] n903_O_6_0_1; // @[Top.scala 1058:22]
  wire [31:0] n903_O_6_0_2; // @[Top.scala 1058:22]
  wire [31:0] n903_O_7_0_0; // @[Top.scala 1058:22]
  wire [31:0] n903_O_7_0_1; // @[Top.scala 1058:22]
  wire [31:0] n903_O_7_0_2; // @[Top.scala 1058:22]
  wire  n910_valid_up; // @[Top.scala 1061:22]
  wire  n910_valid_down; // @[Top.scala 1061:22]
  wire [31:0] n910_I_0_0_0; // @[Top.scala 1061:22]
  wire [31:0] n910_I_0_0_1; // @[Top.scala 1061:22]
  wire [31:0] n910_I_0_0_2; // @[Top.scala 1061:22]
  wire [31:0] n910_I_1_0_0; // @[Top.scala 1061:22]
  wire [31:0] n910_I_1_0_1; // @[Top.scala 1061:22]
  wire [31:0] n910_I_1_0_2; // @[Top.scala 1061:22]
  wire [31:0] n910_I_2_0_0; // @[Top.scala 1061:22]
  wire [31:0] n910_I_2_0_1; // @[Top.scala 1061:22]
  wire [31:0] n910_I_2_0_2; // @[Top.scala 1061:22]
  wire [31:0] n910_I_3_0_0; // @[Top.scala 1061:22]
  wire [31:0] n910_I_3_0_1; // @[Top.scala 1061:22]
  wire [31:0] n910_I_3_0_2; // @[Top.scala 1061:22]
  wire [31:0] n910_I_4_0_0; // @[Top.scala 1061:22]
  wire [31:0] n910_I_4_0_1; // @[Top.scala 1061:22]
  wire [31:0] n910_I_4_0_2; // @[Top.scala 1061:22]
  wire [31:0] n910_I_5_0_0; // @[Top.scala 1061:22]
  wire [31:0] n910_I_5_0_1; // @[Top.scala 1061:22]
  wire [31:0] n910_I_5_0_2; // @[Top.scala 1061:22]
  wire [31:0] n910_I_6_0_0; // @[Top.scala 1061:22]
  wire [31:0] n910_I_6_0_1; // @[Top.scala 1061:22]
  wire [31:0] n910_I_6_0_2; // @[Top.scala 1061:22]
  wire [31:0] n910_I_7_0_0; // @[Top.scala 1061:22]
  wire [31:0] n910_I_7_0_1; // @[Top.scala 1061:22]
  wire [31:0] n910_I_7_0_2; // @[Top.scala 1061:22]
  wire [31:0] n910_O_0_0; // @[Top.scala 1061:22]
  wire [31:0] n910_O_0_1; // @[Top.scala 1061:22]
  wire [31:0] n910_O_0_2; // @[Top.scala 1061:22]
  wire [31:0] n910_O_1_0; // @[Top.scala 1061:22]
  wire [31:0] n910_O_1_1; // @[Top.scala 1061:22]
  wire [31:0] n910_O_1_2; // @[Top.scala 1061:22]
  wire [31:0] n910_O_2_0; // @[Top.scala 1061:22]
  wire [31:0] n910_O_2_1; // @[Top.scala 1061:22]
  wire [31:0] n910_O_2_2; // @[Top.scala 1061:22]
  wire [31:0] n910_O_3_0; // @[Top.scala 1061:22]
  wire [31:0] n910_O_3_1; // @[Top.scala 1061:22]
  wire [31:0] n910_O_3_2; // @[Top.scala 1061:22]
  wire [31:0] n910_O_4_0; // @[Top.scala 1061:22]
  wire [31:0] n910_O_4_1; // @[Top.scala 1061:22]
  wire [31:0] n910_O_4_2; // @[Top.scala 1061:22]
  wire [31:0] n910_O_5_0; // @[Top.scala 1061:22]
  wire [31:0] n910_O_5_1; // @[Top.scala 1061:22]
  wire [31:0] n910_O_5_2; // @[Top.scala 1061:22]
  wire [31:0] n910_O_6_0; // @[Top.scala 1061:22]
  wire [31:0] n910_O_6_1; // @[Top.scala 1061:22]
  wire [31:0] n910_O_6_2; // @[Top.scala 1061:22]
  wire [31:0] n910_O_7_0; // @[Top.scala 1061:22]
  wire [31:0] n910_O_7_1; // @[Top.scala 1061:22]
  wire [31:0] n910_O_7_2; // @[Top.scala 1061:22]
  wire  n911_valid_up; // @[Top.scala 1064:22]
  wire  n911_valid_down; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_0_0_0; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_0_0_1; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_0_0_2; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_0_1_0; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_0_1_1; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_0_1_2; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_1_0_0; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_1_0_1; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_1_0_2; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_1_1_0; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_1_1_1; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_1_1_2; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_2_0_0; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_2_0_1; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_2_0_2; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_2_1_0; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_2_1_1; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_2_1_2; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_3_0_0; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_3_0_1; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_3_0_2; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_3_1_0; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_3_1_1; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_3_1_2; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_4_0_0; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_4_0_1; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_4_0_2; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_4_1_0; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_4_1_1; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_4_1_2; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_5_0_0; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_5_0_1; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_5_0_2; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_5_1_0; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_5_1_1; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_5_1_2; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_6_0_0; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_6_0_1; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_6_0_2; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_6_1_0; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_6_1_1; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_6_1_2; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_7_0_0; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_7_0_1; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_7_0_2; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_7_1_0; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_7_1_1; // @[Top.scala 1064:22]
  wire [31:0] n911_I0_7_1_2; // @[Top.scala 1064:22]
  wire [31:0] n911_I1_0_0; // @[Top.scala 1064:22]
  wire [31:0] n911_I1_0_1; // @[Top.scala 1064:22]
  wire [31:0] n911_I1_0_2; // @[Top.scala 1064:22]
  wire [31:0] n911_I1_1_0; // @[Top.scala 1064:22]
  wire [31:0] n911_I1_1_1; // @[Top.scala 1064:22]
  wire [31:0] n911_I1_1_2; // @[Top.scala 1064:22]
  wire [31:0] n911_I1_2_0; // @[Top.scala 1064:22]
  wire [31:0] n911_I1_2_1; // @[Top.scala 1064:22]
  wire [31:0] n911_I1_2_2; // @[Top.scala 1064:22]
  wire [31:0] n911_I1_3_0; // @[Top.scala 1064:22]
  wire [31:0] n911_I1_3_1; // @[Top.scala 1064:22]
  wire [31:0] n911_I1_3_2; // @[Top.scala 1064:22]
  wire [31:0] n911_I1_4_0; // @[Top.scala 1064:22]
  wire [31:0] n911_I1_4_1; // @[Top.scala 1064:22]
  wire [31:0] n911_I1_4_2; // @[Top.scala 1064:22]
  wire [31:0] n911_I1_5_0; // @[Top.scala 1064:22]
  wire [31:0] n911_I1_5_1; // @[Top.scala 1064:22]
  wire [31:0] n911_I1_5_2; // @[Top.scala 1064:22]
  wire [31:0] n911_I1_6_0; // @[Top.scala 1064:22]
  wire [31:0] n911_I1_6_1; // @[Top.scala 1064:22]
  wire [31:0] n911_I1_6_2; // @[Top.scala 1064:22]
  wire [31:0] n911_I1_7_0; // @[Top.scala 1064:22]
  wire [31:0] n911_I1_7_1; // @[Top.scala 1064:22]
  wire [31:0] n911_I1_7_2; // @[Top.scala 1064:22]
  wire [31:0] n911_O_0_0_0; // @[Top.scala 1064:22]
  wire [31:0] n911_O_0_0_1; // @[Top.scala 1064:22]
  wire [31:0] n911_O_0_0_2; // @[Top.scala 1064:22]
  wire [31:0] n911_O_0_1_0; // @[Top.scala 1064:22]
  wire [31:0] n911_O_0_1_1; // @[Top.scala 1064:22]
  wire [31:0] n911_O_0_1_2; // @[Top.scala 1064:22]
  wire [31:0] n911_O_0_2_0; // @[Top.scala 1064:22]
  wire [31:0] n911_O_0_2_1; // @[Top.scala 1064:22]
  wire [31:0] n911_O_0_2_2; // @[Top.scala 1064:22]
  wire [31:0] n911_O_1_0_0; // @[Top.scala 1064:22]
  wire [31:0] n911_O_1_0_1; // @[Top.scala 1064:22]
  wire [31:0] n911_O_1_0_2; // @[Top.scala 1064:22]
  wire [31:0] n911_O_1_1_0; // @[Top.scala 1064:22]
  wire [31:0] n911_O_1_1_1; // @[Top.scala 1064:22]
  wire [31:0] n911_O_1_1_2; // @[Top.scala 1064:22]
  wire [31:0] n911_O_1_2_0; // @[Top.scala 1064:22]
  wire [31:0] n911_O_1_2_1; // @[Top.scala 1064:22]
  wire [31:0] n911_O_1_2_2; // @[Top.scala 1064:22]
  wire [31:0] n911_O_2_0_0; // @[Top.scala 1064:22]
  wire [31:0] n911_O_2_0_1; // @[Top.scala 1064:22]
  wire [31:0] n911_O_2_0_2; // @[Top.scala 1064:22]
  wire [31:0] n911_O_2_1_0; // @[Top.scala 1064:22]
  wire [31:0] n911_O_2_1_1; // @[Top.scala 1064:22]
  wire [31:0] n911_O_2_1_2; // @[Top.scala 1064:22]
  wire [31:0] n911_O_2_2_0; // @[Top.scala 1064:22]
  wire [31:0] n911_O_2_2_1; // @[Top.scala 1064:22]
  wire [31:0] n911_O_2_2_2; // @[Top.scala 1064:22]
  wire [31:0] n911_O_3_0_0; // @[Top.scala 1064:22]
  wire [31:0] n911_O_3_0_1; // @[Top.scala 1064:22]
  wire [31:0] n911_O_3_0_2; // @[Top.scala 1064:22]
  wire [31:0] n911_O_3_1_0; // @[Top.scala 1064:22]
  wire [31:0] n911_O_3_1_1; // @[Top.scala 1064:22]
  wire [31:0] n911_O_3_1_2; // @[Top.scala 1064:22]
  wire [31:0] n911_O_3_2_0; // @[Top.scala 1064:22]
  wire [31:0] n911_O_3_2_1; // @[Top.scala 1064:22]
  wire [31:0] n911_O_3_2_2; // @[Top.scala 1064:22]
  wire [31:0] n911_O_4_0_0; // @[Top.scala 1064:22]
  wire [31:0] n911_O_4_0_1; // @[Top.scala 1064:22]
  wire [31:0] n911_O_4_0_2; // @[Top.scala 1064:22]
  wire [31:0] n911_O_4_1_0; // @[Top.scala 1064:22]
  wire [31:0] n911_O_4_1_1; // @[Top.scala 1064:22]
  wire [31:0] n911_O_4_1_2; // @[Top.scala 1064:22]
  wire [31:0] n911_O_4_2_0; // @[Top.scala 1064:22]
  wire [31:0] n911_O_4_2_1; // @[Top.scala 1064:22]
  wire [31:0] n911_O_4_2_2; // @[Top.scala 1064:22]
  wire [31:0] n911_O_5_0_0; // @[Top.scala 1064:22]
  wire [31:0] n911_O_5_0_1; // @[Top.scala 1064:22]
  wire [31:0] n911_O_5_0_2; // @[Top.scala 1064:22]
  wire [31:0] n911_O_5_1_0; // @[Top.scala 1064:22]
  wire [31:0] n911_O_5_1_1; // @[Top.scala 1064:22]
  wire [31:0] n911_O_5_1_2; // @[Top.scala 1064:22]
  wire [31:0] n911_O_5_2_0; // @[Top.scala 1064:22]
  wire [31:0] n911_O_5_2_1; // @[Top.scala 1064:22]
  wire [31:0] n911_O_5_2_2; // @[Top.scala 1064:22]
  wire [31:0] n911_O_6_0_0; // @[Top.scala 1064:22]
  wire [31:0] n911_O_6_0_1; // @[Top.scala 1064:22]
  wire [31:0] n911_O_6_0_2; // @[Top.scala 1064:22]
  wire [31:0] n911_O_6_1_0; // @[Top.scala 1064:22]
  wire [31:0] n911_O_6_1_1; // @[Top.scala 1064:22]
  wire [31:0] n911_O_6_1_2; // @[Top.scala 1064:22]
  wire [31:0] n911_O_6_2_0; // @[Top.scala 1064:22]
  wire [31:0] n911_O_6_2_1; // @[Top.scala 1064:22]
  wire [31:0] n911_O_6_2_2; // @[Top.scala 1064:22]
  wire [31:0] n911_O_7_0_0; // @[Top.scala 1064:22]
  wire [31:0] n911_O_7_0_1; // @[Top.scala 1064:22]
  wire [31:0] n911_O_7_0_2; // @[Top.scala 1064:22]
  wire [31:0] n911_O_7_1_0; // @[Top.scala 1064:22]
  wire [31:0] n911_O_7_1_1; // @[Top.scala 1064:22]
  wire [31:0] n911_O_7_1_2; // @[Top.scala 1064:22]
  wire [31:0] n911_O_7_2_0; // @[Top.scala 1064:22]
  wire [31:0] n911_O_7_2_1; // @[Top.scala 1064:22]
  wire [31:0] n911_O_7_2_2; // @[Top.scala 1064:22]
  wire  n920_valid_up; // @[Top.scala 1068:22]
  wire  n920_valid_down; // @[Top.scala 1068:22]
  wire [31:0] n920_I_0_0_0; // @[Top.scala 1068:22]
  wire [31:0] n920_I_0_0_1; // @[Top.scala 1068:22]
  wire [31:0] n920_I_0_0_2; // @[Top.scala 1068:22]
  wire [31:0] n920_I_0_1_0; // @[Top.scala 1068:22]
  wire [31:0] n920_I_0_1_1; // @[Top.scala 1068:22]
  wire [31:0] n920_I_0_1_2; // @[Top.scala 1068:22]
  wire [31:0] n920_I_0_2_0; // @[Top.scala 1068:22]
  wire [31:0] n920_I_0_2_1; // @[Top.scala 1068:22]
  wire [31:0] n920_I_0_2_2; // @[Top.scala 1068:22]
  wire [31:0] n920_I_1_0_0; // @[Top.scala 1068:22]
  wire [31:0] n920_I_1_0_1; // @[Top.scala 1068:22]
  wire [31:0] n920_I_1_0_2; // @[Top.scala 1068:22]
  wire [31:0] n920_I_1_1_0; // @[Top.scala 1068:22]
  wire [31:0] n920_I_1_1_1; // @[Top.scala 1068:22]
  wire [31:0] n920_I_1_1_2; // @[Top.scala 1068:22]
  wire [31:0] n920_I_1_2_0; // @[Top.scala 1068:22]
  wire [31:0] n920_I_1_2_1; // @[Top.scala 1068:22]
  wire [31:0] n920_I_1_2_2; // @[Top.scala 1068:22]
  wire [31:0] n920_I_2_0_0; // @[Top.scala 1068:22]
  wire [31:0] n920_I_2_0_1; // @[Top.scala 1068:22]
  wire [31:0] n920_I_2_0_2; // @[Top.scala 1068:22]
  wire [31:0] n920_I_2_1_0; // @[Top.scala 1068:22]
  wire [31:0] n920_I_2_1_1; // @[Top.scala 1068:22]
  wire [31:0] n920_I_2_1_2; // @[Top.scala 1068:22]
  wire [31:0] n920_I_2_2_0; // @[Top.scala 1068:22]
  wire [31:0] n920_I_2_2_1; // @[Top.scala 1068:22]
  wire [31:0] n920_I_2_2_2; // @[Top.scala 1068:22]
  wire [31:0] n920_I_3_0_0; // @[Top.scala 1068:22]
  wire [31:0] n920_I_3_0_1; // @[Top.scala 1068:22]
  wire [31:0] n920_I_3_0_2; // @[Top.scala 1068:22]
  wire [31:0] n920_I_3_1_0; // @[Top.scala 1068:22]
  wire [31:0] n920_I_3_1_1; // @[Top.scala 1068:22]
  wire [31:0] n920_I_3_1_2; // @[Top.scala 1068:22]
  wire [31:0] n920_I_3_2_0; // @[Top.scala 1068:22]
  wire [31:0] n920_I_3_2_1; // @[Top.scala 1068:22]
  wire [31:0] n920_I_3_2_2; // @[Top.scala 1068:22]
  wire [31:0] n920_I_4_0_0; // @[Top.scala 1068:22]
  wire [31:0] n920_I_4_0_1; // @[Top.scala 1068:22]
  wire [31:0] n920_I_4_0_2; // @[Top.scala 1068:22]
  wire [31:0] n920_I_4_1_0; // @[Top.scala 1068:22]
  wire [31:0] n920_I_4_1_1; // @[Top.scala 1068:22]
  wire [31:0] n920_I_4_1_2; // @[Top.scala 1068:22]
  wire [31:0] n920_I_4_2_0; // @[Top.scala 1068:22]
  wire [31:0] n920_I_4_2_1; // @[Top.scala 1068:22]
  wire [31:0] n920_I_4_2_2; // @[Top.scala 1068:22]
  wire [31:0] n920_I_5_0_0; // @[Top.scala 1068:22]
  wire [31:0] n920_I_5_0_1; // @[Top.scala 1068:22]
  wire [31:0] n920_I_5_0_2; // @[Top.scala 1068:22]
  wire [31:0] n920_I_5_1_0; // @[Top.scala 1068:22]
  wire [31:0] n920_I_5_1_1; // @[Top.scala 1068:22]
  wire [31:0] n920_I_5_1_2; // @[Top.scala 1068:22]
  wire [31:0] n920_I_5_2_0; // @[Top.scala 1068:22]
  wire [31:0] n920_I_5_2_1; // @[Top.scala 1068:22]
  wire [31:0] n920_I_5_2_2; // @[Top.scala 1068:22]
  wire [31:0] n920_I_6_0_0; // @[Top.scala 1068:22]
  wire [31:0] n920_I_6_0_1; // @[Top.scala 1068:22]
  wire [31:0] n920_I_6_0_2; // @[Top.scala 1068:22]
  wire [31:0] n920_I_6_1_0; // @[Top.scala 1068:22]
  wire [31:0] n920_I_6_1_1; // @[Top.scala 1068:22]
  wire [31:0] n920_I_6_1_2; // @[Top.scala 1068:22]
  wire [31:0] n920_I_6_2_0; // @[Top.scala 1068:22]
  wire [31:0] n920_I_6_2_1; // @[Top.scala 1068:22]
  wire [31:0] n920_I_6_2_2; // @[Top.scala 1068:22]
  wire [31:0] n920_I_7_0_0; // @[Top.scala 1068:22]
  wire [31:0] n920_I_7_0_1; // @[Top.scala 1068:22]
  wire [31:0] n920_I_7_0_2; // @[Top.scala 1068:22]
  wire [31:0] n920_I_7_1_0; // @[Top.scala 1068:22]
  wire [31:0] n920_I_7_1_1; // @[Top.scala 1068:22]
  wire [31:0] n920_I_7_1_2; // @[Top.scala 1068:22]
  wire [31:0] n920_I_7_2_0; // @[Top.scala 1068:22]
  wire [31:0] n920_I_7_2_1; // @[Top.scala 1068:22]
  wire [31:0] n920_I_7_2_2; // @[Top.scala 1068:22]
  wire [31:0] n920_O_0_0_0_0; // @[Top.scala 1068:22]
  wire [31:0] n920_O_0_0_0_1; // @[Top.scala 1068:22]
  wire [31:0] n920_O_0_0_0_2; // @[Top.scala 1068:22]
  wire [31:0] n920_O_0_0_1_0; // @[Top.scala 1068:22]
  wire [31:0] n920_O_0_0_1_1; // @[Top.scala 1068:22]
  wire [31:0] n920_O_0_0_1_2; // @[Top.scala 1068:22]
  wire [31:0] n920_O_0_0_2_0; // @[Top.scala 1068:22]
  wire [31:0] n920_O_0_0_2_1; // @[Top.scala 1068:22]
  wire [31:0] n920_O_0_0_2_2; // @[Top.scala 1068:22]
  wire [31:0] n920_O_1_0_0_0; // @[Top.scala 1068:22]
  wire [31:0] n920_O_1_0_0_1; // @[Top.scala 1068:22]
  wire [31:0] n920_O_1_0_0_2; // @[Top.scala 1068:22]
  wire [31:0] n920_O_1_0_1_0; // @[Top.scala 1068:22]
  wire [31:0] n920_O_1_0_1_1; // @[Top.scala 1068:22]
  wire [31:0] n920_O_1_0_1_2; // @[Top.scala 1068:22]
  wire [31:0] n920_O_1_0_2_0; // @[Top.scala 1068:22]
  wire [31:0] n920_O_1_0_2_1; // @[Top.scala 1068:22]
  wire [31:0] n920_O_1_0_2_2; // @[Top.scala 1068:22]
  wire [31:0] n920_O_2_0_0_0; // @[Top.scala 1068:22]
  wire [31:0] n920_O_2_0_0_1; // @[Top.scala 1068:22]
  wire [31:0] n920_O_2_0_0_2; // @[Top.scala 1068:22]
  wire [31:0] n920_O_2_0_1_0; // @[Top.scala 1068:22]
  wire [31:0] n920_O_2_0_1_1; // @[Top.scala 1068:22]
  wire [31:0] n920_O_2_0_1_2; // @[Top.scala 1068:22]
  wire [31:0] n920_O_2_0_2_0; // @[Top.scala 1068:22]
  wire [31:0] n920_O_2_0_2_1; // @[Top.scala 1068:22]
  wire [31:0] n920_O_2_0_2_2; // @[Top.scala 1068:22]
  wire [31:0] n920_O_3_0_0_0; // @[Top.scala 1068:22]
  wire [31:0] n920_O_3_0_0_1; // @[Top.scala 1068:22]
  wire [31:0] n920_O_3_0_0_2; // @[Top.scala 1068:22]
  wire [31:0] n920_O_3_0_1_0; // @[Top.scala 1068:22]
  wire [31:0] n920_O_3_0_1_1; // @[Top.scala 1068:22]
  wire [31:0] n920_O_3_0_1_2; // @[Top.scala 1068:22]
  wire [31:0] n920_O_3_0_2_0; // @[Top.scala 1068:22]
  wire [31:0] n920_O_3_0_2_1; // @[Top.scala 1068:22]
  wire [31:0] n920_O_3_0_2_2; // @[Top.scala 1068:22]
  wire [31:0] n920_O_4_0_0_0; // @[Top.scala 1068:22]
  wire [31:0] n920_O_4_0_0_1; // @[Top.scala 1068:22]
  wire [31:0] n920_O_4_0_0_2; // @[Top.scala 1068:22]
  wire [31:0] n920_O_4_0_1_0; // @[Top.scala 1068:22]
  wire [31:0] n920_O_4_0_1_1; // @[Top.scala 1068:22]
  wire [31:0] n920_O_4_0_1_2; // @[Top.scala 1068:22]
  wire [31:0] n920_O_4_0_2_0; // @[Top.scala 1068:22]
  wire [31:0] n920_O_4_0_2_1; // @[Top.scala 1068:22]
  wire [31:0] n920_O_4_0_2_2; // @[Top.scala 1068:22]
  wire [31:0] n920_O_5_0_0_0; // @[Top.scala 1068:22]
  wire [31:0] n920_O_5_0_0_1; // @[Top.scala 1068:22]
  wire [31:0] n920_O_5_0_0_2; // @[Top.scala 1068:22]
  wire [31:0] n920_O_5_0_1_0; // @[Top.scala 1068:22]
  wire [31:0] n920_O_5_0_1_1; // @[Top.scala 1068:22]
  wire [31:0] n920_O_5_0_1_2; // @[Top.scala 1068:22]
  wire [31:0] n920_O_5_0_2_0; // @[Top.scala 1068:22]
  wire [31:0] n920_O_5_0_2_1; // @[Top.scala 1068:22]
  wire [31:0] n920_O_5_0_2_2; // @[Top.scala 1068:22]
  wire [31:0] n920_O_6_0_0_0; // @[Top.scala 1068:22]
  wire [31:0] n920_O_6_0_0_1; // @[Top.scala 1068:22]
  wire [31:0] n920_O_6_0_0_2; // @[Top.scala 1068:22]
  wire [31:0] n920_O_6_0_1_0; // @[Top.scala 1068:22]
  wire [31:0] n920_O_6_0_1_1; // @[Top.scala 1068:22]
  wire [31:0] n920_O_6_0_1_2; // @[Top.scala 1068:22]
  wire [31:0] n920_O_6_0_2_0; // @[Top.scala 1068:22]
  wire [31:0] n920_O_6_0_2_1; // @[Top.scala 1068:22]
  wire [31:0] n920_O_6_0_2_2; // @[Top.scala 1068:22]
  wire [31:0] n920_O_7_0_0_0; // @[Top.scala 1068:22]
  wire [31:0] n920_O_7_0_0_1; // @[Top.scala 1068:22]
  wire [31:0] n920_O_7_0_0_2; // @[Top.scala 1068:22]
  wire [31:0] n920_O_7_0_1_0; // @[Top.scala 1068:22]
  wire [31:0] n920_O_7_0_1_1; // @[Top.scala 1068:22]
  wire [31:0] n920_O_7_0_1_2; // @[Top.scala 1068:22]
  wire [31:0] n920_O_7_0_2_0; // @[Top.scala 1068:22]
  wire [31:0] n920_O_7_0_2_1; // @[Top.scala 1068:22]
  wire [31:0] n920_O_7_0_2_2; // @[Top.scala 1068:22]
  wire  n927_valid_up; // @[Top.scala 1071:22]
  wire  n927_valid_down; // @[Top.scala 1071:22]
  wire [31:0] n927_I_0_0_0_0; // @[Top.scala 1071:22]
  wire [31:0] n927_I_0_0_0_1; // @[Top.scala 1071:22]
  wire [31:0] n927_I_0_0_0_2; // @[Top.scala 1071:22]
  wire [31:0] n927_I_0_0_1_0; // @[Top.scala 1071:22]
  wire [31:0] n927_I_0_0_1_1; // @[Top.scala 1071:22]
  wire [31:0] n927_I_0_0_1_2; // @[Top.scala 1071:22]
  wire [31:0] n927_I_0_0_2_0; // @[Top.scala 1071:22]
  wire [31:0] n927_I_0_0_2_1; // @[Top.scala 1071:22]
  wire [31:0] n927_I_0_0_2_2; // @[Top.scala 1071:22]
  wire [31:0] n927_I_1_0_0_0; // @[Top.scala 1071:22]
  wire [31:0] n927_I_1_0_0_1; // @[Top.scala 1071:22]
  wire [31:0] n927_I_1_0_0_2; // @[Top.scala 1071:22]
  wire [31:0] n927_I_1_0_1_0; // @[Top.scala 1071:22]
  wire [31:0] n927_I_1_0_1_1; // @[Top.scala 1071:22]
  wire [31:0] n927_I_1_0_1_2; // @[Top.scala 1071:22]
  wire [31:0] n927_I_1_0_2_0; // @[Top.scala 1071:22]
  wire [31:0] n927_I_1_0_2_1; // @[Top.scala 1071:22]
  wire [31:0] n927_I_1_0_2_2; // @[Top.scala 1071:22]
  wire [31:0] n927_I_2_0_0_0; // @[Top.scala 1071:22]
  wire [31:0] n927_I_2_0_0_1; // @[Top.scala 1071:22]
  wire [31:0] n927_I_2_0_0_2; // @[Top.scala 1071:22]
  wire [31:0] n927_I_2_0_1_0; // @[Top.scala 1071:22]
  wire [31:0] n927_I_2_0_1_1; // @[Top.scala 1071:22]
  wire [31:0] n927_I_2_0_1_2; // @[Top.scala 1071:22]
  wire [31:0] n927_I_2_0_2_0; // @[Top.scala 1071:22]
  wire [31:0] n927_I_2_0_2_1; // @[Top.scala 1071:22]
  wire [31:0] n927_I_2_0_2_2; // @[Top.scala 1071:22]
  wire [31:0] n927_I_3_0_0_0; // @[Top.scala 1071:22]
  wire [31:0] n927_I_3_0_0_1; // @[Top.scala 1071:22]
  wire [31:0] n927_I_3_0_0_2; // @[Top.scala 1071:22]
  wire [31:0] n927_I_3_0_1_0; // @[Top.scala 1071:22]
  wire [31:0] n927_I_3_0_1_1; // @[Top.scala 1071:22]
  wire [31:0] n927_I_3_0_1_2; // @[Top.scala 1071:22]
  wire [31:0] n927_I_3_0_2_0; // @[Top.scala 1071:22]
  wire [31:0] n927_I_3_0_2_1; // @[Top.scala 1071:22]
  wire [31:0] n927_I_3_0_2_2; // @[Top.scala 1071:22]
  wire [31:0] n927_I_4_0_0_0; // @[Top.scala 1071:22]
  wire [31:0] n927_I_4_0_0_1; // @[Top.scala 1071:22]
  wire [31:0] n927_I_4_0_0_2; // @[Top.scala 1071:22]
  wire [31:0] n927_I_4_0_1_0; // @[Top.scala 1071:22]
  wire [31:0] n927_I_4_0_1_1; // @[Top.scala 1071:22]
  wire [31:0] n927_I_4_0_1_2; // @[Top.scala 1071:22]
  wire [31:0] n927_I_4_0_2_0; // @[Top.scala 1071:22]
  wire [31:0] n927_I_4_0_2_1; // @[Top.scala 1071:22]
  wire [31:0] n927_I_4_0_2_2; // @[Top.scala 1071:22]
  wire [31:0] n927_I_5_0_0_0; // @[Top.scala 1071:22]
  wire [31:0] n927_I_5_0_0_1; // @[Top.scala 1071:22]
  wire [31:0] n927_I_5_0_0_2; // @[Top.scala 1071:22]
  wire [31:0] n927_I_5_0_1_0; // @[Top.scala 1071:22]
  wire [31:0] n927_I_5_0_1_1; // @[Top.scala 1071:22]
  wire [31:0] n927_I_5_0_1_2; // @[Top.scala 1071:22]
  wire [31:0] n927_I_5_0_2_0; // @[Top.scala 1071:22]
  wire [31:0] n927_I_5_0_2_1; // @[Top.scala 1071:22]
  wire [31:0] n927_I_5_0_2_2; // @[Top.scala 1071:22]
  wire [31:0] n927_I_6_0_0_0; // @[Top.scala 1071:22]
  wire [31:0] n927_I_6_0_0_1; // @[Top.scala 1071:22]
  wire [31:0] n927_I_6_0_0_2; // @[Top.scala 1071:22]
  wire [31:0] n927_I_6_0_1_0; // @[Top.scala 1071:22]
  wire [31:0] n927_I_6_0_1_1; // @[Top.scala 1071:22]
  wire [31:0] n927_I_6_0_1_2; // @[Top.scala 1071:22]
  wire [31:0] n927_I_6_0_2_0; // @[Top.scala 1071:22]
  wire [31:0] n927_I_6_0_2_1; // @[Top.scala 1071:22]
  wire [31:0] n927_I_6_0_2_2; // @[Top.scala 1071:22]
  wire [31:0] n927_I_7_0_0_0; // @[Top.scala 1071:22]
  wire [31:0] n927_I_7_0_0_1; // @[Top.scala 1071:22]
  wire [31:0] n927_I_7_0_0_2; // @[Top.scala 1071:22]
  wire [31:0] n927_I_7_0_1_0; // @[Top.scala 1071:22]
  wire [31:0] n927_I_7_0_1_1; // @[Top.scala 1071:22]
  wire [31:0] n927_I_7_0_1_2; // @[Top.scala 1071:22]
  wire [31:0] n927_I_7_0_2_0; // @[Top.scala 1071:22]
  wire [31:0] n927_I_7_0_2_1; // @[Top.scala 1071:22]
  wire [31:0] n927_I_7_0_2_2; // @[Top.scala 1071:22]
  wire [31:0] n927_O_0_0_0; // @[Top.scala 1071:22]
  wire [31:0] n927_O_0_0_1; // @[Top.scala 1071:22]
  wire [31:0] n927_O_0_0_2; // @[Top.scala 1071:22]
  wire [31:0] n927_O_0_1_0; // @[Top.scala 1071:22]
  wire [31:0] n927_O_0_1_1; // @[Top.scala 1071:22]
  wire [31:0] n927_O_0_1_2; // @[Top.scala 1071:22]
  wire [31:0] n927_O_0_2_0; // @[Top.scala 1071:22]
  wire [31:0] n927_O_0_2_1; // @[Top.scala 1071:22]
  wire [31:0] n927_O_0_2_2; // @[Top.scala 1071:22]
  wire [31:0] n927_O_1_0_0; // @[Top.scala 1071:22]
  wire [31:0] n927_O_1_0_1; // @[Top.scala 1071:22]
  wire [31:0] n927_O_1_0_2; // @[Top.scala 1071:22]
  wire [31:0] n927_O_1_1_0; // @[Top.scala 1071:22]
  wire [31:0] n927_O_1_1_1; // @[Top.scala 1071:22]
  wire [31:0] n927_O_1_1_2; // @[Top.scala 1071:22]
  wire [31:0] n927_O_1_2_0; // @[Top.scala 1071:22]
  wire [31:0] n927_O_1_2_1; // @[Top.scala 1071:22]
  wire [31:0] n927_O_1_2_2; // @[Top.scala 1071:22]
  wire [31:0] n927_O_2_0_0; // @[Top.scala 1071:22]
  wire [31:0] n927_O_2_0_1; // @[Top.scala 1071:22]
  wire [31:0] n927_O_2_0_2; // @[Top.scala 1071:22]
  wire [31:0] n927_O_2_1_0; // @[Top.scala 1071:22]
  wire [31:0] n927_O_2_1_1; // @[Top.scala 1071:22]
  wire [31:0] n927_O_2_1_2; // @[Top.scala 1071:22]
  wire [31:0] n927_O_2_2_0; // @[Top.scala 1071:22]
  wire [31:0] n927_O_2_2_1; // @[Top.scala 1071:22]
  wire [31:0] n927_O_2_2_2; // @[Top.scala 1071:22]
  wire [31:0] n927_O_3_0_0; // @[Top.scala 1071:22]
  wire [31:0] n927_O_3_0_1; // @[Top.scala 1071:22]
  wire [31:0] n927_O_3_0_2; // @[Top.scala 1071:22]
  wire [31:0] n927_O_3_1_0; // @[Top.scala 1071:22]
  wire [31:0] n927_O_3_1_1; // @[Top.scala 1071:22]
  wire [31:0] n927_O_3_1_2; // @[Top.scala 1071:22]
  wire [31:0] n927_O_3_2_0; // @[Top.scala 1071:22]
  wire [31:0] n927_O_3_2_1; // @[Top.scala 1071:22]
  wire [31:0] n927_O_3_2_2; // @[Top.scala 1071:22]
  wire [31:0] n927_O_4_0_0; // @[Top.scala 1071:22]
  wire [31:0] n927_O_4_0_1; // @[Top.scala 1071:22]
  wire [31:0] n927_O_4_0_2; // @[Top.scala 1071:22]
  wire [31:0] n927_O_4_1_0; // @[Top.scala 1071:22]
  wire [31:0] n927_O_4_1_1; // @[Top.scala 1071:22]
  wire [31:0] n927_O_4_1_2; // @[Top.scala 1071:22]
  wire [31:0] n927_O_4_2_0; // @[Top.scala 1071:22]
  wire [31:0] n927_O_4_2_1; // @[Top.scala 1071:22]
  wire [31:0] n927_O_4_2_2; // @[Top.scala 1071:22]
  wire [31:0] n927_O_5_0_0; // @[Top.scala 1071:22]
  wire [31:0] n927_O_5_0_1; // @[Top.scala 1071:22]
  wire [31:0] n927_O_5_0_2; // @[Top.scala 1071:22]
  wire [31:0] n927_O_5_1_0; // @[Top.scala 1071:22]
  wire [31:0] n927_O_5_1_1; // @[Top.scala 1071:22]
  wire [31:0] n927_O_5_1_2; // @[Top.scala 1071:22]
  wire [31:0] n927_O_5_2_0; // @[Top.scala 1071:22]
  wire [31:0] n927_O_5_2_1; // @[Top.scala 1071:22]
  wire [31:0] n927_O_5_2_2; // @[Top.scala 1071:22]
  wire [31:0] n927_O_6_0_0; // @[Top.scala 1071:22]
  wire [31:0] n927_O_6_0_1; // @[Top.scala 1071:22]
  wire [31:0] n927_O_6_0_2; // @[Top.scala 1071:22]
  wire [31:0] n927_O_6_1_0; // @[Top.scala 1071:22]
  wire [31:0] n927_O_6_1_1; // @[Top.scala 1071:22]
  wire [31:0] n927_O_6_1_2; // @[Top.scala 1071:22]
  wire [31:0] n927_O_6_2_0; // @[Top.scala 1071:22]
  wire [31:0] n927_O_6_2_1; // @[Top.scala 1071:22]
  wire [31:0] n927_O_6_2_2; // @[Top.scala 1071:22]
  wire [31:0] n927_O_7_0_0; // @[Top.scala 1071:22]
  wire [31:0] n927_O_7_0_1; // @[Top.scala 1071:22]
  wire [31:0] n927_O_7_0_2; // @[Top.scala 1071:22]
  wire [31:0] n927_O_7_1_0; // @[Top.scala 1071:22]
  wire [31:0] n927_O_7_1_1; // @[Top.scala 1071:22]
  wire [31:0] n927_O_7_1_2; // @[Top.scala 1071:22]
  wire [31:0] n927_O_7_2_0; // @[Top.scala 1071:22]
  wire [31:0] n927_O_7_2_1; // @[Top.scala 1071:22]
  wire [31:0] n927_O_7_2_2; // @[Top.scala 1071:22]
  wire  n969_clock; // @[Top.scala 1074:22]
  wire  n969_reset; // @[Top.scala 1074:22]
  wire  n969_valid_up; // @[Top.scala 1074:22]
  wire  n969_valid_down; // @[Top.scala 1074:22]
  wire [31:0] n969_I_0_0_0; // @[Top.scala 1074:22]
  wire [31:0] n969_I_0_0_1; // @[Top.scala 1074:22]
  wire [31:0] n969_I_0_0_2; // @[Top.scala 1074:22]
  wire [31:0] n969_I_0_1_0; // @[Top.scala 1074:22]
  wire [31:0] n969_I_0_1_1; // @[Top.scala 1074:22]
  wire [31:0] n969_I_0_1_2; // @[Top.scala 1074:22]
  wire [31:0] n969_I_0_2_0; // @[Top.scala 1074:22]
  wire [31:0] n969_I_0_2_1; // @[Top.scala 1074:22]
  wire [31:0] n969_I_0_2_2; // @[Top.scala 1074:22]
  wire [31:0] n969_I_1_0_0; // @[Top.scala 1074:22]
  wire [31:0] n969_I_1_0_1; // @[Top.scala 1074:22]
  wire [31:0] n969_I_1_0_2; // @[Top.scala 1074:22]
  wire [31:0] n969_I_1_1_0; // @[Top.scala 1074:22]
  wire [31:0] n969_I_1_1_1; // @[Top.scala 1074:22]
  wire [31:0] n969_I_1_1_2; // @[Top.scala 1074:22]
  wire [31:0] n969_I_1_2_0; // @[Top.scala 1074:22]
  wire [31:0] n969_I_1_2_1; // @[Top.scala 1074:22]
  wire [31:0] n969_I_1_2_2; // @[Top.scala 1074:22]
  wire [31:0] n969_I_2_0_0; // @[Top.scala 1074:22]
  wire [31:0] n969_I_2_0_1; // @[Top.scala 1074:22]
  wire [31:0] n969_I_2_0_2; // @[Top.scala 1074:22]
  wire [31:0] n969_I_2_1_0; // @[Top.scala 1074:22]
  wire [31:0] n969_I_2_1_1; // @[Top.scala 1074:22]
  wire [31:0] n969_I_2_1_2; // @[Top.scala 1074:22]
  wire [31:0] n969_I_2_2_0; // @[Top.scala 1074:22]
  wire [31:0] n969_I_2_2_1; // @[Top.scala 1074:22]
  wire [31:0] n969_I_2_2_2; // @[Top.scala 1074:22]
  wire [31:0] n969_I_3_0_0; // @[Top.scala 1074:22]
  wire [31:0] n969_I_3_0_1; // @[Top.scala 1074:22]
  wire [31:0] n969_I_3_0_2; // @[Top.scala 1074:22]
  wire [31:0] n969_I_3_1_0; // @[Top.scala 1074:22]
  wire [31:0] n969_I_3_1_1; // @[Top.scala 1074:22]
  wire [31:0] n969_I_3_1_2; // @[Top.scala 1074:22]
  wire [31:0] n969_I_3_2_0; // @[Top.scala 1074:22]
  wire [31:0] n969_I_3_2_1; // @[Top.scala 1074:22]
  wire [31:0] n969_I_3_2_2; // @[Top.scala 1074:22]
  wire [31:0] n969_I_4_0_0; // @[Top.scala 1074:22]
  wire [31:0] n969_I_4_0_1; // @[Top.scala 1074:22]
  wire [31:0] n969_I_4_0_2; // @[Top.scala 1074:22]
  wire [31:0] n969_I_4_1_0; // @[Top.scala 1074:22]
  wire [31:0] n969_I_4_1_1; // @[Top.scala 1074:22]
  wire [31:0] n969_I_4_1_2; // @[Top.scala 1074:22]
  wire [31:0] n969_I_4_2_0; // @[Top.scala 1074:22]
  wire [31:0] n969_I_4_2_1; // @[Top.scala 1074:22]
  wire [31:0] n969_I_4_2_2; // @[Top.scala 1074:22]
  wire [31:0] n969_I_5_0_0; // @[Top.scala 1074:22]
  wire [31:0] n969_I_5_0_1; // @[Top.scala 1074:22]
  wire [31:0] n969_I_5_0_2; // @[Top.scala 1074:22]
  wire [31:0] n969_I_5_1_0; // @[Top.scala 1074:22]
  wire [31:0] n969_I_5_1_1; // @[Top.scala 1074:22]
  wire [31:0] n969_I_5_1_2; // @[Top.scala 1074:22]
  wire [31:0] n969_I_5_2_0; // @[Top.scala 1074:22]
  wire [31:0] n969_I_5_2_1; // @[Top.scala 1074:22]
  wire [31:0] n969_I_5_2_2; // @[Top.scala 1074:22]
  wire [31:0] n969_I_6_0_0; // @[Top.scala 1074:22]
  wire [31:0] n969_I_6_0_1; // @[Top.scala 1074:22]
  wire [31:0] n969_I_6_0_2; // @[Top.scala 1074:22]
  wire [31:0] n969_I_6_1_0; // @[Top.scala 1074:22]
  wire [31:0] n969_I_6_1_1; // @[Top.scala 1074:22]
  wire [31:0] n969_I_6_1_2; // @[Top.scala 1074:22]
  wire [31:0] n969_I_6_2_0; // @[Top.scala 1074:22]
  wire [31:0] n969_I_6_2_1; // @[Top.scala 1074:22]
  wire [31:0] n969_I_6_2_2; // @[Top.scala 1074:22]
  wire [31:0] n969_I_7_0_0; // @[Top.scala 1074:22]
  wire [31:0] n969_I_7_0_1; // @[Top.scala 1074:22]
  wire [31:0] n969_I_7_0_2; // @[Top.scala 1074:22]
  wire [31:0] n969_I_7_1_0; // @[Top.scala 1074:22]
  wire [31:0] n969_I_7_1_1; // @[Top.scala 1074:22]
  wire [31:0] n969_I_7_1_2; // @[Top.scala 1074:22]
  wire [31:0] n969_I_7_2_0; // @[Top.scala 1074:22]
  wire [31:0] n969_I_7_2_1; // @[Top.scala 1074:22]
  wire [31:0] n969_I_7_2_2; // @[Top.scala 1074:22]
  wire [31:0] n969_O_0_0_0; // @[Top.scala 1074:22]
  wire [31:0] n969_O_1_0_0; // @[Top.scala 1074:22]
  wire [31:0] n969_O_2_0_0; // @[Top.scala 1074:22]
  wire [31:0] n969_O_3_0_0; // @[Top.scala 1074:22]
  wire [31:0] n969_O_4_0_0; // @[Top.scala 1074:22]
  wire [31:0] n969_O_5_0_0; // @[Top.scala 1074:22]
  wire [31:0] n969_O_6_0_0; // @[Top.scala 1074:22]
  wire [31:0] n969_O_7_0_0; // @[Top.scala 1074:22]
  wire  n970_valid_up; // @[Top.scala 1077:22]
  wire  n970_valid_down; // @[Top.scala 1077:22]
  wire [31:0] n970_I_0_0_0; // @[Top.scala 1077:22]
  wire [31:0] n970_I_1_0_0; // @[Top.scala 1077:22]
  wire [31:0] n970_I_2_0_0; // @[Top.scala 1077:22]
  wire [31:0] n970_I_3_0_0; // @[Top.scala 1077:22]
  wire [31:0] n970_I_4_0_0; // @[Top.scala 1077:22]
  wire [31:0] n970_I_5_0_0; // @[Top.scala 1077:22]
  wire [31:0] n970_I_6_0_0; // @[Top.scala 1077:22]
  wire [31:0] n970_I_7_0_0; // @[Top.scala 1077:22]
  wire [31:0] n970_O_0_0; // @[Top.scala 1077:22]
  wire [31:0] n970_O_1_0; // @[Top.scala 1077:22]
  wire [31:0] n970_O_2_0; // @[Top.scala 1077:22]
  wire [31:0] n970_O_3_0; // @[Top.scala 1077:22]
  wire [31:0] n970_O_4_0; // @[Top.scala 1077:22]
  wire [31:0] n970_O_5_0; // @[Top.scala 1077:22]
  wire [31:0] n970_O_6_0; // @[Top.scala 1077:22]
  wire [31:0] n970_O_7_0; // @[Top.scala 1077:22]
  wire  n971_valid_up; // @[Top.scala 1080:22]
  wire  n971_valid_down; // @[Top.scala 1080:22]
  wire [31:0] n971_I_0_0; // @[Top.scala 1080:22]
  wire [31:0] n971_I_1_0; // @[Top.scala 1080:22]
  wire [31:0] n971_I_2_0; // @[Top.scala 1080:22]
  wire [31:0] n971_I_3_0; // @[Top.scala 1080:22]
  wire [31:0] n971_I_4_0; // @[Top.scala 1080:22]
  wire [31:0] n971_I_5_0; // @[Top.scala 1080:22]
  wire [31:0] n971_I_6_0; // @[Top.scala 1080:22]
  wire [31:0] n971_I_7_0; // @[Top.scala 1080:22]
  wire [31:0] n971_O_0; // @[Top.scala 1080:22]
  wire [31:0] n971_O_1; // @[Top.scala 1080:22]
  wire [31:0] n971_O_2; // @[Top.scala 1080:22]
  wire [31:0] n971_O_3; // @[Top.scala 1080:22]
  wire [31:0] n971_O_4; // @[Top.scala 1080:22]
  wire [31:0] n971_O_5; // @[Top.scala 1080:22]
  wire [31:0] n971_O_6; // @[Top.scala 1080:22]
  wire [31:0] n971_O_7; // @[Top.scala 1080:22]
  wire  n972_clock; // @[Top.scala 1083:22]
  wire  n972_reset; // @[Top.scala 1083:22]
  wire  n972_valid_up; // @[Top.scala 1083:22]
  wire  n972_valid_down; // @[Top.scala 1083:22]
  wire [31:0] n972_I_0; // @[Top.scala 1083:22]
  wire [31:0] n972_I_1; // @[Top.scala 1083:22]
  wire [31:0] n972_I_2; // @[Top.scala 1083:22]
  wire [31:0] n972_I_3; // @[Top.scala 1083:22]
  wire [31:0] n972_I_4; // @[Top.scala 1083:22]
  wire [31:0] n972_I_5; // @[Top.scala 1083:22]
  wire [31:0] n972_I_6; // @[Top.scala 1083:22]
  wire [31:0] n972_I_7; // @[Top.scala 1083:22]
  wire [31:0] n972_O_0; // @[Top.scala 1083:22]
  wire [31:0] n972_O_1; // @[Top.scala 1083:22]
  wire [31:0] n972_O_2; // @[Top.scala 1083:22]
  wire [31:0] n972_O_3; // @[Top.scala 1083:22]
  wire [31:0] n972_O_4; // @[Top.scala 1083:22]
  wire [31:0] n972_O_5; // @[Top.scala 1083:22]
  wire [31:0] n972_O_6; // @[Top.scala 1083:22]
  wire [31:0] n972_O_7; // @[Top.scala 1083:22]
  wire  n973_clock; // @[Top.scala 1086:22]
  wire  n973_reset; // @[Top.scala 1086:22]
  wire  n973_valid_up; // @[Top.scala 1086:22]
  wire  n973_valid_down; // @[Top.scala 1086:22]
  wire [31:0] n973_I0_0; // @[Top.scala 1086:22]
  wire [31:0] n973_I0_1; // @[Top.scala 1086:22]
  wire [31:0] n973_I0_2; // @[Top.scala 1086:22]
  wire [31:0] n973_I0_3; // @[Top.scala 1086:22]
  wire [31:0] n973_I0_4; // @[Top.scala 1086:22]
  wire [31:0] n973_I0_5; // @[Top.scala 1086:22]
  wire [31:0] n973_I0_6; // @[Top.scala 1086:22]
  wire [31:0] n973_I0_7; // @[Top.scala 1086:22]
  wire [31:0] n973_I1_0; // @[Top.scala 1086:22]
  wire [31:0] n973_I1_1; // @[Top.scala 1086:22]
  wire [31:0] n973_I1_2; // @[Top.scala 1086:22]
  wire [31:0] n973_I1_3; // @[Top.scala 1086:22]
  wire [31:0] n973_I1_4; // @[Top.scala 1086:22]
  wire [31:0] n973_I1_5; // @[Top.scala 1086:22]
  wire [31:0] n973_I1_6; // @[Top.scala 1086:22]
  wire [31:0] n973_I1_7; // @[Top.scala 1086:22]
  wire [31:0] n973_O_0; // @[Top.scala 1086:22]
  wire [31:0] n973_O_1; // @[Top.scala 1086:22]
  wire [31:0] n973_O_2; // @[Top.scala 1086:22]
  wire [31:0] n973_O_3; // @[Top.scala 1086:22]
  wire [31:0] n973_O_4; // @[Top.scala 1086:22]
  wire [31:0] n973_O_5; // @[Top.scala 1086:22]
  wire [31:0] n973_O_6; // @[Top.scala 1086:22]
  wire [31:0] n973_O_7; // @[Top.scala 1086:22]
  wire  n1004_valid_up; // @[Top.scala 1090:23]
  wire  n1004_valid_down; // @[Top.scala 1090:23]
  wire [31:0] n1004_I0_0; // @[Top.scala 1090:23]
  wire [31:0] n1004_I0_1; // @[Top.scala 1090:23]
  wire [31:0] n1004_I0_2; // @[Top.scala 1090:23]
  wire [31:0] n1004_I0_3; // @[Top.scala 1090:23]
  wire [31:0] n1004_I0_4; // @[Top.scala 1090:23]
  wire [31:0] n1004_I0_5; // @[Top.scala 1090:23]
  wire [31:0] n1004_I0_6; // @[Top.scala 1090:23]
  wire [31:0] n1004_I0_7; // @[Top.scala 1090:23]
  wire [31:0] n1004_I1_0; // @[Top.scala 1090:23]
  wire [31:0] n1004_I1_1; // @[Top.scala 1090:23]
  wire [31:0] n1004_I1_2; // @[Top.scala 1090:23]
  wire [31:0] n1004_I1_3; // @[Top.scala 1090:23]
  wire [31:0] n1004_I1_4; // @[Top.scala 1090:23]
  wire [31:0] n1004_I1_5; // @[Top.scala 1090:23]
  wire [31:0] n1004_I1_6; // @[Top.scala 1090:23]
  wire [31:0] n1004_I1_7; // @[Top.scala 1090:23]
  wire [31:0] n1004_O_0_t0b; // @[Top.scala 1090:23]
  wire [31:0] n1004_O_0_t1b; // @[Top.scala 1090:23]
  wire [31:0] n1004_O_1_t0b; // @[Top.scala 1090:23]
  wire [31:0] n1004_O_1_t1b; // @[Top.scala 1090:23]
  wire [31:0] n1004_O_2_t0b; // @[Top.scala 1090:23]
  wire [31:0] n1004_O_2_t1b; // @[Top.scala 1090:23]
  wire [31:0] n1004_O_3_t0b; // @[Top.scala 1090:23]
  wire [31:0] n1004_O_3_t1b; // @[Top.scala 1090:23]
  wire [31:0] n1004_O_4_t0b; // @[Top.scala 1090:23]
  wire [31:0] n1004_O_4_t1b; // @[Top.scala 1090:23]
  wire [31:0] n1004_O_5_t0b; // @[Top.scala 1090:23]
  wire [31:0] n1004_O_5_t1b; // @[Top.scala 1090:23]
  wire [31:0] n1004_O_6_t0b; // @[Top.scala 1090:23]
  wire [31:0] n1004_O_6_t1b; // @[Top.scala 1090:23]
  wire [31:0] n1004_O_7_t0b; // @[Top.scala 1090:23]
  wire [31:0] n1004_O_7_t1b; // @[Top.scala 1090:23]
  wire  n1011_valid_up; // @[Top.scala 1094:23]
  wire  n1011_valid_down; // @[Top.scala 1094:23]
  wire [31:0] n1011_I0_0; // @[Top.scala 1094:23]
  wire [31:0] n1011_I0_1; // @[Top.scala 1094:23]
  wire [31:0] n1011_I0_2; // @[Top.scala 1094:23]
  wire [31:0] n1011_I0_3; // @[Top.scala 1094:23]
  wire [31:0] n1011_I0_4; // @[Top.scala 1094:23]
  wire [31:0] n1011_I0_5; // @[Top.scala 1094:23]
  wire [31:0] n1011_I0_6; // @[Top.scala 1094:23]
  wire [31:0] n1011_I0_7; // @[Top.scala 1094:23]
  wire [31:0] n1011_I1_0_t0b; // @[Top.scala 1094:23]
  wire [31:0] n1011_I1_0_t1b; // @[Top.scala 1094:23]
  wire [31:0] n1011_I1_1_t0b; // @[Top.scala 1094:23]
  wire [31:0] n1011_I1_1_t1b; // @[Top.scala 1094:23]
  wire [31:0] n1011_I1_2_t0b; // @[Top.scala 1094:23]
  wire [31:0] n1011_I1_2_t1b; // @[Top.scala 1094:23]
  wire [31:0] n1011_I1_3_t0b; // @[Top.scala 1094:23]
  wire [31:0] n1011_I1_3_t1b; // @[Top.scala 1094:23]
  wire [31:0] n1011_I1_4_t0b; // @[Top.scala 1094:23]
  wire [31:0] n1011_I1_4_t1b; // @[Top.scala 1094:23]
  wire [31:0] n1011_I1_5_t0b; // @[Top.scala 1094:23]
  wire [31:0] n1011_I1_5_t1b; // @[Top.scala 1094:23]
  wire [31:0] n1011_I1_6_t0b; // @[Top.scala 1094:23]
  wire [31:0] n1011_I1_6_t1b; // @[Top.scala 1094:23]
  wire [31:0] n1011_I1_7_t0b; // @[Top.scala 1094:23]
  wire [31:0] n1011_I1_7_t1b; // @[Top.scala 1094:23]
  wire [31:0] n1011_O_0_t0b; // @[Top.scala 1094:23]
  wire [31:0] n1011_O_0_t1b_t0b; // @[Top.scala 1094:23]
  wire [31:0] n1011_O_0_t1b_t1b; // @[Top.scala 1094:23]
  wire [31:0] n1011_O_1_t0b; // @[Top.scala 1094:23]
  wire [31:0] n1011_O_1_t1b_t0b; // @[Top.scala 1094:23]
  wire [31:0] n1011_O_1_t1b_t1b; // @[Top.scala 1094:23]
  wire [31:0] n1011_O_2_t0b; // @[Top.scala 1094:23]
  wire [31:0] n1011_O_2_t1b_t0b; // @[Top.scala 1094:23]
  wire [31:0] n1011_O_2_t1b_t1b; // @[Top.scala 1094:23]
  wire [31:0] n1011_O_3_t0b; // @[Top.scala 1094:23]
  wire [31:0] n1011_O_3_t1b_t0b; // @[Top.scala 1094:23]
  wire [31:0] n1011_O_3_t1b_t1b; // @[Top.scala 1094:23]
  wire [31:0] n1011_O_4_t0b; // @[Top.scala 1094:23]
  wire [31:0] n1011_O_4_t1b_t0b; // @[Top.scala 1094:23]
  wire [31:0] n1011_O_4_t1b_t1b; // @[Top.scala 1094:23]
  wire [31:0] n1011_O_5_t0b; // @[Top.scala 1094:23]
  wire [31:0] n1011_O_5_t1b_t0b; // @[Top.scala 1094:23]
  wire [31:0] n1011_O_5_t1b_t1b; // @[Top.scala 1094:23]
  wire [31:0] n1011_O_6_t0b; // @[Top.scala 1094:23]
  wire [31:0] n1011_O_6_t1b_t0b; // @[Top.scala 1094:23]
  wire [31:0] n1011_O_6_t1b_t1b; // @[Top.scala 1094:23]
  wire [31:0] n1011_O_7_t0b; // @[Top.scala 1094:23]
  wire [31:0] n1011_O_7_t1b_t0b; // @[Top.scala 1094:23]
  wire [31:0] n1011_O_7_t1b_t1b; // @[Top.scala 1094:23]
  wire  n1018_clock; // @[Top.scala 1098:23]
  wire  n1018_reset; // @[Top.scala 1098:23]
  wire  n1018_valid_up; // @[Top.scala 1098:23]
  wire  n1018_valid_down; // @[Top.scala 1098:23]
  wire [31:0] n1018_I_0_t0b; // @[Top.scala 1098:23]
  wire [31:0] n1018_I_0_t1b_t0b; // @[Top.scala 1098:23]
  wire [31:0] n1018_I_0_t1b_t1b; // @[Top.scala 1098:23]
  wire [31:0] n1018_I_1_t0b; // @[Top.scala 1098:23]
  wire [31:0] n1018_I_1_t1b_t0b; // @[Top.scala 1098:23]
  wire [31:0] n1018_I_1_t1b_t1b; // @[Top.scala 1098:23]
  wire [31:0] n1018_I_2_t0b; // @[Top.scala 1098:23]
  wire [31:0] n1018_I_2_t1b_t0b; // @[Top.scala 1098:23]
  wire [31:0] n1018_I_2_t1b_t1b; // @[Top.scala 1098:23]
  wire [31:0] n1018_I_3_t0b; // @[Top.scala 1098:23]
  wire [31:0] n1018_I_3_t1b_t0b; // @[Top.scala 1098:23]
  wire [31:0] n1018_I_3_t1b_t1b; // @[Top.scala 1098:23]
  wire [31:0] n1018_I_4_t0b; // @[Top.scala 1098:23]
  wire [31:0] n1018_I_4_t1b_t0b; // @[Top.scala 1098:23]
  wire [31:0] n1018_I_4_t1b_t1b; // @[Top.scala 1098:23]
  wire [31:0] n1018_I_5_t0b; // @[Top.scala 1098:23]
  wire [31:0] n1018_I_5_t1b_t0b; // @[Top.scala 1098:23]
  wire [31:0] n1018_I_5_t1b_t1b; // @[Top.scala 1098:23]
  wire [31:0] n1018_I_6_t0b; // @[Top.scala 1098:23]
  wire [31:0] n1018_I_6_t1b_t0b; // @[Top.scala 1098:23]
  wire [31:0] n1018_I_6_t1b_t1b; // @[Top.scala 1098:23]
  wire [31:0] n1018_I_7_t0b; // @[Top.scala 1098:23]
  wire [31:0] n1018_I_7_t1b_t0b; // @[Top.scala 1098:23]
  wire [31:0] n1018_I_7_t1b_t1b; // @[Top.scala 1098:23]
  wire [31:0] n1018_O_0_t0b; // @[Top.scala 1098:23]
  wire [31:0] n1018_O_0_t1b_t0b; // @[Top.scala 1098:23]
  wire [31:0] n1018_O_0_t1b_t1b; // @[Top.scala 1098:23]
  wire [31:0] n1018_O_1_t0b; // @[Top.scala 1098:23]
  wire [31:0] n1018_O_1_t1b_t0b; // @[Top.scala 1098:23]
  wire [31:0] n1018_O_1_t1b_t1b; // @[Top.scala 1098:23]
  wire [31:0] n1018_O_2_t0b; // @[Top.scala 1098:23]
  wire [31:0] n1018_O_2_t1b_t0b; // @[Top.scala 1098:23]
  wire [31:0] n1018_O_2_t1b_t1b; // @[Top.scala 1098:23]
  wire [31:0] n1018_O_3_t0b; // @[Top.scala 1098:23]
  wire [31:0] n1018_O_3_t1b_t0b; // @[Top.scala 1098:23]
  wire [31:0] n1018_O_3_t1b_t1b; // @[Top.scala 1098:23]
  wire [31:0] n1018_O_4_t0b; // @[Top.scala 1098:23]
  wire [31:0] n1018_O_4_t1b_t0b; // @[Top.scala 1098:23]
  wire [31:0] n1018_O_4_t1b_t1b; // @[Top.scala 1098:23]
  wire [31:0] n1018_O_5_t0b; // @[Top.scala 1098:23]
  wire [31:0] n1018_O_5_t1b_t0b; // @[Top.scala 1098:23]
  wire [31:0] n1018_O_5_t1b_t1b; // @[Top.scala 1098:23]
  wire [31:0] n1018_O_6_t0b; // @[Top.scala 1098:23]
  wire [31:0] n1018_O_6_t1b_t0b; // @[Top.scala 1098:23]
  wire [31:0] n1018_O_6_t1b_t1b; // @[Top.scala 1098:23]
  wire [31:0] n1018_O_7_t0b; // @[Top.scala 1098:23]
  wire [31:0] n1018_O_7_t1b_t0b; // @[Top.scala 1098:23]
  wire [31:0] n1018_O_7_t1b_t1b; // @[Top.scala 1098:23]
  wire  n1019_clock; // @[Top.scala 1101:23]
  wire  n1019_reset; // @[Top.scala 1101:23]
  wire  n1019_valid_up; // @[Top.scala 1101:23]
  wire  n1019_valid_down; // @[Top.scala 1101:23]
  wire [31:0] n1019_I_0_t0b; // @[Top.scala 1101:23]
  wire [31:0] n1019_I_0_t1b_t0b; // @[Top.scala 1101:23]
  wire [31:0] n1019_I_0_t1b_t1b; // @[Top.scala 1101:23]
  wire [31:0] n1019_I_1_t0b; // @[Top.scala 1101:23]
  wire [31:0] n1019_I_1_t1b_t0b; // @[Top.scala 1101:23]
  wire [31:0] n1019_I_1_t1b_t1b; // @[Top.scala 1101:23]
  wire [31:0] n1019_I_2_t0b; // @[Top.scala 1101:23]
  wire [31:0] n1019_I_2_t1b_t0b; // @[Top.scala 1101:23]
  wire [31:0] n1019_I_2_t1b_t1b; // @[Top.scala 1101:23]
  wire [31:0] n1019_I_3_t0b; // @[Top.scala 1101:23]
  wire [31:0] n1019_I_3_t1b_t0b; // @[Top.scala 1101:23]
  wire [31:0] n1019_I_3_t1b_t1b; // @[Top.scala 1101:23]
  wire [31:0] n1019_I_4_t0b; // @[Top.scala 1101:23]
  wire [31:0] n1019_I_4_t1b_t0b; // @[Top.scala 1101:23]
  wire [31:0] n1019_I_4_t1b_t1b; // @[Top.scala 1101:23]
  wire [31:0] n1019_I_5_t0b; // @[Top.scala 1101:23]
  wire [31:0] n1019_I_5_t1b_t0b; // @[Top.scala 1101:23]
  wire [31:0] n1019_I_5_t1b_t1b; // @[Top.scala 1101:23]
  wire [31:0] n1019_I_6_t0b; // @[Top.scala 1101:23]
  wire [31:0] n1019_I_6_t1b_t0b; // @[Top.scala 1101:23]
  wire [31:0] n1019_I_6_t1b_t1b; // @[Top.scala 1101:23]
  wire [31:0] n1019_I_7_t0b; // @[Top.scala 1101:23]
  wire [31:0] n1019_I_7_t1b_t0b; // @[Top.scala 1101:23]
  wire [31:0] n1019_I_7_t1b_t1b; // @[Top.scala 1101:23]
  wire [31:0] n1019_O_0_t0b; // @[Top.scala 1101:23]
  wire [31:0] n1019_O_0_t1b_t0b; // @[Top.scala 1101:23]
  wire [31:0] n1019_O_0_t1b_t1b; // @[Top.scala 1101:23]
  wire [31:0] n1019_O_1_t0b; // @[Top.scala 1101:23]
  wire [31:0] n1019_O_1_t1b_t0b; // @[Top.scala 1101:23]
  wire [31:0] n1019_O_1_t1b_t1b; // @[Top.scala 1101:23]
  wire [31:0] n1019_O_2_t0b; // @[Top.scala 1101:23]
  wire [31:0] n1019_O_2_t1b_t0b; // @[Top.scala 1101:23]
  wire [31:0] n1019_O_2_t1b_t1b; // @[Top.scala 1101:23]
  wire [31:0] n1019_O_3_t0b; // @[Top.scala 1101:23]
  wire [31:0] n1019_O_3_t1b_t0b; // @[Top.scala 1101:23]
  wire [31:0] n1019_O_3_t1b_t1b; // @[Top.scala 1101:23]
  wire [31:0] n1019_O_4_t0b; // @[Top.scala 1101:23]
  wire [31:0] n1019_O_4_t1b_t0b; // @[Top.scala 1101:23]
  wire [31:0] n1019_O_4_t1b_t1b; // @[Top.scala 1101:23]
  wire [31:0] n1019_O_5_t0b; // @[Top.scala 1101:23]
  wire [31:0] n1019_O_5_t1b_t0b; // @[Top.scala 1101:23]
  wire [31:0] n1019_O_5_t1b_t1b; // @[Top.scala 1101:23]
  wire [31:0] n1019_O_6_t0b; // @[Top.scala 1101:23]
  wire [31:0] n1019_O_6_t1b_t0b; // @[Top.scala 1101:23]
  wire [31:0] n1019_O_6_t1b_t1b; // @[Top.scala 1101:23]
  wire [31:0] n1019_O_7_t0b; // @[Top.scala 1101:23]
  wire [31:0] n1019_O_7_t1b_t0b; // @[Top.scala 1101:23]
  wire [31:0] n1019_O_7_t1b_t1b; // @[Top.scala 1101:23]
  wire  n1020_clock; // @[Top.scala 1104:23]
  wire  n1020_reset; // @[Top.scala 1104:23]
  wire  n1020_valid_up; // @[Top.scala 1104:23]
  wire  n1020_valid_down; // @[Top.scala 1104:23]
  wire [31:0] n1020_I_0_t0b; // @[Top.scala 1104:23]
  wire [31:0] n1020_I_0_t1b_t0b; // @[Top.scala 1104:23]
  wire [31:0] n1020_I_0_t1b_t1b; // @[Top.scala 1104:23]
  wire [31:0] n1020_I_1_t0b; // @[Top.scala 1104:23]
  wire [31:0] n1020_I_1_t1b_t0b; // @[Top.scala 1104:23]
  wire [31:0] n1020_I_1_t1b_t1b; // @[Top.scala 1104:23]
  wire [31:0] n1020_I_2_t0b; // @[Top.scala 1104:23]
  wire [31:0] n1020_I_2_t1b_t0b; // @[Top.scala 1104:23]
  wire [31:0] n1020_I_2_t1b_t1b; // @[Top.scala 1104:23]
  wire [31:0] n1020_I_3_t0b; // @[Top.scala 1104:23]
  wire [31:0] n1020_I_3_t1b_t0b; // @[Top.scala 1104:23]
  wire [31:0] n1020_I_3_t1b_t1b; // @[Top.scala 1104:23]
  wire [31:0] n1020_I_4_t0b; // @[Top.scala 1104:23]
  wire [31:0] n1020_I_4_t1b_t0b; // @[Top.scala 1104:23]
  wire [31:0] n1020_I_4_t1b_t1b; // @[Top.scala 1104:23]
  wire [31:0] n1020_I_5_t0b; // @[Top.scala 1104:23]
  wire [31:0] n1020_I_5_t1b_t0b; // @[Top.scala 1104:23]
  wire [31:0] n1020_I_5_t1b_t1b; // @[Top.scala 1104:23]
  wire [31:0] n1020_I_6_t0b; // @[Top.scala 1104:23]
  wire [31:0] n1020_I_6_t1b_t0b; // @[Top.scala 1104:23]
  wire [31:0] n1020_I_6_t1b_t1b; // @[Top.scala 1104:23]
  wire [31:0] n1020_I_7_t0b; // @[Top.scala 1104:23]
  wire [31:0] n1020_I_7_t1b_t0b; // @[Top.scala 1104:23]
  wire [31:0] n1020_I_7_t1b_t1b; // @[Top.scala 1104:23]
  wire [31:0] n1020_O_0_t0b; // @[Top.scala 1104:23]
  wire [31:0] n1020_O_0_t1b_t0b; // @[Top.scala 1104:23]
  wire [31:0] n1020_O_0_t1b_t1b; // @[Top.scala 1104:23]
  wire [31:0] n1020_O_1_t0b; // @[Top.scala 1104:23]
  wire [31:0] n1020_O_1_t1b_t0b; // @[Top.scala 1104:23]
  wire [31:0] n1020_O_1_t1b_t1b; // @[Top.scala 1104:23]
  wire [31:0] n1020_O_2_t0b; // @[Top.scala 1104:23]
  wire [31:0] n1020_O_2_t1b_t0b; // @[Top.scala 1104:23]
  wire [31:0] n1020_O_2_t1b_t1b; // @[Top.scala 1104:23]
  wire [31:0] n1020_O_3_t0b; // @[Top.scala 1104:23]
  wire [31:0] n1020_O_3_t1b_t0b; // @[Top.scala 1104:23]
  wire [31:0] n1020_O_3_t1b_t1b; // @[Top.scala 1104:23]
  wire [31:0] n1020_O_4_t0b; // @[Top.scala 1104:23]
  wire [31:0] n1020_O_4_t1b_t0b; // @[Top.scala 1104:23]
  wire [31:0] n1020_O_4_t1b_t1b; // @[Top.scala 1104:23]
  wire [31:0] n1020_O_5_t0b; // @[Top.scala 1104:23]
  wire [31:0] n1020_O_5_t1b_t0b; // @[Top.scala 1104:23]
  wire [31:0] n1020_O_5_t1b_t1b; // @[Top.scala 1104:23]
  wire [31:0] n1020_O_6_t0b; // @[Top.scala 1104:23]
  wire [31:0] n1020_O_6_t1b_t0b; // @[Top.scala 1104:23]
  wire [31:0] n1020_O_6_t1b_t1b; // @[Top.scala 1104:23]
  wire [31:0] n1020_O_7_t0b; // @[Top.scala 1104:23]
  wire [31:0] n1020_O_7_t1b_t0b; // @[Top.scala 1104:23]
  wire [31:0] n1020_O_7_t1b_t1b; // @[Top.scala 1104:23]
  FIFO n1 ( // @[Top.scala 695:20]
    .clock(n1_clock),
    .reset(n1_reset),
    .valid_up(n1_valid_up),
    .valid_down(n1_valid_down),
    .I_0(n1_I_0),
    .I_1(n1_I_1),
    .I_2(n1_I_2),
    .I_3(n1_I_3),
    .I_4(n1_I_4),
    .I_5(n1_I_5),
    .I_6(n1_I_6),
    .I_7(n1_I_7),
    .O_0(n1_O_0),
    .O_1(n1_O_1),
    .O_2(n1_O_2),
    .O_3(n1_O_3),
    .O_4(n1_O_4),
    .O_5(n1_O_5),
    .O_6(n1_O_6),
    .O_7(n1_O_7)
  );
  ShiftTS n2 ( // @[Top.scala 698:20]
    .clock(n2_clock),
    .reset(n2_reset),
    .valid_up(n2_valid_up),
    .valid_down(n2_valid_down),
    .I_0(n2_I_0),
    .I_1(n2_I_1),
    .I_2(n2_I_2),
    .I_3(n2_I_3),
    .I_4(n2_I_4),
    .I_5(n2_I_5),
    .I_6(n2_I_6),
    .I_7(n2_I_7),
    .O_0(n2_O_0),
    .O_1(n2_O_1),
    .O_2(n2_O_2),
    .O_3(n2_O_3),
    .O_4(n2_O_4),
    .O_5(n2_O_5),
    .O_6(n2_O_6),
    .O_7(n2_O_7)
  );
  ShiftTS n3 ( // @[Top.scala 701:20]
    .clock(n3_clock),
    .reset(n3_reset),
    .valid_up(n3_valid_up),
    .valid_down(n3_valid_down),
    .I_0(n3_I_0),
    .I_1(n3_I_1),
    .I_2(n3_I_2),
    .I_3(n3_I_3),
    .I_4(n3_I_4),
    .I_5(n3_I_5),
    .I_6(n3_I_6),
    .I_7(n3_I_7),
    .O_0(n3_O_0),
    .O_1(n3_O_1),
    .O_2(n3_O_2),
    .O_3(n3_O_3),
    .O_4(n3_O_4),
    .O_5(n3_O_5),
    .O_6(n3_O_6),
    .O_7(n3_O_7)
  );
  ShiftTS_2 n4 ( // @[Top.scala 704:20]
    .clock(n4_clock),
    .valid_up(n4_valid_up),
    .valid_down(n4_valid_down),
    .I_0(n4_I_0),
    .I_1(n4_I_1),
    .I_2(n4_I_2),
    .I_3(n4_I_3),
    .I_4(n4_I_4),
    .I_5(n4_I_5),
    .I_6(n4_I_6),
    .I_7(n4_I_7),
    .O_0(n4_O_0),
    .O_1(n4_O_1),
    .O_2(n4_O_2),
    .O_3(n4_O_3),
    .O_4(n4_O_4),
    .O_5(n4_O_5),
    .O_6(n4_O_6),
    .O_7(n4_O_7)
  );
  ShiftTS_2 n5 ( // @[Top.scala 707:20]
    .clock(n5_clock),
    .valid_up(n5_valid_up),
    .valid_down(n5_valid_down),
    .I_0(n5_I_0),
    .I_1(n5_I_1),
    .I_2(n5_I_2),
    .I_3(n5_I_3),
    .I_4(n5_I_4),
    .I_5(n5_I_5),
    .I_6(n5_I_6),
    .I_7(n5_I_7),
    .O_0(n5_O_0),
    .O_1(n5_O_1),
    .O_2(n5_O_2),
    .O_3(n5_O_3),
    .O_4(n5_O_4),
    .O_5(n5_O_5),
    .O_6(n5_O_6),
    .O_7(n5_O_7)
  );
  Map2T n6 ( // @[Top.scala 710:20]
    .valid_up(n6_valid_up),
    .valid_down(n6_valid_down),
    .I0_0(n6_I0_0),
    .I0_1(n6_I0_1),
    .I0_2(n6_I0_2),
    .I0_3(n6_I0_3),
    .I0_4(n6_I0_4),
    .I0_5(n6_I0_5),
    .I0_6(n6_I0_6),
    .I0_7(n6_I0_7),
    .I1_0(n6_I1_0),
    .I1_1(n6_I1_1),
    .I1_2(n6_I1_2),
    .I1_3(n6_I1_3),
    .I1_4(n6_I1_4),
    .I1_5(n6_I1_5),
    .I1_6(n6_I1_6),
    .I1_7(n6_I1_7),
    .O_0_0(n6_O_0_0),
    .O_0_1(n6_O_0_1),
    .O_1_0(n6_O_1_0),
    .O_1_1(n6_O_1_1),
    .O_2_0(n6_O_2_0),
    .O_2_1(n6_O_2_1),
    .O_3_0(n6_O_3_0),
    .O_3_1(n6_O_3_1),
    .O_4_0(n6_O_4_0),
    .O_4_1(n6_O_4_1),
    .O_5_0(n6_O_5_0),
    .O_5_1(n6_O_5_1),
    .O_6_0(n6_O_6_0),
    .O_6_1(n6_O_6_1),
    .O_7_0(n6_O_7_0),
    .O_7_1(n6_O_7_1)
  );
  Map2T_1 n13 ( // @[Top.scala 714:21]
    .valid_up(n13_valid_up),
    .valid_down(n13_valid_down),
    .I0_0_0(n13_I0_0_0),
    .I0_0_1(n13_I0_0_1),
    .I0_1_0(n13_I0_1_0),
    .I0_1_1(n13_I0_1_1),
    .I0_2_0(n13_I0_2_0),
    .I0_2_1(n13_I0_2_1),
    .I0_3_0(n13_I0_3_0),
    .I0_3_1(n13_I0_3_1),
    .I0_4_0(n13_I0_4_0),
    .I0_4_1(n13_I0_4_1),
    .I0_5_0(n13_I0_5_0),
    .I0_5_1(n13_I0_5_1),
    .I0_6_0(n13_I0_6_0),
    .I0_6_1(n13_I0_6_1),
    .I0_7_0(n13_I0_7_0),
    .I0_7_1(n13_I0_7_1),
    .I1_0(n13_I1_0),
    .I1_1(n13_I1_1),
    .I1_2(n13_I1_2),
    .I1_3(n13_I1_3),
    .I1_4(n13_I1_4),
    .I1_5(n13_I1_5),
    .I1_6(n13_I1_6),
    .I1_7(n13_I1_7),
    .O_0_0(n13_O_0_0),
    .O_0_1(n13_O_0_1),
    .O_0_2(n13_O_0_2),
    .O_1_0(n13_O_1_0),
    .O_1_1(n13_O_1_1),
    .O_1_2(n13_O_1_2),
    .O_2_0(n13_O_2_0),
    .O_2_1(n13_O_2_1),
    .O_2_2(n13_O_2_2),
    .O_3_0(n13_O_3_0),
    .O_3_1(n13_O_3_1),
    .O_3_2(n13_O_3_2),
    .O_4_0(n13_O_4_0),
    .O_4_1(n13_O_4_1),
    .O_4_2(n13_O_4_2),
    .O_5_0(n13_O_5_0),
    .O_5_1(n13_O_5_1),
    .O_5_2(n13_O_5_2),
    .O_6_0(n13_O_6_0),
    .O_6_1(n13_O_6_1),
    .O_6_2(n13_O_6_2),
    .O_7_0(n13_O_7_0),
    .O_7_1(n13_O_7_1),
    .O_7_2(n13_O_7_2)
  );
  MapT n22 ( // @[Top.scala 718:21]
    .valid_up(n22_valid_up),
    .valid_down(n22_valid_down),
    .I_0_0(n22_I_0_0),
    .I_0_1(n22_I_0_1),
    .I_0_2(n22_I_0_2),
    .I_1_0(n22_I_1_0),
    .I_1_1(n22_I_1_1),
    .I_1_2(n22_I_1_2),
    .I_2_0(n22_I_2_0),
    .I_2_1(n22_I_2_1),
    .I_2_2(n22_I_2_2),
    .I_3_0(n22_I_3_0),
    .I_3_1(n22_I_3_1),
    .I_3_2(n22_I_3_2),
    .I_4_0(n22_I_4_0),
    .I_4_1(n22_I_4_1),
    .I_4_2(n22_I_4_2),
    .I_5_0(n22_I_5_0),
    .I_5_1(n22_I_5_1),
    .I_5_2(n22_I_5_2),
    .I_6_0(n22_I_6_0),
    .I_6_1(n22_I_6_1),
    .I_6_2(n22_I_6_2),
    .I_7_0(n22_I_7_0),
    .I_7_1(n22_I_7_1),
    .I_7_2(n22_I_7_2),
    .O_0_0_0(n22_O_0_0_0),
    .O_0_0_1(n22_O_0_0_1),
    .O_0_0_2(n22_O_0_0_2),
    .O_1_0_0(n22_O_1_0_0),
    .O_1_0_1(n22_O_1_0_1),
    .O_1_0_2(n22_O_1_0_2),
    .O_2_0_0(n22_O_2_0_0),
    .O_2_0_1(n22_O_2_0_1),
    .O_2_0_2(n22_O_2_0_2),
    .O_3_0_0(n22_O_3_0_0),
    .O_3_0_1(n22_O_3_0_1),
    .O_3_0_2(n22_O_3_0_2),
    .O_4_0_0(n22_O_4_0_0),
    .O_4_0_1(n22_O_4_0_1),
    .O_4_0_2(n22_O_4_0_2),
    .O_5_0_0(n22_O_5_0_0),
    .O_5_0_1(n22_O_5_0_1),
    .O_5_0_2(n22_O_5_0_2),
    .O_6_0_0(n22_O_6_0_0),
    .O_6_0_1(n22_O_6_0_1),
    .O_6_0_2(n22_O_6_0_2),
    .O_7_0_0(n22_O_7_0_0),
    .O_7_0_1(n22_O_7_0_1),
    .O_7_0_2(n22_O_7_0_2)
  );
  MapT_1 n29 ( // @[Top.scala 721:21]
    .valid_up(n29_valid_up),
    .valid_down(n29_valid_down),
    .I_0_0_0(n29_I_0_0_0),
    .I_0_0_1(n29_I_0_0_1),
    .I_0_0_2(n29_I_0_0_2),
    .I_1_0_0(n29_I_1_0_0),
    .I_1_0_1(n29_I_1_0_1),
    .I_1_0_2(n29_I_1_0_2),
    .I_2_0_0(n29_I_2_0_0),
    .I_2_0_1(n29_I_2_0_1),
    .I_2_0_2(n29_I_2_0_2),
    .I_3_0_0(n29_I_3_0_0),
    .I_3_0_1(n29_I_3_0_1),
    .I_3_0_2(n29_I_3_0_2),
    .I_4_0_0(n29_I_4_0_0),
    .I_4_0_1(n29_I_4_0_1),
    .I_4_0_2(n29_I_4_0_2),
    .I_5_0_0(n29_I_5_0_0),
    .I_5_0_1(n29_I_5_0_1),
    .I_5_0_2(n29_I_5_0_2),
    .I_6_0_0(n29_I_6_0_0),
    .I_6_0_1(n29_I_6_0_1),
    .I_6_0_2(n29_I_6_0_2),
    .I_7_0_0(n29_I_7_0_0),
    .I_7_0_1(n29_I_7_0_1),
    .I_7_0_2(n29_I_7_0_2),
    .O_0_0(n29_O_0_0),
    .O_0_1(n29_O_0_1),
    .O_0_2(n29_O_0_2),
    .O_1_0(n29_O_1_0),
    .O_1_1(n29_O_1_1),
    .O_1_2(n29_O_1_2),
    .O_2_0(n29_O_2_0),
    .O_2_1(n29_O_2_1),
    .O_2_2(n29_O_2_2),
    .O_3_0(n29_O_3_0),
    .O_3_1(n29_O_3_1),
    .O_3_2(n29_O_3_2),
    .O_4_0(n29_O_4_0),
    .O_4_1(n29_O_4_1),
    .O_4_2(n29_O_4_2),
    .O_5_0(n29_O_5_0),
    .O_5_1(n29_O_5_1),
    .O_5_2(n29_O_5_2),
    .O_6_0(n29_O_6_0),
    .O_6_1(n29_O_6_1),
    .O_6_2(n29_O_6_2),
    .O_7_0(n29_O_7_0),
    .O_7_1(n29_O_7_1),
    .O_7_2(n29_O_7_2)
  );
  ShiftTS_2 n30 ( // @[Top.scala 724:21]
    .clock(n30_clock),
    .valid_up(n30_valid_up),
    .valid_down(n30_valid_down),
    .I_0(n30_I_0),
    .I_1(n30_I_1),
    .I_2(n30_I_2),
    .I_3(n30_I_3),
    .I_4(n30_I_4),
    .I_5(n30_I_5),
    .I_6(n30_I_6),
    .I_7(n30_I_7),
    .O_0(n30_O_0),
    .O_1(n30_O_1),
    .O_2(n30_O_2),
    .O_3(n30_O_3),
    .O_4(n30_O_4),
    .O_5(n30_O_5),
    .O_6(n30_O_6),
    .O_7(n30_O_7)
  );
  ShiftTS_2 n31 ( // @[Top.scala 727:21]
    .clock(n31_clock),
    .valid_up(n31_valid_up),
    .valid_down(n31_valid_down),
    .I_0(n31_I_0),
    .I_1(n31_I_1),
    .I_2(n31_I_2),
    .I_3(n31_I_3),
    .I_4(n31_I_4),
    .I_5(n31_I_5),
    .I_6(n31_I_6),
    .I_7(n31_I_7),
    .O_0(n31_O_0),
    .O_1(n31_O_1),
    .O_2(n31_O_2),
    .O_3(n31_O_3),
    .O_4(n31_O_4),
    .O_5(n31_O_5),
    .O_6(n31_O_6),
    .O_7(n31_O_7)
  );
  Map2T n32 ( // @[Top.scala 730:21]
    .valid_up(n32_valid_up),
    .valid_down(n32_valid_down),
    .I0_0(n32_I0_0),
    .I0_1(n32_I0_1),
    .I0_2(n32_I0_2),
    .I0_3(n32_I0_3),
    .I0_4(n32_I0_4),
    .I0_5(n32_I0_5),
    .I0_6(n32_I0_6),
    .I0_7(n32_I0_7),
    .I1_0(n32_I1_0),
    .I1_1(n32_I1_1),
    .I1_2(n32_I1_2),
    .I1_3(n32_I1_3),
    .I1_4(n32_I1_4),
    .I1_5(n32_I1_5),
    .I1_6(n32_I1_6),
    .I1_7(n32_I1_7),
    .O_0_0(n32_O_0_0),
    .O_0_1(n32_O_0_1),
    .O_1_0(n32_O_1_0),
    .O_1_1(n32_O_1_1),
    .O_2_0(n32_O_2_0),
    .O_2_1(n32_O_2_1),
    .O_3_0(n32_O_3_0),
    .O_3_1(n32_O_3_1),
    .O_4_0(n32_O_4_0),
    .O_4_1(n32_O_4_1),
    .O_5_0(n32_O_5_0),
    .O_5_1(n32_O_5_1),
    .O_6_0(n32_O_6_0),
    .O_6_1(n32_O_6_1),
    .O_7_0(n32_O_7_0),
    .O_7_1(n32_O_7_1)
  );
  Map2T_1 n39 ( // @[Top.scala 734:21]
    .valid_up(n39_valid_up),
    .valid_down(n39_valid_down),
    .I0_0_0(n39_I0_0_0),
    .I0_0_1(n39_I0_0_1),
    .I0_1_0(n39_I0_1_0),
    .I0_1_1(n39_I0_1_1),
    .I0_2_0(n39_I0_2_0),
    .I0_2_1(n39_I0_2_1),
    .I0_3_0(n39_I0_3_0),
    .I0_3_1(n39_I0_3_1),
    .I0_4_0(n39_I0_4_0),
    .I0_4_1(n39_I0_4_1),
    .I0_5_0(n39_I0_5_0),
    .I0_5_1(n39_I0_5_1),
    .I0_6_0(n39_I0_6_0),
    .I0_6_1(n39_I0_6_1),
    .I0_7_0(n39_I0_7_0),
    .I0_7_1(n39_I0_7_1),
    .I1_0(n39_I1_0),
    .I1_1(n39_I1_1),
    .I1_2(n39_I1_2),
    .I1_3(n39_I1_3),
    .I1_4(n39_I1_4),
    .I1_5(n39_I1_5),
    .I1_6(n39_I1_6),
    .I1_7(n39_I1_7),
    .O_0_0(n39_O_0_0),
    .O_0_1(n39_O_0_1),
    .O_0_2(n39_O_0_2),
    .O_1_0(n39_O_1_0),
    .O_1_1(n39_O_1_1),
    .O_1_2(n39_O_1_2),
    .O_2_0(n39_O_2_0),
    .O_2_1(n39_O_2_1),
    .O_2_2(n39_O_2_2),
    .O_3_0(n39_O_3_0),
    .O_3_1(n39_O_3_1),
    .O_3_2(n39_O_3_2),
    .O_4_0(n39_O_4_0),
    .O_4_1(n39_O_4_1),
    .O_4_2(n39_O_4_2),
    .O_5_0(n39_O_5_0),
    .O_5_1(n39_O_5_1),
    .O_5_2(n39_O_5_2),
    .O_6_0(n39_O_6_0),
    .O_6_1(n39_O_6_1),
    .O_6_2(n39_O_6_2),
    .O_7_0(n39_O_7_0),
    .O_7_1(n39_O_7_1),
    .O_7_2(n39_O_7_2)
  );
  MapT n48 ( // @[Top.scala 738:21]
    .valid_up(n48_valid_up),
    .valid_down(n48_valid_down),
    .I_0_0(n48_I_0_0),
    .I_0_1(n48_I_0_1),
    .I_0_2(n48_I_0_2),
    .I_1_0(n48_I_1_0),
    .I_1_1(n48_I_1_1),
    .I_1_2(n48_I_1_2),
    .I_2_0(n48_I_2_0),
    .I_2_1(n48_I_2_1),
    .I_2_2(n48_I_2_2),
    .I_3_0(n48_I_3_0),
    .I_3_1(n48_I_3_1),
    .I_3_2(n48_I_3_2),
    .I_4_0(n48_I_4_0),
    .I_4_1(n48_I_4_1),
    .I_4_2(n48_I_4_2),
    .I_5_0(n48_I_5_0),
    .I_5_1(n48_I_5_1),
    .I_5_2(n48_I_5_2),
    .I_6_0(n48_I_6_0),
    .I_6_1(n48_I_6_1),
    .I_6_2(n48_I_6_2),
    .I_7_0(n48_I_7_0),
    .I_7_1(n48_I_7_1),
    .I_7_2(n48_I_7_2),
    .O_0_0_0(n48_O_0_0_0),
    .O_0_0_1(n48_O_0_0_1),
    .O_0_0_2(n48_O_0_0_2),
    .O_1_0_0(n48_O_1_0_0),
    .O_1_0_1(n48_O_1_0_1),
    .O_1_0_2(n48_O_1_0_2),
    .O_2_0_0(n48_O_2_0_0),
    .O_2_0_1(n48_O_2_0_1),
    .O_2_0_2(n48_O_2_0_2),
    .O_3_0_0(n48_O_3_0_0),
    .O_3_0_1(n48_O_3_0_1),
    .O_3_0_2(n48_O_3_0_2),
    .O_4_0_0(n48_O_4_0_0),
    .O_4_0_1(n48_O_4_0_1),
    .O_4_0_2(n48_O_4_0_2),
    .O_5_0_0(n48_O_5_0_0),
    .O_5_0_1(n48_O_5_0_1),
    .O_5_0_2(n48_O_5_0_2),
    .O_6_0_0(n48_O_6_0_0),
    .O_6_0_1(n48_O_6_0_1),
    .O_6_0_2(n48_O_6_0_2),
    .O_7_0_0(n48_O_7_0_0),
    .O_7_0_1(n48_O_7_0_1),
    .O_7_0_2(n48_O_7_0_2)
  );
  MapT_1 n55 ( // @[Top.scala 741:21]
    .valid_up(n55_valid_up),
    .valid_down(n55_valid_down),
    .I_0_0_0(n55_I_0_0_0),
    .I_0_0_1(n55_I_0_0_1),
    .I_0_0_2(n55_I_0_0_2),
    .I_1_0_0(n55_I_1_0_0),
    .I_1_0_1(n55_I_1_0_1),
    .I_1_0_2(n55_I_1_0_2),
    .I_2_0_0(n55_I_2_0_0),
    .I_2_0_1(n55_I_2_0_1),
    .I_2_0_2(n55_I_2_0_2),
    .I_3_0_0(n55_I_3_0_0),
    .I_3_0_1(n55_I_3_0_1),
    .I_3_0_2(n55_I_3_0_2),
    .I_4_0_0(n55_I_4_0_0),
    .I_4_0_1(n55_I_4_0_1),
    .I_4_0_2(n55_I_4_0_2),
    .I_5_0_0(n55_I_5_0_0),
    .I_5_0_1(n55_I_5_0_1),
    .I_5_0_2(n55_I_5_0_2),
    .I_6_0_0(n55_I_6_0_0),
    .I_6_0_1(n55_I_6_0_1),
    .I_6_0_2(n55_I_6_0_2),
    .I_7_0_0(n55_I_7_0_0),
    .I_7_0_1(n55_I_7_0_1),
    .I_7_0_2(n55_I_7_0_2),
    .O_0_0(n55_O_0_0),
    .O_0_1(n55_O_0_1),
    .O_0_2(n55_O_0_2),
    .O_1_0(n55_O_1_0),
    .O_1_1(n55_O_1_1),
    .O_1_2(n55_O_1_2),
    .O_2_0(n55_O_2_0),
    .O_2_1(n55_O_2_1),
    .O_2_2(n55_O_2_2),
    .O_3_0(n55_O_3_0),
    .O_3_1(n55_O_3_1),
    .O_3_2(n55_O_3_2),
    .O_4_0(n55_O_4_0),
    .O_4_1(n55_O_4_1),
    .O_4_2(n55_O_4_2),
    .O_5_0(n55_O_5_0),
    .O_5_1(n55_O_5_1),
    .O_5_2(n55_O_5_2),
    .O_6_0(n55_O_6_0),
    .O_6_1(n55_O_6_1),
    .O_6_2(n55_O_6_2),
    .O_7_0(n55_O_7_0),
    .O_7_1(n55_O_7_1),
    .O_7_2(n55_O_7_2)
  );
  Map2T_4 n56 ( // @[Top.scala 744:21]
    .valid_up(n56_valid_up),
    .valid_down(n56_valid_down),
    .I0_0_0(n56_I0_0_0),
    .I0_0_1(n56_I0_0_1),
    .I0_0_2(n56_I0_0_2),
    .I0_1_0(n56_I0_1_0),
    .I0_1_1(n56_I0_1_1),
    .I0_1_2(n56_I0_1_2),
    .I0_2_0(n56_I0_2_0),
    .I0_2_1(n56_I0_2_1),
    .I0_2_2(n56_I0_2_2),
    .I0_3_0(n56_I0_3_0),
    .I0_3_1(n56_I0_3_1),
    .I0_3_2(n56_I0_3_2),
    .I0_4_0(n56_I0_4_0),
    .I0_4_1(n56_I0_4_1),
    .I0_4_2(n56_I0_4_2),
    .I0_5_0(n56_I0_5_0),
    .I0_5_1(n56_I0_5_1),
    .I0_5_2(n56_I0_5_2),
    .I0_6_0(n56_I0_6_0),
    .I0_6_1(n56_I0_6_1),
    .I0_6_2(n56_I0_6_2),
    .I0_7_0(n56_I0_7_0),
    .I0_7_1(n56_I0_7_1),
    .I0_7_2(n56_I0_7_2),
    .I1_0_0(n56_I1_0_0),
    .I1_0_1(n56_I1_0_1),
    .I1_0_2(n56_I1_0_2),
    .I1_1_0(n56_I1_1_0),
    .I1_1_1(n56_I1_1_1),
    .I1_1_2(n56_I1_1_2),
    .I1_2_0(n56_I1_2_0),
    .I1_2_1(n56_I1_2_1),
    .I1_2_2(n56_I1_2_2),
    .I1_3_0(n56_I1_3_0),
    .I1_3_1(n56_I1_3_1),
    .I1_3_2(n56_I1_3_2),
    .I1_4_0(n56_I1_4_0),
    .I1_4_1(n56_I1_4_1),
    .I1_4_2(n56_I1_4_2),
    .I1_5_0(n56_I1_5_0),
    .I1_5_1(n56_I1_5_1),
    .I1_5_2(n56_I1_5_2),
    .I1_6_0(n56_I1_6_0),
    .I1_6_1(n56_I1_6_1),
    .I1_6_2(n56_I1_6_2),
    .I1_7_0(n56_I1_7_0),
    .I1_7_1(n56_I1_7_1),
    .I1_7_2(n56_I1_7_2),
    .O_0_0_0(n56_O_0_0_0),
    .O_0_0_1(n56_O_0_0_1),
    .O_0_0_2(n56_O_0_0_2),
    .O_0_1_0(n56_O_0_1_0),
    .O_0_1_1(n56_O_0_1_1),
    .O_0_1_2(n56_O_0_1_2),
    .O_1_0_0(n56_O_1_0_0),
    .O_1_0_1(n56_O_1_0_1),
    .O_1_0_2(n56_O_1_0_2),
    .O_1_1_0(n56_O_1_1_0),
    .O_1_1_1(n56_O_1_1_1),
    .O_1_1_2(n56_O_1_1_2),
    .O_2_0_0(n56_O_2_0_0),
    .O_2_0_1(n56_O_2_0_1),
    .O_2_0_2(n56_O_2_0_2),
    .O_2_1_0(n56_O_2_1_0),
    .O_2_1_1(n56_O_2_1_1),
    .O_2_1_2(n56_O_2_1_2),
    .O_3_0_0(n56_O_3_0_0),
    .O_3_0_1(n56_O_3_0_1),
    .O_3_0_2(n56_O_3_0_2),
    .O_3_1_0(n56_O_3_1_0),
    .O_3_1_1(n56_O_3_1_1),
    .O_3_1_2(n56_O_3_1_2),
    .O_4_0_0(n56_O_4_0_0),
    .O_4_0_1(n56_O_4_0_1),
    .O_4_0_2(n56_O_4_0_2),
    .O_4_1_0(n56_O_4_1_0),
    .O_4_1_1(n56_O_4_1_1),
    .O_4_1_2(n56_O_4_1_2),
    .O_5_0_0(n56_O_5_0_0),
    .O_5_0_1(n56_O_5_0_1),
    .O_5_0_2(n56_O_5_0_2),
    .O_5_1_0(n56_O_5_1_0),
    .O_5_1_1(n56_O_5_1_1),
    .O_5_1_2(n56_O_5_1_2),
    .O_6_0_0(n56_O_6_0_0),
    .O_6_0_1(n56_O_6_0_1),
    .O_6_0_2(n56_O_6_0_2),
    .O_6_1_0(n56_O_6_1_0),
    .O_6_1_1(n56_O_6_1_1),
    .O_6_1_2(n56_O_6_1_2),
    .O_7_0_0(n56_O_7_0_0),
    .O_7_0_1(n56_O_7_0_1),
    .O_7_0_2(n56_O_7_0_2),
    .O_7_1_0(n56_O_7_1_0),
    .O_7_1_1(n56_O_7_1_1),
    .O_7_1_2(n56_O_7_1_2)
  );
  ShiftTS_2 n63 ( // @[Top.scala 748:21]
    .clock(n63_clock),
    .valid_up(n63_valid_up),
    .valid_down(n63_valid_down),
    .I_0(n63_I_0),
    .I_1(n63_I_1),
    .I_2(n63_I_2),
    .I_3(n63_I_3),
    .I_4(n63_I_4),
    .I_5(n63_I_5),
    .I_6(n63_I_6),
    .I_7(n63_I_7),
    .O_0(n63_O_0),
    .O_1(n63_O_1),
    .O_2(n63_O_2),
    .O_3(n63_O_3),
    .O_4(n63_O_4),
    .O_5(n63_O_5),
    .O_6(n63_O_6),
    .O_7(n63_O_7)
  );
  ShiftTS_2 n64 ( // @[Top.scala 751:21]
    .clock(n64_clock),
    .valid_up(n64_valid_up),
    .valid_down(n64_valid_down),
    .I_0(n64_I_0),
    .I_1(n64_I_1),
    .I_2(n64_I_2),
    .I_3(n64_I_3),
    .I_4(n64_I_4),
    .I_5(n64_I_5),
    .I_6(n64_I_6),
    .I_7(n64_I_7),
    .O_0(n64_O_0),
    .O_1(n64_O_1),
    .O_2(n64_O_2),
    .O_3(n64_O_3),
    .O_4(n64_O_4),
    .O_5(n64_O_5),
    .O_6(n64_O_6),
    .O_7(n64_O_7)
  );
  Map2T n65 ( // @[Top.scala 754:21]
    .valid_up(n65_valid_up),
    .valid_down(n65_valid_down),
    .I0_0(n65_I0_0),
    .I0_1(n65_I0_1),
    .I0_2(n65_I0_2),
    .I0_3(n65_I0_3),
    .I0_4(n65_I0_4),
    .I0_5(n65_I0_5),
    .I0_6(n65_I0_6),
    .I0_7(n65_I0_7),
    .I1_0(n65_I1_0),
    .I1_1(n65_I1_1),
    .I1_2(n65_I1_2),
    .I1_3(n65_I1_3),
    .I1_4(n65_I1_4),
    .I1_5(n65_I1_5),
    .I1_6(n65_I1_6),
    .I1_7(n65_I1_7),
    .O_0_0(n65_O_0_0),
    .O_0_1(n65_O_0_1),
    .O_1_0(n65_O_1_0),
    .O_1_1(n65_O_1_1),
    .O_2_0(n65_O_2_0),
    .O_2_1(n65_O_2_1),
    .O_3_0(n65_O_3_0),
    .O_3_1(n65_O_3_1),
    .O_4_0(n65_O_4_0),
    .O_4_1(n65_O_4_1),
    .O_5_0(n65_O_5_0),
    .O_5_1(n65_O_5_1),
    .O_6_0(n65_O_6_0),
    .O_6_1(n65_O_6_1),
    .O_7_0(n65_O_7_0),
    .O_7_1(n65_O_7_1)
  );
  Map2T_1 n72 ( // @[Top.scala 758:21]
    .valid_up(n72_valid_up),
    .valid_down(n72_valid_down),
    .I0_0_0(n72_I0_0_0),
    .I0_0_1(n72_I0_0_1),
    .I0_1_0(n72_I0_1_0),
    .I0_1_1(n72_I0_1_1),
    .I0_2_0(n72_I0_2_0),
    .I0_2_1(n72_I0_2_1),
    .I0_3_0(n72_I0_3_0),
    .I0_3_1(n72_I0_3_1),
    .I0_4_0(n72_I0_4_0),
    .I0_4_1(n72_I0_4_1),
    .I0_5_0(n72_I0_5_0),
    .I0_5_1(n72_I0_5_1),
    .I0_6_0(n72_I0_6_0),
    .I0_6_1(n72_I0_6_1),
    .I0_7_0(n72_I0_7_0),
    .I0_7_1(n72_I0_7_1),
    .I1_0(n72_I1_0),
    .I1_1(n72_I1_1),
    .I1_2(n72_I1_2),
    .I1_3(n72_I1_3),
    .I1_4(n72_I1_4),
    .I1_5(n72_I1_5),
    .I1_6(n72_I1_6),
    .I1_7(n72_I1_7),
    .O_0_0(n72_O_0_0),
    .O_0_1(n72_O_0_1),
    .O_0_2(n72_O_0_2),
    .O_1_0(n72_O_1_0),
    .O_1_1(n72_O_1_1),
    .O_1_2(n72_O_1_2),
    .O_2_0(n72_O_2_0),
    .O_2_1(n72_O_2_1),
    .O_2_2(n72_O_2_2),
    .O_3_0(n72_O_3_0),
    .O_3_1(n72_O_3_1),
    .O_3_2(n72_O_3_2),
    .O_4_0(n72_O_4_0),
    .O_4_1(n72_O_4_1),
    .O_4_2(n72_O_4_2),
    .O_5_0(n72_O_5_0),
    .O_5_1(n72_O_5_1),
    .O_5_2(n72_O_5_2),
    .O_6_0(n72_O_6_0),
    .O_6_1(n72_O_6_1),
    .O_6_2(n72_O_6_2),
    .O_7_0(n72_O_7_0),
    .O_7_1(n72_O_7_1),
    .O_7_2(n72_O_7_2)
  );
  MapT n81 ( // @[Top.scala 762:21]
    .valid_up(n81_valid_up),
    .valid_down(n81_valid_down),
    .I_0_0(n81_I_0_0),
    .I_0_1(n81_I_0_1),
    .I_0_2(n81_I_0_2),
    .I_1_0(n81_I_1_0),
    .I_1_1(n81_I_1_1),
    .I_1_2(n81_I_1_2),
    .I_2_0(n81_I_2_0),
    .I_2_1(n81_I_2_1),
    .I_2_2(n81_I_2_2),
    .I_3_0(n81_I_3_0),
    .I_3_1(n81_I_3_1),
    .I_3_2(n81_I_3_2),
    .I_4_0(n81_I_4_0),
    .I_4_1(n81_I_4_1),
    .I_4_2(n81_I_4_2),
    .I_5_0(n81_I_5_0),
    .I_5_1(n81_I_5_1),
    .I_5_2(n81_I_5_2),
    .I_6_0(n81_I_6_0),
    .I_6_1(n81_I_6_1),
    .I_6_2(n81_I_6_2),
    .I_7_0(n81_I_7_0),
    .I_7_1(n81_I_7_1),
    .I_7_2(n81_I_7_2),
    .O_0_0_0(n81_O_0_0_0),
    .O_0_0_1(n81_O_0_0_1),
    .O_0_0_2(n81_O_0_0_2),
    .O_1_0_0(n81_O_1_0_0),
    .O_1_0_1(n81_O_1_0_1),
    .O_1_0_2(n81_O_1_0_2),
    .O_2_0_0(n81_O_2_0_0),
    .O_2_0_1(n81_O_2_0_1),
    .O_2_0_2(n81_O_2_0_2),
    .O_3_0_0(n81_O_3_0_0),
    .O_3_0_1(n81_O_3_0_1),
    .O_3_0_2(n81_O_3_0_2),
    .O_4_0_0(n81_O_4_0_0),
    .O_4_0_1(n81_O_4_0_1),
    .O_4_0_2(n81_O_4_0_2),
    .O_5_0_0(n81_O_5_0_0),
    .O_5_0_1(n81_O_5_0_1),
    .O_5_0_2(n81_O_5_0_2),
    .O_6_0_0(n81_O_6_0_0),
    .O_6_0_1(n81_O_6_0_1),
    .O_6_0_2(n81_O_6_0_2),
    .O_7_0_0(n81_O_7_0_0),
    .O_7_0_1(n81_O_7_0_1),
    .O_7_0_2(n81_O_7_0_2)
  );
  MapT_1 n88 ( // @[Top.scala 765:21]
    .valid_up(n88_valid_up),
    .valid_down(n88_valid_down),
    .I_0_0_0(n88_I_0_0_0),
    .I_0_0_1(n88_I_0_0_1),
    .I_0_0_2(n88_I_0_0_2),
    .I_1_0_0(n88_I_1_0_0),
    .I_1_0_1(n88_I_1_0_1),
    .I_1_0_2(n88_I_1_0_2),
    .I_2_0_0(n88_I_2_0_0),
    .I_2_0_1(n88_I_2_0_1),
    .I_2_0_2(n88_I_2_0_2),
    .I_3_0_0(n88_I_3_0_0),
    .I_3_0_1(n88_I_3_0_1),
    .I_3_0_2(n88_I_3_0_2),
    .I_4_0_0(n88_I_4_0_0),
    .I_4_0_1(n88_I_4_0_1),
    .I_4_0_2(n88_I_4_0_2),
    .I_5_0_0(n88_I_5_0_0),
    .I_5_0_1(n88_I_5_0_1),
    .I_5_0_2(n88_I_5_0_2),
    .I_6_0_0(n88_I_6_0_0),
    .I_6_0_1(n88_I_6_0_1),
    .I_6_0_2(n88_I_6_0_2),
    .I_7_0_0(n88_I_7_0_0),
    .I_7_0_1(n88_I_7_0_1),
    .I_7_0_2(n88_I_7_0_2),
    .O_0_0(n88_O_0_0),
    .O_0_1(n88_O_0_1),
    .O_0_2(n88_O_0_2),
    .O_1_0(n88_O_1_0),
    .O_1_1(n88_O_1_1),
    .O_1_2(n88_O_1_2),
    .O_2_0(n88_O_2_0),
    .O_2_1(n88_O_2_1),
    .O_2_2(n88_O_2_2),
    .O_3_0(n88_O_3_0),
    .O_3_1(n88_O_3_1),
    .O_3_2(n88_O_3_2),
    .O_4_0(n88_O_4_0),
    .O_4_1(n88_O_4_1),
    .O_4_2(n88_O_4_2),
    .O_5_0(n88_O_5_0),
    .O_5_1(n88_O_5_1),
    .O_5_2(n88_O_5_2),
    .O_6_0(n88_O_6_0),
    .O_6_1(n88_O_6_1),
    .O_6_2(n88_O_6_2),
    .O_7_0(n88_O_7_0),
    .O_7_1(n88_O_7_1),
    .O_7_2(n88_O_7_2)
  );
  Map2T_7 n89 ( // @[Top.scala 768:21]
    .valid_up(n89_valid_up),
    .valid_down(n89_valid_down),
    .I0_0_0_0(n89_I0_0_0_0),
    .I0_0_0_1(n89_I0_0_0_1),
    .I0_0_0_2(n89_I0_0_0_2),
    .I0_0_1_0(n89_I0_0_1_0),
    .I0_0_1_1(n89_I0_0_1_1),
    .I0_0_1_2(n89_I0_0_1_2),
    .I0_1_0_0(n89_I0_1_0_0),
    .I0_1_0_1(n89_I0_1_0_1),
    .I0_1_0_2(n89_I0_1_0_2),
    .I0_1_1_0(n89_I0_1_1_0),
    .I0_1_1_1(n89_I0_1_1_1),
    .I0_1_1_2(n89_I0_1_1_2),
    .I0_2_0_0(n89_I0_2_0_0),
    .I0_2_0_1(n89_I0_2_0_1),
    .I0_2_0_2(n89_I0_2_0_2),
    .I0_2_1_0(n89_I0_2_1_0),
    .I0_2_1_1(n89_I0_2_1_1),
    .I0_2_1_2(n89_I0_2_1_2),
    .I0_3_0_0(n89_I0_3_0_0),
    .I0_3_0_1(n89_I0_3_0_1),
    .I0_3_0_2(n89_I0_3_0_2),
    .I0_3_1_0(n89_I0_3_1_0),
    .I0_3_1_1(n89_I0_3_1_1),
    .I0_3_1_2(n89_I0_3_1_2),
    .I0_4_0_0(n89_I0_4_0_0),
    .I0_4_0_1(n89_I0_4_0_1),
    .I0_4_0_2(n89_I0_4_0_2),
    .I0_4_1_0(n89_I0_4_1_0),
    .I0_4_1_1(n89_I0_4_1_1),
    .I0_4_1_2(n89_I0_4_1_2),
    .I0_5_0_0(n89_I0_5_0_0),
    .I0_5_0_1(n89_I0_5_0_1),
    .I0_5_0_2(n89_I0_5_0_2),
    .I0_5_1_0(n89_I0_5_1_0),
    .I0_5_1_1(n89_I0_5_1_1),
    .I0_5_1_2(n89_I0_5_1_2),
    .I0_6_0_0(n89_I0_6_0_0),
    .I0_6_0_1(n89_I0_6_0_1),
    .I0_6_0_2(n89_I0_6_0_2),
    .I0_6_1_0(n89_I0_6_1_0),
    .I0_6_1_1(n89_I0_6_1_1),
    .I0_6_1_2(n89_I0_6_1_2),
    .I0_7_0_0(n89_I0_7_0_0),
    .I0_7_0_1(n89_I0_7_0_1),
    .I0_7_0_2(n89_I0_7_0_2),
    .I0_7_1_0(n89_I0_7_1_0),
    .I0_7_1_1(n89_I0_7_1_1),
    .I0_7_1_2(n89_I0_7_1_2),
    .I1_0_0(n89_I1_0_0),
    .I1_0_1(n89_I1_0_1),
    .I1_0_2(n89_I1_0_2),
    .I1_1_0(n89_I1_1_0),
    .I1_1_1(n89_I1_1_1),
    .I1_1_2(n89_I1_1_2),
    .I1_2_0(n89_I1_2_0),
    .I1_2_1(n89_I1_2_1),
    .I1_2_2(n89_I1_2_2),
    .I1_3_0(n89_I1_3_0),
    .I1_3_1(n89_I1_3_1),
    .I1_3_2(n89_I1_3_2),
    .I1_4_0(n89_I1_4_0),
    .I1_4_1(n89_I1_4_1),
    .I1_4_2(n89_I1_4_2),
    .I1_5_0(n89_I1_5_0),
    .I1_5_1(n89_I1_5_1),
    .I1_5_2(n89_I1_5_2),
    .I1_6_0(n89_I1_6_0),
    .I1_6_1(n89_I1_6_1),
    .I1_6_2(n89_I1_6_2),
    .I1_7_0(n89_I1_7_0),
    .I1_7_1(n89_I1_7_1),
    .I1_7_2(n89_I1_7_2),
    .O_0_0_0(n89_O_0_0_0),
    .O_0_0_1(n89_O_0_0_1),
    .O_0_0_2(n89_O_0_0_2),
    .O_0_1_0(n89_O_0_1_0),
    .O_0_1_1(n89_O_0_1_1),
    .O_0_1_2(n89_O_0_1_2),
    .O_0_2_0(n89_O_0_2_0),
    .O_0_2_1(n89_O_0_2_1),
    .O_0_2_2(n89_O_0_2_2),
    .O_1_0_0(n89_O_1_0_0),
    .O_1_0_1(n89_O_1_0_1),
    .O_1_0_2(n89_O_1_0_2),
    .O_1_1_0(n89_O_1_1_0),
    .O_1_1_1(n89_O_1_1_1),
    .O_1_1_2(n89_O_1_1_2),
    .O_1_2_0(n89_O_1_2_0),
    .O_1_2_1(n89_O_1_2_1),
    .O_1_2_2(n89_O_1_2_2),
    .O_2_0_0(n89_O_2_0_0),
    .O_2_0_1(n89_O_2_0_1),
    .O_2_0_2(n89_O_2_0_2),
    .O_2_1_0(n89_O_2_1_0),
    .O_2_1_1(n89_O_2_1_1),
    .O_2_1_2(n89_O_2_1_2),
    .O_2_2_0(n89_O_2_2_0),
    .O_2_2_1(n89_O_2_2_1),
    .O_2_2_2(n89_O_2_2_2),
    .O_3_0_0(n89_O_3_0_0),
    .O_3_0_1(n89_O_3_0_1),
    .O_3_0_2(n89_O_3_0_2),
    .O_3_1_0(n89_O_3_1_0),
    .O_3_1_1(n89_O_3_1_1),
    .O_3_1_2(n89_O_3_1_2),
    .O_3_2_0(n89_O_3_2_0),
    .O_3_2_1(n89_O_3_2_1),
    .O_3_2_2(n89_O_3_2_2),
    .O_4_0_0(n89_O_4_0_0),
    .O_4_0_1(n89_O_4_0_1),
    .O_4_0_2(n89_O_4_0_2),
    .O_4_1_0(n89_O_4_1_0),
    .O_4_1_1(n89_O_4_1_1),
    .O_4_1_2(n89_O_4_1_2),
    .O_4_2_0(n89_O_4_2_0),
    .O_4_2_1(n89_O_4_2_1),
    .O_4_2_2(n89_O_4_2_2),
    .O_5_0_0(n89_O_5_0_0),
    .O_5_0_1(n89_O_5_0_1),
    .O_5_0_2(n89_O_5_0_2),
    .O_5_1_0(n89_O_5_1_0),
    .O_5_1_1(n89_O_5_1_1),
    .O_5_1_2(n89_O_5_1_2),
    .O_5_2_0(n89_O_5_2_0),
    .O_5_2_1(n89_O_5_2_1),
    .O_5_2_2(n89_O_5_2_2),
    .O_6_0_0(n89_O_6_0_0),
    .O_6_0_1(n89_O_6_0_1),
    .O_6_0_2(n89_O_6_0_2),
    .O_6_1_0(n89_O_6_1_0),
    .O_6_1_1(n89_O_6_1_1),
    .O_6_1_2(n89_O_6_1_2),
    .O_6_2_0(n89_O_6_2_0),
    .O_6_2_1(n89_O_6_2_1),
    .O_6_2_2(n89_O_6_2_2),
    .O_7_0_0(n89_O_7_0_0),
    .O_7_0_1(n89_O_7_0_1),
    .O_7_0_2(n89_O_7_0_2),
    .O_7_1_0(n89_O_7_1_0),
    .O_7_1_1(n89_O_7_1_1),
    .O_7_1_2(n89_O_7_1_2),
    .O_7_2_0(n89_O_7_2_0),
    .O_7_2_1(n89_O_7_2_1),
    .O_7_2_2(n89_O_7_2_2)
  );
  MapT_6 n98 ( // @[Top.scala 772:21]
    .valid_up(n98_valid_up),
    .valid_down(n98_valid_down),
    .I_0_0_0(n98_I_0_0_0),
    .I_0_0_1(n98_I_0_0_1),
    .I_0_0_2(n98_I_0_0_2),
    .I_0_1_0(n98_I_0_1_0),
    .I_0_1_1(n98_I_0_1_1),
    .I_0_1_2(n98_I_0_1_2),
    .I_0_2_0(n98_I_0_2_0),
    .I_0_2_1(n98_I_0_2_1),
    .I_0_2_2(n98_I_0_2_2),
    .I_1_0_0(n98_I_1_0_0),
    .I_1_0_1(n98_I_1_0_1),
    .I_1_0_2(n98_I_1_0_2),
    .I_1_1_0(n98_I_1_1_0),
    .I_1_1_1(n98_I_1_1_1),
    .I_1_1_2(n98_I_1_1_2),
    .I_1_2_0(n98_I_1_2_0),
    .I_1_2_1(n98_I_1_2_1),
    .I_1_2_2(n98_I_1_2_2),
    .I_2_0_0(n98_I_2_0_0),
    .I_2_0_1(n98_I_2_0_1),
    .I_2_0_2(n98_I_2_0_2),
    .I_2_1_0(n98_I_2_1_0),
    .I_2_1_1(n98_I_2_1_1),
    .I_2_1_2(n98_I_2_1_2),
    .I_2_2_0(n98_I_2_2_0),
    .I_2_2_1(n98_I_2_2_1),
    .I_2_2_2(n98_I_2_2_2),
    .I_3_0_0(n98_I_3_0_0),
    .I_3_0_1(n98_I_3_0_1),
    .I_3_0_2(n98_I_3_0_2),
    .I_3_1_0(n98_I_3_1_0),
    .I_3_1_1(n98_I_3_1_1),
    .I_3_1_2(n98_I_3_1_2),
    .I_3_2_0(n98_I_3_2_0),
    .I_3_2_1(n98_I_3_2_1),
    .I_3_2_2(n98_I_3_2_2),
    .I_4_0_0(n98_I_4_0_0),
    .I_4_0_1(n98_I_4_0_1),
    .I_4_0_2(n98_I_4_0_2),
    .I_4_1_0(n98_I_4_1_0),
    .I_4_1_1(n98_I_4_1_1),
    .I_4_1_2(n98_I_4_1_2),
    .I_4_2_0(n98_I_4_2_0),
    .I_4_2_1(n98_I_4_2_1),
    .I_4_2_2(n98_I_4_2_2),
    .I_5_0_0(n98_I_5_0_0),
    .I_5_0_1(n98_I_5_0_1),
    .I_5_0_2(n98_I_5_0_2),
    .I_5_1_0(n98_I_5_1_0),
    .I_5_1_1(n98_I_5_1_1),
    .I_5_1_2(n98_I_5_1_2),
    .I_5_2_0(n98_I_5_2_0),
    .I_5_2_1(n98_I_5_2_1),
    .I_5_2_2(n98_I_5_2_2),
    .I_6_0_0(n98_I_6_0_0),
    .I_6_0_1(n98_I_6_0_1),
    .I_6_0_2(n98_I_6_0_2),
    .I_6_1_0(n98_I_6_1_0),
    .I_6_1_1(n98_I_6_1_1),
    .I_6_1_2(n98_I_6_1_2),
    .I_6_2_0(n98_I_6_2_0),
    .I_6_2_1(n98_I_6_2_1),
    .I_6_2_2(n98_I_6_2_2),
    .I_7_0_0(n98_I_7_0_0),
    .I_7_0_1(n98_I_7_0_1),
    .I_7_0_2(n98_I_7_0_2),
    .I_7_1_0(n98_I_7_1_0),
    .I_7_1_1(n98_I_7_1_1),
    .I_7_1_2(n98_I_7_1_2),
    .I_7_2_0(n98_I_7_2_0),
    .I_7_2_1(n98_I_7_2_1),
    .I_7_2_2(n98_I_7_2_2),
    .O_0_0_0_0(n98_O_0_0_0_0),
    .O_0_0_0_1(n98_O_0_0_0_1),
    .O_0_0_0_2(n98_O_0_0_0_2),
    .O_0_0_1_0(n98_O_0_0_1_0),
    .O_0_0_1_1(n98_O_0_0_1_1),
    .O_0_0_1_2(n98_O_0_0_1_2),
    .O_0_0_2_0(n98_O_0_0_2_0),
    .O_0_0_2_1(n98_O_0_0_2_1),
    .O_0_0_2_2(n98_O_0_0_2_2),
    .O_1_0_0_0(n98_O_1_0_0_0),
    .O_1_0_0_1(n98_O_1_0_0_1),
    .O_1_0_0_2(n98_O_1_0_0_2),
    .O_1_0_1_0(n98_O_1_0_1_0),
    .O_1_0_1_1(n98_O_1_0_1_1),
    .O_1_0_1_2(n98_O_1_0_1_2),
    .O_1_0_2_0(n98_O_1_0_2_0),
    .O_1_0_2_1(n98_O_1_0_2_1),
    .O_1_0_2_2(n98_O_1_0_2_2),
    .O_2_0_0_0(n98_O_2_0_0_0),
    .O_2_0_0_1(n98_O_2_0_0_1),
    .O_2_0_0_2(n98_O_2_0_0_2),
    .O_2_0_1_0(n98_O_2_0_1_0),
    .O_2_0_1_1(n98_O_2_0_1_1),
    .O_2_0_1_2(n98_O_2_0_1_2),
    .O_2_0_2_0(n98_O_2_0_2_0),
    .O_2_0_2_1(n98_O_2_0_2_1),
    .O_2_0_2_2(n98_O_2_0_2_2),
    .O_3_0_0_0(n98_O_3_0_0_0),
    .O_3_0_0_1(n98_O_3_0_0_1),
    .O_3_0_0_2(n98_O_3_0_0_2),
    .O_3_0_1_0(n98_O_3_0_1_0),
    .O_3_0_1_1(n98_O_3_0_1_1),
    .O_3_0_1_2(n98_O_3_0_1_2),
    .O_3_0_2_0(n98_O_3_0_2_0),
    .O_3_0_2_1(n98_O_3_0_2_1),
    .O_3_0_2_2(n98_O_3_0_2_2),
    .O_4_0_0_0(n98_O_4_0_0_0),
    .O_4_0_0_1(n98_O_4_0_0_1),
    .O_4_0_0_2(n98_O_4_0_0_2),
    .O_4_0_1_0(n98_O_4_0_1_0),
    .O_4_0_1_1(n98_O_4_0_1_1),
    .O_4_0_1_2(n98_O_4_0_1_2),
    .O_4_0_2_0(n98_O_4_0_2_0),
    .O_4_0_2_1(n98_O_4_0_2_1),
    .O_4_0_2_2(n98_O_4_0_2_2),
    .O_5_0_0_0(n98_O_5_0_0_0),
    .O_5_0_0_1(n98_O_5_0_0_1),
    .O_5_0_0_2(n98_O_5_0_0_2),
    .O_5_0_1_0(n98_O_5_0_1_0),
    .O_5_0_1_1(n98_O_5_0_1_1),
    .O_5_0_1_2(n98_O_5_0_1_2),
    .O_5_0_2_0(n98_O_5_0_2_0),
    .O_5_0_2_1(n98_O_5_0_2_1),
    .O_5_0_2_2(n98_O_5_0_2_2),
    .O_6_0_0_0(n98_O_6_0_0_0),
    .O_6_0_0_1(n98_O_6_0_0_1),
    .O_6_0_0_2(n98_O_6_0_0_2),
    .O_6_0_1_0(n98_O_6_0_1_0),
    .O_6_0_1_1(n98_O_6_0_1_1),
    .O_6_0_1_2(n98_O_6_0_1_2),
    .O_6_0_2_0(n98_O_6_0_2_0),
    .O_6_0_2_1(n98_O_6_0_2_1),
    .O_6_0_2_2(n98_O_6_0_2_2),
    .O_7_0_0_0(n98_O_7_0_0_0),
    .O_7_0_0_1(n98_O_7_0_0_1),
    .O_7_0_0_2(n98_O_7_0_0_2),
    .O_7_0_1_0(n98_O_7_0_1_0),
    .O_7_0_1_1(n98_O_7_0_1_1),
    .O_7_0_1_2(n98_O_7_0_1_2),
    .O_7_0_2_0(n98_O_7_0_2_0),
    .O_7_0_2_1(n98_O_7_0_2_1),
    .O_7_0_2_2(n98_O_7_0_2_2)
  );
  MapT_7 n105 ( // @[Top.scala 775:22]
    .valid_up(n105_valid_up),
    .valid_down(n105_valid_down),
    .I_0_0_0_0(n105_I_0_0_0_0),
    .I_0_0_0_1(n105_I_0_0_0_1),
    .I_0_0_0_2(n105_I_0_0_0_2),
    .I_0_0_1_0(n105_I_0_0_1_0),
    .I_0_0_1_1(n105_I_0_0_1_1),
    .I_0_0_1_2(n105_I_0_0_1_2),
    .I_0_0_2_0(n105_I_0_0_2_0),
    .I_0_0_2_1(n105_I_0_0_2_1),
    .I_0_0_2_2(n105_I_0_0_2_2),
    .I_1_0_0_0(n105_I_1_0_0_0),
    .I_1_0_0_1(n105_I_1_0_0_1),
    .I_1_0_0_2(n105_I_1_0_0_2),
    .I_1_0_1_0(n105_I_1_0_1_0),
    .I_1_0_1_1(n105_I_1_0_1_1),
    .I_1_0_1_2(n105_I_1_0_1_2),
    .I_1_0_2_0(n105_I_1_0_2_0),
    .I_1_0_2_1(n105_I_1_0_2_1),
    .I_1_0_2_2(n105_I_1_0_2_2),
    .I_2_0_0_0(n105_I_2_0_0_0),
    .I_2_0_0_1(n105_I_2_0_0_1),
    .I_2_0_0_2(n105_I_2_0_0_2),
    .I_2_0_1_0(n105_I_2_0_1_0),
    .I_2_0_1_1(n105_I_2_0_1_1),
    .I_2_0_1_2(n105_I_2_0_1_2),
    .I_2_0_2_0(n105_I_2_0_2_0),
    .I_2_0_2_1(n105_I_2_0_2_1),
    .I_2_0_2_2(n105_I_2_0_2_2),
    .I_3_0_0_0(n105_I_3_0_0_0),
    .I_3_0_0_1(n105_I_3_0_0_1),
    .I_3_0_0_2(n105_I_3_0_0_2),
    .I_3_0_1_0(n105_I_3_0_1_0),
    .I_3_0_1_1(n105_I_3_0_1_1),
    .I_3_0_1_2(n105_I_3_0_1_2),
    .I_3_0_2_0(n105_I_3_0_2_0),
    .I_3_0_2_1(n105_I_3_0_2_1),
    .I_3_0_2_2(n105_I_3_0_2_2),
    .I_4_0_0_0(n105_I_4_0_0_0),
    .I_4_0_0_1(n105_I_4_0_0_1),
    .I_4_0_0_2(n105_I_4_0_0_2),
    .I_4_0_1_0(n105_I_4_0_1_0),
    .I_4_0_1_1(n105_I_4_0_1_1),
    .I_4_0_1_2(n105_I_4_0_1_2),
    .I_4_0_2_0(n105_I_4_0_2_0),
    .I_4_0_2_1(n105_I_4_0_2_1),
    .I_4_0_2_2(n105_I_4_0_2_2),
    .I_5_0_0_0(n105_I_5_0_0_0),
    .I_5_0_0_1(n105_I_5_0_0_1),
    .I_5_0_0_2(n105_I_5_0_0_2),
    .I_5_0_1_0(n105_I_5_0_1_0),
    .I_5_0_1_1(n105_I_5_0_1_1),
    .I_5_0_1_2(n105_I_5_0_1_2),
    .I_5_0_2_0(n105_I_5_0_2_0),
    .I_5_0_2_1(n105_I_5_0_2_1),
    .I_5_0_2_2(n105_I_5_0_2_2),
    .I_6_0_0_0(n105_I_6_0_0_0),
    .I_6_0_0_1(n105_I_6_0_0_1),
    .I_6_0_0_2(n105_I_6_0_0_2),
    .I_6_0_1_0(n105_I_6_0_1_0),
    .I_6_0_1_1(n105_I_6_0_1_1),
    .I_6_0_1_2(n105_I_6_0_1_2),
    .I_6_0_2_0(n105_I_6_0_2_0),
    .I_6_0_2_1(n105_I_6_0_2_1),
    .I_6_0_2_2(n105_I_6_0_2_2),
    .I_7_0_0_0(n105_I_7_0_0_0),
    .I_7_0_0_1(n105_I_7_0_0_1),
    .I_7_0_0_2(n105_I_7_0_0_2),
    .I_7_0_1_0(n105_I_7_0_1_0),
    .I_7_0_1_1(n105_I_7_0_1_1),
    .I_7_0_1_2(n105_I_7_0_1_2),
    .I_7_0_2_0(n105_I_7_0_2_0),
    .I_7_0_2_1(n105_I_7_0_2_1),
    .I_7_0_2_2(n105_I_7_0_2_2),
    .O_0_0_0(n105_O_0_0_0),
    .O_0_0_1(n105_O_0_0_1),
    .O_0_0_2(n105_O_0_0_2),
    .O_0_1_0(n105_O_0_1_0),
    .O_0_1_1(n105_O_0_1_1),
    .O_0_1_2(n105_O_0_1_2),
    .O_0_2_0(n105_O_0_2_0),
    .O_0_2_1(n105_O_0_2_1),
    .O_0_2_2(n105_O_0_2_2),
    .O_1_0_0(n105_O_1_0_0),
    .O_1_0_1(n105_O_1_0_1),
    .O_1_0_2(n105_O_1_0_2),
    .O_1_1_0(n105_O_1_1_0),
    .O_1_1_1(n105_O_1_1_1),
    .O_1_1_2(n105_O_1_1_2),
    .O_1_2_0(n105_O_1_2_0),
    .O_1_2_1(n105_O_1_2_1),
    .O_1_2_2(n105_O_1_2_2),
    .O_2_0_0(n105_O_2_0_0),
    .O_2_0_1(n105_O_2_0_1),
    .O_2_0_2(n105_O_2_0_2),
    .O_2_1_0(n105_O_2_1_0),
    .O_2_1_1(n105_O_2_1_1),
    .O_2_1_2(n105_O_2_1_2),
    .O_2_2_0(n105_O_2_2_0),
    .O_2_2_1(n105_O_2_2_1),
    .O_2_2_2(n105_O_2_2_2),
    .O_3_0_0(n105_O_3_0_0),
    .O_3_0_1(n105_O_3_0_1),
    .O_3_0_2(n105_O_3_0_2),
    .O_3_1_0(n105_O_3_1_0),
    .O_3_1_1(n105_O_3_1_1),
    .O_3_1_2(n105_O_3_1_2),
    .O_3_2_0(n105_O_3_2_0),
    .O_3_2_1(n105_O_3_2_1),
    .O_3_2_2(n105_O_3_2_2),
    .O_4_0_0(n105_O_4_0_0),
    .O_4_0_1(n105_O_4_0_1),
    .O_4_0_2(n105_O_4_0_2),
    .O_4_1_0(n105_O_4_1_0),
    .O_4_1_1(n105_O_4_1_1),
    .O_4_1_2(n105_O_4_1_2),
    .O_4_2_0(n105_O_4_2_0),
    .O_4_2_1(n105_O_4_2_1),
    .O_4_2_2(n105_O_4_2_2),
    .O_5_0_0(n105_O_5_0_0),
    .O_5_0_1(n105_O_5_0_1),
    .O_5_0_2(n105_O_5_0_2),
    .O_5_1_0(n105_O_5_1_0),
    .O_5_1_1(n105_O_5_1_1),
    .O_5_1_2(n105_O_5_1_2),
    .O_5_2_0(n105_O_5_2_0),
    .O_5_2_1(n105_O_5_2_1),
    .O_5_2_2(n105_O_5_2_2),
    .O_6_0_0(n105_O_6_0_0),
    .O_6_0_1(n105_O_6_0_1),
    .O_6_0_2(n105_O_6_0_2),
    .O_6_1_0(n105_O_6_1_0),
    .O_6_1_1(n105_O_6_1_1),
    .O_6_1_2(n105_O_6_1_2),
    .O_6_2_0(n105_O_6_2_0),
    .O_6_2_1(n105_O_6_2_1),
    .O_6_2_2(n105_O_6_2_2),
    .O_7_0_0(n105_O_7_0_0),
    .O_7_0_1(n105_O_7_0_1),
    .O_7_0_2(n105_O_7_0_2),
    .O_7_1_0(n105_O_7_1_0),
    .O_7_1_1(n105_O_7_1_1),
    .O_7_1_2(n105_O_7_1_2),
    .O_7_2_0(n105_O_7_2_0),
    .O_7_2_1(n105_O_7_2_1),
    .O_7_2_2(n105_O_7_2_2)
  );
  Passthrough n106 ( // @[Top.scala 778:22]
    .valid_up(n106_valid_up),
    .valid_down(n106_valid_down),
    .I_0_0_0(n106_I_0_0_0),
    .I_0_0_1(n106_I_0_0_1),
    .I_0_0_2(n106_I_0_0_2),
    .I_0_1_0(n106_I_0_1_0),
    .I_0_1_1(n106_I_0_1_1),
    .I_0_1_2(n106_I_0_1_2),
    .I_0_2_0(n106_I_0_2_0),
    .I_0_2_1(n106_I_0_2_1),
    .I_0_2_2(n106_I_0_2_2),
    .I_1_0_0(n106_I_1_0_0),
    .I_1_0_1(n106_I_1_0_1),
    .I_1_0_2(n106_I_1_0_2),
    .I_1_1_0(n106_I_1_1_0),
    .I_1_1_1(n106_I_1_1_1),
    .I_1_1_2(n106_I_1_1_2),
    .I_1_2_0(n106_I_1_2_0),
    .I_1_2_1(n106_I_1_2_1),
    .I_1_2_2(n106_I_1_2_2),
    .I_2_0_0(n106_I_2_0_0),
    .I_2_0_1(n106_I_2_0_1),
    .I_2_0_2(n106_I_2_0_2),
    .I_2_1_0(n106_I_2_1_0),
    .I_2_1_1(n106_I_2_1_1),
    .I_2_1_2(n106_I_2_1_2),
    .I_2_2_0(n106_I_2_2_0),
    .I_2_2_1(n106_I_2_2_1),
    .I_2_2_2(n106_I_2_2_2),
    .I_3_0_0(n106_I_3_0_0),
    .I_3_0_1(n106_I_3_0_1),
    .I_3_0_2(n106_I_3_0_2),
    .I_3_1_0(n106_I_3_1_0),
    .I_3_1_1(n106_I_3_1_1),
    .I_3_1_2(n106_I_3_1_2),
    .I_3_2_0(n106_I_3_2_0),
    .I_3_2_1(n106_I_3_2_1),
    .I_3_2_2(n106_I_3_2_2),
    .I_4_0_0(n106_I_4_0_0),
    .I_4_0_1(n106_I_4_0_1),
    .I_4_0_2(n106_I_4_0_2),
    .I_4_1_0(n106_I_4_1_0),
    .I_4_1_1(n106_I_4_1_1),
    .I_4_1_2(n106_I_4_1_2),
    .I_4_2_0(n106_I_4_2_0),
    .I_4_2_1(n106_I_4_2_1),
    .I_4_2_2(n106_I_4_2_2),
    .I_5_0_0(n106_I_5_0_0),
    .I_5_0_1(n106_I_5_0_1),
    .I_5_0_2(n106_I_5_0_2),
    .I_5_1_0(n106_I_5_1_0),
    .I_5_1_1(n106_I_5_1_1),
    .I_5_1_2(n106_I_5_1_2),
    .I_5_2_0(n106_I_5_2_0),
    .I_5_2_1(n106_I_5_2_1),
    .I_5_2_2(n106_I_5_2_2),
    .I_6_0_0(n106_I_6_0_0),
    .I_6_0_1(n106_I_6_0_1),
    .I_6_0_2(n106_I_6_0_2),
    .I_6_1_0(n106_I_6_1_0),
    .I_6_1_1(n106_I_6_1_1),
    .I_6_1_2(n106_I_6_1_2),
    .I_6_2_0(n106_I_6_2_0),
    .I_6_2_1(n106_I_6_2_1),
    .I_6_2_2(n106_I_6_2_2),
    .I_7_0_0(n106_I_7_0_0),
    .I_7_0_1(n106_I_7_0_1),
    .I_7_0_2(n106_I_7_0_2),
    .I_7_1_0(n106_I_7_1_0),
    .I_7_1_1(n106_I_7_1_1),
    .I_7_1_2(n106_I_7_1_2),
    .I_7_2_0(n106_I_7_2_0),
    .I_7_2_1(n106_I_7_2_1),
    .I_7_2_2(n106_I_7_2_2),
    .O_0_0_0(n106_O_0_0_0),
    .O_0_0_1(n106_O_0_0_1),
    .O_0_0_2(n106_O_0_0_2),
    .O_0_1_0(n106_O_0_1_0),
    .O_0_1_1(n106_O_0_1_1),
    .O_0_1_2(n106_O_0_1_2),
    .O_0_2_0(n106_O_0_2_0),
    .O_0_2_1(n106_O_0_2_1),
    .O_0_2_2(n106_O_0_2_2),
    .O_1_0_0(n106_O_1_0_0),
    .O_1_0_1(n106_O_1_0_1),
    .O_1_0_2(n106_O_1_0_2),
    .O_1_1_0(n106_O_1_1_0),
    .O_1_1_1(n106_O_1_1_1),
    .O_1_1_2(n106_O_1_1_2),
    .O_1_2_0(n106_O_1_2_0),
    .O_1_2_1(n106_O_1_2_1),
    .O_1_2_2(n106_O_1_2_2),
    .O_2_0_0(n106_O_2_0_0),
    .O_2_0_1(n106_O_2_0_1),
    .O_2_0_2(n106_O_2_0_2),
    .O_2_1_0(n106_O_2_1_0),
    .O_2_1_1(n106_O_2_1_1),
    .O_2_1_2(n106_O_2_1_2),
    .O_2_2_0(n106_O_2_2_0),
    .O_2_2_1(n106_O_2_2_1),
    .O_2_2_2(n106_O_2_2_2),
    .O_3_0_0(n106_O_3_0_0),
    .O_3_0_1(n106_O_3_0_1),
    .O_3_0_2(n106_O_3_0_2),
    .O_3_1_0(n106_O_3_1_0),
    .O_3_1_1(n106_O_3_1_1),
    .O_3_1_2(n106_O_3_1_2),
    .O_3_2_0(n106_O_3_2_0),
    .O_3_2_1(n106_O_3_2_1),
    .O_3_2_2(n106_O_3_2_2),
    .O_4_0_0(n106_O_4_0_0),
    .O_4_0_1(n106_O_4_0_1),
    .O_4_0_2(n106_O_4_0_2),
    .O_4_1_0(n106_O_4_1_0),
    .O_4_1_1(n106_O_4_1_1),
    .O_4_1_2(n106_O_4_1_2),
    .O_4_2_0(n106_O_4_2_0),
    .O_4_2_1(n106_O_4_2_1),
    .O_4_2_2(n106_O_4_2_2),
    .O_5_0_0(n106_O_5_0_0),
    .O_5_0_1(n106_O_5_0_1),
    .O_5_0_2(n106_O_5_0_2),
    .O_5_1_0(n106_O_5_1_0),
    .O_5_1_1(n106_O_5_1_1),
    .O_5_1_2(n106_O_5_1_2),
    .O_5_2_0(n106_O_5_2_0),
    .O_5_2_1(n106_O_5_2_1),
    .O_5_2_2(n106_O_5_2_2),
    .O_6_0_0(n106_O_6_0_0),
    .O_6_0_1(n106_O_6_0_1),
    .O_6_0_2(n106_O_6_0_2),
    .O_6_1_0(n106_O_6_1_0),
    .O_6_1_1(n106_O_6_1_1),
    .O_6_1_2(n106_O_6_1_2),
    .O_6_2_0(n106_O_6_2_0),
    .O_6_2_1(n106_O_6_2_1),
    .O_6_2_2(n106_O_6_2_2),
    .O_7_0_0(n106_O_7_0_0),
    .O_7_0_1(n106_O_7_0_1),
    .O_7_0_2(n106_O_7_0_2),
    .O_7_1_0(n106_O_7_1_0),
    .O_7_1_1(n106_O_7_1_1),
    .O_7_1_2(n106_O_7_1_2),
    .O_7_2_0(n106_O_7_2_0),
    .O_7_2_1(n106_O_7_2_1),
    .O_7_2_2(n106_O_7_2_2)
  );
  MapT_12 n443 ( // @[Top.scala 781:22]
    .clock(n443_clock),
    .reset(n443_reset),
    .valid_up(n443_valid_up),
    .valid_down(n443_valid_down),
    .I_0_0_0(n443_I_0_0_0),
    .I_0_0_1(n443_I_0_0_1),
    .I_0_0_2(n443_I_0_0_2),
    .I_0_1_0(n443_I_0_1_0),
    .I_0_1_1(n443_I_0_1_1),
    .I_0_1_2(n443_I_0_1_2),
    .I_0_2_0(n443_I_0_2_0),
    .I_0_2_1(n443_I_0_2_1),
    .I_0_2_2(n443_I_0_2_2),
    .I_1_0_0(n443_I_1_0_0),
    .I_1_0_1(n443_I_1_0_1),
    .I_1_0_2(n443_I_1_0_2),
    .I_1_1_0(n443_I_1_1_0),
    .I_1_1_1(n443_I_1_1_1),
    .I_1_1_2(n443_I_1_1_2),
    .I_1_2_0(n443_I_1_2_0),
    .I_1_2_1(n443_I_1_2_1),
    .I_1_2_2(n443_I_1_2_2),
    .I_2_0_0(n443_I_2_0_0),
    .I_2_0_1(n443_I_2_0_1),
    .I_2_0_2(n443_I_2_0_2),
    .I_2_1_0(n443_I_2_1_0),
    .I_2_1_1(n443_I_2_1_1),
    .I_2_1_2(n443_I_2_1_2),
    .I_2_2_0(n443_I_2_2_0),
    .I_2_2_1(n443_I_2_2_1),
    .I_2_2_2(n443_I_2_2_2),
    .I_3_0_0(n443_I_3_0_0),
    .I_3_0_1(n443_I_3_0_1),
    .I_3_0_2(n443_I_3_0_2),
    .I_3_1_0(n443_I_3_1_0),
    .I_3_1_1(n443_I_3_1_1),
    .I_3_1_2(n443_I_3_1_2),
    .I_3_2_0(n443_I_3_2_0),
    .I_3_2_1(n443_I_3_2_1),
    .I_3_2_2(n443_I_3_2_2),
    .I_4_0_0(n443_I_4_0_0),
    .I_4_0_1(n443_I_4_0_1),
    .I_4_0_2(n443_I_4_0_2),
    .I_4_1_0(n443_I_4_1_0),
    .I_4_1_1(n443_I_4_1_1),
    .I_4_1_2(n443_I_4_1_2),
    .I_4_2_0(n443_I_4_2_0),
    .I_4_2_1(n443_I_4_2_1),
    .I_4_2_2(n443_I_4_2_2),
    .I_5_0_0(n443_I_5_0_0),
    .I_5_0_1(n443_I_5_0_1),
    .I_5_0_2(n443_I_5_0_2),
    .I_5_1_0(n443_I_5_1_0),
    .I_5_1_1(n443_I_5_1_1),
    .I_5_1_2(n443_I_5_1_2),
    .I_5_2_0(n443_I_5_2_0),
    .I_5_2_1(n443_I_5_2_1),
    .I_5_2_2(n443_I_5_2_2),
    .I_6_0_0(n443_I_6_0_0),
    .I_6_0_1(n443_I_6_0_1),
    .I_6_0_2(n443_I_6_0_2),
    .I_6_1_0(n443_I_6_1_0),
    .I_6_1_1(n443_I_6_1_1),
    .I_6_1_2(n443_I_6_1_2),
    .I_6_2_0(n443_I_6_2_0),
    .I_6_2_1(n443_I_6_2_1),
    .I_6_2_2(n443_I_6_2_2),
    .I_7_0_0(n443_I_7_0_0),
    .I_7_0_1(n443_I_7_0_1),
    .I_7_0_2(n443_I_7_0_2),
    .I_7_1_0(n443_I_7_1_0),
    .I_7_1_1(n443_I_7_1_1),
    .I_7_1_2(n443_I_7_1_2),
    .I_7_2_0(n443_I_7_2_0),
    .I_7_2_1(n443_I_7_2_1),
    .I_7_2_2(n443_I_7_2_2),
    .O_0_0_0_t0b(n443_O_0_0_0_t0b),
    .O_0_0_0_t1b_t0b(n443_O_0_0_0_t1b_t0b),
    .O_0_0_0_t1b_t1b(n443_O_0_0_0_t1b_t1b),
    .O_1_0_0_t0b(n443_O_1_0_0_t0b),
    .O_1_0_0_t1b_t0b(n443_O_1_0_0_t1b_t0b),
    .O_1_0_0_t1b_t1b(n443_O_1_0_0_t1b_t1b),
    .O_2_0_0_t0b(n443_O_2_0_0_t0b),
    .O_2_0_0_t1b_t0b(n443_O_2_0_0_t1b_t0b),
    .O_2_0_0_t1b_t1b(n443_O_2_0_0_t1b_t1b),
    .O_3_0_0_t0b(n443_O_3_0_0_t0b),
    .O_3_0_0_t1b_t0b(n443_O_3_0_0_t1b_t0b),
    .O_3_0_0_t1b_t1b(n443_O_3_0_0_t1b_t1b),
    .O_4_0_0_t0b(n443_O_4_0_0_t0b),
    .O_4_0_0_t1b_t0b(n443_O_4_0_0_t1b_t0b),
    .O_4_0_0_t1b_t1b(n443_O_4_0_0_t1b_t1b),
    .O_5_0_0_t0b(n443_O_5_0_0_t0b),
    .O_5_0_0_t1b_t0b(n443_O_5_0_0_t1b_t0b),
    .O_5_0_0_t1b_t1b(n443_O_5_0_0_t1b_t1b),
    .O_6_0_0_t0b(n443_O_6_0_0_t0b),
    .O_6_0_0_t1b_t0b(n443_O_6_0_0_t1b_t0b),
    .O_6_0_0_t1b_t1b(n443_O_6_0_0_t1b_t1b),
    .O_7_0_0_t0b(n443_O_7_0_0_t0b),
    .O_7_0_0_t1b_t0b(n443_O_7_0_0_t1b_t0b),
    .O_7_0_0_t1b_t1b(n443_O_7_0_0_t1b_t1b)
  );
  Passthrough_1 n444 ( // @[Top.scala 784:22]
    .valid_up(n444_valid_up),
    .valid_down(n444_valid_down),
    .I_0_0_0_t0b(n444_I_0_0_0_t0b),
    .I_0_0_0_t1b_t0b(n444_I_0_0_0_t1b_t0b),
    .I_0_0_0_t1b_t1b(n444_I_0_0_0_t1b_t1b),
    .I_1_0_0_t0b(n444_I_1_0_0_t0b),
    .I_1_0_0_t1b_t0b(n444_I_1_0_0_t1b_t0b),
    .I_1_0_0_t1b_t1b(n444_I_1_0_0_t1b_t1b),
    .I_2_0_0_t0b(n444_I_2_0_0_t0b),
    .I_2_0_0_t1b_t0b(n444_I_2_0_0_t1b_t0b),
    .I_2_0_0_t1b_t1b(n444_I_2_0_0_t1b_t1b),
    .I_3_0_0_t0b(n444_I_3_0_0_t0b),
    .I_3_0_0_t1b_t0b(n444_I_3_0_0_t1b_t0b),
    .I_3_0_0_t1b_t1b(n444_I_3_0_0_t1b_t1b),
    .I_4_0_0_t0b(n444_I_4_0_0_t0b),
    .I_4_0_0_t1b_t0b(n444_I_4_0_0_t1b_t0b),
    .I_4_0_0_t1b_t1b(n444_I_4_0_0_t1b_t1b),
    .I_5_0_0_t0b(n444_I_5_0_0_t0b),
    .I_5_0_0_t1b_t0b(n444_I_5_0_0_t1b_t0b),
    .I_5_0_0_t1b_t1b(n444_I_5_0_0_t1b_t1b),
    .I_6_0_0_t0b(n444_I_6_0_0_t0b),
    .I_6_0_0_t1b_t0b(n444_I_6_0_0_t1b_t0b),
    .I_6_0_0_t1b_t1b(n444_I_6_0_0_t1b_t1b),
    .I_7_0_0_t0b(n444_I_7_0_0_t0b),
    .I_7_0_0_t1b_t0b(n444_I_7_0_0_t1b_t0b),
    .I_7_0_0_t1b_t1b(n444_I_7_0_0_t1b_t1b),
    .O_0_0_0_t0b(n444_O_0_0_0_t0b),
    .O_0_0_0_t1b_t0b(n444_O_0_0_0_t1b_t0b),
    .O_0_0_0_t1b_t1b(n444_O_0_0_0_t1b_t1b),
    .O_1_0_0_t0b(n444_O_1_0_0_t0b),
    .O_1_0_0_t1b_t0b(n444_O_1_0_0_t1b_t0b),
    .O_1_0_0_t1b_t1b(n444_O_1_0_0_t1b_t1b),
    .O_2_0_0_t0b(n444_O_2_0_0_t0b),
    .O_2_0_0_t1b_t0b(n444_O_2_0_0_t1b_t0b),
    .O_2_0_0_t1b_t1b(n444_O_2_0_0_t1b_t1b),
    .O_3_0_0_t0b(n444_O_3_0_0_t0b),
    .O_3_0_0_t1b_t0b(n444_O_3_0_0_t1b_t0b),
    .O_3_0_0_t1b_t1b(n444_O_3_0_0_t1b_t1b),
    .O_4_0_0_t0b(n444_O_4_0_0_t0b),
    .O_4_0_0_t1b_t0b(n444_O_4_0_0_t1b_t0b),
    .O_4_0_0_t1b_t1b(n444_O_4_0_0_t1b_t1b),
    .O_5_0_0_t0b(n444_O_5_0_0_t0b),
    .O_5_0_0_t1b_t0b(n444_O_5_0_0_t1b_t0b),
    .O_5_0_0_t1b_t1b(n444_O_5_0_0_t1b_t1b),
    .O_6_0_0_t0b(n444_O_6_0_0_t0b),
    .O_6_0_0_t1b_t0b(n444_O_6_0_0_t1b_t0b),
    .O_6_0_0_t1b_t1b(n444_O_6_0_0_t1b_t1b),
    .O_7_0_0_t0b(n444_O_7_0_0_t0b),
    .O_7_0_0_t1b_t0b(n444_O_7_0_0_t1b_t0b),
    .O_7_0_0_t1b_t1b(n444_O_7_0_0_t1b_t1b)
  );
  Passthrough_2 n445 ( // @[Top.scala 787:22]
    .valid_up(n445_valid_up),
    .valid_down(n445_valid_down),
    .I_0_0_0_t0b(n445_I_0_0_0_t0b),
    .I_0_0_0_t1b_t0b(n445_I_0_0_0_t1b_t0b),
    .I_0_0_0_t1b_t1b(n445_I_0_0_0_t1b_t1b),
    .I_1_0_0_t0b(n445_I_1_0_0_t0b),
    .I_1_0_0_t1b_t0b(n445_I_1_0_0_t1b_t0b),
    .I_1_0_0_t1b_t1b(n445_I_1_0_0_t1b_t1b),
    .I_2_0_0_t0b(n445_I_2_0_0_t0b),
    .I_2_0_0_t1b_t0b(n445_I_2_0_0_t1b_t0b),
    .I_2_0_0_t1b_t1b(n445_I_2_0_0_t1b_t1b),
    .I_3_0_0_t0b(n445_I_3_0_0_t0b),
    .I_3_0_0_t1b_t0b(n445_I_3_0_0_t1b_t0b),
    .I_3_0_0_t1b_t1b(n445_I_3_0_0_t1b_t1b),
    .I_4_0_0_t0b(n445_I_4_0_0_t0b),
    .I_4_0_0_t1b_t0b(n445_I_4_0_0_t1b_t0b),
    .I_4_0_0_t1b_t1b(n445_I_4_0_0_t1b_t1b),
    .I_5_0_0_t0b(n445_I_5_0_0_t0b),
    .I_5_0_0_t1b_t0b(n445_I_5_0_0_t1b_t0b),
    .I_5_0_0_t1b_t1b(n445_I_5_0_0_t1b_t1b),
    .I_6_0_0_t0b(n445_I_6_0_0_t0b),
    .I_6_0_0_t1b_t0b(n445_I_6_0_0_t1b_t0b),
    .I_6_0_0_t1b_t1b(n445_I_6_0_0_t1b_t1b),
    .I_7_0_0_t0b(n445_I_7_0_0_t0b),
    .I_7_0_0_t1b_t0b(n445_I_7_0_0_t1b_t0b),
    .I_7_0_0_t1b_t1b(n445_I_7_0_0_t1b_t1b),
    .O_0_0_t0b(n445_O_0_0_t0b),
    .O_0_0_t1b_t0b(n445_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(n445_O_0_0_t1b_t1b),
    .O_1_0_t0b(n445_O_1_0_t0b),
    .O_1_0_t1b_t0b(n445_O_1_0_t1b_t0b),
    .O_1_0_t1b_t1b(n445_O_1_0_t1b_t1b),
    .O_2_0_t0b(n445_O_2_0_t0b),
    .O_2_0_t1b_t0b(n445_O_2_0_t1b_t0b),
    .O_2_0_t1b_t1b(n445_O_2_0_t1b_t1b),
    .O_3_0_t0b(n445_O_3_0_t0b),
    .O_3_0_t1b_t0b(n445_O_3_0_t1b_t0b),
    .O_3_0_t1b_t1b(n445_O_3_0_t1b_t1b),
    .O_4_0_t0b(n445_O_4_0_t0b),
    .O_4_0_t1b_t0b(n445_O_4_0_t1b_t0b),
    .O_4_0_t1b_t1b(n445_O_4_0_t1b_t1b),
    .O_5_0_t0b(n445_O_5_0_t0b),
    .O_5_0_t1b_t0b(n445_O_5_0_t1b_t0b),
    .O_5_0_t1b_t1b(n445_O_5_0_t1b_t1b),
    .O_6_0_t0b(n445_O_6_0_t0b),
    .O_6_0_t1b_t0b(n445_O_6_0_t1b_t0b),
    .O_6_0_t1b_t1b(n445_O_6_0_t1b_t1b),
    .O_7_0_t0b(n445_O_7_0_t0b),
    .O_7_0_t1b_t0b(n445_O_7_0_t1b_t0b),
    .O_7_0_t1b_t1b(n445_O_7_0_t1b_t1b)
  );
  Passthrough_3 n446 ( // @[Top.scala 790:22]
    .valid_up(n446_valid_up),
    .valid_down(n446_valid_down),
    .I_0_0_t0b(n446_I_0_0_t0b),
    .I_0_0_t1b_t0b(n446_I_0_0_t1b_t0b),
    .I_0_0_t1b_t1b(n446_I_0_0_t1b_t1b),
    .I_1_0_t0b(n446_I_1_0_t0b),
    .I_1_0_t1b_t0b(n446_I_1_0_t1b_t0b),
    .I_1_0_t1b_t1b(n446_I_1_0_t1b_t1b),
    .I_2_0_t0b(n446_I_2_0_t0b),
    .I_2_0_t1b_t0b(n446_I_2_0_t1b_t0b),
    .I_2_0_t1b_t1b(n446_I_2_0_t1b_t1b),
    .I_3_0_t0b(n446_I_3_0_t0b),
    .I_3_0_t1b_t0b(n446_I_3_0_t1b_t0b),
    .I_3_0_t1b_t1b(n446_I_3_0_t1b_t1b),
    .I_4_0_t0b(n446_I_4_0_t0b),
    .I_4_0_t1b_t0b(n446_I_4_0_t1b_t0b),
    .I_4_0_t1b_t1b(n446_I_4_0_t1b_t1b),
    .I_5_0_t0b(n446_I_5_0_t0b),
    .I_5_0_t1b_t0b(n446_I_5_0_t1b_t0b),
    .I_5_0_t1b_t1b(n446_I_5_0_t1b_t1b),
    .I_6_0_t0b(n446_I_6_0_t0b),
    .I_6_0_t1b_t0b(n446_I_6_0_t1b_t0b),
    .I_6_0_t1b_t1b(n446_I_6_0_t1b_t1b),
    .I_7_0_t0b(n446_I_7_0_t0b),
    .I_7_0_t1b_t0b(n446_I_7_0_t1b_t0b),
    .I_7_0_t1b_t1b(n446_I_7_0_t1b_t1b),
    .O_0_t0b(n446_O_0_t0b),
    .O_0_t1b_t0b(n446_O_0_t1b_t0b),
    .O_0_t1b_t1b(n446_O_0_t1b_t1b),
    .O_1_t0b(n446_O_1_t0b),
    .O_1_t1b_t0b(n446_O_1_t1b_t0b),
    .O_1_t1b_t1b(n446_O_1_t1b_t1b),
    .O_2_t0b(n446_O_2_t0b),
    .O_2_t1b_t0b(n446_O_2_t1b_t0b),
    .O_2_t1b_t1b(n446_O_2_t1b_t1b),
    .O_3_t0b(n446_O_3_t0b),
    .O_3_t1b_t0b(n446_O_3_t1b_t0b),
    .O_3_t1b_t1b(n446_O_3_t1b_t1b),
    .O_4_t0b(n446_O_4_t0b),
    .O_4_t1b_t0b(n446_O_4_t1b_t0b),
    .O_4_t1b_t1b(n446_O_4_t1b_t1b),
    .O_5_t0b(n446_O_5_t0b),
    .O_5_t1b_t0b(n446_O_5_t1b_t0b),
    .O_5_t1b_t1b(n446_O_5_t1b_t1b),
    .O_6_t0b(n446_O_6_t0b),
    .O_6_t1b_t0b(n446_O_6_t1b_t0b),
    .O_6_t1b_t1b(n446_O_6_t1b_t1b),
    .O_7_t0b(n446_O_7_t0b),
    .O_7_t1b_t0b(n446_O_7_t1b_t0b),
    .O_7_t1b_t1b(n446_O_7_t1b_t1b)
  );
  MapT_13 n451 ( // @[Top.scala 793:22]
    .valid_up(n451_valid_up),
    .valid_down(n451_valid_down),
    .I_0_t0b(n451_I_0_t0b),
    .I_1_t0b(n451_I_1_t0b),
    .I_2_t0b(n451_I_2_t0b),
    .I_3_t0b(n451_I_3_t0b),
    .I_4_t0b(n451_I_4_t0b),
    .I_5_t0b(n451_I_5_t0b),
    .I_6_t0b(n451_I_6_t0b),
    .I_7_t0b(n451_I_7_t0b),
    .O_0(n451_O_0),
    .O_1(n451_O_1),
    .O_2(n451_O_2),
    .O_3(n451_O_3),
    .O_4(n451_O_4),
    .O_5(n451_O_5),
    .O_6(n451_O_6),
    .O_7(n451_O_7)
  );
  ShiftTS n452 ( // @[Top.scala 796:22]
    .clock(n452_clock),
    .reset(n452_reset),
    .valid_up(n452_valid_up),
    .valid_down(n452_valid_down),
    .I_0(n452_I_0),
    .I_1(n452_I_1),
    .I_2(n452_I_2),
    .I_3(n452_I_3),
    .I_4(n452_I_4),
    .I_5(n452_I_5),
    .I_6(n452_I_6),
    .I_7(n452_I_7),
    .O_0(n452_O_0),
    .O_1(n452_O_1),
    .O_2(n452_O_2),
    .O_3(n452_O_3),
    .O_4(n452_O_4),
    .O_5(n452_O_5),
    .O_6(n452_O_6),
    .O_7(n452_O_7)
  );
  ShiftTS n453 ( // @[Top.scala 799:22]
    .clock(n453_clock),
    .reset(n453_reset),
    .valid_up(n453_valid_up),
    .valid_down(n453_valid_down),
    .I_0(n453_I_0),
    .I_1(n453_I_1),
    .I_2(n453_I_2),
    .I_3(n453_I_3),
    .I_4(n453_I_4),
    .I_5(n453_I_5),
    .I_6(n453_I_6),
    .I_7(n453_I_7),
    .O_0(n453_O_0),
    .O_1(n453_O_1),
    .O_2(n453_O_2),
    .O_3(n453_O_3),
    .O_4(n453_O_4),
    .O_5(n453_O_5),
    .O_6(n453_O_6),
    .O_7(n453_O_7)
  );
  ShiftTS_2 n454 ( // @[Top.scala 802:22]
    .clock(n454_clock),
    .valid_up(n454_valid_up),
    .valid_down(n454_valid_down),
    .I_0(n454_I_0),
    .I_1(n454_I_1),
    .I_2(n454_I_2),
    .I_3(n454_I_3),
    .I_4(n454_I_4),
    .I_5(n454_I_5),
    .I_6(n454_I_6),
    .I_7(n454_I_7),
    .O_0(n454_O_0),
    .O_1(n454_O_1),
    .O_2(n454_O_2),
    .O_3(n454_O_3),
    .O_4(n454_O_4),
    .O_5(n454_O_5),
    .O_6(n454_O_6),
    .O_7(n454_O_7)
  );
  ShiftTS_2 n455 ( // @[Top.scala 805:22]
    .clock(n455_clock),
    .valid_up(n455_valid_up),
    .valid_down(n455_valid_down),
    .I_0(n455_I_0),
    .I_1(n455_I_1),
    .I_2(n455_I_2),
    .I_3(n455_I_3),
    .I_4(n455_I_4),
    .I_5(n455_I_5),
    .I_6(n455_I_6),
    .I_7(n455_I_7),
    .O_0(n455_O_0),
    .O_1(n455_O_1),
    .O_2(n455_O_2),
    .O_3(n455_O_3),
    .O_4(n455_O_4),
    .O_5(n455_O_5),
    .O_6(n455_O_6),
    .O_7(n455_O_7)
  );
  Map2T n456 ( // @[Top.scala 808:22]
    .valid_up(n456_valid_up),
    .valid_down(n456_valid_down),
    .I0_0(n456_I0_0),
    .I0_1(n456_I0_1),
    .I0_2(n456_I0_2),
    .I0_3(n456_I0_3),
    .I0_4(n456_I0_4),
    .I0_5(n456_I0_5),
    .I0_6(n456_I0_6),
    .I0_7(n456_I0_7),
    .I1_0(n456_I1_0),
    .I1_1(n456_I1_1),
    .I1_2(n456_I1_2),
    .I1_3(n456_I1_3),
    .I1_4(n456_I1_4),
    .I1_5(n456_I1_5),
    .I1_6(n456_I1_6),
    .I1_7(n456_I1_7),
    .O_0_0(n456_O_0_0),
    .O_0_1(n456_O_0_1),
    .O_1_0(n456_O_1_0),
    .O_1_1(n456_O_1_1),
    .O_2_0(n456_O_2_0),
    .O_2_1(n456_O_2_1),
    .O_3_0(n456_O_3_0),
    .O_3_1(n456_O_3_1),
    .O_4_0(n456_O_4_0),
    .O_4_1(n456_O_4_1),
    .O_5_0(n456_O_5_0),
    .O_5_1(n456_O_5_1),
    .O_6_0(n456_O_6_0),
    .O_6_1(n456_O_6_1),
    .O_7_0(n456_O_7_0),
    .O_7_1(n456_O_7_1)
  );
  Map2T_1 n463 ( // @[Top.scala 812:22]
    .valid_up(n463_valid_up),
    .valid_down(n463_valid_down),
    .I0_0_0(n463_I0_0_0),
    .I0_0_1(n463_I0_0_1),
    .I0_1_0(n463_I0_1_0),
    .I0_1_1(n463_I0_1_1),
    .I0_2_0(n463_I0_2_0),
    .I0_2_1(n463_I0_2_1),
    .I0_3_0(n463_I0_3_0),
    .I0_3_1(n463_I0_3_1),
    .I0_4_0(n463_I0_4_0),
    .I0_4_1(n463_I0_4_1),
    .I0_5_0(n463_I0_5_0),
    .I0_5_1(n463_I0_5_1),
    .I0_6_0(n463_I0_6_0),
    .I0_6_1(n463_I0_6_1),
    .I0_7_0(n463_I0_7_0),
    .I0_7_1(n463_I0_7_1),
    .I1_0(n463_I1_0),
    .I1_1(n463_I1_1),
    .I1_2(n463_I1_2),
    .I1_3(n463_I1_3),
    .I1_4(n463_I1_4),
    .I1_5(n463_I1_5),
    .I1_6(n463_I1_6),
    .I1_7(n463_I1_7),
    .O_0_0(n463_O_0_0),
    .O_0_1(n463_O_0_1),
    .O_0_2(n463_O_0_2),
    .O_1_0(n463_O_1_0),
    .O_1_1(n463_O_1_1),
    .O_1_2(n463_O_1_2),
    .O_2_0(n463_O_2_0),
    .O_2_1(n463_O_2_1),
    .O_2_2(n463_O_2_2),
    .O_3_0(n463_O_3_0),
    .O_3_1(n463_O_3_1),
    .O_3_2(n463_O_3_2),
    .O_4_0(n463_O_4_0),
    .O_4_1(n463_O_4_1),
    .O_4_2(n463_O_4_2),
    .O_5_0(n463_O_5_0),
    .O_5_1(n463_O_5_1),
    .O_5_2(n463_O_5_2),
    .O_6_0(n463_O_6_0),
    .O_6_1(n463_O_6_1),
    .O_6_2(n463_O_6_2),
    .O_7_0(n463_O_7_0),
    .O_7_1(n463_O_7_1),
    .O_7_2(n463_O_7_2)
  );
  MapT n472 ( // @[Top.scala 816:22]
    .valid_up(n472_valid_up),
    .valid_down(n472_valid_down),
    .I_0_0(n472_I_0_0),
    .I_0_1(n472_I_0_1),
    .I_0_2(n472_I_0_2),
    .I_1_0(n472_I_1_0),
    .I_1_1(n472_I_1_1),
    .I_1_2(n472_I_1_2),
    .I_2_0(n472_I_2_0),
    .I_2_1(n472_I_2_1),
    .I_2_2(n472_I_2_2),
    .I_3_0(n472_I_3_0),
    .I_3_1(n472_I_3_1),
    .I_3_2(n472_I_3_2),
    .I_4_0(n472_I_4_0),
    .I_4_1(n472_I_4_1),
    .I_4_2(n472_I_4_2),
    .I_5_0(n472_I_5_0),
    .I_5_1(n472_I_5_1),
    .I_5_2(n472_I_5_2),
    .I_6_0(n472_I_6_0),
    .I_6_1(n472_I_6_1),
    .I_6_2(n472_I_6_2),
    .I_7_0(n472_I_7_0),
    .I_7_1(n472_I_7_1),
    .I_7_2(n472_I_7_2),
    .O_0_0_0(n472_O_0_0_0),
    .O_0_0_1(n472_O_0_0_1),
    .O_0_0_2(n472_O_0_0_2),
    .O_1_0_0(n472_O_1_0_0),
    .O_1_0_1(n472_O_1_0_1),
    .O_1_0_2(n472_O_1_0_2),
    .O_2_0_0(n472_O_2_0_0),
    .O_2_0_1(n472_O_2_0_1),
    .O_2_0_2(n472_O_2_0_2),
    .O_3_0_0(n472_O_3_0_0),
    .O_3_0_1(n472_O_3_0_1),
    .O_3_0_2(n472_O_3_0_2),
    .O_4_0_0(n472_O_4_0_0),
    .O_4_0_1(n472_O_4_0_1),
    .O_4_0_2(n472_O_4_0_2),
    .O_5_0_0(n472_O_5_0_0),
    .O_5_0_1(n472_O_5_0_1),
    .O_5_0_2(n472_O_5_0_2),
    .O_6_0_0(n472_O_6_0_0),
    .O_6_0_1(n472_O_6_0_1),
    .O_6_0_2(n472_O_6_0_2),
    .O_7_0_0(n472_O_7_0_0),
    .O_7_0_1(n472_O_7_0_1),
    .O_7_0_2(n472_O_7_0_2)
  );
  MapT_1 n479 ( // @[Top.scala 819:22]
    .valid_up(n479_valid_up),
    .valid_down(n479_valid_down),
    .I_0_0_0(n479_I_0_0_0),
    .I_0_0_1(n479_I_0_0_1),
    .I_0_0_2(n479_I_0_0_2),
    .I_1_0_0(n479_I_1_0_0),
    .I_1_0_1(n479_I_1_0_1),
    .I_1_0_2(n479_I_1_0_2),
    .I_2_0_0(n479_I_2_0_0),
    .I_2_0_1(n479_I_2_0_1),
    .I_2_0_2(n479_I_2_0_2),
    .I_3_0_0(n479_I_3_0_0),
    .I_3_0_1(n479_I_3_0_1),
    .I_3_0_2(n479_I_3_0_2),
    .I_4_0_0(n479_I_4_0_0),
    .I_4_0_1(n479_I_4_0_1),
    .I_4_0_2(n479_I_4_0_2),
    .I_5_0_0(n479_I_5_0_0),
    .I_5_0_1(n479_I_5_0_1),
    .I_5_0_2(n479_I_5_0_2),
    .I_6_0_0(n479_I_6_0_0),
    .I_6_0_1(n479_I_6_0_1),
    .I_6_0_2(n479_I_6_0_2),
    .I_7_0_0(n479_I_7_0_0),
    .I_7_0_1(n479_I_7_0_1),
    .I_7_0_2(n479_I_7_0_2),
    .O_0_0(n479_O_0_0),
    .O_0_1(n479_O_0_1),
    .O_0_2(n479_O_0_2),
    .O_1_0(n479_O_1_0),
    .O_1_1(n479_O_1_1),
    .O_1_2(n479_O_1_2),
    .O_2_0(n479_O_2_0),
    .O_2_1(n479_O_2_1),
    .O_2_2(n479_O_2_2),
    .O_3_0(n479_O_3_0),
    .O_3_1(n479_O_3_1),
    .O_3_2(n479_O_3_2),
    .O_4_0(n479_O_4_0),
    .O_4_1(n479_O_4_1),
    .O_4_2(n479_O_4_2),
    .O_5_0(n479_O_5_0),
    .O_5_1(n479_O_5_1),
    .O_5_2(n479_O_5_2),
    .O_6_0(n479_O_6_0),
    .O_6_1(n479_O_6_1),
    .O_6_2(n479_O_6_2),
    .O_7_0(n479_O_7_0),
    .O_7_1(n479_O_7_1),
    .O_7_2(n479_O_7_2)
  );
  ShiftTS_2 n480 ( // @[Top.scala 822:22]
    .clock(n480_clock),
    .valid_up(n480_valid_up),
    .valid_down(n480_valid_down),
    .I_0(n480_I_0),
    .I_1(n480_I_1),
    .I_2(n480_I_2),
    .I_3(n480_I_3),
    .I_4(n480_I_4),
    .I_5(n480_I_5),
    .I_6(n480_I_6),
    .I_7(n480_I_7),
    .O_0(n480_O_0),
    .O_1(n480_O_1),
    .O_2(n480_O_2),
    .O_3(n480_O_3),
    .O_4(n480_O_4),
    .O_5(n480_O_5),
    .O_6(n480_O_6),
    .O_7(n480_O_7)
  );
  ShiftTS_2 n481 ( // @[Top.scala 825:22]
    .clock(n481_clock),
    .valid_up(n481_valid_up),
    .valid_down(n481_valid_down),
    .I_0(n481_I_0),
    .I_1(n481_I_1),
    .I_2(n481_I_2),
    .I_3(n481_I_3),
    .I_4(n481_I_4),
    .I_5(n481_I_5),
    .I_6(n481_I_6),
    .I_7(n481_I_7),
    .O_0(n481_O_0),
    .O_1(n481_O_1),
    .O_2(n481_O_2),
    .O_3(n481_O_3),
    .O_4(n481_O_4),
    .O_5(n481_O_5),
    .O_6(n481_O_6),
    .O_7(n481_O_7)
  );
  Map2T n482 ( // @[Top.scala 828:22]
    .valid_up(n482_valid_up),
    .valid_down(n482_valid_down),
    .I0_0(n482_I0_0),
    .I0_1(n482_I0_1),
    .I0_2(n482_I0_2),
    .I0_3(n482_I0_3),
    .I0_4(n482_I0_4),
    .I0_5(n482_I0_5),
    .I0_6(n482_I0_6),
    .I0_7(n482_I0_7),
    .I1_0(n482_I1_0),
    .I1_1(n482_I1_1),
    .I1_2(n482_I1_2),
    .I1_3(n482_I1_3),
    .I1_4(n482_I1_4),
    .I1_5(n482_I1_5),
    .I1_6(n482_I1_6),
    .I1_7(n482_I1_7),
    .O_0_0(n482_O_0_0),
    .O_0_1(n482_O_0_1),
    .O_1_0(n482_O_1_0),
    .O_1_1(n482_O_1_1),
    .O_2_0(n482_O_2_0),
    .O_2_1(n482_O_2_1),
    .O_3_0(n482_O_3_0),
    .O_3_1(n482_O_3_1),
    .O_4_0(n482_O_4_0),
    .O_4_1(n482_O_4_1),
    .O_5_0(n482_O_5_0),
    .O_5_1(n482_O_5_1),
    .O_6_0(n482_O_6_0),
    .O_6_1(n482_O_6_1),
    .O_7_0(n482_O_7_0),
    .O_7_1(n482_O_7_1)
  );
  Map2T_1 n489 ( // @[Top.scala 832:22]
    .valid_up(n489_valid_up),
    .valid_down(n489_valid_down),
    .I0_0_0(n489_I0_0_0),
    .I0_0_1(n489_I0_0_1),
    .I0_1_0(n489_I0_1_0),
    .I0_1_1(n489_I0_1_1),
    .I0_2_0(n489_I0_2_0),
    .I0_2_1(n489_I0_2_1),
    .I0_3_0(n489_I0_3_0),
    .I0_3_1(n489_I0_3_1),
    .I0_4_0(n489_I0_4_0),
    .I0_4_1(n489_I0_4_1),
    .I0_5_0(n489_I0_5_0),
    .I0_5_1(n489_I0_5_1),
    .I0_6_0(n489_I0_6_0),
    .I0_6_1(n489_I0_6_1),
    .I0_7_0(n489_I0_7_0),
    .I0_7_1(n489_I0_7_1),
    .I1_0(n489_I1_0),
    .I1_1(n489_I1_1),
    .I1_2(n489_I1_2),
    .I1_3(n489_I1_3),
    .I1_4(n489_I1_4),
    .I1_5(n489_I1_5),
    .I1_6(n489_I1_6),
    .I1_7(n489_I1_7),
    .O_0_0(n489_O_0_0),
    .O_0_1(n489_O_0_1),
    .O_0_2(n489_O_0_2),
    .O_1_0(n489_O_1_0),
    .O_1_1(n489_O_1_1),
    .O_1_2(n489_O_1_2),
    .O_2_0(n489_O_2_0),
    .O_2_1(n489_O_2_1),
    .O_2_2(n489_O_2_2),
    .O_3_0(n489_O_3_0),
    .O_3_1(n489_O_3_1),
    .O_3_2(n489_O_3_2),
    .O_4_0(n489_O_4_0),
    .O_4_1(n489_O_4_1),
    .O_4_2(n489_O_4_2),
    .O_5_0(n489_O_5_0),
    .O_5_1(n489_O_5_1),
    .O_5_2(n489_O_5_2),
    .O_6_0(n489_O_6_0),
    .O_6_1(n489_O_6_1),
    .O_6_2(n489_O_6_2),
    .O_7_0(n489_O_7_0),
    .O_7_1(n489_O_7_1),
    .O_7_2(n489_O_7_2)
  );
  MapT n498 ( // @[Top.scala 836:22]
    .valid_up(n498_valid_up),
    .valid_down(n498_valid_down),
    .I_0_0(n498_I_0_0),
    .I_0_1(n498_I_0_1),
    .I_0_2(n498_I_0_2),
    .I_1_0(n498_I_1_0),
    .I_1_1(n498_I_1_1),
    .I_1_2(n498_I_1_2),
    .I_2_0(n498_I_2_0),
    .I_2_1(n498_I_2_1),
    .I_2_2(n498_I_2_2),
    .I_3_0(n498_I_3_0),
    .I_3_1(n498_I_3_1),
    .I_3_2(n498_I_3_2),
    .I_4_0(n498_I_4_0),
    .I_4_1(n498_I_4_1),
    .I_4_2(n498_I_4_2),
    .I_5_0(n498_I_5_0),
    .I_5_1(n498_I_5_1),
    .I_5_2(n498_I_5_2),
    .I_6_0(n498_I_6_0),
    .I_6_1(n498_I_6_1),
    .I_6_2(n498_I_6_2),
    .I_7_0(n498_I_7_0),
    .I_7_1(n498_I_7_1),
    .I_7_2(n498_I_7_2),
    .O_0_0_0(n498_O_0_0_0),
    .O_0_0_1(n498_O_0_0_1),
    .O_0_0_2(n498_O_0_0_2),
    .O_1_0_0(n498_O_1_0_0),
    .O_1_0_1(n498_O_1_0_1),
    .O_1_0_2(n498_O_1_0_2),
    .O_2_0_0(n498_O_2_0_0),
    .O_2_0_1(n498_O_2_0_1),
    .O_2_0_2(n498_O_2_0_2),
    .O_3_0_0(n498_O_3_0_0),
    .O_3_0_1(n498_O_3_0_1),
    .O_3_0_2(n498_O_3_0_2),
    .O_4_0_0(n498_O_4_0_0),
    .O_4_0_1(n498_O_4_0_1),
    .O_4_0_2(n498_O_4_0_2),
    .O_5_0_0(n498_O_5_0_0),
    .O_5_0_1(n498_O_5_0_1),
    .O_5_0_2(n498_O_5_0_2),
    .O_6_0_0(n498_O_6_0_0),
    .O_6_0_1(n498_O_6_0_1),
    .O_6_0_2(n498_O_6_0_2),
    .O_7_0_0(n498_O_7_0_0),
    .O_7_0_1(n498_O_7_0_1),
    .O_7_0_2(n498_O_7_0_2)
  );
  MapT_1 n505 ( // @[Top.scala 839:22]
    .valid_up(n505_valid_up),
    .valid_down(n505_valid_down),
    .I_0_0_0(n505_I_0_0_0),
    .I_0_0_1(n505_I_0_0_1),
    .I_0_0_2(n505_I_0_0_2),
    .I_1_0_0(n505_I_1_0_0),
    .I_1_0_1(n505_I_1_0_1),
    .I_1_0_2(n505_I_1_0_2),
    .I_2_0_0(n505_I_2_0_0),
    .I_2_0_1(n505_I_2_0_1),
    .I_2_0_2(n505_I_2_0_2),
    .I_3_0_0(n505_I_3_0_0),
    .I_3_0_1(n505_I_3_0_1),
    .I_3_0_2(n505_I_3_0_2),
    .I_4_0_0(n505_I_4_0_0),
    .I_4_0_1(n505_I_4_0_1),
    .I_4_0_2(n505_I_4_0_2),
    .I_5_0_0(n505_I_5_0_0),
    .I_5_0_1(n505_I_5_0_1),
    .I_5_0_2(n505_I_5_0_2),
    .I_6_0_0(n505_I_6_0_0),
    .I_6_0_1(n505_I_6_0_1),
    .I_6_0_2(n505_I_6_0_2),
    .I_7_0_0(n505_I_7_0_0),
    .I_7_0_1(n505_I_7_0_1),
    .I_7_0_2(n505_I_7_0_2),
    .O_0_0(n505_O_0_0),
    .O_0_1(n505_O_0_1),
    .O_0_2(n505_O_0_2),
    .O_1_0(n505_O_1_0),
    .O_1_1(n505_O_1_1),
    .O_1_2(n505_O_1_2),
    .O_2_0(n505_O_2_0),
    .O_2_1(n505_O_2_1),
    .O_2_2(n505_O_2_2),
    .O_3_0(n505_O_3_0),
    .O_3_1(n505_O_3_1),
    .O_3_2(n505_O_3_2),
    .O_4_0(n505_O_4_0),
    .O_4_1(n505_O_4_1),
    .O_4_2(n505_O_4_2),
    .O_5_0(n505_O_5_0),
    .O_5_1(n505_O_5_1),
    .O_5_2(n505_O_5_2),
    .O_6_0(n505_O_6_0),
    .O_6_1(n505_O_6_1),
    .O_6_2(n505_O_6_2),
    .O_7_0(n505_O_7_0),
    .O_7_1(n505_O_7_1),
    .O_7_2(n505_O_7_2)
  );
  Map2T_4 n506 ( // @[Top.scala 842:22]
    .valid_up(n506_valid_up),
    .valid_down(n506_valid_down),
    .I0_0_0(n506_I0_0_0),
    .I0_0_1(n506_I0_0_1),
    .I0_0_2(n506_I0_0_2),
    .I0_1_0(n506_I0_1_0),
    .I0_1_1(n506_I0_1_1),
    .I0_1_2(n506_I0_1_2),
    .I0_2_0(n506_I0_2_0),
    .I0_2_1(n506_I0_2_1),
    .I0_2_2(n506_I0_2_2),
    .I0_3_0(n506_I0_3_0),
    .I0_3_1(n506_I0_3_1),
    .I0_3_2(n506_I0_3_2),
    .I0_4_0(n506_I0_4_0),
    .I0_4_1(n506_I0_4_1),
    .I0_4_2(n506_I0_4_2),
    .I0_5_0(n506_I0_5_0),
    .I0_5_1(n506_I0_5_1),
    .I0_5_2(n506_I0_5_2),
    .I0_6_0(n506_I0_6_0),
    .I0_6_1(n506_I0_6_1),
    .I0_6_2(n506_I0_6_2),
    .I0_7_0(n506_I0_7_0),
    .I0_7_1(n506_I0_7_1),
    .I0_7_2(n506_I0_7_2),
    .I1_0_0(n506_I1_0_0),
    .I1_0_1(n506_I1_0_1),
    .I1_0_2(n506_I1_0_2),
    .I1_1_0(n506_I1_1_0),
    .I1_1_1(n506_I1_1_1),
    .I1_1_2(n506_I1_1_2),
    .I1_2_0(n506_I1_2_0),
    .I1_2_1(n506_I1_2_1),
    .I1_2_2(n506_I1_2_2),
    .I1_3_0(n506_I1_3_0),
    .I1_3_1(n506_I1_3_1),
    .I1_3_2(n506_I1_3_2),
    .I1_4_0(n506_I1_4_0),
    .I1_4_1(n506_I1_4_1),
    .I1_4_2(n506_I1_4_2),
    .I1_5_0(n506_I1_5_0),
    .I1_5_1(n506_I1_5_1),
    .I1_5_2(n506_I1_5_2),
    .I1_6_0(n506_I1_6_0),
    .I1_6_1(n506_I1_6_1),
    .I1_6_2(n506_I1_6_2),
    .I1_7_0(n506_I1_7_0),
    .I1_7_1(n506_I1_7_1),
    .I1_7_2(n506_I1_7_2),
    .O_0_0_0(n506_O_0_0_0),
    .O_0_0_1(n506_O_0_0_1),
    .O_0_0_2(n506_O_0_0_2),
    .O_0_1_0(n506_O_0_1_0),
    .O_0_1_1(n506_O_0_1_1),
    .O_0_1_2(n506_O_0_1_2),
    .O_1_0_0(n506_O_1_0_0),
    .O_1_0_1(n506_O_1_0_1),
    .O_1_0_2(n506_O_1_0_2),
    .O_1_1_0(n506_O_1_1_0),
    .O_1_1_1(n506_O_1_1_1),
    .O_1_1_2(n506_O_1_1_2),
    .O_2_0_0(n506_O_2_0_0),
    .O_2_0_1(n506_O_2_0_1),
    .O_2_0_2(n506_O_2_0_2),
    .O_2_1_0(n506_O_2_1_0),
    .O_2_1_1(n506_O_2_1_1),
    .O_2_1_2(n506_O_2_1_2),
    .O_3_0_0(n506_O_3_0_0),
    .O_3_0_1(n506_O_3_0_1),
    .O_3_0_2(n506_O_3_0_2),
    .O_3_1_0(n506_O_3_1_0),
    .O_3_1_1(n506_O_3_1_1),
    .O_3_1_2(n506_O_3_1_2),
    .O_4_0_0(n506_O_4_0_0),
    .O_4_0_1(n506_O_4_0_1),
    .O_4_0_2(n506_O_4_0_2),
    .O_4_1_0(n506_O_4_1_0),
    .O_4_1_1(n506_O_4_1_1),
    .O_4_1_2(n506_O_4_1_2),
    .O_5_0_0(n506_O_5_0_0),
    .O_5_0_1(n506_O_5_0_1),
    .O_5_0_2(n506_O_5_0_2),
    .O_5_1_0(n506_O_5_1_0),
    .O_5_1_1(n506_O_5_1_1),
    .O_5_1_2(n506_O_5_1_2),
    .O_6_0_0(n506_O_6_0_0),
    .O_6_0_1(n506_O_6_0_1),
    .O_6_0_2(n506_O_6_0_2),
    .O_6_1_0(n506_O_6_1_0),
    .O_6_1_1(n506_O_6_1_1),
    .O_6_1_2(n506_O_6_1_2),
    .O_7_0_0(n506_O_7_0_0),
    .O_7_0_1(n506_O_7_0_1),
    .O_7_0_2(n506_O_7_0_2),
    .O_7_1_0(n506_O_7_1_0),
    .O_7_1_1(n506_O_7_1_1),
    .O_7_1_2(n506_O_7_1_2)
  );
  ShiftTS_2 n513 ( // @[Top.scala 846:22]
    .clock(n513_clock),
    .valid_up(n513_valid_up),
    .valid_down(n513_valid_down),
    .I_0(n513_I_0),
    .I_1(n513_I_1),
    .I_2(n513_I_2),
    .I_3(n513_I_3),
    .I_4(n513_I_4),
    .I_5(n513_I_5),
    .I_6(n513_I_6),
    .I_7(n513_I_7),
    .O_0(n513_O_0),
    .O_1(n513_O_1),
    .O_2(n513_O_2),
    .O_3(n513_O_3),
    .O_4(n513_O_4),
    .O_5(n513_O_5),
    .O_6(n513_O_6),
    .O_7(n513_O_7)
  );
  ShiftTS_2 n514 ( // @[Top.scala 849:22]
    .clock(n514_clock),
    .valid_up(n514_valid_up),
    .valid_down(n514_valid_down),
    .I_0(n514_I_0),
    .I_1(n514_I_1),
    .I_2(n514_I_2),
    .I_3(n514_I_3),
    .I_4(n514_I_4),
    .I_5(n514_I_5),
    .I_6(n514_I_6),
    .I_7(n514_I_7),
    .O_0(n514_O_0),
    .O_1(n514_O_1),
    .O_2(n514_O_2),
    .O_3(n514_O_3),
    .O_4(n514_O_4),
    .O_5(n514_O_5),
    .O_6(n514_O_6),
    .O_7(n514_O_7)
  );
  Map2T n515 ( // @[Top.scala 852:22]
    .valid_up(n515_valid_up),
    .valid_down(n515_valid_down),
    .I0_0(n515_I0_0),
    .I0_1(n515_I0_1),
    .I0_2(n515_I0_2),
    .I0_3(n515_I0_3),
    .I0_4(n515_I0_4),
    .I0_5(n515_I0_5),
    .I0_6(n515_I0_6),
    .I0_7(n515_I0_7),
    .I1_0(n515_I1_0),
    .I1_1(n515_I1_1),
    .I1_2(n515_I1_2),
    .I1_3(n515_I1_3),
    .I1_4(n515_I1_4),
    .I1_5(n515_I1_5),
    .I1_6(n515_I1_6),
    .I1_7(n515_I1_7),
    .O_0_0(n515_O_0_0),
    .O_0_1(n515_O_0_1),
    .O_1_0(n515_O_1_0),
    .O_1_1(n515_O_1_1),
    .O_2_0(n515_O_2_0),
    .O_2_1(n515_O_2_1),
    .O_3_0(n515_O_3_0),
    .O_3_1(n515_O_3_1),
    .O_4_0(n515_O_4_0),
    .O_4_1(n515_O_4_1),
    .O_5_0(n515_O_5_0),
    .O_5_1(n515_O_5_1),
    .O_6_0(n515_O_6_0),
    .O_6_1(n515_O_6_1),
    .O_7_0(n515_O_7_0),
    .O_7_1(n515_O_7_1)
  );
  Map2T_1 n522 ( // @[Top.scala 856:22]
    .valid_up(n522_valid_up),
    .valid_down(n522_valid_down),
    .I0_0_0(n522_I0_0_0),
    .I0_0_1(n522_I0_0_1),
    .I0_1_0(n522_I0_1_0),
    .I0_1_1(n522_I0_1_1),
    .I0_2_0(n522_I0_2_0),
    .I0_2_1(n522_I0_2_1),
    .I0_3_0(n522_I0_3_0),
    .I0_3_1(n522_I0_3_1),
    .I0_4_0(n522_I0_4_0),
    .I0_4_1(n522_I0_4_1),
    .I0_5_0(n522_I0_5_0),
    .I0_5_1(n522_I0_5_1),
    .I0_6_0(n522_I0_6_0),
    .I0_6_1(n522_I0_6_1),
    .I0_7_0(n522_I0_7_0),
    .I0_7_1(n522_I0_7_1),
    .I1_0(n522_I1_0),
    .I1_1(n522_I1_1),
    .I1_2(n522_I1_2),
    .I1_3(n522_I1_3),
    .I1_4(n522_I1_4),
    .I1_5(n522_I1_5),
    .I1_6(n522_I1_6),
    .I1_7(n522_I1_7),
    .O_0_0(n522_O_0_0),
    .O_0_1(n522_O_0_1),
    .O_0_2(n522_O_0_2),
    .O_1_0(n522_O_1_0),
    .O_1_1(n522_O_1_1),
    .O_1_2(n522_O_1_2),
    .O_2_0(n522_O_2_0),
    .O_2_1(n522_O_2_1),
    .O_2_2(n522_O_2_2),
    .O_3_0(n522_O_3_0),
    .O_3_1(n522_O_3_1),
    .O_3_2(n522_O_3_2),
    .O_4_0(n522_O_4_0),
    .O_4_1(n522_O_4_1),
    .O_4_2(n522_O_4_2),
    .O_5_0(n522_O_5_0),
    .O_5_1(n522_O_5_1),
    .O_5_2(n522_O_5_2),
    .O_6_0(n522_O_6_0),
    .O_6_1(n522_O_6_1),
    .O_6_2(n522_O_6_2),
    .O_7_0(n522_O_7_0),
    .O_7_1(n522_O_7_1),
    .O_7_2(n522_O_7_2)
  );
  MapT n531 ( // @[Top.scala 860:22]
    .valid_up(n531_valid_up),
    .valid_down(n531_valid_down),
    .I_0_0(n531_I_0_0),
    .I_0_1(n531_I_0_1),
    .I_0_2(n531_I_0_2),
    .I_1_0(n531_I_1_0),
    .I_1_1(n531_I_1_1),
    .I_1_2(n531_I_1_2),
    .I_2_0(n531_I_2_0),
    .I_2_1(n531_I_2_1),
    .I_2_2(n531_I_2_2),
    .I_3_0(n531_I_3_0),
    .I_3_1(n531_I_3_1),
    .I_3_2(n531_I_3_2),
    .I_4_0(n531_I_4_0),
    .I_4_1(n531_I_4_1),
    .I_4_2(n531_I_4_2),
    .I_5_0(n531_I_5_0),
    .I_5_1(n531_I_5_1),
    .I_5_2(n531_I_5_2),
    .I_6_0(n531_I_6_0),
    .I_6_1(n531_I_6_1),
    .I_6_2(n531_I_6_2),
    .I_7_0(n531_I_7_0),
    .I_7_1(n531_I_7_1),
    .I_7_2(n531_I_7_2),
    .O_0_0_0(n531_O_0_0_0),
    .O_0_0_1(n531_O_0_0_1),
    .O_0_0_2(n531_O_0_0_2),
    .O_1_0_0(n531_O_1_0_0),
    .O_1_0_1(n531_O_1_0_1),
    .O_1_0_2(n531_O_1_0_2),
    .O_2_0_0(n531_O_2_0_0),
    .O_2_0_1(n531_O_2_0_1),
    .O_2_0_2(n531_O_2_0_2),
    .O_3_0_0(n531_O_3_0_0),
    .O_3_0_1(n531_O_3_0_1),
    .O_3_0_2(n531_O_3_0_2),
    .O_4_0_0(n531_O_4_0_0),
    .O_4_0_1(n531_O_4_0_1),
    .O_4_0_2(n531_O_4_0_2),
    .O_5_0_0(n531_O_5_0_0),
    .O_5_0_1(n531_O_5_0_1),
    .O_5_0_2(n531_O_5_0_2),
    .O_6_0_0(n531_O_6_0_0),
    .O_6_0_1(n531_O_6_0_1),
    .O_6_0_2(n531_O_6_0_2),
    .O_7_0_0(n531_O_7_0_0),
    .O_7_0_1(n531_O_7_0_1),
    .O_7_0_2(n531_O_7_0_2)
  );
  MapT_1 n538 ( // @[Top.scala 863:22]
    .valid_up(n538_valid_up),
    .valid_down(n538_valid_down),
    .I_0_0_0(n538_I_0_0_0),
    .I_0_0_1(n538_I_0_0_1),
    .I_0_0_2(n538_I_0_0_2),
    .I_1_0_0(n538_I_1_0_0),
    .I_1_0_1(n538_I_1_0_1),
    .I_1_0_2(n538_I_1_0_2),
    .I_2_0_0(n538_I_2_0_0),
    .I_2_0_1(n538_I_2_0_1),
    .I_2_0_2(n538_I_2_0_2),
    .I_3_0_0(n538_I_3_0_0),
    .I_3_0_1(n538_I_3_0_1),
    .I_3_0_2(n538_I_3_0_2),
    .I_4_0_0(n538_I_4_0_0),
    .I_4_0_1(n538_I_4_0_1),
    .I_4_0_2(n538_I_4_0_2),
    .I_5_0_0(n538_I_5_0_0),
    .I_5_0_1(n538_I_5_0_1),
    .I_5_0_2(n538_I_5_0_2),
    .I_6_0_0(n538_I_6_0_0),
    .I_6_0_1(n538_I_6_0_1),
    .I_6_0_2(n538_I_6_0_2),
    .I_7_0_0(n538_I_7_0_0),
    .I_7_0_1(n538_I_7_0_1),
    .I_7_0_2(n538_I_7_0_2),
    .O_0_0(n538_O_0_0),
    .O_0_1(n538_O_0_1),
    .O_0_2(n538_O_0_2),
    .O_1_0(n538_O_1_0),
    .O_1_1(n538_O_1_1),
    .O_1_2(n538_O_1_2),
    .O_2_0(n538_O_2_0),
    .O_2_1(n538_O_2_1),
    .O_2_2(n538_O_2_2),
    .O_3_0(n538_O_3_0),
    .O_3_1(n538_O_3_1),
    .O_3_2(n538_O_3_2),
    .O_4_0(n538_O_4_0),
    .O_4_1(n538_O_4_1),
    .O_4_2(n538_O_4_2),
    .O_5_0(n538_O_5_0),
    .O_5_1(n538_O_5_1),
    .O_5_2(n538_O_5_2),
    .O_6_0(n538_O_6_0),
    .O_6_1(n538_O_6_1),
    .O_6_2(n538_O_6_2),
    .O_7_0(n538_O_7_0),
    .O_7_1(n538_O_7_1),
    .O_7_2(n538_O_7_2)
  );
  Map2T_7 n539 ( // @[Top.scala 866:22]
    .valid_up(n539_valid_up),
    .valid_down(n539_valid_down),
    .I0_0_0_0(n539_I0_0_0_0),
    .I0_0_0_1(n539_I0_0_0_1),
    .I0_0_0_2(n539_I0_0_0_2),
    .I0_0_1_0(n539_I0_0_1_0),
    .I0_0_1_1(n539_I0_0_1_1),
    .I0_0_1_2(n539_I0_0_1_2),
    .I0_1_0_0(n539_I0_1_0_0),
    .I0_1_0_1(n539_I0_1_0_1),
    .I0_1_0_2(n539_I0_1_0_2),
    .I0_1_1_0(n539_I0_1_1_0),
    .I0_1_1_1(n539_I0_1_1_1),
    .I0_1_1_2(n539_I0_1_1_2),
    .I0_2_0_0(n539_I0_2_0_0),
    .I0_2_0_1(n539_I0_2_0_1),
    .I0_2_0_2(n539_I0_2_0_2),
    .I0_2_1_0(n539_I0_2_1_0),
    .I0_2_1_1(n539_I0_2_1_1),
    .I0_2_1_2(n539_I0_2_1_2),
    .I0_3_0_0(n539_I0_3_0_0),
    .I0_3_0_1(n539_I0_3_0_1),
    .I0_3_0_2(n539_I0_3_0_2),
    .I0_3_1_0(n539_I0_3_1_0),
    .I0_3_1_1(n539_I0_3_1_1),
    .I0_3_1_2(n539_I0_3_1_2),
    .I0_4_0_0(n539_I0_4_0_0),
    .I0_4_0_1(n539_I0_4_0_1),
    .I0_4_0_2(n539_I0_4_0_2),
    .I0_4_1_0(n539_I0_4_1_0),
    .I0_4_1_1(n539_I0_4_1_1),
    .I0_4_1_2(n539_I0_4_1_2),
    .I0_5_0_0(n539_I0_5_0_0),
    .I0_5_0_1(n539_I0_5_0_1),
    .I0_5_0_2(n539_I0_5_0_2),
    .I0_5_1_0(n539_I0_5_1_0),
    .I0_5_1_1(n539_I0_5_1_1),
    .I0_5_1_2(n539_I0_5_1_2),
    .I0_6_0_0(n539_I0_6_0_0),
    .I0_6_0_1(n539_I0_6_0_1),
    .I0_6_0_2(n539_I0_6_0_2),
    .I0_6_1_0(n539_I0_6_1_0),
    .I0_6_1_1(n539_I0_6_1_1),
    .I0_6_1_2(n539_I0_6_1_2),
    .I0_7_0_0(n539_I0_7_0_0),
    .I0_7_0_1(n539_I0_7_0_1),
    .I0_7_0_2(n539_I0_7_0_2),
    .I0_7_1_0(n539_I0_7_1_0),
    .I0_7_1_1(n539_I0_7_1_1),
    .I0_7_1_2(n539_I0_7_1_2),
    .I1_0_0(n539_I1_0_0),
    .I1_0_1(n539_I1_0_1),
    .I1_0_2(n539_I1_0_2),
    .I1_1_0(n539_I1_1_0),
    .I1_1_1(n539_I1_1_1),
    .I1_1_2(n539_I1_1_2),
    .I1_2_0(n539_I1_2_0),
    .I1_2_1(n539_I1_2_1),
    .I1_2_2(n539_I1_2_2),
    .I1_3_0(n539_I1_3_0),
    .I1_3_1(n539_I1_3_1),
    .I1_3_2(n539_I1_3_2),
    .I1_4_0(n539_I1_4_0),
    .I1_4_1(n539_I1_4_1),
    .I1_4_2(n539_I1_4_2),
    .I1_5_0(n539_I1_5_0),
    .I1_5_1(n539_I1_5_1),
    .I1_5_2(n539_I1_5_2),
    .I1_6_0(n539_I1_6_0),
    .I1_6_1(n539_I1_6_1),
    .I1_6_2(n539_I1_6_2),
    .I1_7_0(n539_I1_7_0),
    .I1_7_1(n539_I1_7_1),
    .I1_7_2(n539_I1_7_2),
    .O_0_0_0(n539_O_0_0_0),
    .O_0_0_1(n539_O_0_0_1),
    .O_0_0_2(n539_O_0_0_2),
    .O_0_1_0(n539_O_0_1_0),
    .O_0_1_1(n539_O_0_1_1),
    .O_0_1_2(n539_O_0_1_2),
    .O_0_2_0(n539_O_0_2_0),
    .O_0_2_1(n539_O_0_2_1),
    .O_0_2_2(n539_O_0_2_2),
    .O_1_0_0(n539_O_1_0_0),
    .O_1_0_1(n539_O_1_0_1),
    .O_1_0_2(n539_O_1_0_2),
    .O_1_1_0(n539_O_1_1_0),
    .O_1_1_1(n539_O_1_1_1),
    .O_1_1_2(n539_O_1_1_2),
    .O_1_2_0(n539_O_1_2_0),
    .O_1_2_1(n539_O_1_2_1),
    .O_1_2_2(n539_O_1_2_2),
    .O_2_0_0(n539_O_2_0_0),
    .O_2_0_1(n539_O_2_0_1),
    .O_2_0_2(n539_O_2_0_2),
    .O_2_1_0(n539_O_2_1_0),
    .O_2_1_1(n539_O_2_1_1),
    .O_2_1_2(n539_O_2_1_2),
    .O_2_2_0(n539_O_2_2_0),
    .O_2_2_1(n539_O_2_2_1),
    .O_2_2_2(n539_O_2_2_2),
    .O_3_0_0(n539_O_3_0_0),
    .O_3_0_1(n539_O_3_0_1),
    .O_3_0_2(n539_O_3_0_2),
    .O_3_1_0(n539_O_3_1_0),
    .O_3_1_1(n539_O_3_1_1),
    .O_3_1_2(n539_O_3_1_2),
    .O_3_2_0(n539_O_3_2_0),
    .O_3_2_1(n539_O_3_2_1),
    .O_3_2_2(n539_O_3_2_2),
    .O_4_0_0(n539_O_4_0_0),
    .O_4_0_1(n539_O_4_0_1),
    .O_4_0_2(n539_O_4_0_2),
    .O_4_1_0(n539_O_4_1_0),
    .O_4_1_1(n539_O_4_1_1),
    .O_4_1_2(n539_O_4_1_2),
    .O_4_2_0(n539_O_4_2_0),
    .O_4_2_1(n539_O_4_2_1),
    .O_4_2_2(n539_O_4_2_2),
    .O_5_0_0(n539_O_5_0_0),
    .O_5_0_1(n539_O_5_0_1),
    .O_5_0_2(n539_O_5_0_2),
    .O_5_1_0(n539_O_5_1_0),
    .O_5_1_1(n539_O_5_1_1),
    .O_5_1_2(n539_O_5_1_2),
    .O_5_2_0(n539_O_5_2_0),
    .O_5_2_1(n539_O_5_2_1),
    .O_5_2_2(n539_O_5_2_2),
    .O_6_0_0(n539_O_6_0_0),
    .O_6_0_1(n539_O_6_0_1),
    .O_6_0_2(n539_O_6_0_2),
    .O_6_1_0(n539_O_6_1_0),
    .O_6_1_1(n539_O_6_1_1),
    .O_6_1_2(n539_O_6_1_2),
    .O_6_2_0(n539_O_6_2_0),
    .O_6_2_1(n539_O_6_2_1),
    .O_6_2_2(n539_O_6_2_2),
    .O_7_0_0(n539_O_7_0_0),
    .O_7_0_1(n539_O_7_0_1),
    .O_7_0_2(n539_O_7_0_2),
    .O_7_1_0(n539_O_7_1_0),
    .O_7_1_1(n539_O_7_1_1),
    .O_7_1_2(n539_O_7_1_2),
    .O_7_2_0(n539_O_7_2_0),
    .O_7_2_1(n539_O_7_2_1),
    .O_7_2_2(n539_O_7_2_2)
  );
  MapT_6 n548 ( // @[Top.scala 870:22]
    .valid_up(n548_valid_up),
    .valid_down(n548_valid_down),
    .I_0_0_0(n548_I_0_0_0),
    .I_0_0_1(n548_I_0_0_1),
    .I_0_0_2(n548_I_0_0_2),
    .I_0_1_0(n548_I_0_1_0),
    .I_0_1_1(n548_I_0_1_1),
    .I_0_1_2(n548_I_0_1_2),
    .I_0_2_0(n548_I_0_2_0),
    .I_0_2_1(n548_I_0_2_1),
    .I_0_2_2(n548_I_0_2_2),
    .I_1_0_0(n548_I_1_0_0),
    .I_1_0_1(n548_I_1_0_1),
    .I_1_0_2(n548_I_1_0_2),
    .I_1_1_0(n548_I_1_1_0),
    .I_1_1_1(n548_I_1_1_1),
    .I_1_1_2(n548_I_1_1_2),
    .I_1_2_0(n548_I_1_2_0),
    .I_1_2_1(n548_I_1_2_1),
    .I_1_2_2(n548_I_1_2_2),
    .I_2_0_0(n548_I_2_0_0),
    .I_2_0_1(n548_I_2_0_1),
    .I_2_0_2(n548_I_2_0_2),
    .I_2_1_0(n548_I_2_1_0),
    .I_2_1_1(n548_I_2_1_1),
    .I_2_1_2(n548_I_2_1_2),
    .I_2_2_0(n548_I_2_2_0),
    .I_2_2_1(n548_I_2_2_1),
    .I_2_2_2(n548_I_2_2_2),
    .I_3_0_0(n548_I_3_0_0),
    .I_3_0_1(n548_I_3_0_1),
    .I_3_0_2(n548_I_3_0_2),
    .I_3_1_0(n548_I_3_1_0),
    .I_3_1_1(n548_I_3_1_1),
    .I_3_1_2(n548_I_3_1_2),
    .I_3_2_0(n548_I_3_2_0),
    .I_3_2_1(n548_I_3_2_1),
    .I_3_2_2(n548_I_3_2_2),
    .I_4_0_0(n548_I_4_0_0),
    .I_4_0_1(n548_I_4_0_1),
    .I_4_0_2(n548_I_4_0_2),
    .I_4_1_0(n548_I_4_1_0),
    .I_4_1_1(n548_I_4_1_1),
    .I_4_1_2(n548_I_4_1_2),
    .I_4_2_0(n548_I_4_2_0),
    .I_4_2_1(n548_I_4_2_1),
    .I_4_2_2(n548_I_4_2_2),
    .I_5_0_0(n548_I_5_0_0),
    .I_5_0_1(n548_I_5_0_1),
    .I_5_0_2(n548_I_5_0_2),
    .I_5_1_0(n548_I_5_1_0),
    .I_5_1_1(n548_I_5_1_1),
    .I_5_1_2(n548_I_5_1_2),
    .I_5_2_0(n548_I_5_2_0),
    .I_5_2_1(n548_I_5_2_1),
    .I_5_2_2(n548_I_5_2_2),
    .I_6_0_0(n548_I_6_0_0),
    .I_6_0_1(n548_I_6_0_1),
    .I_6_0_2(n548_I_6_0_2),
    .I_6_1_0(n548_I_6_1_0),
    .I_6_1_1(n548_I_6_1_1),
    .I_6_1_2(n548_I_6_1_2),
    .I_6_2_0(n548_I_6_2_0),
    .I_6_2_1(n548_I_6_2_1),
    .I_6_2_2(n548_I_6_2_2),
    .I_7_0_0(n548_I_7_0_0),
    .I_7_0_1(n548_I_7_0_1),
    .I_7_0_2(n548_I_7_0_2),
    .I_7_1_0(n548_I_7_1_0),
    .I_7_1_1(n548_I_7_1_1),
    .I_7_1_2(n548_I_7_1_2),
    .I_7_2_0(n548_I_7_2_0),
    .I_7_2_1(n548_I_7_2_1),
    .I_7_2_2(n548_I_7_2_2),
    .O_0_0_0_0(n548_O_0_0_0_0),
    .O_0_0_0_1(n548_O_0_0_0_1),
    .O_0_0_0_2(n548_O_0_0_0_2),
    .O_0_0_1_0(n548_O_0_0_1_0),
    .O_0_0_1_1(n548_O_0_0_1_1),
    .O_0_0_1_2(n548_O_0_0_1_2),
    .O_0_0_2_0(n548_O_0_0_2_0),
    .O_0_0_2_1(n548_O_0_0_2_1),
    .O_0_0_2_2(n548_O_0_0_2_2),
    .O_1_0_0_0(n548_O_1_0_0_0),
    .O_1_0_0_1(n548_O_1_0_0_1),
    .O_1_0_0_2(n548_O_1_0_0_2),
    .O_1_0_1_0(n548_O_1_0_1_0),
    .O_1_0_1_1(n548_O_1_0_1_1),
    .O_1_0_1_2(n548_O_1_0_1_2),
    .O_1_0_2_0(n548_O_1_0_2_0),
    .O_1_0_2_1(n548_O_1_0_2_1),
    .O_1_0_2_2(n548_O_1_0_2_2),
    .O_2_0_0_0(n548_O_2_0_0_0),
    .O_2_0_0_1(n548_O_2_0_0_1),
    .O_2_0_0_2(n548_O_2_0_0_2),
    .O_2_0_1_0(n548_O_2_0_1_0),
    .O_2_0_1_1(n548_O_2_0_1_1),
    .O_2_0_1_2(n548_O_2_0_1_2),
    .O_2_0_2_0(n548_O_2_0_2_0),
    .O_2_0_2_1(n548_O_2_0_2_1),
    .O_2_0_2_2(n548_O_2_0_2_2),
    .O_3_0_0_0(n548_O_3_0_0_0),
    .O_3_0_0_1(n548_O_3_0_0_1),
    .O_3_0_0_2(n548_O_3_0_0_2),
    .O_3_0_1_0(n548_O_3_0_1_0),
    .O_3_0_1_1(n548_O_3_0_1_1),
    .O_3_0_1_2(n548_O_3_0_1_2),
    .O_3_0_2_0(n548_O_3_0_2_0),
    .O_3_0_2_1(n548_O_3_0_2_1),
    .O_3_0_2_2(n548_O_3_0_2_2),
    .O_4_0_0_0(n548_O_4_0_0_0),
    .O_4_0_0_1(n548_O_4_0_0_1),
    .O_4_0_0_2(n548_O_4_0_0_2),
    .O_4_0_1_0(n548_O_4_0_1_0),
    .O_4_0_1_1(n548_O_4_0_1_1),
    .O_4_0_1_2(n548_O_4_0_1_2),
    .O_4_0_2_0(n548_O_4_0_2_0),
    .O_4_0_2_1(n548_O_4_0_2_1),
    .O_4_0_2_2(n548_O_4_0_2_2),
    .O_5_0_0_0(n548_O_5_0_0_0),
    .O_5_0_0_1(n548_O_5_0_0_1),
    .O_5_0_0_2(n548_O_5_0_0_2),
    .O_5_0_1_0(n548_O_5_0_1_0),
    .O_5_0_1_1(n548_O_5_0_1_1),
    .O_5_0_1_2(n548_O_5_0_1_2),
    .O_5_0_2_0(n548_O_5_0_2_0),
    .O_5_0_2_1(n548_O_5_0_2_1),
    .O_5_0_2_2(n548_O_5_0_2_2),
    .O_6_0_0_0(n548_O_6_0_0_0),
    .O_6_0_0_1(n548_O_6_0_0_1),
    .O_6_0_0_2(n548_O_6_0_0_2),
    .O_6_0_1_0(n548_O_6_0_1_0),
    .O_6_0_1_1(n548_O_6_0_1_1),
    .O_6_0_1_2(n548_O_6_0_1_2),
    .O_6_0_2_0(n548_O_6_0_2_0),
    .O_6_0_2_1(n548_O_6_0_2_1),
    .O_6_0_2_2(n548_O_6_0_2_2),
    .O_7_0_0_0(n548_O_7_0_0_0),
    .O_7_0_0_1(n548_O_7_0_0_1),
    .O_7_0_0_2(n548_O_7_0_0_2),
    .O_7_0_1_0(n548_O_7_0_1_0),
    .O_7_0_1_1(n548_O_7_0_1_1),
    .O_7_0_1_2(n548_O_7_0_1_2),
    .O_7_0_2_0(n548_O_7_0_2_0),
    .O_7_0_2_1(n548_O_7_0_2_1),
    .O_7_0_2_2(n548_O_7_0_2_2)
  );
  MapT_7 n555 ( // @[Top.scala 873:22]
    .valid_up(n555_valid_up),
    .valid_down(n555_valid_down),
    .I_0_0_0_0(n555_I_0_0_0_0),
    .I_0_0_0_1(n555_I_0_0_0_1),
    .I_0_0_0_2(n555_I_0_0_0_2),
    .I_0_0_1_0(n555_I_0_0_1_0),
    .I_0_0_1_1(n555_I_0_0_1_1),
    .I_0_0_1_2(n555_I_0_0_1_2),
    .I_0_0_2_0(n555_I_0_0_2_0),
    .I_0_0_2_1(n555_I_0_0_2_1),
    .I_0_0_2_2(n555_I_0_0_2_2),
    .I_1_0_0_0(n555_I_1_0_0_0),
    .I_1_0_0_1(n555_I_1_0_0_1),
    .I_1_0_0_2(n555_I_1_0_0_2),
    .I_1_0_1_0(n555_I_1_0_1_0),
    .I_1_0_1_1(n555_I_1_0_1_1),
    .I_1_0_1_2(n555_I_1_0_1_2),
    .I_1_0_2_0(n555_I_1_0_2_0),
    .I_1_0_2_1(n555_I_1_0_2_1),
    .I_1_0_2_2(n555_I_1_0_2_2),
    .I_2_0_0_0(n555_I_2_0_0_0),
    .I_2_0_0_1(n555_I_2_0_0_1),
    .I_2_0_0_2(n555_I_2_0_0_2),
    .I_2_0_1_0(n555_I_2_0_1_0),
    .I_2_0_1_1(n555_I_2_0_1_1),
    .I_2_0_1_2(n555_I_2_0_1_2),
    .I_2_0_2_0(n555_I_2_0_2_0),
    .I_2_0_2_1(n555_I_2_0_2_1),
    .I_2_0_2_2(n555_I_2_0_2_2),
    .I_3_0_0_0(n555_I_3_0_0_0),
    .I_3_0_0_1(n555_I_3_0_0_1),
    .I_3_0_0_2(n555_I_3_0_0_2),
    .I_3_0_1_0(n555_I_3_0_1_0),
    .I_3_0_1_1(n555_I_3_0_1_1),
    .I_3_0_1_2(n555_I_3_0_1_2),
    .I_3_0_2_0(n555_I_3_0_2_0),
    .I_3_0_2_1(n555_I_3_0_2_1),
    .I_3_0_2_2(n555_I_3_0_2_2),
    .I_4_0_0_0(n555_I_4_0_0_0),
    .I_4_0_0_1(n555_I_4_0_0_1),
    .I_4_0_0_2(n555_I_4_0_0_2),
    .I_4_0_1_0(n555_I_4_0_1_0),
    .I_4_0_1_1(n555_I_4_0_1_1),
    .I_4_0_1_2(n555_I_4_0_1_2),
    .I_4_0_2_0(n555_I_4_0_2_0),
    .I_4_0_2_1(n555_I_4_0_2_1),
    .I_4_0_2_2(n555_I_4_0_2_2),
    .I_5_0_0_0(n555_I_5_0_0_0),
    .I_5_0_0_1(n555_I_5_0_0_1),
    .I_5_0_0_2(n555_I_5_0_0_2),
    .I_5_0_1_0(n555_I_5_0_1_0),
    .I_5_0_1_1(n555_I_5_0_1_1),
    .I_5_0_1_2(n555_I_5_0_1_2),
    .I_5_0_2_0(n555_I_5_0_2_0),
    .I_5_0_2_1(n555_I_5_0_2_1),
    .I_5_0_2_2(n555_I_5_0_2_2),
    .I_6_0_0_0(n555_I_6_0_0_0),
    .I_6_0_0_1(n555_I_6_0_0_1),
    .I_6_0_0_2(n555_I_6_0_0_2),
    .I_6_0_1_0(n555_I_6_0_1_0),
    .I_6_0_1_1(n555_I_6_0_1_1),
    .I_6_0_1_2(n555_I_6_0_1_2),
    .I_6_0_2_0(n555_I_6_0_2_0),
    .I_6_0_2_1(n555_I_6_0_2_1),
    .I_6_0_2_2(n555_I_6_0_2_2),
    .I_7_0_0_0(n555_I_7_0_0_0),
    .I_7_0_0_1(n555_I_7_0_0_1),
    .I_7_0_0_2(n555_I_7_0_0_2),
    .I_7_0_1_0(n555_I_7_0_1_0),
    .I_7_0_1_1(n555_I_7_0_1_1),
    .I_7_0_1_2(n555_I_7_0_1_2),
    .I_7_0_2_0(n555_I_7_0_2_0),
    .I_7_0_2_1(n555_I_7_0_2_1),
    .I_7_0_2_2(n555_I_7_0_2_2),
    .O_0_0_0(n555_O_0_0_0),
    .O_0_0_1(n555_O_0_0_1),
    .O_0_0_2(n555_O_0_0_2),
    .O_0_1_0(n555_O_0_1_0),
    .O_0_1_1(n555_O_0_1_1),
    .O_0_1_2(n555_O_0_1_2),
    .O_0_2_0(n555_O_0_2_0),
    .O_0_2_1(n555_O_0_2_1),
    .O_0_2_2(n555_O_0_2_2),
    .O_1_0_0(n555_O_1_0_0),
    .O_1_0_1(n555_O_1_0_1),
    .O_1_0_2(n555_O_1_0_2),
    .O_1_1_0(n555_O_1_1_0),
    .O_1_1_1(n555_O_1_1_1),
    .O_1_1_2(n555_O_1_1_2),
    .O_1_2_0(n555_O_1_2_0),
    .O_1_2_1(n555_O_1_2_1),
    .O_1_2_2(n555_O_1_2_2),
    .O_2_0_0(n555_O_2_0_0),
    .O_2_0_1(n555_O_2_0_1),
    .O_2_0_2(n555_O_2_0_2),
    .O_2_1_0(n555_O_2_1_0),
    .O_2_1_1(n555_O_2_1_1),
    .O_2_1_2(n555_O_2_1_2),
    .O_2_2_0(n555_O_2_2_0),
    .O_2_2_1(n555_O_2_2_1),
    .O_2_2_2(n555_O_2_2_2),
    .O_3_0_0(n555_O_3_0_0),
    .O_3_0_1(n555_O_3_0_1),
    .O_3_0_2(n555_O_3_0_2),
    .O_3_1_0(n555_O_3_1_0),
    .O_3_1_1(n555_O_3_1_1),
    .O_3_1_2(n555_O_3_1_2),
    .O_3_2_0(n555_O_3_2_0),
    .O_3_2_1(n555_O_3_2_1),
    .O_3_2_2(n555_O_3_2_2),
    .O_4_0_0(n555_O_4_0_0),
    .O_4_0_1(n555_O_4_0_1),
    .O_4_0_2(n555_O_4_0_2),
    .O_4_1_0(n555_O_4_1_0),
    .O_4_1_1(n555_O_4_1_1),
    .O_4_1_2(n555_O_4_1_2),
    .O_4_2_0(n555_O_4_2_0),
    .O_4_2_1(n555_O_4_2_1),
    .O_4_2_2(n555_O_4_2_2),
    .O_5_0_0(n555_O_5_0_0),
    .O_5_0_1(n555_O_5_0_1),
    .O_5_0_2(n555_O_5_0_2),
    .O_5_1_0(n555_O_5_1_0),
    .O_5_1_1(n555_O_5_1_1),
    .O_5_1_2(n555_O_5_1_2),
    .O_5_2_0(n555_O_5_2_0),
    .O_5_2_1(n555_O_5_2_1),
    .O_5_2_2(n555_O_5_2_2),
    .O_6_0_0(n555_O_6_0_0),
    .O_6_0_1(n555_O_6_0_1),
    .O_6_0_2(n555_O_6_0_2),
    .O_6_1_0(n555_O_6_1_0),
    .O_6_1_1(n555_O_6_1_1),
    .O_6_1_2(n555_O_6_1_2),
    .O_6_2_0(n555_O_6_2_0),
    .O_6_2_1(n555_O_6_2_1),
    .O_6_2_2(n555_O_6_2_2),
    .O_7_0_0(n555_O_7_0_0),
    .O_7_0_1(n555_O_7_0_1),
    .O_7_0_2(n555_O_7_0_2),
    .O_7_1_0(n555_O_7_1_0),
    .O_7_1_1(n555_O_7_1_1),
    .O_7_1_2(n555_O_7_1_2),
    .O_7_2_0(n555_O_7_2_0),
    .O_7_2_1(n555_O_7_2_1),
    .O_7_2_2(n555_O_7_2_2)
  );
  MapT_22 n597 ( // @[Top.scala 876:22]
    .clock(n597_clock),
    .reset(n597_reset),
    .valid_up(n597_valid_up),
    .valid_down(n597_valid_down),
    .I_0_0_0(n597_I_0_0_0),
    .I_0_0_1(n597_I_0_0_1),
    .I_0_0_2(n597_I_0_0_2),
    .I_0_1_0(n597_I_0_1_0),
    .I_0_1_1(n597_I_0_1_1),
    .I_0_1_2(n597_I_0_1_2),
    .I_0_2_0(n597_I_0_2_0),
    .I_0_2_1(n597_I_0_2_1),
    .I_0_2_2(n597_I_0_2_2),
    .I_1_0_0(n597_I_1_0_0),
    .I_1_0_1(n597_I_1_0_1),
    .I_1_0_2(n597_I_1_0_2),
    .I_1_1_0(n597_I_1_1_0),
    .I_1_1_1(n597_I_1_1_1),
    .I_1_1_2(n597_I_1_1_2),
    .I_1_2_0(n597_I_1_2_0),
    .I_1_2_1(n597_I_1_2_1),
    .I_1_2_2(n597_I_1_2_2),
    .I_2_0_0(n597_I_2_0_0),
    .I_2_0_1(n597_I_2_0_1),
    .I_2_0_2(n597_I_2_0_2),
    .I_2_1_0(n597_I_2_1_0),
    .I_2_1_1(n597_I_2_1_1),
    .I_2_1_2(n597_I_2_1_2),
    .I_2_2_0(n597_I_2_2_0),
    .I_2_2_1(n597_I_2_2_1),
    .I_2_2_2(n597_I_2_2_2),
    .I_3_0_0(n597_I_3_0_0),
    .I_3_0_1(n597_I_3_0_1),
    .I_3_0_2(n597_I_3_0_2),
    .I_3_1_0(n597_I_3_1_0),
    .I_3_1_1(n597_I_3_1_1),
    .I_3_1_2(n597_I_3_1_2),
    .I_3_2_0(n597_I_3_2_0),
    .I_3_2_1(n597_I_3_2_1),
    .I_3_2_2(n597_I_3_2_2),
    .I_4_0_0(n597_I_4_0_0),
    .I_4_0_1(n597_I_4_0_1),
    .I_4_0_2(n597_I_4_0_2),
    .I_4_1_0(n597_I_4_1_0),
    .I_4_1_1(n597_I_4_1_1),
    .I_4_1_2(n597_I_4_1_2),
    .I_4_2_0(n597_I_4_2_0),
    .I_4_2_1(n597_I_4_2_1),
    .I_4_2_2(n597_I_4_2_2),
    .I_5_0_0(n597_I_5_0_0),
    .I_5_0_1(n597_I_5_0_1),
    .I_5_0_2(n597_I_5_0_2),
    .I_5_1_0(n597_I_5_1_0),
    .I_5_1_1(n597_I_5_1_1),
    .I_5_1_2(n597_I_5_1_2),
    .I_5_2_0(n597_I_5_2_0),
    .I_5_2_1(n597_I_5_2_1),
    .I_5_2_2(n597_I_5_2_2),
    .I_6_0_0(n597_I_6_0_0),
    .I_6_0_1(n597_I_6_0_1),
    .I_6_0_2(n597_I_6_0_2),
    .I_6_1_0(n597_I_6_1_0),
    .I_6_1_1(n597_I_6_1_1),
    .I_6_1_2(n597_I_6_1_2),
    .I_6_2_0(n597_I_6_2_0),
    .I_6_2_1(n597_I_6_2_1),
    .I_6_2_2(n597_I_6_2_2),
    .I_7_0_0(n597_I_7_0_0),
    .I_7_0_1(n597_I_7_0_1),
    .I_7_0_2(n597_I_7_0_2),
    .I_7_1_0(n597_I_7_1_0),
    .I_7_1_1(n597_I_7_1_1),
    .I_7_1_2(n597_I_7_1_2),
    .I_7_2_0(n597_I_7_2_0),
    .I_7_2_1(n597_I_7_2_1),
    .I_7_2_2(n597_I_7_2_2),
    .O_0_0_0(n597_O_0_0_0),
    .O_1_0_0(n597_O_1_0_0),
    .O_2_0_0(n597_O_2_0_0),
    .O_3_0_0(n597_O_3_0_0),
    .O_4_0_0(n597_O_4_0_0),
    .O_5_0_0(n597_O_5_0_0),
    .O_6_0_0(n597_O_6_0_0),
    .O_7_0_0(n597_O_7_0_0)
  );
  Passthrough_4 n598 ( // @[Top.scala 879:22]
    .valid_up(n598_valid_up),
    .valid_down(n598_valid_down),
    .I_0_0_0(n598_I_0_0_0),
    .I_1_0_0(n598_I_1_0_0),
    .I_2_0_0(n598_I_2_0_0),
    .I_3_0_0(n598_I_3_0_0),
    .I_4_0_0(n598_I_4_0_0),
    .I_5_0_0(n598_I_5_0_0),
    .I_6_0_0(n598_I_6_0_0),
    .I_7_0_0(n598_I_7_0_0),
    .O_0_0(n598_O_0_0),
    .O_1_0(n598_O_1_0),
    .O_2_0(n598_O_2_0),
    .O_3_0(n598_O_3_0),
    .O_4_0(n598_O_4_0),
    .O_5_0(n598_O_5_0),
    .O_6_0(n598_O_6_0),
    .O_7_0(n598_O_7_0)
  );
  Passthrough_5 n599 ( // @[Top.scala 882:22]
    .valid_up(n599_valid_up),
    .valid_down(n599_valid_down),
    .I_0_0(n599_I_0_0),
    .I_1_0(n599_I_1_0),
    .I_2_0(n599_I_2_0),
    .I_3_0(n599_I_3_0),
    .I_4_0(n599_I_4_0),
    .I_5_0(n599_I_5_0),
    .I_6_0(n599_I_6_0),
    .I_7_0(n599_I_7_0),
    .O_0(n599_O_0),
    .O_1(n599_O_1),
    .O_2(n599_O_2),
    .O_3(n599_O_3),
    .O_4(n599_O_4),
    .O_5(n599_O_5),
    .O_6(n599_O_6),
    .O_7(n599_O_7)
  );
  FIFO_9 n600 ( // @[Top.scala 885:22]
    .clock(n600_clock),
    .reset(n600_reset),
    .valid_up(n600_valid_up),
    .valid_down(n600_valid_down),
    .I_0(n600_I_0),
    .I_1(n600_I_1),
    .I_2(n600_I_2),
    .I_3(n600_I_3),
    .I_4(n600_I_4),
    .I_5(n600_I_5),
    .I_6(n600_I_6),
    .I_7(n600_I_7),
    .O_0(n600_O_0),
    .O_1(n600_O_1),
    .O_2(n600_O_2),
    .O_3(n600_O_3),
    .O_4(n600_O_4),
    .O_5(n600_O_5),
    .O_6(n600_O_6),
    .O_7(n600_O_7)
  );
  Map2T_18 n601 ( // @[Top.scala 888:22]
    .clock(n601_clock),
    .reset(n601_reset),
    .valid_up(n601_valid_up),
    .valid_down(n601_valid_down),
    .I0_0(n601_I0_0),
    .I0_1(n601_I0_1),
    .I0_2(n601_I0_2),
    .I0_3(n601_I0_3),
    .I0_4(n601_I0_4),
    .I0_5(n601_I0_5),
    .I0_6(n601_I0_6),
    .I0_7(n601_I0_7),
    .I1_0(n601_I1_0),
    .I1_1(n601_I1_1),
    .I1_2(n601_I1_2),
    .I1_3(n601_I1_3),
    .I1_4(n601_I1_4),
    .I1_5(n601_I1_5),
    .I1_6(n601_I1_6),
    .I1_7(n601_I1_7),
    .O_0(n601_O_0),
    .O_1(n601_O_1),
    .O_2(n601_O_2),
    .O_3(n601_O_3),
    .O_4(n601_O_4),
    .O_5(n601_O_5),
    .O_6(n601_O_6),
    .O_7(n601_O_7)
  );
  MapT_23 n637 ( // @[Top.scala 892:22]
    .valid_up(n637_valid_up),
    .valid_down(n637_valid_down),
    .I_0_t1b_t0b(n637_I_0_t1b_t0b),
    .I_0_t1b_t1b(n637_I_0_t1b_t1b),
    .I_1_t1b_t0b(n637_I_1_t1b_t0b),
    .I_1_t1b_t1b(n637_I_1_t1b_t1b),
    .I_2_t1b_t0b(n637_I_2_t1b_t0b),
    .I_2_t1b_t1b(n637_I_2_t1b_t1b),
    .I_3_t1b_t0b(n637_I_3_t1b_t0b),
    .I_3_t1b_t1b(n637_I_3_t1b_t1b),
    .I_4_t1b_t0b(n637_I_4_t1b_t0b),
    .I_4_t1b_t1b(n637_I_4_t1b_t1b),
    .I_5_t1b_t0b(n637_I_5_t1b_t0b),
    .I_5_t1b_t1b(n637_I_5_t1b_t1b),
    .I_6_t1b_t0b(n637_I_6_t1b_t0b),
    .I_6_t1b_t1b(n637_I_6_t1b_t1b),
    .I_7_t1b_t0b(n637_I_7_t1b_t0b),
    .I_7_t1b_t1b(n637_I_7_t1b_t1b),
    .O_0(n637_O_0),
    .O_1(n637_O_1),
    .O_2(n637_O_2),
    .O_3(n637_O_3),
    .O_4(n637_O_4),
    .O_5(n637_O_5),
    .O_6(n637_O_6),
    .O_7(n637_O_7)
  );
  ShiftTS n638 ( // @[Top.scala 895:22]
    .clock(n638_clock),
    .reset(n638_reset),
    .valid_up(n638_valid_up),
    .valid_down(n638_valid_down),
    .I_0(n638_I_0),
    .I_1(n638_I_1),
    .I_2(n638_I_2),
    .I_3(n638_I_3),
    .I_4(n638_I_4),
    .I_5(n638_I_5),
    .I_6(n638_I_6),
    .I_7(n638_I_7),
    .O_0(n638_O_0),
    .O_1(n638_O_1),
    .O_2(n638_O_2),
    .O_3(n638_O_3),
    .O_4(n638_O_4),
    .O_5(n638_O_5),
    .O_6(n638_O_6),
    .O_7(n638_O_7)
  );
  ShiftTS n639 ( // @[Top.scala 898:22]
    .clock(n639_clock),
    .reset(n639_reset),
    .valid_up(n639_valid_up),
    .valid_down(n639_valid_down),
    .I_0(n639_I_0),
    .I_1(n639_I_1),
    .I_2(n639_I_2),
    .I_3(n639_I_3),
    .I_4(n639_I_4),
    .I_5(n639_I_5),
    .I_6(n639_I_6),
    .I_7(n639_I_7),
    .O_0(n639_O_0),
    .O_1(n639_O_1),
    .O_2(n639_O_2),
    .O_3(n639_O_3),
    .O_4(n639_O_4),
    .O_5(n639_O_5),
    .O_6(n639_O_6),
    .O_7(n639_O_7)
  );
  ShiftTS_2 n640 ( // @[Top.scala 901:22]
    .clock(n640_clock),
    .valid_up(n640_valid_up),
    .valid_down(n640_valid_down),
    .I_0(n640_I_0),
    .I_1(n640_I_1),
    .I_2(n640_I_2),
    .I_3(n640_I_3),
    .I_4(n640_I_4),
    .I_5(n640_I_5),
    .I_6(n640_I_6),
    .I_7(n640_I_7),
    .O_0(n640_O_0),
    .O_1(n640_O_1),
    .O_2(n640_O_2),
    .O_3(n640_O_3),
    .O_4(n640_O_4),
    .O_5(n640_O_5),
    .O_6(n640_O_6),
    .O_7(n640_O_7)
  );
  ShiftTS_2 n641 ( // @[Top.scala 904:22]
    .clock(n641_clock),
    .valid_up(n641_valid_up),
    .valid_down(n641_valid_down),
    .I_0(n641_I_0),
    .I_1(n641_I_1),
    .I_2(n641_I_2),
    .I_3(n641_I_3),
    .I_4(n641_I_4),
    .I_5(n641_I_5),
    .I_6(n641_I_6),
    .I_7(n641_I_7),
    .O_0(n641_O_0),
    .O_1(n641_O_1),
    .O_2(n641_O_2),
    .O_3(n641_O_3),
    .O_4(n641_O_4),
    .O_5(n641_O_5),
    .O_6(n641_O_6),
    .O_7(n641_O_7)
  );
  Map2T n642 ( // @[Top.scala 907:22]
    .valid_up(n642_valid_up),
    .valid_down(n642_valid_down),
    .I0_0(n642_I0_0),
    .I0_1(n642_I0_1),
    .I0_2(n642_I0_2),
    .I0_3(n642_I0_3),
    .I0_4(n642_I0_4),
    .I0_5(n642_I0_5),
    .I0_6(n642_I0_6),
    .I0_7(n642_I0_7),
    .I1_0(n642_I1_0),
    .I1_1(n642_I1_1),
    .I1_2(n642_I1_2),
    .I1_3(n642_I1_3),
    .I1_4(n642_I1_4),
    .I1_5(n642_I1_5),
    .I1_6(n642_I1_6),
    .I1_7(n642_I1_7),
    .O_0_0(n642_O_0_0),
    .O_0_1(n642_O_0_1),
    .O_1_0(n642_O_1_0),
    .O_1_1(n642_O_1_1),
    .O_2_0(n642_O_2_0),
    .O_2_1(n642_O_2_1),
    .O_3_0(n642_O_3_0),
    .O_3_1(n642_O_3_1),
    .O_4_0(n642_O_4_0),
    .O_4_1(n642_O_4_1),
    .O_5_0(n642_O_5_0),
    .O_5_1(n642_O_5_1),
    .O_6_0(n642_O_6_0),
    .O_6_1(n642_O_6_1),
    .O_7_0(n642_O_7_0),
    .O_7_1(n642_O_7_1)
  );
  Map2T_1 n649 ( // @[Top.scala 911:22]
    .valid_up(n649_valid_up),
    .valid_down(n649_valid_down),
    .I0_0_0(n649_I0_0_0),
    .I0_0_1(n649_I0_0_1),
    .I0_1_0(n649_I0_1_0),
    .I0_1_1(n649_I0_1_1),
    .I0_2_0(n649_I0_2_0),
    .I0_2_1(n649_I0_2_1),
    .I0_3_0(n649_I0_3_0),
    .I0_3_1(n649_I0_3_1),
    .I0_4_0(n649_I0_4_0),
    .I0_4_1(n649_I0_4_1),
    .I0_5_0(n649_I0_5_0),
    .I0_5_1(n649_I0_5_1),
    .I0_6_0(n649_I0_6_0),
    .I0_6_1(n649_I0_6_1),
    .I0_7_0(n649_I0_7_0),
    .I0_7_1(n649_I0_7_1),
    .I1_0(n649_I1_0),
    .I1_1(n649_I1_1),
    .I1_2(n649_I1_2),
    .I1_3(n649_I1_3),
    .I1_4(n649_I1_4),
    .I1_5(n649_I1_5),
    .I1_6(n649_I1_6),
    .I1_7(n649_I1_7),
    .O_0_0(n649_O_0_0),
    .O_0_1(n649_O_0_1),
    .O_0_2(n649_O_0_2),
    .O_1_0(n649_O_1_0),
    .O_1_1(n649_O_1_1),
    .O_1_2(n649_O_1_2),
    .O_2_0(n649_O_2_0),
    .O_2_1(n649_O_2_1),
    .O_2_2(n649_O_2_2),
    .O_3_0(n649_O_3_0),
    .O_3_1(n649_O_3_1),
    .O_3_2(n649_O_3_2),
    .O_4_0(n649_O_4_0),
    .O_4_1(n649_O_4_1),
    .O_4_2(n649_O_4_2),
    .O_5_0(n649_O_5_0),
    .O_5_1(n649_O_5_1),
    .O_5_2(n649_O_5_2),
    .O_6_0(n649_O_6_0),
    .O_6_1(n649_O_6_1),
    .O_6_2(n649_O_6_2),
    .O_7_0(n649_O_7_0),
    .O_7_1(n649_O_7_1),
    .O_7_2(n649_O_7_2)
  );
  MapT n658 ( // @[Top.scala 915:22]
    .valid_up(n658_valid_up),
    .valid_down(n658_valid_down),
    .I_0_0(n658_I_0_0),
    .I_0_1(n658_I_0_1),
    .I_0_2(n658_I_0_2),
    .I_1_0(n658_I_1_0),
    .I_1_1(n658_I_1_1),
    .I_1_2(n658_I_1_2),
    .I_2_0(n658_I_2_0),
    .I_2_1(n658_I_2_1),
    .I_2_2(n658_I_2_2),
    .I_3_0(n658_I_3_0),
    .I_3_1(n658_I_3_1),
    .I_3_2(n658_I_3_2),
    .I_4_0(n658_I_4_0),
    .I_4_1(n658_I_4_1),
    .I_4_2(n658_I_4_2),
    .I_5_0(n658_I_5_0),
    .I_5_1(n658_I_5_1),
    .I_5_2(n658_I_5_2),
    .I_6_0(n658_I_6_0),
    .I_6_1(n658_I_6_1),
    .I_6_2(n658_I_6_2),
    .I_7_0(n658_I_7_0),
    .I_7_1(n658_I_7_1),
    .I_7_2(n658_I_7_2),
    .O_0_0_0(n658_O_0_0_0),
    .O_0_0_1(n658_O_0_0_1),
    .O_0_0_2(n658_O_0_0_2),
    .O_1_0_0(n658_O_1_0_0),
    .O_1_0_1(n658_O_1_0_1),
    .O_1_0_2(n658_O_1_0_2),
    .O_2_0_0(n658_O_2_0_0),
    .O_2_0_1(n658_O_2_0_1),
    .O_2_0_2(n658_O_2_0_2),
    .O_3_0_0(n658_O_3_0_0),
    .O_3_0_1(n658_O_3_0_1),
    .O_3_0_2(n658_O_3_0_2),
    .O_4_0_0(n658_O_4_0_0),
    .O_4_0_1(n658_O_4_0_1),
    .O_4_0_2(n658_O_4_0_2),
    .O_5_0_0(n658_O_5_0_0),
    .O_5_0_1(n658_O_5_0_1),
    .O_5_0_2(n658_O_5_0_2),
    .O_6_0_0(n658_O_6_0_0),
    .O_6_0_1(n658_O_6_0_1),
    .O_6_0_2(n658_O_6_0_2),
    .O_7_0_0(n658_O_7_0_0),
    .O_7_0_1(n658_O_7_0_1),
    .O_7_0_2(n658_O_7_0_2)
  );
  MapT_1 n665 ( // @[Top.scala 918:22]
    .valid_up(n665_valid_up),
    .valid_down(n665_valid_down),
    .I_0_0_0(n665_I_0_0_0),
    .I_0_0_1(n665_I_0_0_1),
    .I_0_0_2(n665_I_0_0_2),
    .I_1_0_0(n665_I_1_0_0),
    .I_1_0_1(n665_I_1_0_1),
    .I_1_0_2(n665_I_1_0_2),
    .I_2_0_0(n665_I_2_0_0),
    .I_2_0_1(n665_I_2_0_1),
    .I_2_0_2(n665_I_2_0_2),
    .I_3_0_0(n665_I_3_0_0),
    .I_3_0_1(n665_I_3_0_1),
    .I_3_0_2(n665_I_3_0_2),
    .I_4_0_0(n665_I_4_0_0),
    .I_4_0_1(n665_I_4_0_1),
    .I_4_0_2(n665_I_4_0_2),
    .I_5_0_0(n665_I_5_0_0),
    .I_5_0_1(n665_I_5_0_1),
    .I_5_0_2(n665_I_5_0_2),
    .I_6_0_0(n665_I_6_0_0),
    .I_6_0_1(n665_I_6_0_1),
    .I_6_0_2(n665_I_6_0_2),
    .I_7_0_0(n665_I_7_0_0),
    .I_7_0_1(n665_I_7_0_1),
    .I_7_0_2(n665_I_7_0_2),
    .O_0_0(n665_O_0_0),
    .O_0_1(n665_O_0_1),
    .O_0_2(n665_O_0_2),
    .O_1_0(n665_O_1_0),
    .O_1_1(n665_O_1_1),
    .O_1_2(n665_O_1_2),
    .O_2_0(n665_O_2_0),
    .O_2_1(n665_O_2_1),
    .O_2_2(n665_O_2_2),
    .O_3_0(n665_O_3_0),
    .O_3_1(n665_O_3_1),
    .O_3_2(n665_O_3_2),
    .O_4_0(n665_O_4_0),
    .O_4_1(n665_O_4_1),
    .O_4_2(n665_O_4_2),
    .O_5_0(n665_O_5_0),
    .O_5_1(n665_O_5_1),
    .O_5_2(n665_O_5_2),
    .O_6_0(n665_O_6_0),
    .O_6_1(n665_O_6_1),
    .O_6_2(n665_O_6_2),
    .O_7_0(n665_O_7_0),
    .O_7_1(n665_O_7_1),
    .O_7_2(n665_O_7_2)
  );
  ShiftTS_2 n666 ( // @[Top.scala 921:22]
    .clock(n666_clock),
    .valid_up(n666_valid_up),
    .valid_down(n666_valid_down),
    .I_0(n666_I_0),
    .I_1(n666_I_1),
    .I_2(n666_I_2),
    .I_3(n666_I_3),
    .I_4(n666_I_4),
    .I_5(n666_I_5),
    .I_6(n666_I_6),
    .I_7(n666_I_7),
    .O_0(n666_O_0),
    .O_1(n666_O_1),
    .O_2(n666_O_2),
    .O_3(n666_O_3),
    .O_4(n666_O_4),
    .O_5(n666_O_5),
    .O_6(n666_O_6),
    .O_7(n666_O_7)
  );
  ShiftTS_2 n667 ( // @[Top.scala 924:22]
    .clock(n667_clock),
    .valid_up(n667_valid_up),
    .valid_down(n667_valid_down),
    .I_0(n667_I_0),
    .I_1(n667_I_1),
    .I_2(n667_I_2),
    .I_3(n667_I_3),
    .I_4(n667_I_4),
    .I_5(n667_I_5),
    .I_6(n667_I_6),
    .I_7(n667_I_7),
    .O_0(n667_O_0),
    .O_1(n667_O_1),
    .O_2(n667_O_2),
    .O_3(n667_O_3),
    .O_4(n667_O_4),
    .O_5(n667_O_5),
    .O_6(n667_O_6),
    .O_7(n667_O_7)
  );
  Map2T n668 ( // @[Top.scala 927:22]
    .valid_up(n668_valid_up),
    .valid_down(n668_valid_down),
    .I0_0(n668_I0_0),
    .I0_1(n668_I0_1),
    .I0_2(n668_I0_2),
    .I0_3(n668_I0_3),
    .I0_4(n668_I0_4),
    .I0_5(n668_I0_5),
    .I0_6(n668_I0_6),
    .I0_7(n668_I0_7),
    .I1_0(n668_I1_0),
    .I1_1(n668_I1_1),
    .I1_2(n668_I1_2),
    .I1_3(n668_I1_3),
    .I1_4(n668_I1_4),
    .I1_5(n668_I1_5),
    .I1_6(n668_I1_6),
    .I1_7(n668_I1_7),
    .O_0_0(n668_O_0_0),
    .O_0_1(n668_O_0_1),
    .O_1_0(n668_O_1_0),
    .O_1_1(n668_O_1_1),
    .O_2_0(n668_O_2_0),
    .O_2_1(n668_O_2_1),
    .O_3_0(n668_O_3_0),
    .O_3_1(n668_O_3_1),
    .O_4_0(n668_O_4_0),
    .O_4_1(n668_O_4_1),
    .O_5_0(n668_O_5_0),
    .O_5_1(n668_O_5_1),
    .O_6_0(n668_O_6_0),
    .O_6_1(n668_O_6_1),
    .O_7_0(n668_O_7_0),
    .O_7_1(n668_O_7_1)
  );
  Map2T_1 n675 ( // @[Top.scala 931:22]
    .valid_up(n675_valid_up),
    .valid_down(n675_valid_down),
    .I0_0_0(n675_I0_0_0),
    .I0_0_1(n675_I0_0_1),
    .I0_1_0(n675_I0_1_0),
    .I0_1_1(n675_I0_1_1),
    .I0_2_0(n675_I0_2_0),
    .I0_2_1(n675_I0_2_1),
    .I0_3_0(n675_I0_3_0),
    .I0_3_1(n675_I0_3_1),
    .I0_4_0(n675_I0_4_0),
    .I0_4_1(n675_I0_4_1),
    .I0_5_0(n675_I0_5_0),
    .I0_5_1(n675_I0_5_1),
    .I0_6_0(n675_I0_6_0),
    .I0_6_1(n675_I0_6_1),
    .I0_7_0(n675_I0_7_0),
    .I0_7_1(n675_I0_7_1),
    .I1_0(n675_I1_0),
    .I1_1(n675_I1_1),
    .I1_2(n675_I1_2),
    .I1_3(n675_I1_3),
    .I1_4(n675_I1_4),
    .I1_5(n675_I1_5),
    .I1_6(n675_I1_6),
    .I1_7(n675_I1_7),
    .O_0_0(n675_O_0_0),
    .O_0_1(n675_O_0_1),
    .O_0_2(n675_O_0_2),
    .O_1_0(n675_O_1_0),
    .O_1_1(n675_O_1_1),
    .O_1_2(n675_O_1_2),
    .O_2_0(n675_O_2_0),
    .O_2_1(n675_O_2_1),
    .O_2_2(n675_O_2_2),
    .O_3_0(n675_O_3_0),
    .O_3_1(n675_O_3_1),
    .O_3_2(n675_O_3_2),
    .O_4_0(n675_O_4_0),
    .O_4_1(n675_O_4_1),
    .O_4_2(n675_O_4_2),
    .O_5_0(n675_O_5_0),
    .O_5_1(n675_O_5_1),
    .O_5_2(n675_O_5_2),
    .O_6_0(n675_O_6_0),
    .O_6_1(n675_O_6_1),
    .O_6_2(n675_O_6_2),
    .O_7_0(n675_O_7_0),
    .O_7_1(n675_O_7_1),
    .O_7_2(n675_O_7_2)
  );
  MapT n684 ( // @[Top.scala 935:22]
    .valid_up(n684_valid_up),
    .valid_down(n684_valid_down),
    .I_0_0(n684_I_0_0),
    .I_0_1(n684_I_0_1),
    .I_0_2(n684_I_0_2),
    .I_1_0(n684_I_1_0),
    .I_1_1(n684_I_1_1),
    .I_1_2(n684_I_1_2),
    .I_2_0(n684_I_2_0),
    .I_2_1(n684_I_2_1),
    .I_2_2(n684_I_2_2),
    .I_3_0(n684_I_3_0),
    .I_3_1(n684_I_3_1),
    .I_3_2(n684_I_3_2),
    .I_4_0(n684_I_4_0),
    .I_4_1(n684_I_4_1),
    .I_4_2(n684_I_4_2),
    .I_5_0(n684_I_5_0),
    .I_5_1(n684_I_5_1),
    .I_5_2(n684_I_5_2),
    .I_6_0(n684_I_6_0),
    .I_6_1(n684_I_6_1),
    .I_6_2(n684_I_6_2),
    .I_7_0(n684_I_7_0),
    .I_7_1(n684_I_7_1),
    .I_7_2(n684_I_7_2),
    .O_0_0_0(n684_O_0_0_0),
    .O_0_0_1(n684_O_0_0_1),
    .O_0_0_2(n684_O_0_0_2),
    .O_1_0_0(n684_O_1_0_0),
    .O_1_0_1(n684_O_1_0_1),
    .O_1_0_2(n684_O_1_0_2),
    .O_2_0_0(n684_O_2_0_0),
    .O_2_0_1(n684_O_2_0_1),
    .O_2_0_2(n684_O_2_0_2),
    .O_3_0_0(n684_O_3_0_0),
    .O_3_0_1(n684_O_3_0_1),
    .O_3_0_2(n684_O_3_0_2),
    .O_4_0_0(n684_O_4_0_0),
    .O_4_0_1(n684_O_4_0_1),
    .O_4_0_2(n684_O_4_0_2),
    .O_5_0_0(n684_O_5_0_0),
    .O_5_0_1(n684_O_5_0_1),
    .O_5_0_2(n684_O_5_0_2),
    .O_6_0_0(n684_O_6_0_0),
    .O_6_0_1(n684_O_6_0_1),
    .O_6_0_2(n684_O_6_0_2),
    .O_7_0_0(n684_O_7_0_0),
    .O_7_0_1(n684_O_7_0_1),
    .O_7_0_2(n684_O_7_0_2)
  );
  MapT_1 n691 ( // @[Top.scala 938:22]
    .valid_up(n691_valid_up),
    .valid_down(n691_valid_down),
    .I_0_0_0(n691_I_0_0_0),
    .I_0_0_1(n691_I_0_0_1),
    .I_0_0_2(n691_I_0_0_2),
    .I_1_0_0(n691_I_1_0_0),
    .I_1_0_1(n691_I_1_0_1),
    .I_1_0_2(n691_I_1_0_2),
    .I_2_0_0(n691_I_2_0_0),
    .I_2_0_1(n691_I_2_0_1),
    .I_2_0_2(n691_I_2_0_2),
    .I_3_0_0(n691_I_3_0_0),
    .I_3_0_1(n691_I_3_0_1),
    .I_3_0_2(n691_I_3_0_2),
    .I_4_0_0(n691_I_4_0_0),
    .I_4_0_1(n691_I_4_0_1),
    .I_4_0_2(n691_I_4_0_2),
    .I_5_0_0(n691_I_5_0_0),
    .I_5_0_1(n691_I_5_0_1),
    .I_5_0_2(n691_I_5_0_2),
    .I_6_0_0(n691_I_6_0_0),
    .I_6_0_1(n691_I_6_0_1),
    .I_6_0_2(n691_I_6_0_2),
    .I_7_0_0(n691_I_7_0_0),
    .I_7_0_1(n691_I_7_0_1),
    .I_7_0_2(n691_I_7_0_2),
    .O_0_0(n691_O_0_0),
    .O_0_1(n691_O_0_1),
    .O_0_2(n691_O_0_2),
    .O_1_0(n691_O_1_0),
    .O_1_1(n691_O_1_1),
    .O_1_2(n691_O_1_2),
    .O_2_0(n691_O_2_0),
    .O_2_1(n691_O_2_1),
    .O_2_2(n691_O_2_2),
    .O_3_0(n691_O_3_0),
    .O_3_1(n691_O_3_1),
    .O_3_2(n691_O_3_2),
    .O_4_0(n691_O_4_0),
    .O_4_1(n691_O_4_1),
    .O_4_2(n691_O_4_2),
    .O_5_0(n691_O_5_0),
    .O_5_1(n691_O_5_1),
    .O_5_2(n691_O_5_2),
    .O_6_0(n691_O_6_0),
    .O_6_1(n691_O_6_1),
    .O_6_2(n691_O_6_2),
    .O_7_0(n691_O_7_0),
    .O_7_1(n691_O_7_1),
    .O_7_2(n691_O_7_2)
  );
  Map2T_4 n692 ( // @[Top.scala 941:22]
    .valid_up(n692_valid_up),
    .valid_down(n692_valid_down),
    .I0_0_0(n692_I0_0_0),
    .I0_0_1(n692_I0_0_1),
    .I0_0_2(n692_I0_0_2),
    .I0_1_0(n692_I0_1_0),
    .I0_1_1(n692_I0_1_1),
    .I0_1_2(n692_I0_1_2),
    .I0_2_0(n692_I0_2_0),
    .I0_2_1(n692_I0_2_1),
    .I0_2_2(n692_I0_2_2),
    .I0_3_0(n692_I0_3_0),
    .I0_3_1(n692_I0_3_1),
    .I0_3_2(n692_I0_3_2),
    .I0_4_0(n692_I0_4_0),
    .I0_4_1(n692_I0_4_1),
    .I0_4_2(n692_I0_4_2),
    .I0_5_0(n692_I0_5_0),
    .I0_5_1(n692_I0_5_1),
    .I0_5_2(n692_I0_5_2),
    .I0_6_0(n692_I0_6_0),
    .I0_6_1(n692_I0_6_1),
    .I0_6_2(n692_I0_6_2),
    .I0_7_0(n692_I0_7_0),
    .I0_7_1(n692_I0_7_1),
    .I0_7_2(n692_I0_7_2),
    .I1_0_0(n692_I1_0_0),
    .I1_0_1(n692_I1_0_1),
    .I1_0_2(n692_I1_0_2),
    .I1_1_0(n692_I1_1_0),
    .I1_1_1(n692_I1_1_1),
    .I1_1_2(n692_I1_1_2),
    .I1_2_0(n692_I1_2_0),
    .I1_2_1(n692_I1_2_1),
    .I1_2_2(n692_I1_2_2),
    .I1_3_0(n692_I1_3_0),
    .I1_3_1(n692_I1_3_1),
    .I1_3_2(n692_I1_3_2),
    .I1_4_0(n692_I1_4_0),
    .I1_4_1(n692_I1_4_1),
    .I1_4_2(n692_I1_4_2),
    .I1_5_0(n692_I1_5_0),
    .I1_5_1(n692_I1_5_1),
    .I1_5_2(n692_I1_5_2),
    .I1_6_0(n692_I1_6_0),
    .I1_6_1(n692_I1_6_1),
    .I1_6_2(n692_I1_6_2),
    .I1_7_0(n692_I1_7_0),
    .I1_7_1(n692_I1_7_1),
    .I1_7_2(n692_I1_7_2),
    .O_0_0_0(n692_O_0_0_0),
    .O_0_0_1(n692_O_0_0_1),
    .O_0_0_2(n692_O_0_0_2),
    .O_0_1_0(n692_O_0_1_0),
    .O_0_1_1(n692_O_0_1_1),
    .O_0_1_2(n692_O_0_1_2),
    .O_1_0_0(n692_O_1_0_0),
    .O_1_0_1(n692_O_1_0_1),
    .O_1_0_2(n692_O_1_0_2),
    .O_1_1_0(n692_O_1_1_0),
    .O_1_1_1(n692_O_1_1_1),
    .O_1_1_2(n692_O_1_1_2),
    .O_2_0_0(n692_O_2_0_0),
    .O_2_0_1(n692_O_2_0_1),
    .O_2_0_2(n692_O_2_0_2),
    .O_2_1_0(n692_O_2_1_0),
    .O_2_1_1(n692_O_2_1_1),
    .O_2_1_2(n692_O_2_1_2),
    .O_3_0_0(n692_O_3_0_0),
    .O_3_0_1(n692_O_3_0_1),
    .O_3_0_2(n692_O_3_0_2),
    .O_3_1_0(n692_O_3_1_0),
    .O_3_1_1(n692_O_3_1_1),
    .O_3_1_2(n692_O_3_1_2),
    .O_4_0_0(n692_O_4_0_0),
    .O_4_0_1(n692_O_4_0_1),
    .O_4_0_2(n692_O_4_0_2),
    .O_4_1_0(n692_O_4_1_0),
    .O_4_1_1(n692_O_4_1_1),
    .O_4_1_2(n692_O_4_1_2),
    .O_5_0_0(n692_O_5_0_0),
    .O_5_0_1(n692_O_5_0_1),
    .O_5_0_2(n692_O_5_0_2),
    .O_5_1_0(n692_O_5_1_0),
    .O_5_1_1(n692_O_5_1_1),
    .O_5_1_2(n692_O_5_1_2),
    .O_6_0_0(n692_O_6_0_0),
    .O_6_0_1(n692_O_6_0_1),
    .O_6_0_2(n692_O_6_0_2),
    .O_6_1_0(n692_O_6_1_0),
    .O_6_1_1(n692_O_6_1_1),
    .O_6_1_2(n692_O_6_1_2),
    .O_7_0_0(n692_O_7_0_0),
    .O_7_0_1(n692_O_7_0_1),
    .O_7_0_2(n692_O_7_0_2),
    .O_7_1_0(n692_O_7_1_0),
    .O_7_1_1(n692_O_7_1_1),
    .O_7_1_2(n692_O_7_1_2)
  );
  ShiftTS_2 n699 ( // @[Top.scala 945:22]
    .clock(n699_clock),
    .valid_up(n699_valid_up),
    .valid_down(n699_valid_down),
    .I_0(n699_I_0),
    .I_1(n699_I_1),
    .I_2(n699_I_2),
    .I_3(n699_I_3),
    .I_4(n699_I_4),
    .I_5(n699_I_5),
    .I_6(n699_I_6),
    .I_7(n699_I_7),
    .O_0(n699_O_0),
    .O_1(n699_O_1),
    .O_2(n699_O_2),
    .O_3(n699_O_3),
    .O_4(n699_O_4),
    .O_5(n699_O_5),
    .O_6(n699_O_6),
    .O_7(n699_O_7)
  );
  ShiftTS_2 n700 ( // @[Top.scala 948:22]
    .clock(n700_clock),
    .valid_up(n700_valid_up),
    .valid_down(n700_valid_down),
    .I_0(n700_I_0),
    .I_1(n700_I_1),
    .I_2(n700_I_2),
    .I_3(n700_I_3),
    .I_4(n700_I_4),
    .I_5(n700_I_5),
    .I_6(n700_I_6),
    .I_7(n700_I_7),
    .O_0(n700_O_0),
    .O_1(n700_O_1),
    .O_2(n700_O_2),
    .O_3(n700_O_3),
    .O_4(n700_O_4),
    .O_5(n700_O_5),
    .O_6(n700_O_6),
    .O_7(n700_O_7)
  );
  Map2T n701 ( // @[Top.scala 951:22]
    .valid_up(n701_valid_up),
    .valid_down(n701_valid_down),
    .I0_0(n701_I0_0),
    .I0_1(n701_I0_1),
    .I0_2(n701_I0_2),
    .I0_3(n701_I0_3),
    .I0_4(n701_I0_4),
    .I0_5(n701_I0_5),
    .I0_6(n701_I0_6),
    .I0_7(n701_I0_7),
    .I1_0(n701_I1_0),
    .I1_1(n701_I1_1),
    .I1_2(n701_I1_2),
    .I1_3(n701_I1_3),
    .I1_4(n701_I1_4),
    .I1_5(n701_I1_5),
    .I1_6(n701_I1_6),
    .I1_7(n701_I1_7),
    .O_0_0(n701_O_0_0),
    .O_0_1(n701_O_0_1),
    .O_1_0(n701_O_1_0),
    .O_1_1(n701_O_1_1),
    .O_2_0(n701_O_2_0),
    .O_2_1(n701_O_2_1),
    .O_3_0(n701_O_3_0),
    .O_3_1(n701_O_3_1),
    .O_4_0(n701_O_4_0),
    .O_4_1(n701_O_4_1),
    .O_5_0(n701_O_5_0),
    .O_5_1(n701_O_5_1),
    .O_6_0(n701_O_6_0),
    .O_6_1(n701_O_6_1),
    .O_7_0(n701_O_7_0),
    .O_7_1(n701_O_7_1)
  );
  Map2T_1 n708 ( // @[Top.scala 955:22]
    .valid_up(n708_valid_up),
    .valid_down(n708_valid_down),
    .I0_0_0(n708_I0_0_0),
    .I0_0_1(n708_I0_0_1),
    .I0_1_0(n708_I0_1_0),
    .I0_1_1(n708_I0_1_1),
    .I0_2_0(n708_I0_2_0),
    .I0_2_1(n708_I0_2_1),
    .I0_3_0(n708_I0_3_0),
    .I0_3_1(n708_I0_3_1),
    .I0_4_0(n708_I0_4_0),
    .I0_4_1(n708_I0_4_1),
    .I0_5_0(n708_I0_5_0),
    .I0_5_1(n708_I0_5_1),
    .I0_6_0(n708_I0_6_0),
    .I0_6_1(n708_I0_6_1),
    .I0_7_0(n708_I0_7_0),
    .I0_7_1(n708_I0_7_1),
    .I1_0(n708_I1_0),
    .I1_1(n708_I1_1),
    .I1_2(n708_I1_2),
    .I1_3(n708_I1_3),
    .I1_4(n708_I1_4),
    .I1_5(n708_I1_5),
    .I1_6(n708_I1_6),
    .I1_7(n708_I1_7),
    .O_0_0(n708_O_0_0),
    .O_0_1(n708_O_0_1),
    .O_0_2(n708_O_0_2),
    .O_1_0(n708_O_1_0),
    .O_1_1(n708_O_1_1),
    .O_1_2(n708_O_1_2),
    .O_2_0(n708_O_2_0),
    .O_2_1(n708_O_2_1),
    .O_2_2(n708_O_2_2),
    .O_3_0(n708_O_3_0),
    .O_3_1(n708_O_3_1),
    .O_3_2(n708_O_3_2),
    .O_4_0(n708_O_4_0),
    .O_4_1(n708_O_4_1),
    .O_4_2(n708_O_4_2),
    .O_5_0(n708_O_5_0),
    .O_5_1(n708_O_5_1),
    .O_5_2(n708_O_5_2),
    .O_6_0(n708_O_6_0),
    .O_6_1(n708_O_6_1),
    .O_6_2(n708_O_6_2),
    .O_7_0(n708_O_7_0),
    .O_7_1(n708_O_7_1),
    .O_7_2(n708_O_7_2)
  );
  MapT n717 ( // @[Top.scala 959:22]
    .valid_up(n717_valid_up),
    .valid_down(n717_valid_down),
    .I_0_0(n717_I_0_0),
    .I_0_1(n717_I_0_1),
    .I_0_2(n717_I_0_2),
    .I_1_0(n717_I_1_0),
    .I_1_1(n717_I_1_1),
    .I_1_2(n717_I_1_2),
    .I_2_0(n717_I_2_0),
    .I_2_1(n717_I_2_1),
    .I_2_2(n717_I_2_2),
    .I_3_0(n717_I_3_0),
    .I_3_1(n717_I_3_1),
    .I_3_2(n717_I_3_2),
    .I_4_0(n717_I_4_0),
    .I_4_1(n717_I_4_1),
    .I_4_2(n717_I_4_2),
    .I_5_0(n717_I_5_0),
    .I_5_1(n717_I_5_1),
    .I_5_2(n717_I_5_2),
    .I_6_0(n717_I_6_0),
    .I_6_1(n717_I_6_1),
    .I_6_2(n717_I_6_2),
    .I_7_0(n717_I_7_0),
    .I_7_1(n717_I_7_1),
    .I_7_2(n717_I_7_2),
    .O_0_0_0(n717_O_0_0_0),
    .O_0_0_1(n717_O_0_0_1),
    .O_0_0_2(n717_O_0_0_2),
    .O_1_0_0(n717_O_1_0_0),
    .O_1_0_1(n717_O_1_0_1),
    .O_1_0_2(n717_O_1_0_2),
    .O_2_0_0(n717_O_2_0_0),
    .O_2_0_1(n717_O_2_0_1),
    .O_2_0_2(n717_O_2_0_2),
    .O_3_0_0(n717_O_3_0_0),
    .O_3_0_1(n717_O_3_0_1),
    .O_3_0_2(n717_O_3_0_2),
    .O_4_0_0(n717_O_4_0_0),
    .O_4_0_1(n717_O_4_0_1),
    .O_4_0_2(n717_O_4_0_2),
    .O_5_0_0(n717_O_5_0_0),
    .O_5_0_1(n717_O_5_0_1),
    .O_5_0_2(n717_O_5_0_2),
    .O_6_0_0(n717_O_6_0_0),
    .O_6_0_1(n717_O_6_0_1),
    .O_6_0_2(n717_O_6_0_2),
    .O_7_0_0(n717_O_7_0_0),
    .O_7_0_1(n717_O_7_0_1),
    .O_7_0_2(n717_O_7_0_2)
  );
  MapT_1 n724 ( // @[Top.scala 962:22]
    .valid_up(n724_valid_up),
    .valid_down(n724_valid_down),
    .I_0_0_0(n724_I_0_0_0),
    .I_0_0_1(n724_I_0_0_1),
    .I_0_0_2(n724_I_0_0_2),
    .I_1_0_0(n724_I_1_0_0),
    .I_1_0_1(n724_I_1_0_1),
    .I_1_0_2(n724_I_1_0_2),
    .I_2_0_0(n724_I_2_0_0),
    .I_2_0_1(n724_I_2_0_1),
    .I_2_0_2(n724_I_2_0_2),
    .I_3_0_0(n724_I_3_0_0),
    .I_3_0_1(n724_I_3_0_1),
    .I_3_0_2(n724_I_3_0_2),
    .I_4_0_0(n724_I_4_0_0),
    .I_4_0_1(n724_I_4_0_1),
    .I_4_0_2(n724_I_4_0_2),
    .I_5_0_0(n724_I_5_0_0),
    .I_5_0_1(n724_I_5_0_1),
    .I_5_0_2(n724_I_5_0_2),
    .I_6_0_0(n724_I_6_0_0),
    .I_6_0_1(n724_I_6_0_1),
    .I_6_0_2(n724_I_6_0_2),
    .I_7_0_0(n724_I_7_0_0),
    .I_7_0_1(n724_I_7_0_1),
    .I_7_0_2(n724_I_7_0_2),
    .O_0_0(n724_O_0_0),
    .O_0_1(n724_O_0_1),
    .O_0_2(n724_O_0_2),
    .O_1_0(n724_O_1_0),
    .O_1_1(n724_O_1_1),
    .O_1_2(n724_O_1_2),
    .O_2_0(n724_O_2_0),
    .O_2_1(n724_O_2_1),
    .O_2_2(n724_O_2_2),
    .O_3_0(n724_O_3_0),
    .O_3_1(n724_O_3_1),
    .O_3_2(n724_O_3_2),
    .O_4_0(n724_O_4_0),
    .O_4_1(n724_O_4_1),
    .O_4_2(n724_O_4_2),
    .O_5_0(n724_O_5_0),
    .O_5_1(n724_O_5_1),
    .O_5_2(n724_O_5_2),
    .O_6_0(n724_O_6_0),
    .O_6_1(n724_O_6_1),
    .O_6_2(n724_O_6_2),
    .O_7_0(n724_O_7_0),
    .O_7_1(n724_O_7_1),
    .O_7_2(n724_O_7_2)
  );
  Map2T_7 n725 ( // @[Top.scala 965:22]
    .valid_up(n725_valid_up),
    .valid_down(n725_valid_down),
    .I0_0_0_0(n725_I0_0_0_0),
    .I0_0_0_1(n725_I0_0_0_1),
    .I0_0_0_2(n725_I0_0_0_2),
    .I0_0_1_0(n725_I0_0_1_0),
    .I0_0_1_1(n725_I0_0_1_1),
    .I0_0_1_2(n725_I0_0_1_2),
    .I0_1_0_0(n725_I0_1_0_0),
    .I0_1_0_1(n725_I0_1_0_1),
    .I0_1_0_2(n725_I0_1_0_2),
    .I0_1_1_0(n725_I0_1_1_0),
    .I0_1_1_1(n725_I0_1_1_1),
    .I0_1_1_2(n725_I0_1_1_2),
    .I0_2_0_0(n725_I0_2_0_0),
    .I0_2_0_1(n725_I0_2_0_1),
    .I0_2_0_2(n725_I0_2_0_2),
    .I0_2_1_0(n725_I0_2_1_0),
    .I0_2_1_1(n725_I0_2_1_1),
    .I0_2_1_2(n725_I0_2_1_2),
    .I0_3_0_0(n725_I0_3_0_0),
    .I0_3_0_1(n725_I0_3_0_1),
    .I0_3_0_2(n725_I0_3_0_2),
    .I0_3_1_0(n725_I0_3_1_0),
    .I0_3_1_1(n725_I0_3_1_1),
    .I0_3_1_2(n725_I0_3_1_2),
    .I0_4_0_0(n725_I0_4_0_0),
    .I0_4_0_1(n725_I0_4_0_1),
    .I0_4_0_2(n725_I0_4_0_2),
    .I0_4_1_0(n725_I0_4_1_0),
    .I0_4_1_1(n725_I0_4_1_1),
    .I0_4_1_2(n725_I0_4_1_2),
    .I0_5_0_0(n725_I0_5_0_0),
    .I0_5_0_1(n725_I0_5_0_1),
    .I0_5_0_2(n725_I0_5_0_2),
    .I0_5_1_0(n725_I0_5_1_0),
    .I0_5_1_1(n725_I0_5_1_1),
    .I0_5_1_2(n725_I0_5_1_2),
    .I0_6_0_0(n725_I0_6_0_0),
    .I0_6_0_1(n725_I0_6_0_1),
    .I0_6_0_2(n725_I0_6_0_2),
    .I0_6_1_0(n725_I0_6_1_0),
    .I0_6_1_1(n725_I0_6_1_1),
    .I0_6_1_2(n725_I0_6_1_2),
    .I0_7_0_0(n725_I0_7_0_0),
    .I0_7_0_1(n725_I0_7_0_1),
    .I0_7_0_2(n725_I0_7_0_2),
    .I0_7_1_0(n725_I0_7_1_0),
    .I0_7_1_1(n725_I0_7_1_1),
    .I0_7_1_2(n725_I0_7_1_2),
    .I1_0_0(n725_I1_0_0),
    .I1_0_1(n725_I1_0_1),
    .I1_0_2(n725_I1_0_2),
    .I1_1_0(n725_I1_1_0),
    .I1_1_1(n725_I1_1_1),
    .I1_1_2(n725_I1_1_2),
    .I1_2_0(n725_I1_2_0),
    .I1_2_1(n725_I1_2_1),
    .I1_2_2(n725_I1_2_2),
    .I1_3_0(n725_I1_3_0),
    .I1_3_1(n725_I1_3_1),
    .I1_3_2(n725_I1_3_2),
    .I1_4_0(n725_I1_4_0),
    .I1_4_1(n725_I1_4_1),
    .I1_4_2(n725_I1_4_2),
    .I1_5_0(n725_I1_5_0),
    .I1_5_1(n725_I1_5_1),
    .I1_5_2(n725_I1_5_2),
    .I1_6_0(n725_I1_6_0),
    .I1_6_1(n725_I1_6_1),
    .I1_6_2(n725_I1_6_2),
    .I1_7_0(n725_I1_7_0),
    .I1_7_1(n725_I1_7_1),
    .I1_7_2(n725_I1_7_2),
    .O_0_0_0(n725_O_0_0_0),
    .O_0_0_1(n725_O_0_0_1),
    .O_0_0_2(n725_O_0_0_2),
    .O_0_1_0(n725_O_0_1_0),
    .O_0_1_1(n725_O_0_1_1),
    .O_0_1_2(n725_O_0_1_2),
    .O_0_2_0(n725_O_0_2_0),
    .O_0_2_1(n725_O_0_2_1),
    .O_0_2_2(n725_O_0_2_2),
    .O_1_0_0(n725_O_1_0_0),
    .O_1_0_1(n725_O_1_0_1),
    .O_1_0_2(n725_O_1_0_2),
    .O_1_1_0(n725_O_1_1_0),
    .O_1_1_1(n725_O_1_1_1),
    .O_1_1_2(n725_O_1_1_2),
    .O_1_2_0(n725_O_1_2_0),
    .O_1_2_1(n725_O_1_2_1),
    .O_1_2_2(n725_O_1_2_2),
    .O_2_0_0(n725_O_2_0_0),
    .O_2_0_1(n725_O_2_0_1),
    .O_2_0_2(n725_O_2_0_2),
    .O_2_1_0(n725_O_2_1_0),
    .O_2_1_1(n725_O_2_1_1),
    .O_2_1_2(n725_O_2_1_2),
    .O_2_2_0(n725_O_2_2_0),
    .O_2_2_1(n725_O_2_2_1),
    .O_2_2_2(n725_O_2_2_2),
    .O_3_0_0(n725_O_3_0_0),
    .O_3_0_1(n725_O_3_0_1),
    .O_3_0_2(n725_O_3_0_2),
    .O_3_1_0(n725_O_3_1_0),
    .O_3_1_1(n725_O_3_1_1),
    .O_3_1_2(n725_O_3_1_2),
    .O_3_2_0(n725_O_3_2_0),
    .O_3_2_1(n725_O_3_2_1),
    .O_3_2_2(n725_O_3_2_2),
    .O_4_0_0(n725_O_4_0_0),
    .O_4_0_1(n725_O_4_0_1),
    .O_4_0_2(n725_O_4_0_2),
    .O_4_1_0(n725_O_4_1_0),
    .O_4_1_1(n725_O_4_1_1),
    .O_4_1_2(n725_O_4_1_2),
    .O_4_2_0(n725_O_4_2_0),
    .O_4_2_1(n725_O_4_2_1),
    .O_4_2_2(n725_O_4_2_2),
    .O_5_0_0(n725_O_5_0_0),
    .O_5_0_1(n725_O_5_0_1),
    .O_5_0_2(n725_O_5_0_2),
    .O_5_1_0(n725_O_5_1_0),
    .O_5_1_1(n725_O_5_1_1),
    .O_5_1_2(n725_O_5_1_2),
    .O_5_2_0(n725_O_5_2_0),
    .O_5_2_1(n725_O_5_2_1),
    .O_5_2_2(n725_O_5_2_2),
    .O_6_0_0(n725_O_6_0_0),
    .O_6_0_1(n725_O_6_0_1),
    .O_6_0_2(n725_O_6_0_2),
    .O_6_1_0(n725_O_6_1_0),
    .O_6_1_1(n725_O_6_1_1),
    .O_6_1_2(n725_O_6_1_2),
    .O_6_2_0(n725_O_6_2_0),
    .O_6_2_1(n725_O_6_2_1),
    .O_6_2_2(n725_O_6_2_2),
    .O_7_0_0(n725_O_7_0_0),
    .O_7_0_1(n725_O_7_0_1),
    .O_7_0_2(n725_O_7_0_2),
    .O_7_1_0(n725_O_7_1_0),
    .O_7_1_1(n725_O_7_1_1),
    .O_7_1_2(n725_O_7_1_2),
    .O_7_2_0(n725_O_7_2_0),
    .O_7_2_1(n725_O_7_2_1),
    .O_7_2_2(n725_O_7_2_2)
  );
  MapT_6 n734 ( // @[Top.scala 969:22]
    .valid_up(n734_valid_up),
    .valid_down(n734_valid_down),
    .I_0_0_0(n734_I_0_0_0),
    .I_0_0_1(n734_I_0_0_1),
    .I_0_0_2(n734_I_0_0_2),
    .I_0_1_0(n734_I_0_1_0),
    .I_0_1_1(n734_I_0_1_1),
    .I_0_1_2(n734_I_0_1_2),
    .I_0_2_0(n734_I_0_2_0),
    .I_0_2_1(n734_I_0_2_1),
    .I_0_2_2(n734_I_0_2_2),
    .I_1_0_0(n734_I_1_0_0),
    .I_1_0_1(n734_I_1_0_1),
    .I_1_0_2(n734_I_1_0_2),
    .I_1_1_0(n734_I_1_1_0),
    .I_1_1_1(n734_I_1_1_1),
    .I_1_1_2(n734_I_1_1_2),
    .I_1_2_0(n734_I_1_2_0),
    .I_1_2_1(n734_I_1_2_1),
    .I_1_2_2(n734_I_1_2_2),
    .I_2_0_0(n734_I_2_0_0),
    .I_2_0_1(n734_I_2_0_1),
    .I_2_0_2(n734_I_2_0_2),
    .I_2_1_0(n734_I_2_1_0),
    .I_2_1_1(n734_I_2_1_1),
    .I_2_1_2(n734_I_2_1_2),
    .I_2_2_0(n734_I_2_2_0),
    .I_2_2_1(n734_I_2_2_1),
    .I_2_2_2(n734_I_2_2_2),
    .I_3_0_0(n734_I_3_0_0),
    .I_3_0_1(n734_I_3_0_1),
    .I_3_0_2(n734_I_3_0_2),
    .I_3_1_0(n734_I_3_1_0),
    .I_3_1_1(n734_I_3_1_1),
    .I_3_1_2(n734_I_3_1_2),
    .I_3_2_0(n734_I_3_2_0),
    .I_3_2_1(n734_I_3_2_1),
    .I_3_2_2(n734_I_3_2_2),
    .I_4_0_0(n734_I_4_0_0),
    .I_4_0_1(n734_I_4_0_1),
    .I_4_0_2(n734_I_4_0_2),
    .I_4_1_0(n734_I_4_1_0),
    .I_4_1_1(n734_I_4_1_1),
    .I_4_1_2(n734_I_4_1_2),
    .I_4_2_0(n734_I_4_2_0),
    .I_4_2_1(n734_I_4_2_1),
    .I_4_2_2(n734_I_4_2_2),
    .I_5_0_0(n734_I_5_0_0),
    .I_5_0_1(n734_I_5_0_1),
    .I_5_0_2(n734_I_5_0_2),
    .I_5_1_0(n734_I_5_1_0),
    .I_5_1_1(n734_I_5_1_1),
    .I_5_1_2(n734_I_5_1_2),
    .I_5_2_0(n734_I_5_2_0),
    .I_5_2_1(n734_I_5_2_1),
    .I_5_2_2(n734_I_5_2_2),
    .I_6_0_0(n734_I_6_0_0),
    .I_6_0_1(n734_I_6_0_1),
    .I_6_0_2(n734_I_6_0_2),
    .I_6_1_0(n734_I_6_1_0),
    .I_6_1_1(n734_I_6_1_1),
    .I_6_1_2(n734_I_6_1_2),
    .I_6_2_0(n734_I_6_2_0),
    .I_6_2_1(n734_I_6_2_1),
    .I_6_2_2(n734_I_6_2_2),
    .I_7_0_0(n734_I_7_0_0),
    .I_7_0_1(n734_I_7_0_1),
    .I_7_0_2(n734_I_7_0_2),
    .I_7_1_0(n734_I_7_1_0),
    .I_7_1_1(n734_I_7_1_1),
    .I_7_1_2(n734_I_7_1_2),
    .I_7_2_0(n734_I_7_2_0),
    .I_7_2_1(n734_I_7_2_1),
    .I_7_2_2(n734_I_7_2_2),
    .O_0_0_0_0(n734_O_0_0_0_0),
    .O_0_0_0_1(n734_O_0_0_0_1),
    .O_0_0_0_2(n734_O_0_0_0_2),
    .O_0_0_1_0(n734_O_0_0_1_0),
    .O_0_0_1_1(n734_O_0_0_1_1),
    .O_0_0_1_2(n734_O_0_0_1_2),
    .O_0_0_2_0(n734_O_0_0_2_0),
    .O_0_0_2_1(n734_O_0_0_2_1),
    .O_0_0_2_2(n734_O_0_0_2_2),
    .O_1_0_0_0(n734_O_1_0_0_0),
    .O_1_0_0_1(n734_O_1_0_0_1),
    .O_1_0_0_2(n734_O_1_0_0_2),
    .O_1_0_1_0(n734_O_1_0_1_0),
    .O_1_0_1_1(n734_O_1_0_1_1),
    .O_1_0_1_2(n734_O_1_0_1_2),
    .O_1_0_2_0(n734_O_1_0_2_0),
    .O_1_0_2_1(n734_O_1_0_2_1),
    .O_1_0_2_2(n734_O_1_0_2_2),
    .O_2_0_0_0(n734_O_2_0_0_0),
    .O_2_0_0_1(n734_O_2_0_0_1),
    .O_2_0_0_2(n734_O_2_0_0_2),
    .O_2_0_1_0(n734_O_2_0_1_0),
    .O_2_0_1_1(n734_O_2_0_1_1),
    .O_2_0_1_2(n734_O_2_0_1_2),
    .O_2_0_2_0(n734_O_2_0_2_0),
    .O_2_0_2_1(n734_O_2_0_2_1),
    .O_2_0_2_2(n734_O_2_0_2_2),
    .O_3_0_0_0(n734_O_3_0_0_0),
    .O_3_0_0_1(n734_O_3_0_0_1),
    .O_3_0_0_2(n734_O_3_0_0_2),
    .O_3_0_1_0(n734_O_3_0_1_0),
    .O_3_0_1_1(n734_O_3_0_1_1),
    .O_3_0_1_2(n734_O_3_0_1_2),
    .O_3_0_2_0(n734_O_3_0_2_0),
    .O_3_0_2_1(n734_O_3_0_2_1),
    .O_3_0_2_2(n734_O_3_0_2_2),
    .O_4_0_0_0(n734_O_4_0_0_0),
    .O_4_0_0_1(n734_O_4_0_0_1),
    .O_4_0_0_2(n734_O_4_0_0_2),
    .O_4_0_1_0(n734_O_4_0_1_0),
    .O_4_0_1_1(n734_O_4_0_1_1),
    .O_4_0_1_2(n734_O_4_0_1_2),
    .O_4_0_2_0(n734_O_4_0_2_0),
    .O_4_0_2_1(n734_O_4_0_2_1),
    .O_4_0_2_2(n734_O_4_0_2_2),
    .O_5_0_0_0(n734_O_5_0_0_0),
    .O_5_0_0_1(n734_O_5_0_0_1),
    .O_5_0_0_2(n734_O_5_0_0_2),
    .O_5_0_1_0(n734_O_5_0_1_0),
    .O_5_0_1_1(n734_O_5_0_1_1),
    .O_5_0_1_2(n734_O_5_0_1_2),
    .O_5_0_2_0(n734_O_5_0_2_0),
    .O_5_0_2_1(n734_O_5_0_2_1),
    .O_5_0_2_2(n734_O_5_0_2_2),
    .O_6_0_0_0(n734_O_6_0_0_0),
    .O_6_0_0_1(n734_O_6_0_0_1),
    .O_6_0_0_2(n734_O_6_0_0_2),
    .O_6_0_1_0(n734_O_6_0_1_0),
    .O_6_0_1_1(n734_O_6_0_1_1),
    .O_6_0_1_2(n734_O_6_0_1_2),
    .O_6_0_2_0(n734_O_6_0_2_0),
    .O_6_0_2_1(n734_O_6_0_2_1),
    .O_6_0_2_2(n734_O_6_0_2_2),
    .O_7_0_0_0(n734_O_7_0_0_0),
    .O_7_0_0_1(n734_O_7_0_0_1),
    .O_7_0_0_2(n734_O_7_0_0_2),
    .O_7_0_1_0(n734_O_7_0_1_0),
    .O_7_0_1_1(n734_O_7_0_1_1),
    .O_7_0_1_2(n734_O_7_0_1_2),
    .O_7_0_2_0(n734_O_7_0_2_0),
    .O_7_0_2_1(n734_O_7_0_2_1),
    .O_7_0_2_2(n734_O_7_0_2_2)
  );
  MapT_7 n741 ( // @[Top.scala 972:22]
    .valid_up(n741_valid_up),
    .valid_down(n741_valid_down),
    .I_0_0_0_0(n741_I_0_0_0_0),
    .I_0_0_0_1(n741_I_0_0_0_1),
    .I_0_0_0_2(n741_I_0_0_0_2),
    .I_0_0_1_0(n741_I_0_0_1_0),
    .I_0_0_1_1(n741_I_0_0_1_1),
    .I_0_0_1_2(n741_I_0_0_1_2),
    .I_0_0_2_0(n741_I_0_0_2_0),
    .I_0_0_2_1(n741_I_0_0_2_1),
    .I_0_0_2_2(n741_I_0_0_2_2),
    .I_1_0_0_0(n741_I_1_0_0_0),
    .I_1_0_0_1(n741_I_1_0_0_1),
    .I_1_0_0_2(n741_I_1_0_0_2),
    .I_1_0_1_0(n741_I_1_0_1_0),
    .I_1_0_1_1(n741_I_1_0_1_1),
    .I_1_0_1_2(n741_I_1_0_1_2),
    .I_1_0_2_0(n741_I_1_0_2_0),
    .I_1_0_2_1(n741_I_1_0_2_1),
    .I_1_0_2_2(n741_I_1_0_2_2),
    .I_2_0_0_0(n741_I_2_0_0_0),
    .I_2_0_0_1(n741_I_2_0_0_1),
    .I_2_0_0_2(n741_I_2_0_0_2),
    .I_2_0_1_0(n741_I_2_0_1_0),
    .I_2_0_1_1(n741_I_2_0_1_1),
    .I_2_0_1_2(n741_I_2_0_1_2),
    .I_2_0_2_0(n741_I_2_0_2_0),
    .I_2_0_2_1(n741_I_2_0_2_1),
    .I_2_0_2_2(n741_I_2_0_2_2),
    .I_3_0_0_0(n741_I_3_0_0_0),
    .I_3_0_0_1(n741_I_3_0_0_1),
    .I_3_0_0_2(n741_I_3_0_0_2),
    .I_3_0_1_0(n741_I_3_0_1_0),
    .I_3_0_1_1(n741_I_3_0_1_1),
    .I_3_0_1_2(n741_I_3_0_1_2),
    .I_3_0_2_0(n741_I_3_0_2_0),
    .I_3_0_2_1(n741_I_3_0_2_1),
    .I_3_0_2_2(n741_I_3_0_2_2),
    .I_4_0_0_0(n741_I_4_0_0_0),
    .I_4_0_0_1(n741_I_4_0_0_1),
    .I_4_0_0_2(n741_I_4_0_0_2),
    .I_4_0_1_0(n741_I_4_0_1_0),
    .I_4_0_1_1(n741_I_4_0_1_1),
    .I_4_0_1_2(n741_I_4_0_1_2),
    .I_4_0_2_0(n741_I_4_0_2_0),
    .I_4_0_2_1(n741_I_4_0_2_1),
    .I_4_0_2_2(n741_I_4_0_2_2),
    .I_5_0_0_0(n741_I_5_0_0_0),
    .I_5_0_0_1(n741_I_5_0_0_1),
    .I_5_0_0_2(n741_I_5_0_0_2),
    .I_5_0_1_0(n741_I_5_0_1_0),
    .I_5_0_1_1(n741_I_5_0_1_1),
    .I_5_0_1_2(n741_I_5_0_1_2),
    .I_5_0_2_0(n741_I_5_0_2_0),
    .I_5_0_2_1(n741_I_5_0_2_1),
    .I_5_0_2_2(n741_I_5_0_2_2),
    .I_6_0_0_0(n741_I_6_0_0_0),
    .I_6_0_0_1(n741_I_6_0_0_1),
    .I_6_0_0_2(n741_I_6_0_0_2),
    .I_6_0_1_0(n741_I_6_0_1_0),
    .I_6_0_1_1(n741_I_6_0_1_1),
    .I_6_0_1_2(n741_I_6_0_1_2),
    .I_6_0_2_0(n741_I_6_0_2_0),
    .I_6_0_2_1(n741_I_6_0_2_1),
    .I_6_0_2_2(n741_I_6_0_2_2),
    .I_7_0_0_0(n741_I_7_0_0_0),
    .I_7_0_0_1(n741_I_7_0_0_1),
    .I_7_0_0_2(n741_I_7_0_0_2),
    .I_7_0_1_0(n741_I_7_0_1_0),
    .I_7_0_1_1(n741_I_7_0_1_1),
    .I_7_0_1_2(n741_I_7_0_1_2),
    .I_7_0_2_0(n741_I_7_0_2_0),
    .I_7_0_2_1(n741_I_7_0_2_1),
    .I_7_0_2_2(n741_I_7_0_2_2),
    .O_0_0_0(n741_O_0_0_0),
    .O_0_0_1(n741_O_0_0_1),
    .O_0_0_2(n741_O_0_0_2),
    .O_0_1_0(n741_O_0_1_0),
    .O_0_1_1(n741_O_0_1_1),
    .O_0_1_2(n741_O_0_1_2),
    .O_0_2_0(n741_O_0_2_0),
    .O_0_2_1(n741_O_0_2_1),
    .O_0_2_2(n741_O_0_2_2),
    .O_1_0_0(n741_O_1_0_0),
    .O_1_0_1(n741_O_1_0_1),
    .O_1_0_2(n741_O_1_0_2),
    .O_1_1_0(n741_O_1_1_0),
    .O_1_1_1(n741_O_1_1_1),
    .O_1_1_2(n741_O_1_1_2),
    .O_1_2_0(n741_O_1_2_0),
    .O_1_2_1(n741_O_1_2_1),
    .O_1_2_2(n741_O_1_2_2),
    .O_2_0_0(n741_O_2_0_0),
    .O_2_0_1(n741_O_2_0_1),
    .O_2_0_2(n741_O_2_0_2),
    .O_2_1_0(n741_O_2_1_0),
    .O_2_1_1(n741_O_2_1_1),
    .O_2_1_2(n741_O_2_1_2),
    .O_2_2_0(n741_O_2_2_0),
    .O_2_2_1(n741_O_2_2_1),
    .O_2_2_2(n741_O_2_2_2),
    .O_3_0_0(n741_O_3_0_0),
    .O_3_0_1(n741_O_3_0_1),
    .O_3_0_2(n741_O_3_0_2),
    .O_3_1_0(n741_O_3_1_0),
    .O_3_1_1(n741_O_3_1_1),
    .O_3_1_2(n741_O_3_1_2),
    .O_3_2_0(n741_O_3_2_0),
    .O_3_2_1(n741_O_3_2_1),
    .O_3_2_2(n741_O_3_2_2),
    .O_4_0_0(n741_O_4_0_0),
    .O_4_0_1(n741_O_4_0_1),
    .O_4_0_2(n741_O_4_0_2),
    .O_4_1_0(n741_O_4_1_0),
    .O_4_1_1(n741_O_4_1_1),
    .O_4_1_2(n741_O_4_1_2),
    .O_4_2_0(n741_O_4_2_0),
    .O_4_2_1(n741_O_4_2_1),
    .O_4_2_2(n741_O_4_2_2),
    .O_5_0_0(n741_O_5_0_0),
    .O_5_0_1(n741_O_5_0_1),
    .O_5_0_2(n741_O_5_0_2),
    .O_5_1_0(n741_O_5_1_0),
    .O_5_1_1(n741_O_5_1_1),
    .O_5_1_2(n741_O_5_1_2),
    .O_5_2_0(n741_O_5_2_0),
    .O_5_2_1(n741_O_5_2_1),
    .O_5_2_2(n741_O_5_2_2),
    .O_6_0_0(n741_O_6_0_0),
    .O_6_0_1(n741_O_6_0_1),
    .O_6_0_2(n741_O_6_0_2),
    .O_6_1_0(n741_O_6_1_0),
    .O_6_1_1(n741_O_6_1_1),
    .O_6_1_2(n741_O_6_1_2),
    .O_6_2_0(n741_O_6_2_0),
    .O_6_2_1(n741_O_6_2_1),
    .O_6_2_2(n741_O_6_2_2),
    .O_7_0_0(n741_O_7_0_0),
    .O_7_0_1(n741_O_7_0_1),
    .O_7_0_2(n741_O_7_0_2),
    .O_7_1_0(n741_O_7_1_0),
    .O_7_1_1(n741_O_7_1_1),
    .O_7_1_2(n741_O_7_1_2),
    .O_7_2_0(n741_O_7_2_0),
    .O_7_2_1(n741_O_7_2_1),
    .O_7_2_2(n741_O_7_2_2)
  );
  MapT_32 n783 ( // @[Top.scala 975:22]
    .clock(n783_clock),
    .reset(n783_reset),
    .valid_up(n783_valid_up),
    .valid_down(n783_valid_down),
    .I_0_0_0(n783_I_0_0_0),
    .I_0_0_1(n783_I_0_0_1),
    .I_0_0_2(n783_I_0_0_2),
    .I_0_1_0(n783_I_0_1_0),
    .I_0_1_1(n783_I_0_1_1),
    .I_0_1_2(n783_I_0_1_2),
    .I_0_2_0(n783_I_0_2_0),
    .I_0_2_1(n783_I_0_2_1),
    .I_0_2_2(n783_I_0_2_2),
    .I_1_0_0(n783_I_1_0_0),
    .I_1_0_1(n783_I_1_0_1),
    .I_1_0_2(n783_I_1_0_2),
    .I_1_1_0(n783_I_1_1_0),
    .I_1_1_1(n783_I_1_1_1),
    .I_1_1_2(n783_I_1_1_2),
    .I_1_2_0(n783_I_1_2_0),
    .I_1_2_1(n783_I_1_2_1),
    .I_1_2_2(n783_I_1_2_2),
    .I_2_0_0(n783_I_2_0_0),
    .I_2_0_1(n783_I_2_0_1),
    .I_2_0_2(n783_I_2_0_2),
    .I_2_1_0(n783_I_2_1_0),
    .I_2_1_1(n783_I_2_1_1),
    .I_2_1_2(n783_I_2_1_2),
    .I_2_2_0(n783_I_2_2_0),
    .I_2_2_1(n783_I_2_2_1),
    .I_2_2_2(n783_I_2_2_2),
    .I_3_0_0(n783_I_3_0_0),
    .I_3_0_1(n783_I_3_0_1),
    .I_3_0_2(n783_I_3_0_2),
    .I_3_1_0(n783_I_3_1_0),
    .I_3_1_1(n783_I_3_1_1),
    .I_3_1_2(n783_I_3_1_2),
    .I_3_2_0(n783_I_3_2_0),
    .I_3_2_1(n783_I_3_2_1),
    .I_3_2_2(n783_I_3_2_2),
    .I_4_0_0(n783_I_4_0_0),
    .I_4_0_1(n783_I_4_0_1),
    .I_4_0_2(n783_I_4_0_2),
    .I_4_1_0(n783_I_4_1_0),
    .I_4_1_1(n783_I_4_1_1),
    .I_4_1_2(n783_I_4_1_2),
    .I_4_2_0(n783_I_4_2_0),
    .I_4_2_1(n783_I_4_2_1),
    .I_4_2_2(n783_I_4_2_2),
    .I_5_0_0(n783_I_5_0_0),
    .I_5_0_1(n783_I_5_0_1),
    .I_5_0_2(n783_I_5_0_2),
    .I_5_1_0(n783_I_5_1_0),
    .I_5_1_1(n783_I_5_1_1),
    .I_5_1_2(n783_I_5_1_2),
    .I_5_2_0(n783_I_5_2_0),
    .I_5_2_1(n783_I_5_2_1),
    .I_5_2_2(n783_I_5_2_2),
    .I_6_0_0(n783_I_6_0_0),
    .I_6_0_1(n783_I_6_0_1),
    .I_6_0_2(n783_I_6_0_2),
    .I_6_1_0(n783_I_6_1_0),
    .I_6_1_1(n783_I_6_1_1),
    .I_6_1_2(n783_I_6_1_2),
    .I_6_2_0(n783_I_6_2_0),
    .I_6_2_1(n783_I_6_2_1),
    .I_6_2_2(n783_I_6_2_2),
    .I_7_0_0(n783_I_7_0_0),
    .I_7_0_1(n783_I_7_0_1),
    .I_7_0_2(n783_I_7_0_2),
    .I_7_1_0(n783_I_7_1_0),
    .I_7_1_1(n783_I_7_1_1),
    .I_7_1_2(n783_I_7_1_2),
    .I_7_2_0(n783_I_7_2_0),
    .I_7_2_1(n783_I_7_2_1),
    .I_7_2_2(n783_I_7_2_2),
    .O_0_0_0(n783_O_0_0_0),
    .O_1_0_0(n783_O_1_0_0),
    .O_2_0_0(n783_O_2_0_0),
    .O_3_0_0(n783_O_3_0_0),
    .O_4_0_0(n783_O_4_0_0),
    .O_5_0_0(n783_O_5_0_0),
    .O_6_0_0(n783_O_6_0_0),
    .O_7_0_0(n783_O_7_0_0)
  );
  Passthrough_4 n784 ( // @[Top.scala 978:22]
    .valid_up(n784_valid_up),
    .valid_down(n784_valid_down),
    .I_0_0_0(n784_I_0_0_0),
    .I_1_0_0(n784_I_1_0_0),
    .I_2_0_0(n784_I_2_0_0),
    .I_3_0_0(n784_I_3_0_0),
    .I_4_0_0(n784_I_4_0_0),
    .I_5_0_0(n784_I_5_0_0),
    .I_6_0_0(n784_I_6_0_0),
    .I_7_0_0(n784_I_7_0_0),
    .O_0_0(n784_O_0_0),
    .O_1_0(n784_O_1_0),
    .O_2_0(n784_O_2_0),
    .O_3_0(n784_O_3_0),
    .O_4_0(n784_O_4_0),
    .O_5_0(n784_O_5_0),
    .O_6_0(n784_O_6_0),
    .O_7_0(n784_O_7_0)
  );
  Passthrough_5 n785 ( // @[Top.scala 981:22]
    .valid_up(n785_valid_up),
    .valid_down(n785_valid_down),
    .I_0_0(n785_I_0_0),
    .I_1_0(n785_I_1_0),
    .I_2_0(n785_I_2_0),
    .I_3_0(n785_I_3_0),
    .I_4_0(n785_I_4_0),
    .I_5_0(n785_I_5_0),
    .I_6_0(n785_I_6_0),
    .I_7_0(n785_I_7_0),
    .O_0(n785_O_0),
    .O_1(n785_O_1),
    .O_2(n785_O_2),
    .O_3(n785_O_3),
    .O_4(n785_O_4),
    .O_5(n785_O_5),
    .O_6(n785_O_6),
    .O_7(n785_O_7)
  );
  FIFO_9 n786 ( // @[Top.scala 984:22]
    .clock(n786_clock),
    .reset(n786_reset),
    .valid_up(n786_valid_up),
    .valid_down(n786_valid_down),
    .I_0(n786_I_0),
    .I_1(n786_I_1),
    .I_2(n786_I_2),
    .I_3(n786_I_3),
    .I_4(n786_I_4),
    .I_5(n786_I_5),
    .I_6(n786_I_6),
    .I_7(n786_I_7),
    .O_0(n786_O_0),
    .O_1(n786_O_1),
    .O_2(n786_O_2),
    .O_3(n786_O_3),
    .O_4(n786_O_4),
    .O_5(n786_O_5),
    .O_6(n786_O_6),
    .O_7(n786_O_7)
  );
  Map2T_18 n787 ( // @[Top.scala 987:22]
    .clock(n787_clock),
    .reset(n787_reset),
    .valid_up(n787_valid_up),
    .valid_down(n787_valid_down),
    .I0_0(n787_I0_0),
    .I0_1(n787_I0_1),
    .I0_2(n787_I0_2),
    .I0_3(n787_I0_3),
    .I0_4(n787_I0_4),
    .I0_5(n787_I0_5),
    .I0_6(n787_I0_6),
    .I0_7(n787_I0_7),
    .I1_0(n787_I1_0),
    .I1_1(n787_I1_1),
    .I1_2(n787_I1_2),
    .I1_3(n787_I1_3),
    .I1_4(n787_I1_4),
    .I1_5(n787_I1_5),
    .I1_6(n787_I1_6),
    .I1_7(n787_I1_7),
    .O_0(n787_O_0),
    .O_1(n787_O_1),
    .O_2(n787_O_2),
    .O_3(n787_O_3),
    .O_4(n787_O_4),
    .O_5(n787_O_5),
    .O_6(n787_O_6),
    .O_7(n787_O_7)
  );
  MapT_33 n823 ( // @[Top.scala 991:22]
    .valid_up(n823_valid_up),
    .valid_down(n823_valid_down),
    .I_0_t1b_t0b(n823_I_0_t1b_t0b),
    .I_0_t1b_t1b(n823_I_0_t1b_t1b),
    .I_1_t1b_t0b(n823_I_1_t1b_t0b),
    .I_1_t1b_t1b(n823_I_1_t1b_t1b),
    .I_2_t1b_t0b(n823_I_2_t1b_t0b),
    .I_2_t1b_t1b(n823_I_2_t1b_t1b),
    .I_3_t1b_t0b(n823_I_3_t1b_t0b),
    .I_3_t1b_t1b(n823_I_3_t1b_t1b),
    .I_4_t1b_t0b(n823_I_4_t1b_t0b),
    .I_4_t1b_t1b(n823_I_4_t1b_t1b),
    .I_5_t1b_t0b(n823_I_5_t1b_t0b),
    .I_5_t1b_t1b(n823_I_5_t1b_t1b),
    .I_6_t1b_t0b(n823_I_6_t1b_t0b),
    .I_6_t1b_t1b(n823_I_6_t1b_t1b),
    .I_7_t1b_t0b(n823_I_7_t1b_t0b),
    .I_7_t1b_t1b(n823_I_7_t1b_t1b),
    .O_0(n823_O_0),
    .O_1(n823_O_1),
    .O_2(n823_O_2),
    .O_3(n823_O_3),
    .O_4(n823_O_4),
    .O_5(n823_O_5),
    .O_6(n823_O_6),
    .O_7(n823_O_7)
  );
  ShiftTS n824 ( // @[Top.scala 994:22]
    .clock(n824_clock),
    .reset(n824_reset),
    .valid_up(n824_valid_up),
    .valid_down(n824_valid_down),
    .I_0(n824_I_0),
    .I_1(n824_I_1),
    .I_2(n824_I_2),
    .I_3(n824_I_3),
    .I_4(n824_I_4),
    .I_5(n824_I_5),
    .I_6(n824_I_6),
    .I_7(n824_I_7),
    .O_0(n824_O_0),
    .O_1(n824_O_1),
    .O_2(n824_O_2),
    .O_3(n824_O_3),
    .O_4(n824_O_4),
    .O_5(n824_O_5),
    .O_6(n824_O_6),
    .O_7(n824_O_7)
  );
  ShiftTS n825 ( // @[Top.scala 997:22]
    .clock(n825_clock),
    .reset(n825_reset),
    .valid_up(n825_valid_up),
    .valid_down(n825_valid_down),
    .I_0(n825_I_0),
    .I_1(n825_I_1),
    .I_2(n825_I_2),
    .I_3(n825_I_3),
    .I_4(n825_I_4),
    .I_5(n825_I_5),
    .I_6(n825_I_6),
    .I_7(n825_I_7),
    .O_0(n825_O_0),
    .O_1(n825_O_1),
    .O_2(n825_O_2),
    .O_3(n825_O_3),
    .O_4(n825_O_4),
    .O_5(n825_O_5),
    .O_6(n825_O_6),
    .O_7(n825_O_7)
  );
  ShiftTS_2 n826 ( // @[Top.scala 1000:22]
    .clock(n826_clock),
    .valid_up(n826_valid_up),
    .valid_down(n826_valid_down),
    .I_0(n826_I_0),
    .I_1(n826_I_1),
    .I_2(n826_I_2),
    .I_3(n826_I_3),
    .I_4(n826_I_4),
    .I_5(n826_I_5),
    .I_6(n826_I_6),
    .I_7(n826_I_7),
    .O_0(n826_O_0),
    .O_1(n826_O_1),
    .O_2(n826_O_2),
    .O_3(n826_O_3),
    .O_4(n826_O_4),
    .O_5(n826_O_5),
    .O_6(n826_O_6),
    .O_7(n826_O_7)
  );
  ShiftTS_2 n827 ( // @[Top.scala 1003:22]
    .clock(n827_clock),
    .valid_up(n827_valid_up),
    .valid_down(n827_valid_down),
    .I_0(n827_I_0),
    .I_1(n827_I_1),
    .I_2(n827_I_2),
    .I_3(n827_I_3),
    .I_4(n827_I_4),
    .I_5(n827_I_5),
    .I_6(n827_I_6),
    .I_7(n827_I_7),
    .O_0(n827_O_0),
    .O_1(n827_O_1),
    .O_2(n827_O_2),
    .O_3(n827_O_3),
    .O_4(n827_O_4),
    .O_5(n827_O_5),
    .O_6(n827_O_6),
    .O_7(n827_O_7)
  );
  Map2T n828 ( // @[Top.scala 1006:22]
    .valid_up(n828_valid_up),
    .valid_down(n828_valid_down),
    .I0_0(n828_I0_0),
    .I0_1(n828_I0_1),
    .I0_2(n828_I0_2),
    .I0_3(n828_I0_3),
    .I0_4(n828_I0_4),
    .I0_5(n828_I0_5),
    .I0_6(n828_I0_6),
    .I0_7(n828_I0_7),
    .I1_0(n828_I1_0),
    .I1_1(n828_I1_1),
    .I1_2(n828_I1_2),
    .I1_3(n828_I1_3),
    .I1_4(n828_I1_4),
    .I1_5(n828_I1_5),
    .I1_6(n828_I1_6),
    .I1_7(n828_I1_7),
    .O_0_0(n828_O_0_0),
    .O_0_1(n828_O_0_1),
    .O_1_0(n828_O_1_0),
    .O_1_1(n828_O_1_1),
    .O_2_0(n828_O_2_0),
    .O_2_1(n828_O_2_1),
    .O_3_0(n828_O_3_0),
    .O_3_1(n828_O_3_1),
    .O_4_0(n828_O_4_0),
    .O_4_1(n828_O_4_1),
    .O_5_0(n828_O_5_0),
    .O_5_1(n828_O_5_1),
    .O_6_0(n828_O_6_0),
    .O_6_1(n828_O_6_1),
    .O_7_0(n828_O_7_0),
    .O_7_1(n828_O_7_1)
  );
  Map2T_1 n835 ( // @[Top.scala 1010:22]
    .valid_up(n835_valid_up),
    .valid_down(n835_valid_down),
    .I0_0_0(n835_I0_0_0),
    .I0_0_1(n835_I0_0_1),
    .I0_1_0(n835_I0_1_0),
    .I0_1_1(n835_I0_1_1),
    .I0_2_0(n835_I0_2_0),
    .I0_2_1(n835_I0_2_1),
    .I0_3_0(n835_I0_3_0),
    .I0_3_1(n835_I0_3_1),
    .I0_4_0(n835_I0_4_0),
    .I0_4_1(n835_I0_4_1),
    .I0_5_0(n835_I0_5_0),
    .I0_5_1(n835_I0_5_1),
    .I0_6_0(n835_I0_6_0),
    .I0_6_1(n835_I0_6_1),
    .I0_7_0(n835_I0_7_0),
    .I0_7_1(n835_I0_7_1),
    .I1_0(n835_I1_0),
    .I1_1(n835_I1_1),
    .I1_2(n835_I1_2),
    .I1_3(n835_I1_3),
    .I1_4(n835_I1_4),
    .I1_5(n835_I1_5),
    .I1_6(n835_I1_6),
    .I1_7(n835_I1_7),
    .O_0_0(n835_O_0_0),
    .O_0_1(n835_O_0_1),
    .O_0_2(n835_O_0_2),
    .O_1_0(n835_O_1_0),
    .O_1_1(n835_O_1_1),
    .O_1_2(n835_O_1_2),
    .O_2_0(n835_O_2_0),
    .O_2_1(n835_O_2_1),
    .O_2_2(n835_O_2_2),
    .O_3_0(n835_O_3_0),
    .O_3_1(n835_O_3_1),
    .O_3_2(n835_O_3_2),
    .O_4_0(n835_O_4_0),
    .O_4_1(n835_O_4_1),
    .O_4_2(n835_O_4_2),
    .O_5_0(n835_O_5_0),
    .O_5_1(n835_O_5_1),
    .O_5_2(n835_O_5_2),
    .O_6_0(n835_O_6_0),
    .O_6_1(n835_O_6_1),
    .O_6_2(n835_O_6_2),
    .O_7_0(n835_O_7_0),
    .O_7_1(n835_O_7_1),
    .O_7_2(n835_O_7_2)
  );
  MapT n844 ( // @[Top.scala 1014:22]
    .valid_up(n844_valid_up),
    .valid_down(n844_valid_down),
    .I_0_0(n844_I_0_0),
    .I_0_1(n844_I_0_1),
    .I_0_2(n844_I_0_2),
    .I_1_0(n844_I_1_0),
    .I_1_1(n844_I_1_1),
    .I_1_2(n844_I_1_2),
    .I_2_0(n844_I_2_0),
    .I_2_1(n844_I_2_1),
    .I_2_2(n844_I_2_2),
    .I_3_0(n844_I_3_0),
    .I_3_1(n844_I_3_1),
    .I_3_2(n844_I_3_2),
    .I_4_0(n844_I_4_0),
    .I_4_1(n844_I_4_1),
    .I_4_2(n844_I_4_2),
    .I_5_0(n844_I_5_0),
    .I_5_1(n844_I_5_1),
    .I_5_2(n844_I_5_2),
    .I_6_0(n844_I_6_0),
    .I_6_1(n844_I_6_1),
    .I_6_2(n844_I_6_2),
    .I_7_0(n844_I_7_0),
    .I_7_1(n844_I_7_1),
    .I_7_2(n844_I_7_2),
    .O_0_0_0(n844_O_0_0_0),
    .O_0_0_1(n844_O_0_0_1),
    .O_0_0_2(n844_O_0_0_2),
    .O_1_0_0(n844_O_1_0_0),
    .O_1_0_1(n844_O_1_0_1),
    .O_1_0_2(n844_O_1_0_2),
    .O_2_0_0(n844_O_2_0_0),
    .O_2_0_1(n844_O_2_0_1),
    .O_2_0_2(n844_O_2_0_2),
    .O_3_0_0(n844_O_3_0_0),
    .O_3_0_1(n844_O_3_0_1),
    .O_3_0_2(n844_O_3_0_2),
    .O_4_0_0(n844_O_4_0_0),
    .O_4_0_1(n844_O_4_0_1),
    .O_4_0_2(n844_O_4_0_2),
    .O_5_0_0(n844_O_5_0_0),
    .O_5_0_1(n844_O_5_0_1),
    .O_5_0_2(n844_O_5_0_2),
    .O_6_0_0(n844_O_6_0_0),
    .O_6_0_1(n844_O_6_0_1),
    .O_6_0_2(n844_O_6_0_2),
    .O_7_0_0(n844_O_7_0_0),
    .O_7_0_1(n844_O_7_0_1),
    .O_7_0_2(n844_O_7_0_2)
  );
  MapT_1 n851 ( // @[Top.scala 1017:22]
    .valid_up(n851_valid_up),
    .valid_down(n851_valid_down),
    .I_0_0_0(n851_I_0_0_0),
    .I_0_0_1(n851_I_0_0_1),
    .I_0_0_2(n851_I_0_0_2),
    .I_1_0_0(n851_I_1_0_0),
    .I_1_0_1(n851_I_1_0_1),
    .I_1_0_2(n851_I_1_0_2),
    .I_2_0_0(n851_I_2_0_0),
    .I_2_0_1(n851_I_2_0_1),
    .I_2_0_2(n851_I_2_0_2),
    .I_3_0_0(n851_I_3_0_0),
    .I_3_0_1(n851_I_3_0_1),
    .I_3_0_2(n851_I_3_0_2),
    .I_4_0_0(n851_I_4_0_0),
    .I_4_0_1(n851_I_4_0_1),
    .I_4_0_2(n851_I_4_0_2),
    .I_5_0_0(n851_I_5_0_0),
    .I_5_0_1(n851_I_5_0_1),
    .I_5_0_2(n851_I_5_0_2),
    .I_6_0_0(n851_I_6_0_0),
    .I_6_0_1(n851_I_6_0_1),
    .I_6_0_2(n851_I_6_0_2),
    .I_7_0_0(n851_I_7_0_0),
    .I_7_0_1(n851_I_7_0_1),
    .I_7_0_2(n851_I_7_0_2),
    .O_0_0(n851_O_0_0),
    .O_0_1(n851_O_0_1),
    .O_0_2(n851_O_0_2),
    .O_1_0(n851_O_1_0),
    .O_1_1(n851_O_1_1),
    .O_1_2(n851_O_1_2),
    .O_2_0(n851_O_2_0),
    .O_2_1(n851_O_2_1),
    .O_2_2(n851_O_2_2),
    .O_3_0(n851_O_3_0),
    .O_3_1(n851_O_3_1),
    .O_3_2(n851_O_3_2),
    .O_4_0(n851_O_4_0),
    .O_4_1(n851_O_4_1),
    .O_4_2(n851_O_4_2),
    .O_5_0(n851_O_5_0),
    .O_5_1(n851_O_5_1),
    .O_5_2(n851_O_5_2),
    .O_6_0(n851_O_6_0),
    .O_6_1(n851_O_6_1),
    .O_6_2(n851_O_6_2),
    .O_7_0(n851_O_7_0),
    .O_7_1(n851_O_7_1),
    .O_7_2(n851_O_7_2)
  );
  ShiftTS_2 n852 ( // @[Top.scala 1020:22]
    .clock(n852_clock),
    .valid_up(n852_valid_up),
    .valid_down(n852_valid_down),
    .I_0(n852_I_0),
    .I_1(n852_I_1),
    .I_2(n852_I_2),
    .I_3(n852_I_3),
    .I_4(n852_I_4),
    .I_5(n852_I_5),
    .I_6(n852_I_6),
    .I_7(n852_I_7),
    .O_0(n852_O_0),
    .O_1(n852_O_1),
    .O_2(n852_O_2),
    .O_3(n852_O_3),
    .O_4(n852_O_4),
    .O_5(n852_O_5),
    .O_6(n852_O_6),
    .O_7(n852_O_7)
  );
  ShiftTS_2 n853 ( // @[Top.scala 1023:22]
    .clock(n853_clock),
    .valid_up(n853_valid_up),
    .valid_down(n853_valid_down),
    .I_0(n853_I_0),
    .I_1(n853_I_1),
    .I_2(n853_I_2),
    .I_3(n853_I_3),
    .I_4(n853_I_4),
    .I_5(n853_I_5),
    .I_6(n853_I_6),
    .I_7(n853_I_7),
    .O_0(n853_O_0),
    .O_1(n853_O_1),
    .O_2(n853_O_2),
    .O_3(n853_O_3),
    .O_4(n853_O_4),
    .O_5(n853_O_5),
    .O_6(n853_O_6),
    .O_7(n853_O_7)
  );
  Map2T n854 ( // @[Top.scala 1026:22]
    .valid_up(n854_valid_up),
    .valid_down(n854_valid_down),
    .I0_0(n854_I0_0),
    .I0_1(n854_I0_1),
    .I0_2(n854_I0_2),
    .I0_3(n854_I0_3),
    .I0_4(n854_I0_4),
    .I0_5(n854_I0_5),
    .I0_6(n854_I0_6),
    .I0_7(n854_I0_7),
    .I1_0(n854_I1_0),
    .I1_1(n854_I1_1),
    .I1_2(n854_I1_2),
    .I1_3(n854_I1_3),
    .I1_4(n854_I1_4),
    .I1_5(n854_I1_5),
    .I1_6(n854_I1_6),
    .I1_7(n854_I1_7),
    .O_0_0(n854_O_0_0),
    .O_0_1(n854_O_0_1),
    .O_1_0(n854_O_1_0),
    .O_1_1(n854_O_1_1),
    .O_2_0(n854_O_2_0),
    .O_2_1(n854_O_2_1),
    .O_3_0(n854_O_3_0),
    .O_3_1(n854_O_3_1),
    .O_4_0(n854_O_4_0),
    .O_4_1(n854_O_4_1),
    .O_5_0(n854_O_5_0),
    .O_5_1(n854_O_5_1),
    .O_6_0(n854_O_6_0),
    .O_6_1(n854_O_6_1),
    .O_7_0(n854_O_7_0),
    .O_7_1(n854_O_7_1)
  );
  Map2T_1 n861 ( // @[Top.scala 1030:22]
    .valid_up(n861_valid_up),
    .valid_down(n861_valid_down),
    .I0_0_0(n861_I0_0_0),
    .I0_0_1(n861_I0_0_1),
    .I0_1_0(n861_I0_1_0),
    .I0_1_1(n861_I0_1_1),
    .I0_2_0(n861_I0_2_0),
    .I0_2_1(n861_I0_2_1),
    .I0_3_0(n861_I0_3_0),
    .I0_3_1(n861_I0_3_1),
    .I0_4_0(n861_I0_4_0),
    .I0_4_1(n861_I0_4_1),
    .I0_5_0(n861_I0_5_0),
    .I0_5_1(n861_I0_5_1),
    .I0_6_0(n861_I0_6_0),
    .I0_6_1(n861_I0_6_1),
    .I0_7_0(n861_I0_7_0),
    .I0_7_1(n861_I0_7_1),
    .I1_0(n861_I1_0),
    .I1_1(n861_I1_1),
    .I1_2(n861_I1_2),
    .I1_3(n861_I1_3),
    .I1_4(n861_I1_4),
    .I1_5(n861_I1_5),
    .I1_6(n861_I1_6),
    .I1_7(n861_I1_7),
    .O_0_0(n861_O_0_0),
    .O_0_1(n861_O_0_1),
    .O_0_2(n861_O_0_2),
    .O_1_0(n861_O_1_0),
    .O_1_1(n861_O_1_1),
    .O_1_2(n861_O_1_2),
    .O_2_0(n861_O_2_0),
    .O_2_1(n861_O_2_1),
    .O_2_2(n861_O_2_2),
    .O_3_0(n861_O_3_0),
    .O_3_1(n861_O_3_1),
    .O_3_2(n861_O_3_2),
    .O_4_0(n861_O_4_0),
    .O_4_1(n861_O_4_1),
    .O_4_2(n861_O_4_2),
    .O_5_0(n861_O_5_0),
    .O_5_1(n861_O_5_1),
    .O_5_2(n861_O_5_2),
    .O_6_0(n861_O_6_0),
    .O_6_1(n861_O_6_1),
    .O_6_2(n861_O_6_2),
    .O_7_0(n861_O_7_0),
    .O_7_1(n861_O_7_1),
    .O_7_2(n861_O_7_2)
  );
  MapT n870 ( // @[Top.scala 1034:22]
    .valid_up(n870_valid_up),
    .valid_down(n870_valid_down),
    .I_0_0(n870_I_0_0),
    .I_0_1(n870_I_0_1),
    .I_0_2(n870_I_0_2),
    .I_1_0(n870_I_1_0),
    .I_1_1(n870_I_1_1),
    .I_1_2(n870_I_1_2),
    .I_2_0(n870_I_2_0),
    .I_2_1(n870_I_2_1),
    .I_2_2(n870_I_2_2),
    .I_3_0(n870_I_3_0),
    .I_3_1(n870_I_3_1),
    .I_3_2(n870_I_3_2),
    .I_4_0(n870_I_4_0),
    .I_4_1(n870_I_4_1),
    .I_4_2(n870_I_4_2),
    .I_5_0(n870_I_5_0),
    .I_5_1(n870_I_5_1),
    .I_5_2(n870_I_5_2),
    .I_6_0(n870_I_6_0),
    .I_6_1(n870_I_6_1),
    .I_6_2(n870_I_6_2),
    .I_7_0(n870_I_7_0),
    .I_7_1(n870_I_7_1),
    .I_7_2(n870_I_7_2),
    .O_0_0_0(n870_O_0_0_0),
    .O_0_0_1(n870_O_0_0_1),
    .O_0_0_2(n870_O_0_0_2),
    .O_1_0_0(n870_O_1_0_0),
    .O_1_0_1(n870_O_1_0_1),
    .O_1_0_2(n870_O_1_0_2),
    .O_2_0_0(n870_O_2_0_0),
    .O_2_0_1(n870_O_2_0_1),
    .O_2_0_2(n870_O_2_0_2),
    .O_3_0_0(n870_O_3_0_0),
    .O_3_0_1(n870_O_3_0_1),
    .O_3_0_2(n870_O_3_0_2),
    .O_4_0_0(n870_O_4_0_0),
    .O_4_0_1(n870_O_4_0_1),
    .O_4_0_2(n870_O_4_0_2),
    .O_5_0_0(n870_O_5_0_0),
    .O_5_0_1(n870_O_5_0_1),
    .O_5_0_2(n870_O_5_0_2),
    .O_6_0_0(n870_O_6_0_0),
    .O_6_0_1(n870_O_6_0_1),
    .O_6_0_2(n870_O_6_0_2),
    .O_7_0_0(n870_O_7_0_0),
    .O_7_0_1(n870_O_7_0_1),
    .O_7_0_2(n870_O_7_0_2)
  );
  MapT_1 n877 ( // @[Top.scala 1037:22]
    .valid_up(n877_valid_up),
    .valid_down(n877_valid_down),
    .I_0_0_0(n877_I_0_0_0),
    .I_0_0_1(n877_I_0_0_1),
    .I_0_0_2(n877_I_0_0_2),
    .I_1_0_0(n877_I_1_0_0),
    .I_1_0_1(n877_I_1_0_1),
    .I_1_0_2(n877_I_1_0_2),
    .I_2_0_0(n877_I_2_0_0),
    .I_2_0_1(n877_I_2_0_1),
    .I_2_0_2(n877_I_2_0_2),
    .I_3_0_0(n877_I_3_0_0),
    .I_3_0_1(n877_I_3_0_1),
    .I_3_0_2(n877_I_3_0_2),
    .I_4_0_0(n877_I_4_0_0),
    .I_4_0_1(n877_I_4_0_1),
    .I_4_0_2(n877_I_4_0_2),
    .I_5_0_0(n877_I_5_0_0),
    .I_5_0_1(n877_I_5_0_1),
    .I_5_0_2(n877_I_5_0_2),
    .I_6_0_0(n877_I_6_0_0),
    .I_6_0_1(n877_I_6_0_1),
    .I_6_0_2(n877_I_6_0_2),
    .I_7_0_0(n877_I_7_0_0),
    .I_7_0_1(n877_I_7_0_1),
    .I_7_0_2(n877_I_7_0_2),
    .O_0_0(n877_O_0_0),
    .O_0_1(n877_O_0_1),
    .O_0_2(n877_O_0_2),
    .O_1_0(n877_O_1_0),
    .O_1_1(n877_O_1_1),
    .O_1_2(n877_O_1_2),
    .O_2_0(n877_O_2_0),
    .O_2_1(n877_O_2_1),
    .O_2_2(n877_O_2_2),
    .O_3_0(n877_O_3_0),
    .O_3_1(n877_O_3_1),
    .O_3_2(n877_O_3_2),
    .O_4_0(n877_O_4_0),
    .O_4_1(n877_O_4_1),
    .O_4_2(n877_O_4_2),
    .O_5_0(n877_O_5_0),
    .O_5_1(n877_O_5_1),
    .O_5_2(n877_O_5_2),
    .O_6_0(n877_O_6_0),
    .O_6_1(n877_O_6_1),
    .O_6_2(n877_O_6_2),
    .O_7_0(n877_O_7_0),
    .O_7_1(n877_O_7_1),
    .O_7_2(n877_O_7_2)
  );
  Map2T_4 n878 ( // @[Top.scala 1040:22]
    .valid_up(n878_valid_up),
    .valid_down(n878_valid_down),
    .I0_0_0(n878_I0_0_0),
    .I0_0_1(n878_I0_0_1),
    .I0_0_2(n878_I0_0_2),
    .I0_1_0(n878_I0_1_0),
    .I0_1_1(n878_I0_1_1),
    .I0_1_2(n878_I0_1_2),
    .I0_2_0(n878_I0_2_0),
    .I0_2_1(n878_I0_2_1),
    .I0_2_2(n878_I0_2_2),
    .I0_3_0(n878_I0_3_0),
    .I0_3_1(n878_I0_3_1),
    .I0_3_2(n878_I0_3_2),
    .I0_4_0(n878_I0_4_0),
    .I0_4_1(n878_I0_4_1),
    .I0_4_2(n878_I0_4_2),
    .I0_5_0(n878_I0_5_0),
    .I0_5_1(n878_I0_5_1),
    .I0_5_2(n878_I0_5_2),
    .I0_6_0(n878_I0_6_0),
    .I0_6_1(n878_I0_6_1),
    .I0_6_2(n878_I0_6_2),
    .I0_7_0(n878_I0_7_0),
    .I0_7_1(n878_I0_7_1),
    .I0_7_2(n878_I0_7_2),
    .I1_0_0(n878_I1_0_0),
    .I1_0_1(n878_I1_0_1),
    .I1_0_2(n878_I1_0_2),
    .I1_1_0(n878_I1_1_0),
    .I1_1_1(n878_I1_1_1),
    .I1_1_2(n878_I1_1_2),
    .I1_2_0(n878_I1_2_0),
    .I1_2_1(n878_I1_2_1),
    .I1_2_2(n878_I1_2_2),
    .I1_3_0(n878_I1_3_0),
    .I1_3_1(n878_I1_3_1),
    .I1_3_2(n878_I1_3_2),
    .I1_4_0(n878_I1_4_0),
    .I1_4_1(n878_I1_4_1),
    .I1_4_2(n878_I1_4_2),
    .I1_5_0(n878_I1_5_0),
    .I1_5_1(n878_I1_5_1),
    .I1_5_2(n878_I1_5_2),
    .I1_6_0(n878_I1_6_0),
    .I1_6_1(n878_I1_6_1),
    .I1_6_2(n878_I1_6_2),
    .I1_7_0(n878_I1_7_0),
    .I1_7_1(n878_I1_7_1),
    .I1_7_2(n878_I1_7_2),
    .O_0_0_0(n878_O_0_0_0),
    .O_0_0_1(n878_O_0_0_1),
    .O_0_0_2(n878_O_0_0_2),
    .O_0_1_0(n878_O_0_1_0),
    .O_0_1_1(n878_O_0_1_1),
    .O_0_1_2(n878_O_0_1_2),
    .O_1_0_0(n878_O_1_0_0),
    .O_1_0_1(n878_O_1_0_1),
    .O_1_0_2(n878_O_1_0_2),
    .O_1_1_0(n878_O_1_1_0),
    .O_1_1_1(n878_O_1_1_1),
    .O_1_1_2(n878_O_1_1_2),
    .O_2_0_0(n878_O_2_0_0),
    .O_2_0_1(n878_O_2_0_1),
    .O_2_0_2(n878_O_2_0_2),
    .O_2_1_0(n878_O_2_1_0),
    .O_2_1_1(n878_O_2_1_1),
    .O_2_1_2(n878_O_2_1_2),
    .O_3_0_0(n878_O_3_0_0),
    .O_3_0_1(n878_O_3_0_1),
    .O_3_0_2(n878_O_3_0_2),
    .O_3_1_0(n878_O_3_1_0),
    .O_3_1_1(n878_O_3_1_1),
    .O_3_1_2(n878_O_3_1_2),
    .O_4_0_0(n878_O_4_0_0),
    .O_4_0_1(n878_O_4_0_1),
    .O_4_0_2(n878_O_4_0_2),
    .O_4_1_0(n878_O_4_1_0),
    .O_4_1_1(n878_O_4_1_1),
    .O_4_1_2(n878_O_4_1_2),
    .O_5_0_0(n878_O_5_0_0),
    .O_5_0_1(n878_O_5_0_1),
    .O_5_0_2(n878_O_5_0_2),
    .O_5_1_0(n878_O_5_1_0),
    .O_5_1_1(n878_O_5_1_1),
    .O_5_1_2(n878_O_5_1_2),
    .O_6_0_0(n878_O_6_0_0),
    .O_6_0_1(n878_O_6_0_1),
    .O_6_0_2(n878_O_6_0_2),
    .O_6_1_0(n878_O_6_1_0),
    .O_6_1_1(n878_O_6_1_1),
    .O_6_1_2(n878_O_6_1_2),
    .O_7_0_0(n878_O_7_0_0),
    .O_7_0_1(n878_O_7_0_1),
    .O_7_0_2(n878_O_7_0_2),
    .O_7_1_0(n878_O_7_1_0),
    .O_7_1_1(n878_O_7_1_1),
    .O_7_1_2(n878_O_7_1_2)
  );
  ShiftTS_2 n885 ( // @[Top.scala 1044:22]
    .clock(n885_clock),
    .valid_up(n885_valid_up),
    .valid_down(n885_valid_down),
    .I_0(n885_I_0),
    .I_1(n885_I_1),
    .I_2(n885_I_2),
    .I_3(n885_I_3),
    .I_4(n885_I_4),
    .I_5(n885_I_5),
    .I_6(n885_I_6),
    .I_7(n885_I_7),
    .O_0(n885_O_0),
    .O_1(n885_O_1),
    .O_2(n885_O_2),
    .O_3(n885_O_3),
    .O_4(n885_O_4),
    .O_5(n885_O_5),
    .O_6(n885_O_6),
    .O_7(n885_O_7)
  );
  ShiftTS_2 n886 ( // @[Top.scala 1047:22]
    .clock(n886_clock),
    .valid_up(n886_valid_up),
    .valid_down(n886_valid_down),
    .I_0(n886_I_0),
    .I_1(n886_I_1),
    .I_2(n886_I_2),
    .I_3(n886_I_3),
    .I_4(n886_I_4),
    .I_5(n886_I_5),
    .I_6(n886_I_6),
    .I_7(n886_I_7),
    .O_0(n886_O_0),
    .O_1(n886_O_1),
    .O_2(n886_O_2),
    .O_3(n886_O_3),
    .O_4(n886_O_4),
    .O_5(n886_O_5),
    .O_6(n886_O_6),
    .O_7(n886_O_7)
  );
  Map2T n887 ( // @[Top.scala 1050:22]
    .valid_up(n887_valid_up),
    .valid_down(n887_valid_down),
    .I0_0(n887_I0_0),
    .I0_1(n887_I0_1),
    .I0_2(n887_I0_2),
    .I0_3(n887_I0_3),
    .I0_4(n887_I0_4),
    .I0_5(n887_I0_5),
    .I0_6(n887_I0_6),
    .I0_7(n887_I0_7),
    .I1_0(n887_I1_0),
    .I1_1(n887_I1_1),
    .I1_2(n887_I1_2),
    .I1_3(n887_I1_3),
    .I1_4(n887_I1_4),
    .I1_5(n887_I1_5),
    .I1_6(n887_I1_6),
    .I1_7(n887_I1_7),
    .O_0_0(n887_O_0_0),
    .O_0_1(n887_O_0_1),
    .O_1_0(n887_O_1_0),
    .O_1_1(n887_O_1_1),
    .O_2_0(n887_O_2_0),
    .O_2_1(n887_O_2_1),
    .O_3_0(n887_O_3_0),
    .O_3_1(n887_O_3_1),
    .O_4_0(n887_O_4_0),
    .O_4_1(n887_O_4_1),
    .O_5_0(n887_O_5_0),
    .O_5_1(n887_O_5_1),
    .O_6_0(n887_O_6_0),
    .O_6_1(n887_O_6_1),
    .O_7_0(n887_O_7_0),
    .O_7_1(n887_O_7_1)
  );
  Map2T_1 n894 ( // @[Top.scala 1054:22]
    .valid_up(n894_valid_up),
    .valid_down(n894_valid_down),
    .I0_0_0(n894_I0_0_0),
    .I0_0_1(n894_I0_0_1),
    .I0_1_0(n894_I0_1_0),
    .I0_1_1(n894_I0_1_1),
    .I0_2_0(n894_I0_2_0),
    .I0_2_1(n894_I0_2_1),
    .I0_3_0(n894_I0_3_0),
    .I0_3_1(n894_I0_3_1),
    .I0_4_0(n894_I0_4_0),
    .I0_4_1(n894_I0_4_1),
    .I0_5_0(n894_I0_5_0),
    .I0_5_1(n894_I0_5_1),
    .I0_6_0(n894_I0_6_0),
    .I0_6_1(n894_I0_6_1),
    .I0_7_0(n894_I0_7_0),
    .I0_7_1(n894_I0_7_1),
    .I1_0(n894_I1_0),
    .I1_1(n894_I1_1),
    .I1_2(n894_I1_2),
    .I1_3(n894_I1_3),
    .I1_4(n894_I1_4),
    .I1_5(n894_I1_5),
    .I1_6(n894_I1_6),
    .I1_7(n894_I1_7),
    .O_0_0(n894_O_0_0),
    .O_0_1(n894_O_0_1),
    .O_0_2(n894_O_0_2),
    .O_1_0(n894_O_1_0),
    .O_1_1(n894_O_1_1),
    .O_1_2(n894_O_1_2),
    .O_2_0(n894_O_2_0),
    .O_2_1(n894_O_2_1),
    .O_2_2(n894_O_2_2),
    .O_3_0(n894_O_3_0),
    .O_3_1(n894_O_3_1),
    .O_3_2(n894_O_3_2),
    .O_4_0(n894_O_4_0),
    .O_4_1(n894_O_4_1),
    .O_4_2(n894_O_4_2),
    .O_5_0(n894_O_5_0),
    .O_5_1(n894_O_5_1),
    .O_5_2(n894_O_5_2),
    .O_6_0(n894_O_6_0),
    .O_6_1(n894_O_6_1),
    .O_6_2(n894_O_6_2),
    .O_7_0(n894_O_7_0),
    .O_7_1(n894_O_7_1),
    .O_7_2(n894_O_7_2)
  );
  MapT n903 ( // @[Top.scala 1058:22]
    .valid_up(n903_valid_up),
    .valid_down(n903_valid_down),
    .I_0_0(n903_I_0_0),
    .I_0_1(n903_I_0_1),
    .I_0_2(n903_I_0_2),
    .I_1_0(n903_I_1_0),
    .I_1_1(n903_I_1_1),
    .I_1_2(n903_I_1_2),
    .I_2_0(n903_I_2_0),
    .I_2_1(n903_I_2_1),
    .I_2_2(n903_I_2_2),
    .I_3_0(n903_I_3_0),
    .I_3_1(n903_I_3_1),
    .I_3_2(n903_I_3_2),
    .I_4_0(n903_I_4_0),
    .I_4_1(n903_I_4_1),
    .I_4_2(n903_I_4_2),
    .I_5_0(n903_I_5_0),
    .I_5_1(n903_I_5_1),
    .I_5_2(n903_I_5_2),
    .I_6_0(n903_I_6_0),
    .I_6_1(n903_I_6_1),
    .I_6_2(n903_I_6_2),
    .I_7_0(n903_I_7_0),
    .I_7_1(n903_I_7_1),
    .I_7_2(n903_I_7_2),
    .O_0_0_0(n903_O_0_0_0),
    .O_0_0_1(n903_O_0_0_1),
    .O_0_0_2(n903_O_0_0_2),
    .O_1_0_0(n903_O_1_0_0),
    .O_1_0_1(n903_O_1_0_1),
    .O_1_0_2(n903_O_1_0_2),
    .O_2_0_0(n903_O_2_0_0),
    .O_2_0_1(n903_O_2_0_1),
    .O_2_0_2(n903_O_2_0_2),
    .O_3_0_0(n903_O_3_0_0),
    .O_3_0_1(n903_O_3_0_1),
    .O_3_0_2(n903_O_3_0_2),
    .O_4_0_0(n903_O_4_0_0),
    .O_4_0_1(n903_O_4_0_1),
    .O_4_0_2(n903_O_4_0_2),
    .O_5_0_0(n903_O_5_0_0),
    .O_5_0_1(n903_O_5_0_1),
    .O_5_0_2(n903_O_5_0_2),
    .O_6_0_0(n903_O_6_0_0),
    .O_6_0_1(n903_O_6_0_1),
    .O_6_0_2(n903_O_6_0_2),
    .O_7_0_0(n903_O_7_0_0),
    .O_7_0_1(n903_O_7_0_1),
    .O_7_0_2(n903_O_7_0_2)
  );
  MapT_1 n910 ( // @[Top.scala 1061:22]
    .valid_up(n910_valid_up),
    .valid_down(n910_valid_down),
    .I_0_0_0(n910_I_0_0_0),
    .I_0_0_1(n910_I_0_0_1),
    .I_0_0_2(n910_I_0_0_2),
    .I_1_0_0(n910_I_1_0_0),
    .I_1_0_1(n910_I_1_0_1),
    .I_1_0_2(n910_I_1_0_2),
    .I_2_0_0(n910_I_2_0_0),
    .I_2_0_1(n910_I_2_0_1),
    .I_2_0_2(n910_I_2_0_2),
    .I_3_0_0(n910_I_3_0_0),
    .I_3_0_1(n910_I_3_0_1),
    .I_3_0_2(n910_I_3_0_2),
    .I_4_0_0(n910_I_4_0_0),
    .I_4_0_1(n910_I_4_0_1),
    .I_4_0_2(n910_I_4_0_2),
    .I_5_0_0(n910_I_5_0_0),
    .I_5_0_1(n910_I_5_0_1),
    .I_5_0_2(n910_I_5_0_2),
    .I_6_0_0(n910_I_6_0_0),
    .I_6_0_1(n910_I_6_0_1),
    .I_6_0_2(n910_I_6_0_2),
    .I_7_0_0(n910_I_7_0_0),
    .I_7_0_1(n910_I_7_0_1),
    .I_7_0_2(n910_I_7_0_2),
    .O_0_0(n910_O_0_0),
    .O_0_1(n910_O_0_1),
    .O_0_2(n910_O_0_2),
    .O_1_0(n910_O_1_0),
    .O_1_1(n910_O_1_1),
    .O_1_2(n910_O_1_2),
    .O_2_0(n910_O_2_0),
    .O_2_1(n910_O_2_1),
    .O_2_2(n910_O_2_2),
    .O_3_0(n910_O_3_0),
    .O_3_1(n910_O_3_1),
    .O_3_2(n910_O_3_2),
    .O_4_0(n910_O_4_0),
    .O_4_1(n910_O_4_1),
    .O_4_2(n910_O_4_2),
    .O_5_0(n910_O_5_0),
    .O_5_1(n910_O_5_1),
    .O_5_2(n910_O_5_2),
    .O_6_0(n910_O_6_0),
    .O_6_1(n910_O_6_1),
    .O_6_2(n910_O_6_2),
    .O_7_0(n910_O_7_0),
    .O_7_1(n910_O_7_1),
    .O_7_2(n910_O_7_2)
  );
  Map2T_7 n911 ( // @[Top.scala 1064:22]
    .valid_up(n911_valid_up),
    .valid_down(n911_valid_down),
    .I0_0_0_0(n911_I0_0_0_0),
    .I0_0_0_1(n911_I0_0_0_1),
    .I0_0_0_2(n911_I0_0_0_2),
    .I0_0_1_0(n911_I0_0_1_0),
    .I0_0_1_1(n911_I0_0_1_1),
    .I0_0_1_2(n911_I0_0_1_2),
    .I0_1_0_0(n911_I0_1_0_0),
    .I0_1_0_1(n911_I0_1_0_1),
    .I0_1_0_2(n911_I0_1_0_2),
    .I0_1_1_0(n911_I0_1_1_0),
    .I0_1_1_1(n911_I0_1_1_1),
    .I0_1_1_2(n911_I0_1_1_2),
    .I0_2_0_0(n911_I0_2_0_0),
    .I0_2_0_1(n911_I0_2_0_1),
    .I0_2_0_2(n911_I0_2_0_2),
    .I0_2_1_0(n911_I0_2_1_0),
    .I0_2_1_1(n911_I0_2_1_1),
    .I0_2_1_2(n911_I0_2_1_2),
    .I0_3_0_0(n911_I0_3_0_0),
    .I0_3_0_1(n911_I0_3_0_1),
    .I0_3_0_2(n911_I0_3_0_2),
    .I0_3_1_0(n911_I0_3_1_0),
    .I0_3_1_1(n911_I0_3_1_1),
    .I0_3_1_2(n911_I0_3_1_2),
    .I0_4_0_0(n911_I0_4_0_0),
    .I0_4_0_1(n911_I0_4_0_1),
    .I0_4_0_2(n911_I0_4_0_2),
    .I0_4_1_0(n911_I0_4_1_0),
    .I0_4_1_1(n911_I0_4_1_1),
    .I0_4_1_2(n911_I0_4_1_2),
    .I0_5_0_0(n911_I0_5_0_0),
    .I0_5_0_1(n911_I0_5_0_1),
    .I0_5_0_2(n911_I0_5_0_2),
    .I0_5_1_0(n911_I0_5_1_0),
    .I0_5_1_1(n911_I0_5_1_1),
    .I0_5_1_2(n911_I0_5_1_2),
    .I0_6_0_0(n911_I0_6_0_0),
    .I0_6_0_1(n911_I0_6_0_1),
    .I0_6_0_2(n911_I0_6_0_2),
    .I0_6_1_0(n911_I0_6_1_0),
    .I0_6_1_1(n911_I0_6_1_1),
    .I0_6_1_2(n911_I0_6_1_2),
    .I0_7_0_0(n911_I0_7_0_0),
    .I0_7_0_1(n911_I0_7_0_1),
    .I0_7_0_2(n911_I0_7_0_2),
    .I0_7_1_0(n911_I0_7_1_0),
    .I0_7_1_1(n911_I0_7_1_1),
    .I0_7_1_2(n911_I0_7_1_2),
    .I1_0_0(n911_I1_0_0),
    .I1_0_1(n911_I1_0_1),
    .I1_0_2(n911_I1_0_2),
    .I1_1_0(n911_I1_1_0),
    .I1_1_1(n911_I1_1_1),
    .I1_1_2(n911_I1_1_2),
    .I1_2_0(n911_I1_2_0),
    .I1_2_1(n911_I1_2_1),
    .I1_2_2(n911_I1_2_2),
    .I1_3_0(n911_I1_3_0),
    .I1_3_1(n911_I1_3_1),
    .I1_3_2(n911_I1_3_2),
    .I1_4_0(n911_I1_4_0),
    .I1_4_1(n911_I1_4_1),
    .I1_4_2(n911_I1_4_2),
    .I1_5_0(n911_I1_5_0),
    .I1_5_1(n911_I1_5_1),
    .I1_5_2(n911_I1_5_2),
    .I1_6_0(n911_I1_6_0),
    .I1_6_1(n911_I1_6_1),
    .I1_6_2(n911_I1_6_2),
    .I1_7_0(n911_I1_7_0),
    .I1_7_1(n911_I1_7_1),
    .I1_7_2(n911_I1_7_2),
    .O_0_0_0(n911_O_0_0_0),
    .O_0_0_1(n911_O_0_0_1),
    .O_0_0_2(n911_O_0_0_2),
    .O_0_1_0(n911_O_0_1_0),
    .O_0_1_1(n911_O_0_1_1),
    .O_0_1_2(n911_O_0_1_2),
    .O_0_2_0(n911_O_0_2_0),
    .O_0_2_1(n911_O_0_2_1),
    .O_0_2_2(n911_O_0_2_2),
    .O_1_0_0(n911_O_1_0_0),
    .O_1_0_1(n911_O_1_0_1),
    .O_1_0_2(n911_O_1_0_2),
    .O_1_1_0(n911_O_1_1_0),
    .O_1_1_1(n911_O_1_1_1),
    .O_1_1_2(n911_O_1_1_2),
    .O_1_2_0(n911_O_1_2_0),
    .O_1_2_1(n911_O_1_2_1),
    .O_1_2_2(n911_O_1_2_2),
    .O_2_0_0(n911_O_2_0_0),
    .O_2_0_1(n911_O_2_0_1),
    .O_2_0_2(n911_O_2_0_2),
    .O_2_1_0(n911_O_2_1_0),
    .O_2_1_1(n911_O_2_1_1),
    .O_2_1_2(n911_O_2_1_2),
    .O_2_2_0(n911_O_2_2_0),
    .O_2_2_1(n911_O_2_2_1),
    .O_2_2_2(n911_O_2_2_2),
    .O_3_0_0(n911_O_3_0_0),
    .O_3_0_1(n911_O_3_0_1),
    .O_3_0_2(n911_O_3_0_2),
    .O_3_1_0(n911_O_3_1_0),
    .O_3_1_1(n911_O_3_1_1),
    .O_3_1_2(n911_O_3_1_2),
    .O_3_2_0(n911_O_3_2_0),
    .O_3_2_1(n911_O_3_2_1),
    .O_3_2_2(n911_O_3_2_2),
    .O_4_0_0(n911_O_4_0_0),
    .O_4_0_1(n911_O_4_0_1),
    .O_4_0_2(n911_O_4_0_2),
    .O_4_1_0(n911_O_4_1_0),
    .O_4_1_1(n911_O_4_1_1),
    .O_4_1_2(n911_O_4_1_2),
    .O_4_2_0(n911_O_4_2_0),
    .O_4_2_1(n911_O_4_2_1),
    .O_4_2_2(n911_O_4_2_2),
    .O_5_0_0(n911_O_5_0_0),
    .O_5_0_1(n911_O_5_0_1),
    .O_5_0_2(n911_O_5_0_2),
    .O_5_1_0(n911_O_5_1_0),
    .O_5_1_1(n911_O_5_1_1),
    .O_5_1_2(n911_O_5_1_2),
    .O_5_2_0(n911_O_5_2_0),
    .O_5_2_1(n911_O_5_2_1),
    .O_5_2_2(n911_O_5_2_2),
    .O_6_0_0(n911_O_6_0_0),
    .O_6_0_1(n911_O_6_0_1),
    .O_6_0_2(n911_O_6_0_2),
    .O_6_1_0(n911_O_6_1_0),
    .O_6_1_1(n911_O_6_1_1),
    .O_6_1_2(n911_O_6_1_2),
    .O_6_2_0(n911_O_6_2_0),
    .O_6_2_1(n911_O_6_2_1),
    .O_6_2_2(n911_O_6_2_2),
    .O_7_0_0(n911_O_7_0_0),
    .O_7_0_1(n911_O_7_0_1),
    .O_7_0_2(n911_O_7_0_2),
    .O_7_1_0(n911_O_7_1_0),
    .O_7_1_1(n911_O_7_1_1),
    .O_7_1_2(n911_O_7_1_2),
    .O_7_2_0(n911_O_7_2_0),
    .O_7_2_1(n911_O_7_2_1),
    .O_7_2_2(n911_O_7_2_2)
  );
  MapT_6 n920 ( // @[Top.scala 1068:22]
    .valid_up(n920_valid_up),
    .valid_down(n920_valid_down),
    .I_0_0_0(n920_I_0_0_0),
    .I_0_0_1(n920_I_0_0_1),
    .I_0_0_2(n920_I_0_0_2),
    .I_0_1_0(n920_I_0_1_0),
    .I_0_1_1(n920_I_0_1_1),
    .I_0_1_2(n920_I_0_1_2),
    .I_0_2_0(n920_I_0_2_0),
    .I_0_2_1(n920_I_0_2_1),
    .I_0_2_2(n920_I_0_2_2),
    .I_1_0_0(n920_I_1_0_0),
    .I_1_0_1(n920_I_1_0_1),
    .I_1_0_2(n920_I_1_0_2),
    .I_1_1_0(n920_I_1_1_0),
    .I_1_1_1(n920_I_1_1_1),
    .I_1_1_2(n920_I_1_1_2),
    .I_1_2_0(n920_I_1_2_0),
    .I_1_2_1(n920_I_1_2_1),
    .I_1_2_2(n920_I_1_2_2),
    .I_2_0_0(n920_I_2_0_0),
    .I_2_0_1(n920_I_2_0_1),
    .I_2_0_2(n920_I_2_0_2),
    .I_2_1_0(n920_I_2_1_0),
    .I_2_1_1(n920_I_2_1_1),
    .I_2_1_2(n920_I_2_1_2),
    .I_2_2_0(n920_I_2_2_0),
    .I_2_2_1(n920_I_2_2_1),
    .I_2_2_2(n920_I_2_2_2),
    .I_3_0_0(n920_I_3_0_0),
    .I_3_0_1(n920_I_3_0_1),
    .I_3_0_2(n920_I_3_0_2),
    .I_3_1_0(n920_I_3_1_0),
    .I_3_1_1(n920_I_3_1_1),
    .I_3_1_2(n920_I_3_1_2),
    .I_3_2_0(n920_I_3_2_0),
    .I_3_2_1(n920_I_3_2_1),
    .I_3_2_2(n920_I_3_2_2),
    .I_4_0_0(n920_I_4_0_0),
    .I_4_0_1(n920_I_4_0_1),
    .I_4_0_2(n920_I_4_0_2),
    .I_4_1_0(n920_I_4_1_0),
    .I_4_1_1(n920_I_4_1_1),
    .I_4_1_2(n920_I_4_1_2),
    .I_4_2_0(n920_I_4_2_0),
    .I_4_2_1(n920_I_4_2_1),
    .I_4_2_2(n920_I_4_2_2),
    .I_5_0_0(n920_I_5_0_0),
    .I_5_0_1(n920_I_5_0_1),
    .I_5_0_2(n920_I_5_0_2),
    .I_5_1_0(n920_I_5_1_0),
    .I_5_1_1(n920_I_5_1_1),
    .I_5_1_2(n920_I_5_1_2),
    .I_5_2_0(n920_I_5_2_0),
    .I_5_2_1(n920_I_5_2_1),
    .I_5_2_2(n920_I_5_2_2),
    .I_6_0_0(n920_I_6_0_0),
    .I_6_0_1(n920_I_6_0_1),
    .I_6_0_2(n920_I_6_0_2),
    .I_6_1_0(n920_I_6_1_0),
    .I_6_1_1(n920_I_6_1_1),
    .I_6_1_2(n920_I_6_1_2),
    .I_6_2_0(n920_I_6_2_0),
    .I_6_2_1(n920_I_6_2_1),
    .I_6_2_2(n920_I_6_2_2),
    .I_7_0_0(n920_I_7_0_0),
    .I_7_0_1(n920_I_7_0_1),
    .I_7_0_2(n920_I_7_0_2),
    .I_7_1_0(n920_I_7_1_0),
    .I_7_1_1(n920_I_7_1_1),
    .I_7_1_2(n920_I_7_1_2),
    .I_7_2_0(n920_I_7_2_0),
    .I_7_2_1(n920_I_7_2_1),
    .I_7_2_2(n920_I_7_2_2),
    .O_0_0_0_0(n920_O_0_0_0_0),
    .O_0_0_0_1(n920_O_0_0_0_1),
    .O_0_0_0_2(n920_O_0_0_0_2),
    .O_0_0_1_0(n920_O_0_0_1_0),
    .O_0_0_1_1(n920_O_0_0_1_1),
    .O_0_0_1_2(n920_O_0_0_1_2),
    .O_0_0_2_0(n920_O_0_0_2_0),
    .O_0_0_2_1(n920_O_0_0_2_1),
    .O_0_0_2_2(n920_O_0_0_2_2),
    .O_1_0_0_0(n920_O_1_0_0_0),
    .O_1_0_0_1(n920_O_1_0_0_1),
    .O_1_0_0_2(n920_O_1_0_0_2),
    .O_1_0_1_0(n920_O_1_0_1_0),
    .O_1_0_1_1(n920_O_1_0_1_1),
    .O_1_0_1_2(n920_O_1_0_1_2),
    .O_1_0_2_0(n920_O_1_0_2_0),
    .O_1_0_2_1(n920_O_1_0_2_1),
    .O_1_0_2_2(n920_O_1_0_2_2),
    .O_2_0_0_0(n920_O_2_0_0_0),
    .O_2_0_0_1(n920_O_2_0_0_1),
    .O_2_0_0_2(n920_O_2_0_0_2),
    .O_2_0_1_0(n920_O_2_0_1_0),
    .O_2_0_1_1(n920_O_2_0_1_1),
    .O_2_0_1_2(n920_O_2_0_1_2),
    .O_2_0_2_0(n920_O_2_0_2_0),
    .O_2_0_2_1(n920_O_2_0_2_1),
    .O_2_0_2_2(n920_O_2_0_2_2),
    .O_3_0_0_0(n920_O_3_0_0_0),
    .O_3_0_0_1(n920_O_3_0_0_1),
    .O_3_0_0_2(n920_O_3_0_0_2),
    .O_3_0_1_0(n920_O_3_0_1_0),
    .O_3_0_1_1(n920_O_3_0_1_1),
    .O_3_0_1_2(n920_O_3_0_1_2),
    .O_3_0_2_0(n920_O_3_0_2_0),
    .O_3_0_2_1(n920_O_3_0_2_1),
    .O_3_0_2_2(n920_O_3_0_2_2),
    .O_4_0_0_0(n920_O_4_0_0_0),
    .O_4_0_0_1(n920_O_4_0_0_1),
    .O_4_0_0_2(n920_O_4_0_0_2),
    .O_4_0_1_0(n920_O_4_0_1_0),
    .O_4_0_1_1(n920_O_4_0_1_1),
    .O_4_0_1_2(n920_O_4_0_1_2),
    .O_4_0_2_0(n920_O_4_0_2_0),
    .O_4_0_2_1(n920_O_4_0_2_1),
    .O_4_0_2_2(n920_O_4_0_2_2),
    .O_5_0_0_0(n920_O_5_0_0_0),
    .O_5_0_0_1(n920_O_5_0_0_1),
    .O_5_0_0_2(n920_O_5_0_0_2),
    .O_5_0_1_0(n920_O_5_0_1_0),
    .O_5_0_1_1(n920_O_5_0_1_1),
    .O_5_0_1_2(n920_O_5_0_1_2),
    .O_5_0_2_0(n920_O_5_0_2_0),
    .O_5_0_2_1(n920_O_5_0_2_1),
    .O_5_0_2_2(n920_O_5_0_2_2),
    .O_6_0_0_0(n920_O_6_0_0_0),
    .O_6_0_0_1(n920_O_6_0_0_1),
    .O_6_0_0_2(n920_O_6_0_0_2),
    .O_6_0_1_0(n920_O_6_0_1_0),
    .O_6_0_1_1(n920_O_6_0_1_1),
    .O_6_0_1_2(n920_O_6_0_1_2),
    .O_6_0_2_0(n920_O_6_0_2_0),
    .O_6_0_2_1(n920_O_6_0_2_1),
    .O_6_0_2_2(n920_O_6_0_2_2),
    .O_7_0_0_0(n920_O_7_0_0_0),
    .O_7_0_0_1(n920_O_7_0_0_1),
    .O_7_0_0_2(n920_O_7_0_0_2),
    .O_7_0_1_0(n920_O_7_0_1_0),
    .O_7_0_1_1(n920_O_7_0_1_1),
    .O_7_0_1_2(n920_O_7_0_1_2),
    .O_7_0_2_0(n920_O_7_0_2_0),
    .O_7_0_2_1(n920_O_7_0_2_1),
    .O_7_0_2_2(n920_O_7_0_2_2)
  );
  MapT_7 n927 ( // @[Top.scala 1071:22]
    .valid_up(n927_valid_up),
    .valid_down(n927_valid_down),
    .I_0_0_0_0(n927_I_0_0_0_0),
    .I_0_0_0_1(n927_I_0_0_0_1),
    .I_0_0_0_2(n927_I_0_0_0_2),
    .I_0_0_1_0(n927_I_0_0_1_0),
    .I_0_0_1_1(n927_I_0_0_1_1),
    .I_0_0_1_2(n927_I_0_0_1_2),
    .I_0_0_2_0(n927_I_0_0_2_0),
    .I_0_0_2_1(n927_I_0_0_2_1),
    .I_0_0_2_2(n927_I_0_0_2_2),
    .I_1_0_0_0(n927_I_1_0_0_0),
    .I_1_0_0_1(n927_I_1_0_0_1),
    .I_1_0_0_2(n927_I_1_0_0_2),
    .I_1_0_1_0(n927_I_1_0_1_0),
    .I_1_0_1_1(n927_I_1_0_1_1),
    .I_1_0_1_2(n927_I_1_0_1_2),
    .I_1_0_2_0(n927_I_1_0_2_0),
    .I_1_0_2_1(n927_I_1_0_2_1),
    .I_1_0_2_2(n927_I_1_0_2_2),
    .I_2_0_0_0(n927_I_2_0_0_0),
    .I_2_0_0_1(n927_I_2_0_0_1),
    .I_2_0_0_2(n927_I_2_0_0_2),
    .I_2_0_1_0(n927_I_2_0_1_0),
    .I_2_0_1_1(n927_I_2_0_1_1),
    .I_2_0_1_2(n927_I_2_0_1_2),
    .I_2_0_2_0(n927_I_2_0_2_0),
    .I_2_0_2_1(n927_I_2_0_2_1),
    .I_2_0_2_2(n927_I_2_0_2_2),
    .I_3_0_0_0(n927_I_3_0_0_0),
    .I_3_0_0_1(n927_I_3_0_0_1),
    .I_3_0_0_2(n927_I_3_0_0_2),
    .I_3_0_1_0(n927_I_3_0_1_0),
    .I_3_0_1_1(n927_I_3_0_1_1),
    .I_3_0_1_2(n927_I_3_0_1_2),
    .I_3_0_2_0(n927_I_3_0_2_0),
    .I_3_0_2_1(n927_I_3_0_2_1),
    .I_3_0_2_2(n927_I_3_0_2_2),
    .I_4_0_0_0(n927_I_4_0_0_0),
    .I_4_0_0_1(n927_I_4_0_0_1),
    .I_4_0_0_2(n927_I_4_0_0_2),
    .I_4_0_1_0(n927_I_4_0_1_0),
    .I_4_0_1_1(n927_I_4_0_1_1),
    .I_4_0_1_2(n927_I_4_0_1_2),
    .I_4_0_2_0(n927_I_4_0_2_0),
    .I_4_0_2_1(n927_I_4_0_2_1),
    .I_4_0_2_2(n927_I_4_0_2_2),
    .I_5_0_0_0(n927_I_5_0_0_0),
    .I_5_0_0_1(n927_I_5_0_0_1),
    .I_5_0_0_2(n927_I_5_0_0_2),
    .I_5_0_1_0(n927_I_5_0_1_0),
    .I_5_0_1_1(n927_I_5_0_1_1),
    .I_5_0_1_2(n927_I_5_0_1_2),
    .I_5_0_2_0(n927_I_5_0_2_0),
    .I_5_0_2_1(n927_I_5_0_2_1),
    .I_5_0_2_2(n927_I_5_0_2_2),
    .I_6_0_0_0(n927_I_6_0_0_0),
    .I_6_0_0_1(n927_I_6_0_0_1),
    .I_6_0_0_2(n927_I_6_0_0_2),
    .I_6_0_1_0(n927_I_6_0_1_0),
    .I_6_0_1_1(n927_I_6_0_1_1),
    .I_6_0_1_2(n927_I_6_0_1_2),
    .I_6_0_2_0(n927_I_6_0_2_0),
    .I_6_0_2_1(n927_I_6_0_2_1),
    .I_6_0_2_2(n927_I_6_0_2_2),
    .I_7_0_0_0(n927_I_7_0_0_0),
    .I_7_0_0_1(n927_I_7_0_0_1),
    .I_7_0_0_2(n927_I_7_0_0_2),
    .I_7_0_1_0(n927_I_7_0_1_0),
    .I_7_0_1_1(n927_I_7_0_1_1),
    .I_7_0_1_2(n927_I_7_0_1_2),
    .I_7_0_2_0(n927_I_7_0_2_0),
    .I_7_0_2_1(n927_I_7_0_2_1),
    .I_7_0_2_2(n927_I_7_0_2_2),
    .O_0_0_0(n927_O_0_0_0),
    .O_0_0_1(n927_O_0_0_1),
    .O_0_0_2(n927_O_0_0_2),
    .O_0_1_0(n927_O_0_1_0),
    .O_0_1_1(n927_O_0_1_1),
    .O_0_1_2(n927_O_0_1_2),
    .O_0_2_0(n927_O_0_2_0),
    .O_0_2_1(n927_O_0_2_1),
    .O_0_2_2(n927_O_0_2_2),
    .O_1_0_0(n927_O_1_0_0),
    .O_1_0_1(n927_O_1_0_1),
    .O_1_0_2(n927_O_1_0_2),
    .O_1_1_0(n927_O_1_1_0),
    .O_1_1_1(n927_O_1_1_1),
    .O_1_1_2(n927_O_1_1_2),
    .O_1_2_0(n927_O_1_2_0),
    .O_1_2_1(n927_O_1_2_1),
    .O_1_2_2(n927_O_1_2_2),
    .O_2_0_0(n927_O_2_0_0),
    .O_2_0_1(n927_O_2_0_1),
    .O_2_0_2(n927_O_2_0_2),
    .O_2_1_0(n927_O_2_1_0),
    .O_2_1_1(n927_O_2_1_1),
    .O_2_1_2(n927_O_2_1_2),
    .O_2_2_0(n927_O_2_2_0),
    .O_2_2_1(n927_O_2_2_1),
    .O_2_2_2(n927_O_2_2_2),
    .O_3_0_0(n927_O_3_0_0),
    .O_3_0_1(n927_O_3_0_1),
    .O_3_0_2(n927_O_3_0_2),
    .O_3_1_0(n927_O_3_1_0),
    .O_3_1_1(n927_O_3_1_1),
    .O_3_1_2(n927_O_3_1_2),
    .O_3_2_0(n927_O_3_2_0),
    .O_3_2_1(n927_O_3_2_1),
    .O_3_2_2(n927_O_3_2_2),
    .O_4_0_0(n927_O_4_0_0),
    .O_4_0_1(n927_O_4_0_1),
    .O_4_0_2(n927_O_4_0_2),
    .O_4_1_0(n927_O_4_1_0),
    .O_4_1_1(n927_O_4_1_1),
    .O_4_1_2(n927_O_4_1_2),
    .O_4_2_0(n927_O_4_2_0),
    .O_4_2_1(n927_O_4_2_1),
    .O_4_2_2(n927_O_4_2_2),
    .O_5_0_0(n927_O_5_0_0),
    .O_5_0_1(n927_O_5_0_1),
    .O_5_0_2(n927_O_5_0_2),
    .O_5_1_0(n927_O_5_1_0),
    .O_5_1_1(n927_O_5_1_1),
    .O_5_1_2(n927_O_5_1_2),
    .O_5_2_0(n927_O_5_2_0),
    .O_5_2_1(n927_O_5_2_1),
    .O_5_2_2(n927_O_5_2_2),
    .O_6_0_0(n927_O_6_0_0),
    .O_6_0_1(n927_O_6_0_1),
    .O_6_0_2(n927_O_6_0_2),
    .O_6_1_0(n927_O_6_1_0),
    .O_6_1_1(n927_O_6_1_1),
    .O_6_1_2(n927_O_6_1_2),
    .O_6_2_0(n927_O_6_2_0),
    .O_6_2_1(n927_O_6_2_1),
    .O_6_2_2(n927_O_6_2_2),
    .O_7_0_0(n927_O_7_0_0),
    .O_7_0_1(n927_O_7_0_1),
    .O_7_0_2(n927_O_7_0_2),
    .O_7_1_0(n927_O_7_1_0),
    .O_7_1_1(n927_O_7_1_1),
    .O_7_1_2(n927_O_7_1_2),
    .O_7_2_0(n927_O_7_2_0),
    .O_7_2_1(n927_O_7_2_1),
    .O_7_2_2(n927_O_7_2_2)
  );
  MapT_42 n969 ( // @[Top.scala 1074:22]
    .clock(n969_clock),
    .reset(n969_reset),
    .valid_up(n969_valid_up),
    .valid_down(n969_valid_down),
    .I_0_0_0(n969_I_0_0_0),
    .I_0_0_1(n969_I_0_0_1),
    .I_0_0_2(n969_I_0_0_2),
    .I_0_1_0(n969_I_0_1_0),
    .I_0_1_1(n969_I_0_1_1),
    .I_0_1_2(n969_I_0_1_2),
    .I_0_2_0(n969_I_0_2_0),
    .I_0_2_1(n969_I_0_2_1),
    .I_0_2_2(n969_I_0_2_2),
    .I_1_0_0(n969_I_1_0_0),
    .I_1_0_1(n969_I_1_0_1),
    .I_1_0_2(n969_I_1_0_2),
    .I_1_1_0(n969_I_1_1_0),
    .I_1_1_1(n969_I_1_1_1),
    .I_1_1_2(n969_I_1_1_2),
    .I_1_2_0(n969_I_1_2_0),
    .I_1_2_1(n969_I_1_2_1),
    .I_1_2_2(n969_I_1_2_2),
    .I_2_0_0(n969_I_2_0_0),
    .I_2_0_1(n969_I_2_0_1),
    .I_2_0_2(n969_I_2_0_2),
    .I_2_1_0(n969_I_2_1_0),
    .I_2_1_1(n969_I_2_1_1),
    .I_2_1_2(n969_I_2_1_2),
    .I_2_2_0(n969_I_2_2_0),
    .I_2_2_1(n969_I_2_2_1),
    .I_2_2_2(n969_I_2_2_2),
    .I_3_0_0(n969_I_3_0_0),
    .I_3_0_1(n969_I_3_0_1),
    .I_3_0_2(n969_I_3_0_2),
    .I_3_1_0(n969_I_3_1_0),
    .I_3_1_1(n969_I_3_1_1),
    .I_3_1_2(n969_I_3_1_2),
    .I_3_2_0(n969_I_3_2_0),
    .I_3_2_1(n969_I_3_2_1),
    .I_3_2_2(n969_I_3_2_2),
    .I_4_0_0(n969_I_4_0_0),
    .I_4_0_1(n969_I_4_0_1),
    .I_4_0_2(n969_I_4_0_2),
    .I_4_1_0(n969_I_4_1_0),
    .I_4_1_1(n969_I_4_1_1),
    .I_4_1_2(n969_I_4_1_2),
    .I_4_2_0(n969_I_4_2_0),
    .I_4_2_1(n969_I_4_2_1),
    .I_4_2_2(n969_I_4_2_2),
    .I_5_0_0(n969_I_5_0_0),
    .I_5_0_1(n969_I_5_0_1),
    .I_5_0_2(n969_I_5_0_2),
    .I_5_1_0(n969_I_5_1_0),
    .I_5_1_1(n969_I_5_1_1),
    .I_5_1_2(n969_I_5_1_2),
    .I_5_2_0(n969_I_5_2_0),
    .I_5_2_1(n969_I_5_2_1),
    .I_5_2_2(n969_I_5_2_2),
    .I_6_0_0(n969_I_6_0_0),
    .I_6_0_1(n969_I_6_0_1),
    .I_6_0_2(n969_I_6_0_2),
    .I_6_1_0(n969_I_6_1_0),
    .I_6_1_1(n969_I_6_1_1),
    .I_6_1_2(n969_I_6_1_2),
    .I_6_2_0(n969_I_6_2_0),
    .I_6_2_1(n969_I_6_2_1),
    .I_6_2_2(n969_I_6_2_2),
    .I_7_0_0(n969_I_7_0_0),
    .I_7_0_1(n969_I_7_0_1),
    .I_7_0_2(n969_I_7_0_2),
    .I_7_1_0(n969_I_7_1_0),
    .I_7_1_1(n969_I_7_1_1),
    .I_7_1_2(n969_I_7_1_2),
    .I_7_2_0(n969_I_7_2_0),
    .I_7_2_1(n969_I_7_2_1),
    .I_7_2_2(n969_I_7_2_2),
    .O_0_0_0(n969_O_0_0_0),
    .O_1_0_0(n969_O_1_0_0),
    .O_2_0_0(n969_O_2_0_0),
    .O_3_0_0(n969_O_3_0_0),
    .O_4_0_0(n969_O_4_0_0),
    .O_5_0_0(n969_O_5_0_0),
    .O_6_0_0(n969_O_6_0_0),
    .O_7_0_0(n969_O_7_0_0)
  );
  Passthrough_4 n970 ( // @[Top.scala 1077:22]
    .valid_up(n970_valid_up),
    .valid_down(n970_valid_down),
    .I_0_0_0(n970_I_0_0_0),
    .I_1_0_0(n970_I_1_0_0),
    .I_2_0_0(n970_I_2_0_0),
    .I_3_0_0(n970_I_3_0_0),
    .I_4_0_0(n970_I_4_0_0),
    .I_5_0_0(n970_I_5_0_0),
    .I_6_0_0(n970_I_6_0_0),
    .I_7_0_0(n970_I_7_0_0),
    .O_0_0(n970_O_0_0),
    .O_1_0(n970_O_1_0),
    .O_2_0(n970_O_2_0),
    .O_3_0(n970_O_3_0),
    .O_4_0(n970_O_4_0),
    .O_5_0(n970_O_5_0),
    .O_6_0(n970_O_6_0),
    .O_7_0(n970_O_7_0)
  );
  Passthrough_5 n971 ( // @[Top.scala 1080:22]
    .valid_up(n971_valid_up),
    .valid_down(n971_valid_down),
    .I_0_0(n971_I_0_0),
    .I_1_0(n971_I_1_0),
    .I_2_0(n971_I_2_0),
    .I_3_0(n971_I_3_0),
    .I_4_0(n971_I_4_0),
    .I_5_0(n971_I_5_0),
    .I_6_0(n971_I_6_0),
    .I_7_0(n971_I_7_0),
    .O_0(n971_O_0),
    .O_1(n971_O_1),
    .O_2(n971_O_2),
    .O_3(n971_O_3),
    .O_4(n971_O_4),
    .O_5(n971_O_5),
    .O_6(n971_O_6),
    .O_7(n971_O_7)
  );
  FIFO_9 n972 ( // @[Top.scala 1083:22]
    .clock(n972_clock),
    .reset(n972_reset),
    .valid_up(n972_valid_up),
    .valid_down(n972_valid_down),
    .I_0(n972_I_0),
    .I_1(n972_I_1),
    .I_2(n972_I_2),
    .I_3(n972_I_3),
    .I_4(n972_I_4),
    .I_5(n972_I_5),
    .I_6(n972_I_6),
    .I_7(n972_I_7),
    .O_0(n972_O_0),
    .O_1(n972_O_1),
    .O_2(n972_O_2),
    .O_3(n972_O_3),
    .O_4(n972_O_4),
    .O_5(n972_O_5),
    .O_6(n972_O_6),
    .O_7(n972_O_7)
  );
  Map2T_18 n973 ( // @[Top.scala 1086:22]
    .clock(n973_clock),
    .reset(n973_reset),
    .valid_up(n973_valid_up),
    .valid_down(n973_valid_down),
    .I0_0(n973_I0_0),
    .I0_1(n973_I0_1),
    .I0_2(n973_I0_2),
    .I0_3(n973_I0_3),
    .I0_4(n973_I0_4),
    .I0_5(n973_I0_5),
    .I0_6(n973_I0_6),
    .I0_7(n973_I0_7),
    .I1_0(n973_I1_0),
    .I1_1(n973_I1_1),
    .I1_2(n973_I1_2),
    .I1_3(n973_I1_3),
    .I1_4(n973_I1_4),
    .I1_5(n973_I1_5),
    .I1_6(n973_I1_6),
    .I1_7(n973_I1_7),
    .O_0(n973_O_0),
    .O_1(n973_O_1),
    .O_2(n973_O_2),
    .O_3(n973_O_3),
    .O_4(n973_O_4),
    .O_5(n973_O_5),
    .O_6(n973_O_6),
    .O_7(n973_O_7)
  );
  Map2T_37 n1004 ( // @[Top.scala 1090:23]
    .valid_up(n1004_valid_up),
    .valid_down(n1004_valid_down),
    .I0_0(n1004_I0_0),
    .I0_1(n1004_I0_1),
    .I0_2(n1004_I0_2),
    .I0_3(n1004_I0_3),
    .I0_4(n1004_I0_4),
    .I0_5(n1004_I0_5),
    .I0_6(n1004_I0_6),
    .I0_7(n1004_I0_7),
    .I1_0(n1004_I1_0),
    .I1_1(n1004_I1_1),
    .I1_2(n1004_I1_2),
    .I1_3(n1004_I1_3),
    .I1_4(n1004_I1_4),
    .I1_5(n1004_I1_5),
    .I1_6(n1004_I1_6),
    .I1_7(n1004_I1_7),
    .O_0_t0b(n1004_O_0_t0b),
    .O_0_t1b(n1004_O_0_t1b),
    .O_1_t0b(n1004_O_1_t0b),
    .O_1_t1b(n1004_O_1_t1b),
    .O_2_t0b(n1004_O_2_t0b),
    .O_2_t1b(n1004_O_2_t1b),
    .O_3_t0b(n1004_O_3_t0b),
    .O_3_t1b(n1004_O_3_t1b),
    .O_4_t0b(n1004_O_4_t0b),
    .O_4_t1b(n1004_O_4_t1b),
    .O_5_t0b(n1004_O_5_t0b),
    .O_5_t1b(n1004_O_5_t1b),
    .O_6_t0b(n1004_O_6_t0b),
    .O_6_t1b(n1004_O_6_t1b),
    .O_7_t0b(n1004_O_7_t0b),
    .O_7_t1b(n1004_O_7_t1b)
  );
  Map2T_38 n1011 ( // @[Top.scala 1094:23]
    .valid_up(n1011_valid_up),
    .valid_down(n1011_valid_down),
    .I0_0(n1011_I0_0),
    .I0_1(n1011_I0_1),
    .I0_2(n1011_I0_2),
    .I0_3(n1011_I0_3),
    .I0_4(n1011_I0_4),
    .I0_5(n1011_I0_5),
    .I0_6(n1011_I0_6),
    .I0_7(n1011_I0_7),
    .I1_0_t0b(n1011_I1_0_t0b),
    .I1_0_t1b(n1011_I1_0_t1b),
    .I1_1_t0b(n1011_I1_1_t0b),
    .I1_1_t1b(n1011_I1_1_t1b),
    .I1_2_t0b(n1011_I1_2_t0b),
    .I1_2_t1b(n1011_I1_2_t1b),
    .I1_3_t0b(n1011_I1_3_t0b),
    .I1_3_t1b(n1011_I1_3_t1b),
    .I1_4_t0b(n1011_I1_4_t0b),
    .I1_4_t1b(n1011_I1_4_t1b),
    .I1_5_t0b(n1011_I1_5_t0b),
    .I1_5_t1b(n1011_I1_5_t1b),
    .I1_6_t0b(n1011_I1_6_t0b),
    .I1_6_t1b(n1011_I1_6_t1b),
    .I1_7_t0b(n1011_I1_7_t0b),
    .I1_7_t1b(n1011_I1_7_t1b),
    .O_0_t0b(n1011_O_0_t0b),
    .O_0_t1b_t0b(n1011_O_0_t1b_t0b),
    .O_0_t1b_t1b(n1011_O_0_t1b_t1b),
    .O_1_t0b(n1011_O_1_t0b),
    .O_1_t1b_t0b(n1011_O_1_t1b_t0b),
    .O_1_t1b_t1b(n1011_O_1_t1b_t1b),
    .O_2_t0b(n1011_O_2_t0b),
    .O_2_t1b_t0b(n1011_O_2_t1b_t0b),
    .O_2_t1b_t1b(n1011_O_2_t1b_t1b),
    .O_3_t0b(n1011_O_3_t0b),
    .O_3_t1b_t0b(n1011_O_3_t1b_t0b),
    .O_3_t1b_t1b(n1011_O_3_t1b_t1b),
    .O_4_t0b(n1011_O_4_t0b),
    .O_4_t1b_t0b(n1011_O_4_t1b_t0b),
    .O_4_t1b_t1b(n1011_O_4_t1b_t1b),
    .O_5_t0b(n1011_O_5_t0b),
    .O_5_t1b_t0b(n1011_O_5_t1b_t0b),
    .O_5_t1b_t1b(n1011_O_5_t1b_t1b),
    .O_6_t0b(n1011_O_6_t0b),
    .O_6_t1b_t0b(n1011_O_6_t1b_t0b),
    .O_6_t1b_t1b(n1011_O_6_t1b_t1b),
    .O_7_t0b(n1011_O_7_t0b),
    .O_7_t1b_t0b(n1011_O_7_t1b_t0b),
    .O_7_t1b_t1b(n1011_O_7_t1b_t1b)
  );
  FIFO_15 n1018 ( // @[Top.scala 1098:23]
    .clock(n1018_clock),
    .reset(n1018_reset),
    .valid_up(n1018_valid_up),
    .valid_down(n1018_valid_down),
    .I_0_t0b(n1018_I_0_t0b),
    .I_0_t1b_t0b(n1018_I_0_t1b_t0b),
    .I_0_t1b_t1b(n1018_I_0_t1b_t1b),
    .I_1_t0b(n1018_I_1_t0b),
    .I_1_t1b_t0b(n1018_I_1_t1b_t0b),
    .I_1_t1b_t1b(n1018_I_1_t1b_t1b),
    .I_2_t0b(n1018_I_2_t0b),
    .I_2_t1b_t0b(n1018_I_2_t1b_t0b),
    .I_2_t1b_t1b(n1018_I_2_t1b_t1b),
    .I_3_t0b(n1018_I_3_t0b),
    .I_3_t1b_t0b(n1018_I_3_t1b_t0b),
    .I_3_t1b_t1b(n1018_I_3_t1b_t1b),
    .I_4_t0b(n1018_I_4_t0b),
    .I_4_t1b_t0b(n1018_I_4_t1b_t0b),
    .I_4_t1b_t1b(n1018_I_4_t1b_t1b),
    .I_5_t0b(n1018_I_5_t0b),
    .I_5_t1b_t0b(n1018_I_5_t1b_t0b),
    .I_5_t1b_t1b(n1018_I_5_t1b_t1b),
    .I_6_t0b(n1018_I_6_t0b),
    .I_6_t1b_t0b(n1018_I_6_t1b_t0b),
    .I_6_t1b_t1b(n1018_I_6_t1b_t1b),
    .I_7_t0b(n1018_I_7_t0b),
    .I_7_t1b_t0b(n1018_I_7_t1b_t0b),
    .I_7_t1b_t1b(n1018_I_7_t1b_t1b),
    .O_0_t0b(n1018_O_0_t0b),
    .O_0_t1b_t0b(n1018_O_0_t1b_t0b),
    .O_0_t1b_t1b(n1018_O_0_t1b_t1b),
    .O_1_t0b(n1018_O_1_t0b),
    .O_1_t1b_t0b(n1018_O_1_t1b_t0b),
    .O_1_t1b_t1b(n1018_O_1_t1b_t1b),
    .O_2_t0b(n1018_O_2_t0b),
    .O_2_t1b_t0b(n1018_O_2_t1b_t0b),
    .O_2_t1b_t1b(n1018_O_2_t1b_t1b),
    .O_3_t0b(n1018_O_3_t0b),
    .O_3_t1b_t0b(n1018_O_3_t1b_t0b),
    .O_3_t1b_t1b(n1018_O_3_t1b_t1b),
    .O_4_t0b(n1018_O_4_t0b),
    .O_4_t1b_t0b(n1018_O_4_t1b_t0b),
    .O_4_t1b_t1b(n1018_O_4_t1b_t1b),
    .O_5_t0b(n1018_O_5_t0b),
    .O_5_t1b_t0b(n1018_O_5_t1b_t0b),
    .O_5_t1b_t1b(n1018_O_5_t1b_t1b),
    .O_6_t0b(n1018_O_6_t0b),
    .O_6_t1b_t0b(n1018_O_6_t1b_t0b),
    .O_6_t1b_t1b(n1018_O_6_t1b_t1b),
    .O_7_t0b(n1018_O_7_t0b),
    .O_7_t1b_t0b(n1018_O_7_t1b_t0b),
    .O_7_t1b_t1b(n1018_O_7_t1b_t1b)
  );
  FIFO_15 n1019 ( // @[Top.scala 1101:23]
    .clock(n1019_clock),
    .reset(n1019_reset),
    .valid_up(n1019_valid_up),
    .valid_down(n1019_valid_down),
    .I_0_t0b(n1019_I_0_t0b),
    .I_0_t1b_t0b(n1019_I_0_t1b_t0b),
    .I_0_t1b_t1b(n1019_I_0_t1b_t1b),
    .I_1_t0b(n1019_I_1_t0b),
    .I_1_t1b_t0b(n1019_I_1_t1b_t0b),
    .I_1_t1b_t1b(n1019_I_1_t1b_t1b),
    .I_2_t0b(n1019_I_2_t0b),
    .I_2_t1b_t0b(n1019_I_2_t1b_t0b),
    .I_2_t1b_t1b(n1019_I_2_t1b_t1b),
    .I_3_t0b(n1019_I_3_t0b),
    .I_3_t1b_t0b(n1019_I_3_t1b_t0b),
    .I_3_t1b_t1b(n1019_I_3_t1b_t1b),
    .I_4_t0b(n1019_I_4_t0b),
    .I_4_t1b_t0b(n1019_I_4_t1b_t0b),
    .I_4_t1b_t1b(n1019_I_4_t1b_t1b),
    .I_5_t0b(n1019_I_5_t0b),
    .I_5_t1b_t0b(n1019_I_5_t1b_t0b),
    .I_5_t1b_t1b(n1019_I_5_t1b_t1b),
    .I_6_t0b(n1019_I_6_t0b),
    .I_6_t1b_t0b(n1019_I_6_t1b_t0b),
    .I_6_t1b_t1b(n1019_I_6_t1b_t1b),
    .I_7_t0b(n1019_I_7_t0b),
    .I_7_t1b_t0b(n1019_I_7_t1b_t0b),
    .I_7_t1b_t1b(n1019_I_7_t1b_t1b),
    .O_0_t0b(n1019_O_0_t0b),
    .O_0_t1b_t0b(n1019_O_0_t1b_t0b),
    .O_0_t1b_t1b(n1019_O_0_t1b_t1b),
    .O_1_t0b(n1019_O_1_t0b),
    .O_1_t1b_t0b(n1019_O_1_t1b_t0b),
    .O_1_t1b_t1b(n1019_O_1_t1b_t1b),
    .O_2_t0b(n1019_O_2_t0b),
    .O_2_t1b_t0b(n1019_O_2_t1b_t0b),
    .O_2_t1b_t1b(n1019_O_2_t1b_t1b),
    .O_3_t0b(n1019_O_3_t0b),
    .O_3_t1b_t0b(n1019_O_3_t1b_t0b),
    .O_3_t1b_t1b(n1019_O_3_t1b_t1b),
    .O_4_t0b(n1019_O_4_t0b),
    .O_4_t1b_t0b(n1019_O_4_t1b_t0b),
    .O_4_t1b_t1b(n1019_O_4_t1b_t1b),
    .O_5_t0b(n1019_O_5_t0b),
    .O_5_t1b_t0b(n1019_O_5_t1b_t0b),
    .O_5_t1b_t1b(n1019_O_5_t1b_t1b),
    .O_6_t0b(n1019_O_6_t0b),
    .O_6_t1b_t0b(n1019_O_6_t1b_t0b),
    .O_6_t1b_t1b(n1019_O_6_t1b_t1b),
    .O_7_t0b(n1019_O_7_t0b),
    .O_7_t1b_t0b(n1019_O_7_t1b_t0b),
    .O_7_t1b_t1b(n1019_O_7_t1b_t1b)
  );
  FIFO_15 n1020 ( // @[Top.scala 1104:23]
    .clock(n1020_clock),
    .reset(n1020_reset),
    .valid_up(n1020_valid_up),
    .valid_down(n1020_valid_down),
    .I_0_t0b(n1020_I_0_t0b),
    .I_0_t1b_t0b(n1020_I_0_t1b_t0b),
    .I_0_t1b_t1b(n1020_I_0_t1b_t1b),
    .I_1_t0b(n1020_I_1_t0b),
    .I_1_t1b_t0b(n1020_I_1_t1b_t0b),
    .I_1_t1b_t1b(n1020_I_1_t1b_t1b),
    .I_2_t0b(n1020_I_2_t0b),
    .I_2_t1b_t0b(n1020_I_2_t1b_t0b),
    .I_2_t1b_t1b(n1020_I_2_t1b_t1b),
    .I_3_t0b(n1020_I_3_t0b),
    .I_3_t1b_t0b(n1020_I_3_t1b_t0b),
    .I_3_t1b_t1b(n1020_I_3_t1b_t1b),
    .I_4_t0b(n1020_I_4_t0b),
    .I_4_t1b_t0b(n1020_I_4_t1b_t0b),
    .I_4_t1b_t1b(n1020_I_4_t1b_t1b),
    .I_5_t0b(n1020_I_5_t0b),
    .I_5_t1b_t0b(n1020_I_5_t1b_t0b),
    .I_5_t1b_t1b(n1020_I_5_t1b_t1b),
    .I_6_t0b(n1020_I_6_t0b),
    .I_6_t1b_t0b(n1020_I_6_t1b_t0b),
    .I_6_t1b_t1b(n1020_I_6_t1b_t1b),
    .I_7_t0b(n1020_I_7_t0b),
    .I_7_t1b_t0b(n1020_I_7_t1b_t0b),
    .I_7_t1b_t1b(n1020_I_7_t1b_t1b),
    .O_0_t0b(n1020_O_0_t0b),
    .O_0_t1b_t0b(n1020_O_0_t1b_t0b),
    .O_0_t1b_t1b(n1020_O_0_t1b_t1b),
    .O_1_t0b(n1020_O_1_t0b),
    .O_1_t1b_t0b(n1020_O_1_t1b_t0b),
    .O_1_t1b_t1b(n1020_O_1_t1b_t1b),
    .O_2_t0b(n1020_O_2_t0b),
    .O_2_t1b_t0b(n1020_O_2_t1b_t0b),
    .O_2_t1b_t1b(n1020_O_2_t1b_t1b),
    .O_3_t0b(n1020_O_3_t0b),
    .O_3_t1b_t0b(n1020_O_3_t1b_t0b),
    .O_3_t1b_t1b(n1020_O_3_t1b_t1b),
    .O_4_t0b(n1020_O_4_t0b),
    .O_4_t1b_t0b(n1020_O_4_t1b_t0b),
    .O_4_t1b_t1b(n1020_O_4_t1b_t1b),
    .O_5_t0b(n1020_O_5_t0b),
    .O_5_t1b_t0b(n1020_O_5_t1b_t0b),
    .O_5_t1b_t1b(n1020_O_5_t1b_t1b),
    .O_6_t0b(n1020_O_6_t0b),
    .O_6_t1b_t0b(n1020_O_6_t1b_t0b),
    .O_6_t1b_t1b(n1020_O_6_t1b_t1b),
    .O_7_t0b(n1020_O_7_t0b),
    .O_7_t1b_t0b(n1020_O_7_t1b_t0b),
    .O_7_t1b_t1b(n1020_O_7_t1b_t1b)
  );
  assign valid_down = n1020_valid_down; // @[Top.scala 1108:16]
  assign O_0_t0b = n1020_O_0_t0b; // @[Top.scala 1107:7]
  assign O_0_t1b_t0b = n1020_O_0_t1b_t0b; // @[Top.scala 1107:7]
  assign O_0_t1b_t1b = n1020_O_0_t1b_t1b; // @[Top.scala 1107:7]
  assign O_1_t0b = n1020_O_1_t0b; // @[Top.scala 1107:7]
  assign O_1_t1b_t0b = n1020_O_1_t1b_t0b; // @[Top.scala 1107:7]
  assign O_1_t1b_t1b = n1020_O_1_t1b_t1b; // @[Top.scala 1107:7]
  assign O_2_t0b = n1020_O_2_t0b; // @[Top.scala 1107:7]
  assign O_2_t1b_t0b = n1020_O_2_t1b_t0b; // @[Top.scala 1107:7]
  assign O_2_t1b_t1b = n1020_O_2_t1b_t1b; // @[Top.scala 1107:7]
  assign O_3_t0b = n1020_O_3_t0b; // @[Top.scala 1107:7]
  assign O_3_t1b_t0b = n1020_O_3_t1b_t0b; // @[Top.scala 1107:7]
  assign O_3_t1b_t1b = n1020_O_3_t1b_t1b; // @[Top.scala 1107:7]
  assign O_4_t0b = n1020_O_4_t0b; // @[Top.scala 1107:7]
  assign O_4_t1b_t0b = n1020_O_4_t1b_t0b; // @[Top.scala 1107:7]
  assign O_4_t1b_t1b = n1020_O_4_t1b_t1b; // @[Top.scala 1107:7]
  assign O_5_t0b = n1020_O_5_t0b; // @[Top.scala 1107:7]
  assign O_5_t1b_t0b = n1020_O_5_t1b_t0b; // @[Top.scala 1107:7]
  assign O_5_t1b_t1b = n1020_O_5_t1b_t1b; // @[Top.scala 1107:7]
  assign O_6_t0b = n1020_O_6_t0b; // @[Top.scala 1107:7]
  assign O_6_t1b_t0b = n1020_O_6_t1b_t0b; // @[Top.scala 1107:7]
  assign O_6_t1b_t1b = n1020_O_6_t1b_t1b; // @[Top.scala 1107:7]
  assign O_7_t0b = n1020_O_7_t0b; // @[Top.scala 1107:7]
  assign O_7_t1b_t0b = n1020_O_7_t1b_t0b; // @[Top.scala 1107:7]
  assign O_7_t1b_t1b = n1020_O_7_t1b_t1b; // @[Top.scala 1107:7]
  assign n1_clock = clock;
  assign n1_reset = reset;
  assign n1_valid_up = valid_up; // @[Top.scala 697:17]
  assign n1_I_0 = I_0; // @[Top.scala 696:10]
  assign n1_I_1 = I_1; // @[Top.scala 696:10]
  assign n1_I_2 = I_2; // @[Top.scala 696:10]
  assign n1_I_3 = I_3; // @[Top.scala 696:10]
  assign n1_I_4 = I_4; // @[Top.scala 696:10]
  assign n1_I_5 = I_5; // @[Top.scala 696:10]
  assign n1_I_6 = I_6; // @[Top.scala 696:10]
  assign n1_I_7 = I_7; // @[Top.scala 696:10]
  assign n2_clock = clock;
  assign n2_reset = reset;
  assign n2_valid_up = n1_valid_down; // @[Top.scala 700:17]
  assign n2_I_0 = n1_O_0; // @[Top.scala 699:10]
  assign n2_I_1 = n1_O_1; // @[Top.scala 699:10]
  assign n2_I_2 = n1_O_2; // @[Top.scala 699:10]
  assign n2_I_3 = n1_O_3; // @[Top.scala 699:10]
  assign n2_I_4 = n1_O_4; // @[Top.scala 699:10]
  assign n2_I_5 = n1_O_5; // @[Top.scala 699:10]
  assign n2_I_6 = n1_O_6; // @[Top.scala 699:10]
  assign n2_I_7 = n1_O_7; // @[Top.scala 699:10]
  assign n3_clock = clock;
  assign n3_reset = reset;
  assign n3_valid_up = n2_valid_down; // @[Top.scala 703:17]
  assign n3_I_0 = n2_O_0; // @[Top.scala 702:10]
  assign n3_I_1 = n2_O_1; // @[Top.scala 702:10]
  assign n3_I_2 = n2_O_2; // @[Top.scala 702:10]
  assign n3_I_3 = n2_O_3; // @[Top.scala 702:10]
  assign n3_I_4 = n2_O_4; // @[Top.scala 702:10]
  assign n3_I_5 = n2_O_5; // @[Top.scala 702:10]
  assign n3_I_6 = n2_O_6; // @[Top.scala 702:10]
  assign n3_I_7 = n2_O_7; // @[Top.scala 702:10]
  assign n4_clock = clock;
  assign n4_valid_up = n3_valid_down; // @[Top.scala 706:17]
  assign n4_I_0 = n3_O_0; // @[Top.scala 705:10]
  assign n4_I_1 = n3_O_1; // @[Top.scala 705:10]
  assign n4_I_2 = n3_O_2; // @[Top.scala 705:10]
  assign n4_I_3 = n3_O_3; // @[Top.scala 705:10]
  assign n4_I_4 = n3_O_4; // @[Top.scala 705:10]
  assign n4_I_5 = n3_O_5; // @[Top.scala 705:10]
  assign n4_I_6 = n3_O_6; // @[Top.scala 705:10]
  assign n4_I_7 = n3_O_7; // @[Top.scala 705:10]
  assign n5_clock = clock;
  assign n5_valid_up = n4_valid_down; // @[Top.scala 709:17]
  assign n5_I_0 = n4_O_0; // @[Top.scala 708:10]
  assign n5_I_1 = n4_O_1; // @[Top.scala 708:10]
  assign n5_I_2 = n4_O_2; // @[Top.scala 708:10]
  assign n5_I_3 = n4_O_3; // @[Top.scala 708:10]
  assign n5_I_4 = n4_O_4; // @[Top.scala 708:10]
  assign n5_I_5 = n4_O_5; // @[Top.scala 708:10]
  assign n5_I_6 = n4_O_6; // @[Top.scala 708:10]
  assign n5_I_7 = n4_O_7; // @[Top.scala 708:10]
  assign n6_valid_up = n5_valid_down & n4_valid_down; // @[Top.scala 713:17]
  assign n6_I0_0 = n5_O_0; // @[Top.scala 711:11]
  assign n6_I0_1 = n5_O_1; // @[Top.scala 711:11]
  assign n6_I0_2 = n5_O_2; // @[Top.scala 711:11]
  assign n6_I0_3 = n5_O_3; // @[Top.scala 711:11]
  assign n6_I0_4 = n5_O_4; // @[Top.scala 711:11]
  assign n6_I0_5 = n5_O_5; // @[Top.scala 711:11]
  assign n6_I0_6 = n5_O_6; // @[Top.scala 711:11]
  assign n6_I0_7 = n5_O_7; // @[Top.scala 711:11]
  assign n6_I1_0 = n4_O_0; // @[Top.scala 712:11]
  assign n6_I1_1 = n4_O_1; // @[Top.scala 712:11]
  assign n6_I1_2 = n4_O_2; // @[Top.scala 712:11]
  assign n6_I1_3 = n4_O_3; // @[Top.scala 712:11]
  assign n6_I1_4 = n4_O_4; // @[Top.scala 712:11]
  assign n6_I1_5 = n4_O_5; // @[Top.scala 712:11]
  assign n6_I1_6 = n4_O_6; // @[Top.scala 712:11]
  assign n6_I1_7 = n4_O_7; // @[Top.scala 712:11]
  assign n13_valid_up = n6_valid_down & n3_valid_down; // @[Top.scala 717:18]
  assign n13_I0_0_0 = n6_O_0_0; // @[Top.scala 715:12]
  assign n13_I0_0_1 = n6_O_0_1; // @[Top.scala 715:12]
  assign n13_I0_1_0 = n6_O_1_0; // @[Top.scala 715:12]
  assign n13_I0_1_1 = n6_O_1_1; // @[Top.scala 715:12]
  assign n13_I0_2_0 = n6_O_2_0; // @[Top.scala 715:12]
  assign n13_I0_2_1 = n6_O_2_1; // @[Top.scala 715:12]
  assign n13_I0_3_0 = n6_O_3_0; // @[Top.scala 715:12]
  assign n13_I0_3_1 = n6_O_3_1; // @[Top.scala 715:12]
  assign n13_I0_4_0 = n6_O_4_0; // @[Top.scala 715:12]
  assign n13_I0_4_1 = n6_O_4_1; // @[Top.scala 715:12]
  assign n13_I0_5_0 = n6_O_5_0; // @[Top.scala 715:12]
  assign n13_I0_5_1 = n6_O_5_1; // @[Top.scala 715:12]
  assign n13_I0_6_0 = n6_O_6_0; // @[Top.scala 715:12]
  assign n13_I0_6_1 = n6_O_6_1; // @[Top.scala 715:12]
  assign n13_I0_7_0 = n6_O_7_0; // @[Top.scala 715:12]
  assign n13_I0_7_1 = n6_O_7_1; // @[Top.scala 715:12]
  assign n13_I1_0 = n3_O_0; // @[Top.scala 716:12]
  assign n13_I1_1 = n3_O_1; // @[Top.scala 716:12]
  assign n13_I1_2 = n3_O_2; // @[Top.scala 716:12]
  assign n13_I1_3 = n3_O_3; // @[Top.scala 716:12]
  assign n13_I1_4 = n3_O_4; // @[Top.scala 716:12]
  assign n13_I1_5 = n3_O_5; // @[Top.scala 716:12]
  assign n13_I1_6 = n3_O_6; // @[Top.scala 716:12]
  assign n13_I1_7 = n3_O_7; // @[Top.scala 716:12]
  assign n22_valid_up = n13_valid_down; // @[Top.scala 720:18]
  assign n22_I_0_0 = n13_O_0_0; // @[Top.scala 719:11]
  assign n22_I_0_1 = n13_O_0_1; // @[Top.scala 719:11]
  assign n22_I_0_2 = n13_O_0_2; // @[Top.scala 719:11]
  assign n22_I_1_0 = n13_O_1_0; // @[Top.scala 719:11]
  assign n22_I_1_1 = n13_O_1_1; // @[Top.scala 719:11]
  assign n22_I_1_2 = n13_O_1_2; // @[Top.scala 719:11]
  assign n22_I_2_0 = n13_O_2_0; // @[Top.scala 719:11]
  assign n22_I_2_1 = n13_O_2_1; // @[Top.scala 719:11]
  assign n22_I_2_2 = n13_O_2_2; // @[Top.scala 719:11]
  assign n22_I_3_0 = n13_O_3_0; // @[Top.scala 719:11]
  assign n22_I_3_1 = n13_O_3_1; // @[Top.scala 719:11]
  assign n22_I_3_2 = n13_O_3_2; // @[Top.scala 719:11]
  assign n22_I_4_0 = n13_O_4_0; // @[Top.scala 719:11]
  assign n22_I_4_1 = n13_O_4_1; // @[Top.scala 719:11]
  assign n22_I_4_2 = n13_O_4_2; // @[Top.scala 719:11]
  assign n22_I_5_0 = n13_O_5_0; // @[Top.scala 719:11]
  assign n22_I_5_1 = n13_O_5_1; // @[Top.scala 719:11]
  assign n22_I_5_2 = n13_O_5_2; // @[Top.scala 719:11]
  assign n22_I_6_0 = n13_O_6_0; // @[Top.scala 719:11]
  assign n22_I_6_1 = n13_O_6_1; // @[Top.scala 719:11]
  assign n22_I_6_2 = n13_O_6_2; // @[Top.scala 719:11]
  assign n22_I_7_0 = n13_O_7_0; // @[Top.scala 719:11]
  assign n22_I_7_1 = n13_O_7_1; // @[Top.scala 719:11]
  assign n22_I_7_2 = n13_O_7_2; // @[Top.scala 719:11]
  assign n29_valid_up = n22_valid_down; // @[Top.scala 723:18]
  assign n29_I_0_0_0 = n22_O_0_0_0; // @[Top.scala 722:11]
  assign n29_I_0_0_1 = n22_O_0_0_1; // @[Top.scala 722:11]
  assign n29_I_0_0_2 = n22_O_0_0_2; // @[Top.scala 722:11]
  assign n29_I_1_0_0 = n22_O_1_0_0; // @[Top.scala 722:11]
  assign n29_I_1_0_1 = n22_O_1_0_1; // @[Top.scala 722:11]
  assign n29_I_1_0_2 = n22_O_1_0_2; // @[Top.scala 722:11]
  assign n29_I_2_0_0 = n22_O_2_0_0; // @[Top.scala 722:11]
  assign n29_I_2_0_1 = n22_O_2_0_1; // @[Top.scala 722:11]
  assign n29_I_2_0_2 = n22_O_2_0_2; // @[Top.scala 722:11]
  assign n29_I_3_0_0 = n22_O_3_0_0; // @[Top.scala 722:11]
  assign n29_I_3_0_1 = n22_O_3_0_1; // @[Top.scala 722:11]
  assign n29_I_3_0_2 = n22_O_3_0_2; // @[Top.scala 722:11]
  assign n29_I_4_0_0 = n22_O_4_0_0; // @[Top.scala 722:11]
  assign n29_I_4_0_1 = n22_O_4_0_1; // @[Top.scala 722:11]
  assign n29_I_4_0_2 = n22_O_4_0_2; // @[Top.scala 722:11]
  assign n29_I_5_0_0 = n22_O_5_0_0; // @[Top.scala 722:11]
  assign n29_I_5_0_1 = n22_O_5_0_1; // @[Top.scala 722:11]
  assign n29_I_5_0_2 = n22_O_5_0_2; // @[Top.scala 722:11]
  assign n29_I_6_0_0 = n22_O_6_0_0; // @[Top.scala 722:11]
  assign n29_I_6_0_1 = n22_O_6_0_1; // @[Top.scala 722:11]
  assign n29_I_6_0_2 = n22_O_6_0_2; // @[Top.scala 722:11]
  assign n29_I_7_0_0 = n22_O_7_0_0; // @[Top.scala 722:11]
  assign n29_I_7_0_1 = n22_O_7_0_1; // @[Top.scala 722:11]
  assign n29_I_7_0_2 = n22_O_7_0_2; // @[Top.scala 722:11]
  assign n30_clock = clock;
  assign n30_valid_up = n2_valid_down; // @[Top.scala 726:18]
  assign n30_I_0 = n2_O_0; // @[Top.scala 725:11]
  assign n30_I_1 = n2_O_1; // @[Top.scala 725:11]
  assign n30_I_2 = n2_O_2; // @[Top.scala 725:11]
  assign n30_I_3 = n2_O_3; // @[Top.scala 725:11]
  assign n30_I_4 = n2_O_4; // @[Top.scala 725:11]
  assign n30_I_5 = n2_O_5; // @[Top.scala 725:11]
  assign n30_I_6 = n2_O_6; // @[Top.scala 725:11]
  assign n30_I_7 = n2_O_7; // @[Top.scala 725:11]
  assign n31_clock = clock;
  assign n31_valid_up = n30_valid_down; // @[Top.scala 729:18]
  assign n31_I_0 = n30_O_0; // @[Top.scala 728:11]
  assign n31_I_1 = n30_O_1; // @[Top.scala 728:11]
  assign n31_I_2 = n30_O_2; // @[Top.scala 728:11]
  assign n31_I_3 = n30_O_3; // @[Top.scala 728:11]
  assign n31_I_4 = n30_O_4; // @[Top.scala 728:11]
  assign n31_I_5 = n30_O_5; // @[Top.scala 728:11]
  assign n31_I_6 = n30_O_6; // @[Top.scala 728:11]
  assign n31_I_7 = n30_O_7; // @[Top.scala 728:11]
  assign n32_valid_up = n31_valid_down & n30_valid_down; // @[Top.scala 733:18]
  assign n32_I0_0 = n31_O_0; // @[Top.scala 731:12]
  assign n32_I0_1 = n31_O_1; // @[Top.scala 731:12]
  assign n32_I0_2 = n31_O_2; // @[Top.scala 731:12]
  assign n32_I0_3 = n31_O_3; // @[Top.scala 731:12]
  assign n32_I0_4 = n31_O_4; // @[Top.scala 731:12]
  assign n32_I0_5 = n31_O_5; // @[Top.scala 731:12]
  assign n32_I0_6 = n31_O_6; // @[Top.scala 731:12]
  assign n32_I0_7 = n31_O_7; // @[Top.scala 731:12]
  assign n32_I1_0 = n30_O_0; // @[Top.scala 732:12]
  assign n32_I1_1 = n30_O_1; // @[Top.scala 732:12]
  assign n32_I1_2 = n30_O_2; // @[Top.scala 732:12]
  assign n32_I1_3 = n30_O_3; // @[Top.scala 732:12]
  assign n32_I1_4 = n30_O_4; // @[Top.scala 732:12]
  assign n32_I1_5 = n30_O_5; // @[Top.scala 732:12]
  assign n32_I1_6 = n30_O_6; // @[Top.scala 732:12]
  assign n32_I1_7 = n30_O_7; // @[Top.scala 732:12]
  assign n39_valid_up = n32_valid_down & n2_valid_down; // @[Top.scala 737:18]
  assign n39_I0_0_0 = n32_O_0_0; // @[Top.scala 735:12]
  assign n39_I0_0_1 = n32_O_0_1; // @[Top.scala 735:12]
  assign n39_I0_1_0 = n32_O_1_0; // @[Top.scala 735:12]
  assign n39_I0_1_1 = n32_O_1_1; // @[Top.scala 735:12]
  assign n39_I0_2_0 = n32_O_2_0; // @[Top.scala 735:12]
  assign n39_I0_2_1 = n32_O_2_1; // @[Top.scala 735:12]
  assign n39_I0_3_0 = n32_O_3_0; // @[Top.scala 735:12]
  assign n39_I0_3_1 = n32_O_3_1; // @[Top.scala 735:12]
  assign n39_I0_4_0 = n32_O_4_0; // @[Top.scala 735:12]
  assign n39_I0_4_1 = n32_O_4_1; // @[Top.scala 735:12]
  assign n39_I0_5_0 = n32_O_5_0; // @[Top.scala 735:12]
  assign n39_I0_5_1 = n32_O_5_1; // @[Top.scala 735:12]
  assign n39_I0_6_0 = n32_O_6_0; // @[Top.scala 735:12]
  assign n39_I0_6_1 = n32_O_6_1; // @[Top.scala 735:12]
  assign n39_I0_7_0 = n32_O_7_0; // @[Top.scala 735:12]
  assign n39_I0_7_1 = n32_O_7_1; // @[Top.scala 735:12]
  assign n39_I1_0 = n2_O_0; // @[Top.scala 736:12]
  assign n39_I1_1 = n2_O_1; // @[Top.scala 736:12]
  assign n39_I1_2 = n2_O_2; // @[Top.scala 736:12]
  assign n39_I1_3 = n2_O_3; // @[Top.scala 736:12]
  assign n39_I1_4 = n2_O_4; // @[Top.scala 736:12]
  assign n39_I1_5 = n2_O_5; // @[Top.scala 736:12]
  assign n39_I1_6 = n2_O_6; // @[Top.scala 736:12]
  assign n39_I1_7 = n2_O_7; // @[Top.scala 736:12]
  assign n48_valid_up = n39_valid_down; // @[Top.scala 740:18]
  assign n48_I_0_0 = n39_O_0_0; // @[Top.scala 739:11]
  assign n48_I_0_1 = n39_O_0_1; // @[Top.scala 739:11]
  assign n48_I_0_2 = n39_O_0_2; // @[Top.scala 739:11]
  assign n48_I_1_0 = n39_O_1_0; // @[Top.scala 739:11]
  assign n48_I_1_1 = n39_O_1_1; // @[Top.scala 739:11]
  assign n48_I_1_2 = n39_O_1_2; // @[Top.scala 739:11]
  assign n48_I_2_0 = n39_O_2_0; // @[Top.scala 739:11]
  assign n48_I_2_1 = n39_O_2_1; // @[Top.scala 739:11]
  assign n48_I_2_2 = n39_O_2_2; // @[Top.scala 739:11]
  assign n48_I_3_0 = n39_O_3_0; // @[Top.scala 739:11]
  assign n48_I_3_1 = n39_O_3_1; // @[Top.scala 739:11]
  assign n48_I_3_2 = n39_O_3_2; // @[Top.scala 739:11]
  assign n48_I_4_0 = n39_O_4_0; // @[Top.scala 739:11]
  assign n48_I_4_1 = n39_O_4_1; // @[Top.scala 739:11]
  assign n48_I_4_2 = n39_O_4_2; // @[Top.scala 739:11]
  assign n48_I_5_0 = n39_O_5_0; // @[Top.scala 739:11]
  assign n48_I_5_1 = n39_O_5_1; // @[Top.scala 739:11]
  assign n48_I_5_2 = n39_O_5_2; // @[Top.scala 739:11]
  assign n48_I_6_0 = n39_O_6_0; // @[Top.scala 739:11]
  assign n48_I_6_1 = n39_O_6_1; // @[Top.scala 739:11]
  assign n48_I_6_2 = n39_O_6_2; // @[Top.scala 739:11]
  assign n48_I_7_0 = n39_O_7_0; // @[Top.scala 739:11]
  assign n48_I_7_1 = n39_O_7_1; // @[Top.scala 739:11]
  assign n48_I_7_2 = n39_O_7_2; // @[Top.scala 739:11]
  assign n55_valid_up = n48_valid_down; // @[Top.scala 743:18]
  assign n55_I_0_0_0 = n48_O_0_0_0; // @[Top.scala 742:11]
  assign n55_I_0_0_1 = n48_O_0_0_1; // @[Top.scala 742:11]
  assign n55_I_0_0_2 = n48_O_0_0_2; // @[Top.scala 742:11]
  assign n55_I_1_0_0 = n48_O_1_0_0; // @[Top.scala 742:11]
  assign n55_I_1_0_1 = n48_O_1_0_1; // @[Top.scala 742:11]
  assign n55_I_1_0_2 = n48_O_1_0_2; // @[Top.scala 742:11]
  assign n55_I_2_0_0 = n48_O_2_0_0; // @[Top.scala 742:11]
  assign n55_I_2_0_1 = n48_O_2_0_1; // @[Top.scala 742:11]
  assign n55_I_2_0_2 = n48_O_2_0_2; // @[Top.scala 742:11]
  assign n55_I_3_0_0 = n48_O_3_0_0; // @[Top.scala 742:11]
  assign n55_I_3_0_1 = n48_O_3_0_1; // @[Top.scala 742:11]
  assign n55_I_3_0_2 = n48_O_3_0_2; // @[Top.scala 742:11]
  assign n55_I_4_0_0 = n48_O_4_0_0; // @[Top.scala 742:11]
  assign n55_I_4_0_1 = n48_O_4_0_1; // @[Top.scala 742:11]
  assign n55_I_4_0_2 = n48_O_4_0_2; // @[Top.scala 742:11]
  assign n55_I_5_0_0 = n48_O_5_0_0; // @[Top.scala 742:11]
  assign n55_I_5_0_1 = n48_O_5_0_1; // @[Top.scala 742:11]
  assign n55_I_5_0_2 = n48_O_5_0_2; // @[Top.scala 742:11]
  assign n55_I_6_0_0 = n48_O_6_0_0; // @[Top.scala 742:11]
  assign n55_I_6_0_1 = n48_O_6_0_1; // @[Top.scala 742:11]
  assign n55_I_6_0_2 = n48_O_6_0_2; // @[Top.scala 742:11]
  assign n55_I_7_0_0 = n48_O_7_0_0; // @[Top.scala 742:11]
  assign n55_I_7_0_1 = n48_O_7_0_1; // @[Top.scala 742:11]
  assign n55_I_7_0_2 = n48_O_7_0_2; // @[Top.scala 742:11]
  assign n56_valid_up = n29_valid_down & n55_valid_down; // @[Top.scala 747:18]
  assign n56_I0_0_0 = n29_O_0_0; // @[Top.scala 745:12]
  assign n56_I0_0_1 = n29_O_0_1; // @[Top.scala 745:12]
  assign n56_I0_0_2 = n29_O_0_2; // @[Top.scala 745:12]
  assign n56_I0_1_0 = n29_O_1_0; // @[Top.scala 745:12]
  assign n56_I0_1_1 = n29_O_1_1; // @[Top.scala 745:12]
  assign n56_I0_1_2 = n29_O_1_2; // @[Top.scala 745:12]
  assign n56_I0_2_0 = n29_O_2_0; // @[Top.scala 745:12]
  assign n56_I0_2_1 = n29_O_2_1; // @[Top.scala 745:12]
  assign n56_I0_2_2 = n29_O_2_2; // @[Top.scala 745:12]
  assign n56_I0_3_0 = n29_O_3_0; // @[Top.scala 745:12]
  assign n56_I0_3_1 = n29_O_3_1; // @[Top.scala 745:12]
  assign n56_I0_3_2 = n29_O_3_2; // @[Top.scala 745:12]
  assign n56_I0_4_0 = n29_O_4_0; // @[Top.scala 745:12]
  assign n56_I0_4_1 = n29_O_4_1; // @[Top.scala 745:12]
  assign n56_I0_4_2 = n29_O_4_2; // @[Top.scala 745:12]
  assign n56_I0_5_0 = n29_O_5_0; // @[Top.scala 745:12]
  assign n56_I0_5_1 = n29_O_5_1; // @[Top.scala 745:12]
  assign n56_I0_5_2 = n29_O_5_2; // @[Top.scala 745:12]
  assign n56_I0_6_0 = n29_O_6_0; // @[Top.scala 745:12]
  assign n56_I0_6_1 = n29_O_6_1; // @[Top.scala 745:12]
  assign n56_I0_6_2 = n29_O_6_2; // @[Top.scala 745:12]
  assign n56_I0_7_0 = n29_O_7_0; // @[Top.scala 745:12]
  assign n56_I0_7_1 = n29_O_7_1; // @[Top.scala 745:12]
  assign n56_I0_7_2 = n29_O_7_2; // @[Top.scala 745:12]
  assign n56_I1_0_0 = n55_O_0_0; // @[Top.scala 746:12]
  assign n56_I1_0_1 = n55_O_0_1; // @[Top.scala 746:12]
  assign n56_I1_0_2 = n55_O_0_2; // @[Top.scala 746:12]
  assign n56_I1_1_0 = n55_O_1_0; // @[Top.scala 746:12]
  assign n56_I1_1_1 = n55_O_1_1; // @[Top.scala 746:12]
  assign n56_I1_1_2 = n55_O_1_2; // @[Top.scala 746:12]
  assign n56_I1_2_0 = n55_O_2_0; // @[Top.scala 746:12]
  assign n56_I1_2_1 = n55_O_2_1; // @[Top.scala 746:12]
  assign n56_I1_2_2 = n55_O_2_2; // @[Top.scala 746:12]
  assign n56_I1_3_0 = n55_O_3_0; // @[Top.scala 746:12]
  assign n56_I1_3_1 = n55_O_3_1; // @[Top.scala 746:12]
  assign n56_I1_3_2 = n55_O_3_2; // @[Top.scala 746:12]
  assign n56_I1_4_0 = n55_O_4_0; // @[Top.scala 746:12]
  assign n56_I1_4_1 = n55_O_4_1; // @[Top.scala 746:12]
  assign n56_I1_4_2 = n55_O_4_2; // @[Top.scala 746:12]
  assign n56_I1_5_0 = n55_O_5_0; // @[Top.scala 746:12]
  assign n56_I1_5_1 = n55_O_5_1; // @[Top.scala 746:12]
  assign n56_I1_5_2 = n55_O_5_2; // @[Top.scala 746:12]
  assign n56_I1_6_0 = n55_O_6_0; // @[Top.scala 746:12]
  assign n56_I1_6_1 = n55_O_6_1; // @[Top.scala 746:12]
  assign n56_I1_6_2 = n55_O_6_2; // @[Top.scala 746:12]
  assign n56_I1_7_0 = n55_O_7_0; // @[Top.scala 746:12]
  assign n56_I1_7_1 = n55_O_7_1; // @[Top.scala 746:12]
  assign n56_I1_7_2 = n55_O_7_2; // @[Top.scala 746:12]
  assign n63_clock = clock;
  assign n63_valid_up = n1_valid_down; // @[Top.scala 750:18]
  assign n63_I_0 = n1_O_0; // @[Top.scala 749:11]
  assign n63_I_1 = n1_O_1; // @[Top.scala 749:11]
  assign n63_I_2 = n1_O_2; // @[Top.scala 749:11]
  assign n63_I_3 = n1_O_3; // @[Top.scala 749:11]
  assign n63_I_4 = n1_O_4; // @[Top.scala 749:11]
  assign n63_I_5 = n1_O_5; // @[Top.scala 749:11]
  assign n63_I_6 = n1_O_6; // @[Top.scala 749:11]
  assign n63_I_7 = n1_O_7; // @[Top.scala 749:11]
  assign n64_clock = clock;
  assign n64_valid_up = n63_valid_down; // @[Top.scala 753:18]
  assign n64_I_0 = n63_O_0; // @[Top.scala 752:11]
  assign n64_I_1 = n63_O_1; // @[Top.scala 752:11]
  assign n64_I_2 = n63_O_2; // @[Top.scala 752:11]
  assign n64_I_3 = n63_O_3; // @[Top.scala 752:11]
  assign n64_I_4 = n63_O_4; // @[Top.scala 752:11]
  assign n64_I_5 = n63_O_5; // @[Top.scala 752:11]
  assign n64_I_6 = n63_O_6; // @[Top.scala 752:11]
  assign n64_I_7 = n63_O_7; // @[Top.scala 752:11]
  assign n65_valid_up = n64_valid_down & n63_valid_down; // @[Top.scala 757:18]
  assign n65_I0_0 = n64_O_0; // @[Top.scala 755:12]
  assign n65_I0_1 = n64_O_1; // @[Top.scala 755:12]
  assign n65_I0_2 = n64_O_2; // @[Top.scala 755:12]
  assign n65_I0_3 = n64_O_3; // @[Top.scala 755:12]
  assign n65_I0_4 = n64_O_4; // @[Top.scala 755:12]
  assign n65_I0_5 = n64_O_5; // @[Top.scala 755:12]
  assign n65_I0_6 = n64_O_6; // @[Top.scala 755:12]
  assign n65_I0_7 = n64_O_7; // @[Top.scala 755:12]
  assign n65_I1_0 = n63_O_0; // @[Top.scala 756:12]
  assign n65_I1_1 = n63_O_1; // @[Top.scala 756:12]
  assign n65_I1_2 = n63_O_2; // @[Top.scala 756:12]
  assign n65_I1_3 = n63_O_3; // @[Top.scala 756:12]
  assign n65_I1_4 = n63_O_4; // @[Top.scala 756:12]
  assign n65_I1_5 = n63_O_5; // @[Top.scala 756:12]
  assign n65_I1_6 = n63_O_6; // @[Top.scala 756:12]
  assign n65_I1_7 = n63_O_7; // @[Top.scala 756:12]
  assign n72_valid_up = n65_valid_down & n1_valid_down; // @[Top.scala 761:18]
  assign n72_I0_0_0 = n65_O_0_0; // @[Top.scala 759:12]
  assign n72_I0_0_1 = n65_O_0_1; // @[Top.scala 759:12]
  assign n72_I0_1_0 = n65_O_1_0; // @[Top.scala 759:12]
  assign n72_I0_1_1 = n65_O_1_1; // @[Top.scala 759:12]
  assign n72_I0_2_0 = n65_O_2_0; // @[Top.scala 759:12]
  assign n72_I0_2_1 = n65_O_2_1; // @[Top.scala 759:12]
  assign n72_I0_3_0 = n65_O_3_0; // @[Top.scala 759:12]
  assign n72_I0_3_1 = n65_O_3_1; // @[Top.scala 759:12]
  assign n72_I0_4_0 = n65_O_4_0; // @[Top.scala 759:12]
  assign n72_I0_4_1 = n65_O_4_1; // @[Top.scala 759:12]
  assign n72_I0_5_0 = n65_O_5_0; // @[Top.scala 759:12]
  assign n72_I0_5_1 = n65_O_5_1; // @[Top.scala 759:12]
  assign n72_I0_6_0 = n65_O_6_0; // @[Top.scala 759:12]
  assign n72_I0_6_1 = n65_O_6_1; // @[Top.scala 759:12]
  assign n72_I0_7_0 = n65_O_7_0; // @[Top.scala 759:12]
  assign n72_I0_7_1 = n65_O_7_1; // @[Top.scala 759:12]
  assign n72_I1_0 = n1_O_0; // @[Top.scala 760:12]
  assign n72_I1_1 = n1_O_1; // @[Top.scala 760:12]
  assign n72_I1_2 = n1_O_2; // @[Top.scala 760:12]
  assign n72_I1_3 = n1_O_3; // @[Top.scala 760:12]
  assign n72_I1_4 = n1_O_4; // @[Top.scala 760:12]
  assign n72_I1_5 = n1_O_5; // @[Top.scala 760:12]
  assign n72_I1_6 = n1_O_6; // @[Top.scala 760:12]
  assign n72_I1_7 = n1_O_7; // @[Top.scala 760:12]
  assign n81_valid_up = n72_valid_down; // @[Top.scala 764:18]
  assign n81_I_0_0 = n72_O_0_0; // @[Top.scala 763:11]
  assign n81_I_0_1 = n72_O_0_1; // @[Top.scala 763:11]
  assign n81_I_0_2 = n72_O_0_2; // @[Top.scala 763:11]
  assign n81_I_1_0 = n72_O_1_0; // @[Top.scala 763:11]
  assign n81_I_1_1 = n72_O_1_1; // @[Top.scala 763:11]
  assign n81_I_1_2 = n72_O_1_2; // @[Top.scala 763:11]
  assign n81_I_2_0 = n72_O_2_0; // @[Top.scala 763:11]
  assign n81_I_2_1 = n72_O_2_1; // @[Top.scala 763:11]
  assign n81_I_2_2 = n72_O_2_2; // @[Top.scala 763:11]
  assign n81_I_3_0 = n72_O_3_0; // @[Top.scala 763:11]
  assign n81_I_3_1 = n72_O_3_1; // @[Top.scala 763:11]
  assign n81_I_3_2 = n72_O_3_2; // @[Top.scala 763:11]
  assign n81_I_4_0 = n72_O_4_0; // @[Top.scala 763:11]
  assign n81_I_4_1 = n72_O_4_1; // @[Top.scala 763:11]
  assign n81_I_4_2 = n72_O_4_2; // @[Top.scala 763:11]
  assign n81_I_5_0 = n72_O_5_0; // @[Top.scala 763:11]
  assign n81_I_5_1 = n72_O_5_1; // @[Top.scala 763:11]
  assign n81_I_5_2 = n72_O_5_2; // @[Top.scala 763:11]
  assign n81_I_6_0 = n72_O_6_0; // @[Top.scala 763:11]
  assign n81_I_6_1 = n72_O_6_1; // @[Top.scala 763:11]
  assign n81_I_6_2 = n72_O_6_2; // @[Top.scala 763:11]
  assign n81_I_7_0 = n72_O_7_0; // @[Top.scala 763:11]
  assign n81_I_7_1 = n72_O_7_1; // @[Top.scala 763:11]
  assign n81_I_7_2 = n72_O_7_2; // @[Top.scala 763:11]
  assign n88_valid_up = n81_valid_down; // @[Top.scala 767:18]
  assign n88_I_0_0_0 = n81_O_0_0_0; // @[Top.scala 766:11]
  assign n88_I_0_0_1 = n81_O_0_0_1; // @[Top.scala 766:11]
  assign n88_I_0_0_2 = n81_O_0_0_2; // @[Top.scala 766:11]
  assign n88_I_1_0_0 = n81_O_1_0_0; // @[Top.scala 766:11]
  assign n88_I_1_0_1 = n81_O_1_0_1; // @[Top.scala 766:11]
  assign n88_I_1_0_2 = n81_O_1_0_2; // @[Top.scala 766:11]
  assign n88_I_2_0_0 = n81_O_2_0_0; // @[Top.scala 766:11]
  assign n88_I_2_0_1 = n81_O_2_0_1; // @[Top.scala 766:11]
  assign n88_I_2_0_2 = n81_O_2_0_2; // @[Top.scala 766:11]
  assign n88_I_3_0_0 = n81_O_3_0_0; // @[Top.scala 766:11]
  assign n88_I_3_0_1 = n81_O_3_0_1; // @[Top.scala 766:11]
  assign n88_I_3_0_2 = n81_O_3_0_2; // @[Top.scala 766:11]
  assign n88_I_4_0_0 = n81_O_4_0_0; // @[Top.scala 766:11]
  assign n88_I_4_0_1 = n81_O_4_0_1; // @[Top.scala 766:11]
  assign n88_I_4_0_2 = n81_O_4_0_2; // @[Top.scala 766:11]
  assign n88_I_5_0_0 = n81_O_5_0_0; // @[Top.scala 766:11]
  assign n88_I_5_0_1 = n81_O_5_0_1; // @[Top.scala 766:11]
  assign n88_I_5_0_2 = n81_O_5_0_2; // @[Top.scala 766:11]
  assign n88_I_6_0_0 = n81_O_6_0_0; // @[Top.scala 766:11]
  assign n88_I_6_0_1 = n81_O_6_0_1; // @[Top.scala 766:11]
  assign n88_I_6_0_2 = n81_O_6_0_2; // @[Top.scala 766:11]
  assign n88_I_7_0_0 = n81_O_7_0_0; // @[Top.scala 766:11]
  assign n88_I_7_0_1 = n81_O_7_0_1; // @[Top.scala 766:11]
  assign n88_I_7_0_2 = n81_O_7_0_2; // @[Top.scala 766:11]
  assign n89_valid_up = n56_valid_down & n88_valid_down; // @[Top.scala 771:18]
  assign n89_I0_0_0_0 = n56_O_0_0_0; // @[Top.scala 769:12]
  assign n89_I0_0_0_1 = n56_O_0_0_1; // @[Top.scala 769:12]
  assign n89_I0_0_0_2 = n56_O_0_0_2; // @[Top.scala 769:12]
  assign n89_I0_0_1_0 = n56_O_0_1_0; // @[Top.scala 769:12]
  assign n89_I0_0_1_1 = n56_O_0_1_1; // @[Top.scala 769:12]
  assign n89_I0_0_1_2 = n56_O_0_1_2; // @[Top.scala 769:12]
  assign n89_I0_1_0_0 = n56_O_1_0_0; // @[Top.scala 769:12]
  assign n89_I0_1_0_1 = n56_O_1_0_1; // @[Top.scala 769:12]
  assign n89_I0_1_0_2 = n56_O_1_0_2; // @[Top.scala 769:12]
  assign n89_I0_1_1_0 = n56_O_1_1_0; // @[Top.scala 769:12]
  assign n89_I0_1_1_1 = n56_O_1_1_1; // @[Top.scala 769:12]
  assign n89_I0_1_1_2 = n56_O_1_1_2; // @[Top.scala 769:12]
  assign n89_I0_2_0_0 = n56_O_2_0_0; // @[Top.scala 769:12]
  assign n89_I0_2_0_1 = n56_O_2_0_1; // @[Top.scala 769:12]
  assign n89_I0_2_0_2 = n56_O_2_0_2; // @[Top.scala 769:12]
  assign n89_I0_2_1_0 = n56_O_2_1_0; // @[Top.scala 769:12]
  assign n89_I0_2_1_1 = n56_O_2_1_1; // @[Top.scala 769:12]
  assign n89_I0_2_1_2 = n56_O_2_1_2; // @[Top.scala 769:12]
  assign n89_I0_3_0_0 = n56_O_3_0_0; // @[Top.scala 769:12]
  assign n89_I0_3_0_1 = n56_O_3_0_1; // @[Top.scala 769:12]
  assign n89_I0_3_0_2 = n56_O_3_0_2; // @[Top.scala 769:12]
  assign n89_I0_3_1_0 = n56_O_3_1_0; // @[Top.scala 769:12]
  assign n89_I0_3_1_1 = n56_O_3_1_1; // @[Top.scala 769:12]
  assign n89_I0_3_1_2 = n56_O_3_1_2; // @[Top.scala 769:12]
  assign n89_I0_4_0_0 = n56_O_4_0_0; // @[Top.scala 769:12]
  assign n89_I0_4_0_1 = n56_O_4_0_1; // @[Top.scala 769:12]
  assign n89_I0_4_0_2 = n56_O_4_0_2; // @[Top.scala 769:12]
  assign n89_I0_4_1_0 = n56_O_4_1_0; // @[Top.scala 769:12]
  assign n89_I0_4_1_1 = n56_O_4_1_1; // @[Top.scala 769:12]
  assign n89_I0_4_1_2 = n56_O_4_1_2; // @[Top.scala 769:12]
  assign n89_I0_5_0_0 = n56_O_5_0_0; // @[Top.scala 769:12]
  assign n89_I0_5_0_1 = n56_O_5_0_1; // @[Top.scala 769:12]
  assign n89_I0_5_0_2 = n56_O_5_0_2; // @[Top.scala 769:12]
  assign n89_I0_5_1_0 = n56_O_5_1_0; // @[Top.scala 769:12]
  assign n89_I0_5_1_1 = n56_O_5_1_1; // @[Top.scala 769:12]
  assign n89_I0_5_1_2 = n56_O_5_1_2; // @[Top.scala 769:12]
  assign n89_I0_6_0_0 = n56_O_6_0_0; // @[Top.scala 769:12]
  assign n89_I0_6_0_1 = n56_O_6_0_1; // @[Top.scala 769:12]
  assign n89_I0_6_0_2 = n56_O_6_0_2; // @[Top.scala 769:12]
  assign n89_I0_6_1_0 = n56_O_6_1_0; // @[Top.scala 769:12]
  assign n89_I0_6_1_1 = n56_O_6_1_1; // @[Top.scala 769:12]
  assign n89_I0_6_1_2 = n56_O_6_1_2; // @[Top.scala 769:12]
  assign n89_I0_7_0_0 = n56_O_7_0_0; // @[Top.scala 769:12]
  assign n89_I0_7_0_1 = n56_O_7_0_1; // @[Top.scala 769:12]
  assign n89_I0_7_0_2 = n56_O_7_0_2; // @[Top.scala 769:12]
  assign n89_I0_7_1_0 = n56_O_7_1_0; // @[Top.scala 769:12]
  assign n89_I0_7_1_1 = n56_O_7_1_1; // @[Top.scala 769:12]
  assign n89_I0_7_1_2 = n56_O_7_1_2; // @[Top.scala 769:12]
  assign n89_I1_0_0 = n88_O_0_0; // @[Top.scala 770:12]
  assign n89_I1_0_1 = n88_O_0_1; // @[Top.scala 770:12]
  assign n89_I1_0_2 = n88_O_0_2; // @[Top.scala 770:12]
  assign n89_I1_1_0 = n88_O_1_0; // @[Top.scala 770:12]
  assign n89_I1_1_1 = n88_O_1_1; // @[Top.scala 770:12]
  assign n89_I1_1_2 = n88_O_1_2; // @[Top.scala 770:12]
  assign n89_I1_2_0 = n88_O_2_0; // @[Top.scala 770:12]
  assign n89_I1_2_1 = n88_O_2_1; // @[Top.scala 770:12]
  assign n89_I1_2_2 = n88_O_2_2; // @[Top.scala 770:12]
  assign n89_I1_3_0 = n88_O_3_0; // @[Top.scala 770:12]
  assign n89_I1_3_1 = n88_O_3_1; // @[Top.scala 770:12]
  assign n89_I1_3_2 = n88_O_3_2; // @[Top.scala 770:12]
  assign n89_I1_4_0 = n88_O_4_0; // @[Top.scala 770:12]
  assign n89_I1_4_1 = n88_O_4_1; // @[Top.scala 770:12]
  assign n89_I1_4_2 = n88_O_4_2; // @[Top.scala 770:12]
  assign n89_I1_5_0 = n88_O_5_0; // @[Top.scala 770:12]
  assign n89_I1_5_1 = n88_O_5_1; // @[Top.scala 770:12]
  assign n89_I1_5_2 = n88_O_5_2; // @[Top.scala 770:12]
  assign n89_I1_6_0 = n88_O_6_0; // @[Top.scala 770:12]
  assign n89_I1_6_1 = n88_O_6_1; // @[Top.scala 770:12]
  assign n89_I1_6_2 = n88_O_6_2; // @[Top.scala 770:12]
  assign n89_I1_7_0 = n88_O_7_0; // @[Top.scala 770:12]
  assign n89_I1_7_1 = n88_O_7_1; // @[Top.scala 770:12]
  assign n89_I1_7_2 = n88_O_7_2; // @[Top.scala 770:12]
  assign n98_valid_up = n89_valid_down; // @[Top.scala 774:18]
  assign n98_I_0_0_0 = n89_O_0_0_0; // @[Top.scala 773:11]
  assign n98_I_0_0_1 = n89_O_0_0_1; // @[Top.scala 773:11]
  assign n98_I_0_0_2 = n89_O_0_0_2; // @[Top.scala 773:11]
  assign n98_I_0_1_0 = n89_O_0_1_0; // @[Top.scala 773:11]
  assign n98_I_0_1_1 = n89_O_0_1_1; // @[Top.scala 773:11]
  assign n98_I_0_1_2 = n89_O_0_1_2; // @[Top.scala 773:11]
  assign n98_I_0_2_0 = n89_O_0_2_0; // @[Top.scala 773:11]
  assign n98_I_0_2_1 = n89_O_0_2_1; // @[Top.scala 773:11]
  assign n98_I_0_2_2 = n89_O_0_2_2; // @[Top.scala 773:11]
  assign n98_I_1_0_0 = n89_O_1_0_0; // @[Top.scala 773:11]
  assign n98_I_1_0_1 = n89_O_1_0_1; // @[Top.scala 773:11]
  assign n98_I_1_0_2 = n89_O_1_0_2; // @[Top.scala 773:11]
  assign n98_I_1_1_0 = n89_O_1_1_0; // @[Top.scala 773:11]
  assign n98_I_1_1_1 = n89_O_1_1_1; // @[Top.scala 773:11]
  assign n98_I_1_1_2 = n89_O_1_1_2; // @[Top.scala 773:11]
  assign n98_I_1_2_0 = n89_O_1_2_0; // @[Top.scala 773:11]
  assign n98_I_1_2_1 = n89_O_1_2_1; // @[Top.scala 773:11]
  assign n98_I_1_2_2 = n89_O_1_2_2; // @[Top.scala 773:11]
  assign n98_I_2_0_0 = n89_O_2_0_0; // @[Top.scala 773:11]
  assign n98_I_2_0_1 = n89_O_2_0_1; // @[Top.scala 773:11]
  assign n98_I_2_0_2 = n89_O_2_0_2; // @[Top.scala 773:11]
  assign n98_I_2_1_0 = n89_O_2_1_0; // @[Top.scala 773:11]
  assign n98_I_2_1_1 = n89_O_2_1_1; // @[Top.scala 773:11]
  assign n98_I_2_1_2 = n89_O_2_1_2; // @[Top.scala 773:11]
  assign n98_I_2_2_0 = n89_O_2_2_0; // @[Top.scala 773:11]
  assign n98_I_2_2_1 = n89_O_2_2_1; // @[Top.scala 773:11]
  assign n98_I_2_2_2 = n89_O_2_2_2; // @[Top.scala 773:11]
  assign n98_I_3_0_0 = n89_O_3_0_0; // @[Top.scala 773:11]
  assign n98_I_3_0_1 = n89_O_3_0_1; // @[Top.scala 773:11]
  assign n98_I_3_0_2 = n89_O_3_0_2; // @[Top.scala 773:11]
  assign n98_I_3_1_0 = n89_O_3_1_0; // @[Top.scala 773:11]
  assign n98_I_3_1_1 = n89_O_3_1_1; // @[Top.scala 773:11]
  assign n98_I_3_1_2 = n89_O_3_1_2; // @[Top.scala 773:11]
  assign n98_I_3_2_0 = n89_O_3_2_0; // @[Top.scala 773:11]
  assign n98_I_3_2_1 = n89_O_3_2_1; // @[Top.scala 773:11]
  assign n98_I_3_2_2 = n89_O_3_2_2; // @[Top.scala 773:11]
  assign n98_I_4_0_0 = n89_O_4_0_0; // @[Top.scala 773:11]
  assign n98_I_4_0_1 = n89_O_4_0_1; // @[Top.scala 773:11]
  assign n98_I_4_0_2 = n89_O_4_0_2; // @[Top.scala 773:11]
  assign n98_I_4_1_0 = n89_O_4_1_0; // @[Top.scala 773:11]
  assign n98_I_4_1_1 = n89_O_4_1_1; // @[Top.scala 773:11]
  assign n98_I_4_1_2 = n89_O_4_1_2; // @[Top.scala 773:11]
  assign n98_I_4_2_0 = n89_O_4_2_0; // @[Top.scala 773:11]
  assign n98_I_4_2_1 = n89_O_4_2_1; // @[Top.scala 773:11]
  assign n98_I_4_2_2 = n89_O_4_2_2; // @[Top.scala 773:11]
  assign n98_I_5_0_0 = n89_O_5_0_0; // @[Top.scala 773:11]
  assign n98_I_5_0_1 = n89_O_5_0_1; // @[Top.scala 773:11]
  assign n98_I_5_0_2 = n89_O_5_0_2; // @[Top.scala 773:11]
  assign n98_I_5_1_0 = n89_O_5_1_0; // @[Top.scala 773:11]
  assign n98_I_5_1_1 = n89_O_5_1_1; // @[Top.scala 773:11]
  assign n98_I_5_1_2 = n89_O_5_1_2; // @[Top.scala 773:11]
  assign n98_I_5_2_0 = n89_O_5_2_0; // @[Top.scala 773:11]
  assign n98_I_5_2_1 = n89_O_5_2_1; // @[Top.scala 773:11]
  assign n98_I_5_2_2 = n89_O_5_2_2; // @[Top.scala 773:11]
  assign n98_I_6_0_0 = n89_O_6_0_0; // @[Top.scala 773:11]
  assign n98_I_6_0_1 = n89_O_6_0_1; // @[Top.scala 773:11]
  assign n98_I_6_0_2 = n89_O_6_0_2; // @[Top.scala 773:11]
  assign n98_I_6_1_0 = n89_O_6_1_0; // @[Top.scala 773:11]
  assign n98_I_6_1_1 = n89_O_6_1_1; // @[Top.scala 773:11]
  assign n98_I_6_1_2 = n89_O_6_1_2; // @[Top.scala 773:11]
  assign n98_I_6_2_0 = n89_O_6_2_0; // @[Top.scala 773:11]
  assign n98_I_6_2_1 = n89_O_6_2_1; // @[Top.scala 773:11]
  assign n98_I_6_2_2 = n89_O_6_2_2; // @[Top.scala 773:11]
  assign n98_I_7_0_0 = n89_O_7_0_0; // @[Top.scala 773:11]
  assign n98_I_7_0_1 = n89_O_7_0_1; // @[Top.scala 773:11]
  assign n98_I_7_0_2 = n89_O_7_0_2; // @[Top.scala 773:11]
  assign n98_I_7_1_0 = n89_O_7_1_0; // @[Top.scala 773:11]
  assign n98_I_7_1_1 = n89_O_7_1_1; // @[Top.scala 773:11]
  assign n98_I_7_1_2 = n89_O_7_1_2; // @[Top.scala 773:11]
  assign n98_I_7_2_0 = n89_O_7_2_0; // @[Top.scala 773:11]
  assign n98_I_7_2_1 = n89_O_7_2_1; // @[Top.scala 773:11]
  assign n98_I_7_2_2 = n89_O_7_2_2; // @[Top.scala 773:11]
  assign n105_valid_up = n98_valid_down; // @[Top.scala 777:19]
  assign n105_I_0_0_0_0 = n98_O_0_0_0_0; // @[Top.scala 776:12]
  assign n105_I_0_0_0_1 = n98_O_0_0_0_1; // @[Top.scala 776:12]
  assign n105_I_0_0_0_2 = n98_O_0_0_0_2; // @[Top.scala 776:12]
  assign n105_I_0_0_1_0 = n98_O_0_0_1_0; // @[Top.scala 776:12]
  assign n105_I_0_0_1_1 = n98_O_0_0_1_1; // @[Top.scala 776:12]
  assign n105_I_0_0_1_2 = n98_O_0_0_1_2; // @[Top.scala 776:12]
  assign n105_I_0_0_2_0 = n98_O_0_0_2_0; // @[Top.scala 776:12]
  assign n105_I_0_0_2_1 = n98_O_0_0_2_1; // @[Top.scala 776:12]
  assign n105_I_0_0_2_2 = n98_O_0_0_2_2; // @[Top.scala 776:12]
  assign n105_I_1_0_0_0 = n98_O_1_0_0_0; // @[Top.scala 776:12]
  assign n105_I_1_0_0_1 = n98_O_1_0_0_1; // @[Top.scala 776:12]
  assign n105_I_1_0_0_2 = n98_O_1_0_0_2; // @[Top.scala 776:12]
  assign n105_I_1_0_1_0 = n98_O_1_0_1_0; // @[Top.scala 776:12]
  assign n105_I_1_0_1_1 = n98_O_1_0_1_1; // @[Top.scala 776:12]
  assign n105_I_1_0_1_2 = n98_O_1_0_1_2; // @[Top.scala 776:12]
  assign n105_I_1_0_2_0 = n98_O_1_0_2_0; // @[Top.scala 776:12]
  assign n105_I_1_0_2_1 = n98_O_1_0_2_1; // @[Top.scala 776:12]
  assign n105_I_1_0_2_2 = n98_O_1_0_2_2; // @[Top.scala 776:12]
  assign n105_I_2_0_0_0 = n98_O_2_0_0_0; // @[Top.scala 776:12]
  assign n105_I_2_0_0_1 = n98_O_2_0_0_1; // @[Top.scala 776:12]
  assign n105_I_2_0_0_2 = n98_O_2_0_0_2; // @[Top.scala 776:12]
  assign n105_I_2_0_1_0 = n98_O_2_0_1_0; // @[Top.scala 776:12]
  assign n105_I_2_0_1_1 = n98_O_2_0_1_1; // @[Top.scala 776:12]
  assign n105_I_2_0_1_2 = n98_O_2_0_1_2; // @[Top.scala 776:12]
  assign n105_I_2_0_2_0 = n98_O_2_0_2_0; // @[Top.scala 776:12]
  assign n105_I_2_0_2_1 = n98_O_2_0_2_1; // @[Top.scala 776:12]
  assign n105_I_2_0_2_2 = n98_O_2_0_2_2; // @[Top.scala 776:12]
  assign n105_I_3_0_0_0 = n98_O_3_0_0_0; // @[Top.scala 776:12]
  assign n105_I_3_0_0_1 = n98_O_3_0_0_1; // @[Top.scala 776:12]
  assign n105_I_3_0_0_2 = n98_O_3_0_0_2; // @[Top.scala 776:12]
  assign n105_I_3_0_1_0 = n98_O_3_0_1_0; // @[Top.scala 776:12]
  assign n105_I_3_0_1_1 = n98_O_3_0_1_1; // @[Top.scala 776:12]
  assign n105_I_3_0_1_2 = n98_O_3_0_1_2; // @[Top.scala 776:12]
  assign n105_I_3_0_2_0 = n98_O_3_0_2_0; // @[Top.scala 776:12]
  assign n105_I_3_0_2_1 = n98_O_3_0_2_1; // @[Top.scala 776:12]
  assign n105_I_3_0_2_2 = n98_O_3_0_2_2; // @[Top.scala 776:12]
  assign n105_I_4_0_0_0 = n98_O_4_0_0_0; // @[Top.scala 776:12]
  assign n105_I_4_0_0_1 = n98_O_4_0_0_1; // @[Top.scala 776:12]
  assign n105_I_4_0_0_2 = n98_O_4_0_0_2; // @[Top.scala 776:12]
  assign n105_I_4_0_1_0 = n98_O_4_0_1_0; // @[Top.scala 776:12]
  assign n105_I_4_0_1_1 = n98_O_4_0_1_1; // @[Top.scala 776:12]
  assign n105_I_4_0_1_2 = n98_O_4_0_1_2; // @[Top.scala 776:12]
  assign n105_I_4_0_2_0 = n98_O_4_0_2_0; // @[Top.scala 776:12]
  assign n105_I_4_0_2_1 = n98_O_4_0_2_1; // @[Top.scala 776:12]
  assign n105_I_4_0_2_2 = n98_O_4_0_2_2; // @[Top.scala 776:12]
  assign n105_I_5_0_0_0 = n98_O_5_0_0_0; // @[Top.scala 776:12]
  assign n105_I_5_0_0_1 = n98_O_5_0_0_1; // @[Top.scala 776:12]
  assign n105_I_5_0_0_2 = n98_O_5_0_0_2; // @[Top.scala 776:12]
  assign n105_I_5_0_1_0 = n98_O_5_0_1_0; // @[Top.scala 776:12]
  assign n105_I_5_0_1_1 = n98_O_5_0_1_1; // @[Top.scala 776:12]
  assign n105_I_5_0_1_2 = n98_O_5_0_1_2; // @[Top.scala 776:12]
  assign n105_I_5_0_2_0 = n98_O_5_0_2_0; // @[Top.scala 776:12]
  assign n105_I_5_0_2_1 = n98_O_5_0_2_1; // @[Top.scala 776:12]
  assign n105_I_5_0_2_2 = n98_O_5_0_2_2; // @[Top.scala 776:12]
  assign n105_I_6_0_0_0 = n98_O_6_0_0_0; // @[Top.scala 776:12]
  assign n105_I_6_0_0_1 = n98_O_6_0_0_1; // @[Top.scala 776:12]
  assign n105_I_6_0_0_2 = n98_O_6_0_0_2; // @[Top.scala 776:12]
  assign n105_I_6_0_1_0 = n98_O_6_0_1_0; // @[Top.scala 776:12]
  assign n105_I_6_0_1_1 = n98_O_6_0_1_1; // @[Top.scala 776:12]
  assign n105_I_6_0_1_2 = n98_O_6_0_1_2; // @[Top.scala 776:12]
  assign n105_I_6_0_2_0 = n98_O_6_0_2_0; // @[Top.scala 776:12]
  assign n105_I_6_0_2_1 = n98_O_6_0_2_1; // @[Top.scala 776:12]
  assign n105_I_6_0_2_2 = n98_O_6_0_2_2; // @[Top.scala 776:12]
  assign n105_I_7_0_0_0 = n98_O_7_0_0_0; // @[Top.scala 776:12]
  assign n105_I_7_0_0_1 = n98_O_7_0_0_1; // @[Top.scala 776:12]
  assign n105_I_7_0_0_2 = n98_O_7_0_0_2; // @[Top.scala 776:12]
  assign n105_I_7_0_1_0 = n98_O_7_0_1_0; // @[Top.scala 776:12]
  assign n105_I_7_0_1_1 = n98_O_7_0_1_1; // @[Top.scala 776:12]
  assign n105_I_7_0_1_2 = n98_O_7_0_1_2; // @[Top.scala 776:12]
  assign n105_I_7_0_2_0 = n98_O_7_0_2_0; // @[Top.scala 776:12]
  assign n105_I_7_0_2_1 = n98_O_7_0_2_1; // @[Top.scala 776:12]
  assign n105_I_7_0_2_2 = n98_O_7_0_2_2; // @[Top.scala 776:12]
  assign n106_valid_up = n105_valid_down; // @[Top.scala 780:19]
  assign n106_I_0_0_0 = n105_O_0_0_0; // @[Top.scala 779:12]
  assign n106_I_0_0_1 = n105_O_0_0_1; // @[Top.scala 779:12]
  assign n106_I_0_0_2 = n105_O_0_0_2; // @[Top.scala 779:12]
  assign n106_I_0_1_0 = n105_O_0_1_0; // @[Top.scala 779:12]
  assign n106_I_0_1_1 = n105_O_0_1_1; // @[Top.scala 779:12]
  assign n106_I_0_1_2 = n105_O_0_1_2; // @[Top.scala 779:12]
  assign n106_I_0_2_0 = n105_O_0_2_0; // @[Top.scala 779:12]
  assign n106_I_0_2_1 = n105_O_0_2_1; // @[Top.scala 779:12]
  assign n106_I_0_2_2 = n105_O_0_2_2; // @[Top.scala 779:12]
  assign n106_I_1_0_0 = n105_O_1_0_0; // @[Top.scala 779:12]
  assign n106_I_1_0_1 = n105_O_1_0_1; // @[Top.scala 779:12]
  assign n106_I_1_0_2 = n105_O_1_0_2; // @[Top.scala 779:12]
  assign n106_I_1_1_0 = n105_O_1_1_0; // @[Top.scala 779:12]
  assign n106_I_1_1_1 = n105_O_1_1_1; // @[Top.scala 779:12]
  assign n106_I_1_1_2 = n105_O_1_1_2; // @[Top.scala 779:12]
  assign n106_I_1_2_0 = n105_O_1_2_0; // @[Top.scala 779:12]
  assign n106_I_1_2_1 = n105_O_1_2_1; // @[Top.scala 779:12]
  assign n106_I_1_2_2 = n105_O_1_2_2; // @[Top.scala 779:12]
  assign n106_I_2_0_0 = n105_O_2_0_0; // @[Top.scala 779:12]
  assign n106_I_2_0_1 = n105_O_2_0_1; // @[Top.scala 779:12]
  assign n106_I_2_0_2 = n105_O_2_0_2; // @[Top.scala 779:12]
  assign n106_I_2_1_0 = n105_O_2_1_0; // @[Top.scala 779:12]
  assign n106_I_2_1_1 = n105_O_2_1_1; // @[Top.scala 779:12]
  assign n106_I_2_1_2 = n105_O_2_1_2; // @[Top.scala 779:12]
  assign n106_I_2_2_0 = n105_O_2_2_0; // @[Top.scala 779:12]
  assign n106_I_2_2_1 = n105_O_2_2_1; // @[Top.scala 779:12]
  assign n106_I_2_2_2 = n105_O_2_2_2; // @[Top.scala 779:12]
  assign n106_I_3_0_0 = n105_O_3_0_0; // @[Top.scala 779:12]
  assign n106_I_3_0_1 = n105_O_3_0_1; // @[Top.scala 779:12]
  assign n106_I_3_0_2 = n105_O_3_0_2; // @[Top.scala 779:12]
  assign n106_I_3_1_0 = n105_O_3_1_0; // @[Top.scala 779:12]
  assign n106_I_3_1_1 = n105_O_3_1_1; // @[Top.scala 779:12]
  assign n106_I_3_1_2 = n105_O_3_1_2; // @[Top.scala 779:12]
  assign n106_I_3_2_0 = n105_O_3_2_0; // @[Top.scala 779:12]
  assign n106_I_3_2_1 = n105_O_3_2_1; // @[Top.scala 779:12]
  assign n106_I_3_2_2 = n105_O_3_2_2; // @[Top.scala 779:12]
  assign n106_I_4_0_0 = n105_O_4_0_0; // @[Top.scala 779:12]
  assign n106_I_4_0_1 = n105_O_4_0_1; // @[Top.scala 779:12]
  assign n106_I_4_0_2 = n105_O_4_0_2; // @[Top.scala 779:12]
  assign n106_I_4_1_0 = n105_O_4_1_0; // @[Top.scala 779:12]
  assign n106_I_4_1_1 = n105_O_4_1_1; // @[Top.scala 779:12]
  assign n106_I_4_1_2 = n105_O_4_1_2; // @[Top.scala 779:12]
  assign n106_I_4_2_0 = n105_O_4_2_0; // @[Top.scala 779:12]
  assign n106_I_4_2_1 = n105_O_4_2_1; // @[Top.scala 779:12]
  assign n106_I_4_2_2 = n105_O_4_2_2; // @[Top.scala 779:12]
  assign n106_I_5_0_0 = n105_O_5_0_0; // @[Top.scala 779:12]
  assign n106_I_5_0_1 = n105_O_5_0_1; // @[Top.scala 779:12]
  assign n106_I_5_0_2 = n105_O_5_0_2; // @[Top.scala 779:12]
  assign n106_I_5_1_0 = n105_O_5_1_0; // @[Top.scala 779:12]
  assign n106_I_5_1_1 = n105_O_5_1_1; // @[Top.scala 779:12]
  assign n106_I_5_1_2 = n105_O_5_1_2; // @[Top.scala 779:12]
  assign n106_I_5_2_0 = n105_O_5_2_0; // @[Top.scala 779:12]
  assign n106_I_5_2_1 = n105_O_5_2_1; // @[Top.scala 779:12]
  assign n106_I_5_2_2 = n105_O_5_2_2; // @[Top.scala 779:12]
  assign n106_I_6_0_0 = n105_O_6_0_0; // @[Top.scala 779:12]
  assign n106_I_6_0_1 = n105_O_6_0_1; // @[Top.scala 779:12]
  assign n106_I_6_0_2 = n105_O_6_0_2; // @[Top.scala 779:12]
  assign n106_I_6_1_0 = n105_O_6_1_0; // @[Top.scala 779:12]
  assign n106_I_6_1_1 = n105_O_6_1_1; // @[Top.scala 779:12]
  assign n106_I_6_1_2 = n105_O_6_1_2; // @[Top.scala 779:12]
  assign n106_I_6_2_0 = n105_O_6_2_0; // @[Top.scala 779:12]
  assign n106_I_6_2_1 = n105_O_6_2_1; // @[Top.scala 779:12]
  assign n106_I_6_2_2 = n105_O_6_2_2; // @[Top.scala 779:12]
  assign n106_I_7_0_0 = n105_O_7_0_0; // @[Top.scala 779:12]
  assign n106_I_7_0_1 = n105_O_7_0_1; // @[Top.scala 779:12]
  assign n106_I_7_0_2 = n105_O_7_0_2; // @[Top.scala 779:12]
  assign n106_I_7_1_0 = n105_O_7_1_0; // @[Top.scala 779:12]
  assign n106_I_7_1_1 = n105_O_7_1_1; // @[Top.scala 779:12]
  assign n106_I_7_1_2 = n105_O_7_1_2; // @[Top.scala 779:12]
  assign n106_I_7_2_0 = n105_O_7_2_0; // @[Top.scala 779:12]
  assign n106_I_7_2_1 = n105_O_7_2_1; // @[Top.scala 779:12]
  assign n106_I_7_2_2 = n105_O_7_2_2; // @[Top.scala 779:12]
  assign n443_clock = clock;
  assign n443_reset = reset;
  assign n443_valid_up = n106_valid_down; // @[Top.scala 783:19]
  assign n443_I_0_0_0 = n106_O_0_0_0; // @[Top.scala 782:12]
  assign n443_I_0_0_1 = n106_O_0_0_1; // @[Top.scala 782:12]
  assign n443_I_0_0_2 = n106_O_0_0_2; // @[Top.scala 782:12]
  assign n443_I_0_1_0 = n106_O_0_1_0; // @[Top.scala 782:12]
  assign n443_I_0_1_1 = n106_O_0_1_1; // @[Top.scala 782:12]
  assign n443_I_0_1_2 = n106_O_0_1_2; // @[Top.scala 782:12]
  assign n443_I_0_2_0 = n106_O_0_2_0; // @[Top.scala 782:12]
  assign n443_I_0_2_1 = n106_O_0_2_1; // @[Top.scala 782:12]
  assign n443_I_0_2_2 = n106_O_0_2_2; // @[Top.scala 782:12]
  assign n443_I_1_0_0 = n106_O_1_0_0; // @[Top.scala 782:12]
  assign n443_I_1_0_1 = n106_O_1_0_1; // @[Top.scala 782:12]
  assign n443_I_1_0_2 = n106_O_1_0_2; // @[Top.scala 782:12]
  assign n443_I_1_1_0 = n106_O_1_1_0; // @[Top.scala 782:12]
  assign n443_I_1_1_1 = n106_O_1_1_1; // @[Top.scala 782:12]
  assign n443_I_1_1_2 = n106_O_1_1_2; // @[Top.scala 782:12]
  assign n443_I_1_2_0 = n106_O_1_2_0; // @[Top.scala 782:12]
  assign n443_I_1_2_1 = n106_O_1_2_1; // @[Top.scala 782:12]
  assign n443_I_1_2_2 = n106_O_1_2_2; // @[Top.scala 782:12]
  assign n443_I_2_0_0 = n106_O_2_0_0; // @[Top.scala 782:12]
  assign n443_I_2_0_1 = n106_O_2_0_1; // @[Top.scala 782:12]
  assign n443_I_2_0_2 = n106_O_2_0_2; // @[Top.scala 782:12]
  assign n443_I_2_1_0 = n106_O_2_1_0; // @[Top.scala 782:12]
  assign n443_I_2_1_1 = n106_O_2_1_1; // @[Top.scala 782:12]
  assign n443_I_2_1_2 = n106_O_2_1_2; // @[Top.scala 782:12]
  assign n443_I_2_2_0 = n106_O_2_2_0; // @[Top.scala 782:12]
  assign n443_I_2_2_1 = n106_O_2_2_1; // @[Top.scala 782:12]
  assign n443_I_2_2_2 = n106_O_2_2_2; // @[Top.scala 782:12]
  assign n443_I_3_0_0 = n106_O_3_0_0; // @[Top.scala 782:12]
  assign n443_I_3_0_1 = n106_O_3_0_1; // @[Top.scala 782:12]
  assign n443_I_3_0_2 = n106_O_3_0_2; // @[Top.scala 782:12]
  assign n443_I_3_1_0 = n106_O_3_1_0; // @[Top.scala 782:12]
  assign n443_I_3_1_1 = n106_O_3_1_1; // @[Top.scala 782:12]
  assign n443_I_3_1_2 = n106_O_3_1_2; // @[Top.scala 782:12]
  assign n443_I_3_2_0 = n106_O_3_2_0; // @[Top.scala 782:12]
  assign n443_I_3_2_1 = n106_O_3_2_1; // @[Top.scala 782:12]
  assign n443_I_3_2_2 = n106_O_3_2_2; // @[Top.scala 782:12]
  assign n443_I_4_0_0 = n106_O_4_0_0; // @[Top.scala 782:12]
  assign n443_I_4_0_1 = n106_O_4_0_1; // @[Top.scala 782:12]
  assign n443_I_4_0_2 = n106_O_4_0_2; // @[Top.scala 782:12]
  assign n443_I_4_1_0 = n106_O_4_1_0; // @[Top.scala 782:12]
  assign n443_I_4_1_1 = n106_O_4_1_1; // @[Top.scala 782:12]
  assign n443_I_4_1_2 = n106_O_4_1_2; // @[Top.scala 782:12]
  assign n443_I_4_2_0 = n106_O_4_2_0; // @[Top.scala 782:12]
  assign n443_I_4_2_1 = n106_O_4_2_1; // @[Top.scala 782:12]
  assign n443_I_4_2_2 = n106_O_4_2_2; // @[Top.scala 782:12]
  assign n443_I_5_0_0 = n106_O_5_0_0; // @[Top.scala 782:12]
  assign n443_I_5_0_1 = n106_O_5_0_1; // @[Top.scala 782:12]
  assign n443_I_5_0_2 = n106_O_5_0_2; // @[Top.scala 782:12]
  assign n443_I_5_1_0 = n106_O_5_1_0; // @[Top.scala 782:12]
  assign n443_I_5_1_1 = n106_O_5_1_1; // @[Top.scala 782:12]
  assign n443_I_5_1_2 = n106_O_5_1_2; // @[Top.scala 782:12]
  assign n443_I_5_2_0 = n106_O_5_2_0; // @[Top.scala 782:12]
  assign n443_I_5_2_1 = n106_O_5_2_1; // @[Top.scala 782:12]
  assign n443_I_5_2_2 = n106_O_5_2_2; // @[Top.scala 782:12]
  assign n443_I_6_0_0 = n106_O_6_0_0; // @[Top.scala 782:12]
  assign n443_I_6_0_1 = n106_O_6_0_1; // @[Top.scala 782:12]
  assign n443_I_6_0_2 = n106_O_6_0_2; // @[Top.scala 782:12]
  assign n443_I_6_1_0 = n106_O_6_1_0; // @[Top.scala 782:12]
  assign n443_I_6_1_1 = n106_O_6_1_1; // @[Top.scala 782:12]
  assign n443_I_6_1_2 = n106_O_6_1_2; // @[Top.scala 782:12]
  assign n443_I_6_2_0 = n106_O_6_2_0; // @[Top.scala 782:12]
  assign n443_I_6_2_1 = n106_O_6_2_1; // @[Top.scala 782:12]
  assign n443_I_6_2_2 = n106_O_6_2_2; // @[Top.scala 782:12]
  assign n443_I_7_0_0 = n106_O_7_0_0; // @[Top.scala 782:12]
  assign n443_I_7_0_1 = n106_O_7_0_1; // @[Top.scala 782:12]
  assign n443_I_7_0_2 = n106_O_7_0_2; // @[Top.scala 782:12]
  assign n443_I_7_1_0 = n106_O_7_1_0; // @[Top.scala 782:12]
  assign n443_I_7_1_1 = n106_O_7_1_1; // @[Top.scala 782:12]
  assign n443_I_7_1_2 = n106_O_7_1_2; // @[Top.scala 782:12]
  assign n443_I_7_2_0 = n106_O_7_2_0; // @[Top.scala 782:12]
  assign n443_I_7_2_1 = n106_O_7_2_1; // @[Top.scala 782:12]
  assign n443_I_7_2_2 = n106_O_7_2_2; // @[Top.scala 782:12]
  assign n444_valid_up = n443_valid_down; // @[Top.scala 786:19]
  assign n444_I_0_0_0_t0b = n443_O_0_0_0_t0b; // @[Top.scala 785:12]
  assign n444_I_0_0_0_t1b_t0b = n443_O_0_0_0_t1b_t0b; // @[Top.scala 785:12]
  assign n444_I_0_0_0_t1b_t1b = n443_O_0_0_0_t1b_t1b; // @[Top.scala 785:12]
  assign n444_I_1_0_0_t0b = n443_O_1_0_0_t0b; // @[Top.scala 785:12]
  assign n444_I_1_0_0_t1b_t0b = n443_O_1_0_0_t1b_t0b; // @[Top.scala 785:12]
  assign n444_I_1_0_0_t1b_t1b = n443_O_1_0_0_t1b_t1b; // @[Top.scala 785:12]
  assign n444_I_2_0_0_t0b = n443_O_2_0_0_t0b; // @[Top.scala 785:12]
  assign n444_I_2_0_0_t1b_t0b = n443_O_2_0_0_t1b_t0b; // @[Top.scala 785:12]
  assign n444_I_2_0_0_t1b_t1b = n443_O_2_0_0_t1b_t1b; // @[Top.scala 785:12]
  assign n444_I_3_0_0_t0b = n443_O_3_0_0_t0b; // @[Top.scala 785:12]
  assign n444_I_3_0_0_t1b_t0b = n443_O_3_0_0_t1b_t0b; // @[Top.scala 785:12]
  assign n444_I_3_0_0_t1b_t1b = n443_O_3_0_0_t1b_t1b; // @[Top.scala 785:12]
  assign n444_I_4_0_0_t0b = n443_O_4_0_0_t0b; // @[Top.scala 785:12]
  assign n444_I_4_0_0_t1b_t0b = n443_O_4_0_0_t1b_t0b; // @[Top.scala 785:12]
  assign n444_I_4_0_0_t1b_t1b = n443_O_4_0_0_t1b_t1b; // @[Top.scala 785:12]
  assign n444_I_5_0_0_t0b = n443_O_5_0_0_t0b; // @[Top.scala 785:12]
  assign n444_I_5_0_0_t1b_t0b = n443_O_5_0_0_t1b_t0b; // @[Top.scala 785:12]
  assign n444_I_5_0_0_t1b_t1b = n443_O_5_0_0_t1b_t1b; // @[Top.scala 785:12]
  assign n444_I_6_0_0_t0b = n443_O_6_0_0_t0b; // @[Top.scala 785:12]
  assign n444_I_6_0_0_t1b_t0b = n443_O_6_0_0_t1b_t0b; // @[Top.scala 785:12]
  assign n444_I_6_0_0_t1b_t1b = n443_O_6_0_0_t1b_t1b; // @[Top.scala 785:12]
  assign n444_I_7_0_0_t0b = n443_O_7_0_0_t0b; // @[Top.scala 785:12]
  assign n444_I_7_0_0_t1b_t0b = n443_O_7_0_0_t1b_t0b; // @[Top.scala 785:12]
  assign n444_I_7_0_0_t1b_t1b = n443_O_7_0_0_t1b_t1b; // @[Top.scala 785:12]
  assign n445_valid_up = n444_valid_down; // @[Top.scala 789:19]
  assign n445_I_0_0_0_t0b = n444_O_0_0_0_t0b; // @[Top.scala 788:12]
  assign n445_I_0_0_0_t1b_t0b = n444_O_0_0_0_t1b_t0b; // @[Top.scala 788:12]
  assign n445_I_0_0_0_t1b_t1b = n444_O_0_0_0_t1b_t1b; // @[Top.scala 788:12]
  assign n445_I_1_0_0_t0b = n444_O_1_0_0_t0b; // @[Top.scala 788:12]
  assign n445_I_1_0_0_t1b_t0b = n444_O_1_0_0_t1b_t0b; // @[Top.scala 788:12]
  assign n445_I_1_0_0_t1b_t1b = n444_O_1_0_0_t1b_t1b; // @[Top.scala 788:12]
  assign n445_I_2_0_0_t0b = n444_O_2_0_0_t0b; // @[Top.scala 788:12]
  assign n445_I_2_0_0_t1b_t0b = n444_O_2_0_0_t1b_t0b; // @[Top.scala 788:12]
  assign n445_I_2_0_0_t1b_t1b = n444_O_2_0_0_t1b_t1b; // @[Top.scala 788:12]
  assign n445_I_3_0_0_t0b = n444_O_3_0_0_t0b; // @[Top.scala 788:12]
  assign n445_I_3_0_0_t1b_t0b = n444_O_3_0_0_t1b_t0b; // @[Top.scala 788:12]
  assign n445_I_3_0_0_t1b_t1b = n444_O_3_0_0_t1b_t1b; // @[Top.scala 788:12]
  assign n445_I_4_0_0_t0b = n444_O_4_0_0_t0b; // @[Top.scala 788:12]
  assign n445_I_4_0_0_t1b_t0b = n444_O_4_0_0_t1b_t0b; // @[Top.scala 788:12]
  assign n445_I_4_0_0_t1b_t1b = n444_O_4_0_0_t1b_t1b; // @[Top.scala 788:12]
  assign n445_I_5_0_0_t0b = n444_O_5_0_0_t0b; // @[Top.scala 788:12]
  assign n445_I_5_0_0_t1b_t0b = n444_O_5_0_0_t1b_t0b; // @[Top.scala 788:12]
  assign n445_I_5_0_0_t1b_t1b = n444_O_5_0_0_t1b_t1b; // @[Top.scala 788:12]
  assign n445_I_6_0_0_t0b = n444_O_6_0_0_t0b; // @[Top.scala 788:12]
  assign n445_I_6_0_0_t1b_t0b = n444_O_6_0_0_t1b_t0b; // @[Top.scala 788:12]
  assign n445_I_6_0_0_t1b_t1b = n444_O_6_0_0_t1b_t1b; // @[Top.scala 788:12]
  assign n445_I_7_0_0_t0b = n444_O_7_0_0_t0b; // @[Top.scala 788:12]
  assign n445_I_7_0_0_t1b_t0b = n444_O_7_0_0_t1b_t0b; // @[Top.scala 788:12]
  assign n445_I_7_0_0_t1b_t1b = n444_O_7_0_0_t1b_t1b; // @[Top.scala 788:12]
  assign n446_valid_up = n445_valid_down; // @[Top.scala 792:19]
  assign n446_I_0_0_t0b = n445_O_0_0_t0b; // @[Top.scala 791:12]
  assign n446_I_0_0_t1b_t0b = n445_O_0_0_t1b_t0b; // @[Top.scala 791:12]
  assign n446_I_0_0_t1b_t1b = n445_O_0_0_t1b_t1b; // @[Top.scala 791:12]
  assign n446_I_1_0_t0b = n445_O_1_0_t0b; // @[Top.scala 791:12]
  assign n446_I_1_0_t1b_t0b = n445_O_1_0_t1b_t0b; // @[Top.scala 791:12]
  assign n446_I_1_0_t1b_t1b = n445_O_1_0_t1b_t1b; // @[Top.scala 791:12]
  assign n446_I_2_0_t0b = n445_O_2_0_t0b; // @[Top.scala 791:12]
  assign n446_I_2_0_t1b_t0b = n445_O_2_0_t1b_t0b; // @[Top.scala 791:12]
  assign n446_I_2_0_t1b_t1b = n445_O_2_0_t1b_t1b; // @[Top.scala 791:12]
  assign n446_I_3_0_t0b = n445_O_3_0_t0b; // @[Top.scala 791:12]
  assign n446_I_3_0_t1b_t0b = n445_O_3_0_t1b_t0b; // @[Top.scala 791:12]
  assign n446_I_3_0_t1b_t1b = n445_O_3_0_t1b_t1b; // @[Top.scala 791:12]
  assign n446_I_4_0_t0b = n445_O_4_0_t0b; // @[Top.scala 791:12]
  assign n446_I_4_0_t1b_t0b = n445_O_4_0_t1b_t0b; // @[Top.scala 791:12]
  assign n446_I_4_0_t1b_t1b = n445_O_4_0_t1b_t1b; // @[Top.scala 791:12]
  assign n446_I_5_0_t0b = n445_O_5_0_t0b; // @[Top.scala 791:12]
  assign n446_I_5_0_t1b_t0b = n445_O_5_0_t1b_t0b; // @[Top.scala 791:12]
  assign n446_I_5_0_t1b_t1b = n445_O_5_0_t1b_t1b; // @[Top.scala 791:12]
  assign n446_I_6_0_t0b = n445_O_6_0_t0b; // @[Top.scala 791:12]
  assign n446_I_6_0_t1b_t0b = n445_O_6_0_t1b_t0b; // @[Top.scala 791:12]
  assign n446_I_6_0_t1b_t1b = n445_O_6_0_t1b_t1b; // @[Top.scala 791:12]
  assign n446_I_7_0_t0b = n445_O_7_0_t0b; // @[Top.scala 791:12]
  assign n446_I_7_0_t1b_t0b = n445_O_7_0_t1b_t0b; // @[Top.scala 791:12]
  assign n446_I_7_0_t1b_t1b = n445_O_7_0_t1b_t1b; // @[Top.scala 791:12]
  assign n451_valid_up = n446_valid_down; // @[Top.scala 795:19]
  assign n451_I_0_t0b = n446_O_0_t0b; // @[Top.scala 794:12]
  assign n451_I_1_t0b = n446_O_1_t0b; // @[Top.scala 794:12]
  assign n451_I_2_t0b = n446_O_2_t0b; // @[Top.scala 794:12]
  assign n451_I_3_t0b = n446_O_3_t0b; // @[Top.scala 794:12]
  assign n451_I_4_t0b = n446_O_4_t0b; // @[Top.scala 794:12]
  assign n451_I_5_t0b = n446_O_5_t0b; // @[Top.scala 794:12]
  assign n451_I_6_t0b = n446_O_6_t0b; // @[Top.scala 794:12]
  assign n451_I_7_t0b = n446_O_7_t0b; // @[Top.scala 794:12]
  assign n452_clock = clock;
  assign n452_reset = reset;
  assign n452_valid_up = n451_valid_down; // @[Top.scala 798:19]
  assign n452_I_0 = n451_O_0; // @[Top.scala 797:12]
  assign n452_I_1 = n451_O_1; // @[Top.scala 797:12]
  assign n452_I_2 = n451_O_2; // @[Top.scala 797:12]
  assign n452_I_3 = n451_O_3; // @[Top.scala 797:12]
  assign n452_I_4 = n451_O_4; // @[Top.scala 797:12]
  assign n452_I_5 = n451_O_5; // @[Top.scala 797:12]
  assign n452_I_6 = n451_O_6; // @[Top.scala 797:12]
  assign n452_I_7 = n451_O_7; // @[Top.scala 797:12]
  assign n453_clock = clock;
  assign n453_reset = reset;
  assign n453_valid_up = n452_valid_down; // @[Top.scala 801:19]
  assign n453_I_0 = n452_O_0; // @[Top.scala 800:12]
  assign n453_I_1 = n452_O_1; // @[Top.scala 800:12]
  assign n453_I_2 = n452_O_2; // @[Top.scala 800:12]
  assign n453_I_3 = n452_O_3; // @[Top.scala 800:12]
  assign n453_I_4 = n452_O_4; // @[Top.scala 800:12]
  assign n453_I_5 = n452_O_5; // @[Top.scala 800:12]
  assign n453_I_6 = n452_O_6; // @[Top.scala 800:12]
  assign n453_I_7 = n452_O_7; // @[Top.scala 800:12]
  assign n454_clock = clock;
  assign n454_valid_up = n453_valid_down; // @[Top.scala 804:19]
  assign n454_I_0 = n453_O_0; // @[Top.scala 803:12]
  assign n454_I_1 = n453_O_1; // @[Top.scala 803:12]
  assign n454_I_2 = n453_O_2; // @[Top.scala 803:12]
  assign n454_I_3 = n453_O_3; // @[Top.scala 803:12]
  assign n454_I_4 = n453_O_4; // @[Top.scala 803:12]
  assign n454_I_5 = n453_O_5; // @[Top.scala 803:12]
  assign n454_I_6 = n453_O_6; // @[Top.scala 803:12]
  assign n454_I_7 = n453_O_7; // @[Top.scala 803:12]
  assign n455_clock = clock;
  assign n455_valid_up = n454_valid_down; // @[Top.scala 807:19]
  assign n455_I_0 = n454_O_0; // @[Top.scala 806:12]
  assign n455_I_1 = n454_O_1; // @[Top.scala 806:12]
  assign n455_I_2 = n454_O_2; // @[Top.scala 806:12]
  assign n455_I_3 = n454_O_3; // @[Top.scala 806:12]
  assign n455_I_4 = n454_O_4; // @[Top.scala 806:12]
  assign n455_I_5 = n454_O_5; // @[Top.scala 806:12]
  assign n455_I_6 = n454_O_6; // @[Top.scala 806:12]
  assign n455_I_7 = n454_O_7; // @[Top.scala 806:12]
  assign n456_valid_up = n455_valid_down & n454_valid_down; // @[Top.scala 811:19]
  assign n456_I0_0 = n455_O_0; // @[Top.scala 809:13]
  assign n456_I0_1 = n455_O_1; // @[Top.scala 809:13]
  assign n456_I0_2 = n455_O_2; // @[Top.scala 809:13]
  assign n456_I0_3 = n455_O_3; // @[Top.scala 809:13]
  assign n456_I0_4 = n455_O_4; // @[Top.scala 809:13]
  assign n456_I0_5 = n455_O_5; // @[Top.scala 809:13]
  assign n456_I0_6 = n455_O_6; // @[Top.scala 809:13]
  assign n456_I0_7 = n455_O_7; // @[Top.scala 809:13]
  assign n456_I1_0 = n454_O_0; // @[Top.scala 810:13]
  assign n456_I1_1 = n454_O_1; // @[Top.scala 810:13]
  assign n456_I1_2 = n454_O_2; // @[Top.scala 810:13]
  assign n456_I1_3 = n454_O_3; // @[Top.scala 810:13]
  assign n456_I1_4 = n454_O_4; // @[Top.scala 810:13]
  assign n456_I1_5 = n454_O_5; // @[Top.scala 810:13]
  assign n456_I1_6 = n454_O_6; // @[Top.scala 810:13]
  assign n456_I1_7 = n454_O_7; // @[Top.scala 810:13]
  assign n463_valid_up = n456_valid_down & n453_valid_down; // @[Top.scala 815:19]
  assign n463_I0_0_0 = n456_O_0_0; // @[Top.scala 813:13]
  assign n463_I0_0_1 = n456_O_0_1; // @[Top.scala 813:13]
  assign n463_I0_1_0 = n456_O_1_0; // @[Top.scala 813:13]
  assign n463_I0_1_1 = n456_O_1_1; // @[Top.scala 813:13]
  assign n463_I0_2_0 = n456_O_2_0; // @[Top.scala 813:13]
  assign n463_I0_2_1 = n456_O_2_1; // @[Top.scala 813:13]
  assign n463_I0_3_0 = n456_O_3_0; // @[Top.scala 813:13]
  assign n463_I0_3_1 = n456_O_3_1; // @[Top.scala 813:13]
  assign n463_I0_4_0 = n456_O_4_0; // @[Top.scala 813:13]
  assign n463_I0_4_1 = n456_O_4_1; // @[Top.scala 813:13]
  assign n463_I0_5_0 = n456_O_5_0; // @[Top.scala 813:13]
  assign n463_I0_5_1 = n456_O_5_1; // @[Top.scala 813:13]
  assign n463_I0_6_0 = n456_O_6_0; // @[Top.scala 813:13]
  assign n463_I0_6_1 = n456_O_6_1; // @[Top.scala 813:13]
  assign n463_I0_7_0 = n456_O_7_0; // @[Top.scala 813:13]
  assign n463_I0_7_1 = n456_O_7_1; // @[Top.scala 813:13]
  assign n463_I1_0 = n453_O_0; // @[Top.scala 814:13]
  assign n463_I1_1 = n453_O_1; // @[Top.scala 814:13]
  assign n463_I1_2 = n453_O_2; // @[Top.scala 814:13]
  assign n463_I1_3 = n453_O_3; // @[Top.scala 814:13]
  assign n463_I1_4 = n453_O_4; // @[Top.scala 814:13]
  assign n463_I1_5 = n453_O_5; // @[Top.scala 814:13]
  assign n463_I1_6 = n453_O_6; // @[Top.scala 814:13]
  assign n463_I1_7 = n453_O_7; // @[Top.scala 814:13]
  assign n472_valid_up = n463_valid_down; // @[Top.scala 818:19]
  assign n472_I_0_0 = n463_O_0_0; // @[Top.scala 817:12]
  assign n472_I_0_1 = n463_O_0_1; // @[Top.scala 817:12]
  assign n472_I_0_2 = n463_O_0_2; // @[Top.scala 817:12]
  assign n472_I_1_0 = n463_O_1_0; // @[Top.scala 817:12]
  assign n472_I_1_1 = n463_O_1_1; // @[Top.scala 817:12]
  assign n472_I_1_2 = n463_O_1_2; // @[Top.scala 817:12]
  assign n472_I_2_0 = n463_O_2_0; // @[Top.scala 817:12]
  assign n472_I_2_1 = n463_O_2_1; // @[Top.scala 817:12]
  assign n472_I_2_2 = n463_O_2_2; // @[Top.scala 817:12]
  assign n472_I_3_0 = n463_O_3_0; // @[Top.scala 817:12]
  assign n472_I_3_1 = n463_O_3_1; // @[Top.scala 817:12]
  assign n472_I_3_2 = n463_O_3_2; // @[Top.scala 817:12]
  assign n472_I_4_0 = n463_O_4_0; // @[Top.scala 817:12]
  assign n472_I_4_1 = n463_O_4_1; // @[Top.scala 817:12]
  assign n472_I_4_2 = n463_O_4_2; // @[Top.scala 817:12]
  assign n472_I_5_0 = n463_O_5_0; // @[Top.scala 817:12]
  assign n472_I_5_1 = n463_O_5_1; // @[Top.scala 817:12]
  assign n472_I_5_2 = n463_O_5_2; // @[Top.scala 817:12]
  assign n472_I_6_0 = n463_O_6_0; // @[Top.scala 817:12]
  assign n472_I_6_1 = n463_O_6_1; // @[Top.scala 817:12]
  assign n472_I_6_2 = n463_O_6_2; // @[Top.scala 817:12]
  assign n472_I_7_0 = n463_O_7_0; // @[Top.scala 817:12]
  assign n472_I_7_1 = n463_O_7_1; // @[Top.scala 817:12]
  assign n472_I_7_2 = n463_O_7_2; // @[Top.scala 817:12]
  assign n479_valid_up = n472_valid_down; // @[Top.scala 821:19]
  assign n479_I_0_0_0 = n472_O_0_0_0; // @[Top.scala 820:12]
  assign n479_I_0_0_1 = n472_O_0_0_1; // @[Top.scala 820:12]
  assign n479_I_0_0_2 = n472_O_0_0_2; // @[Top.scala 820:12]
  assign n479_I_1_0_0 = n472_O_1_0_0; // @[Top.scala 820:12]
  assign n479_I_1_0_1 = n472_O_1_0_1; // @[Top.scala 820:12]
  assign n479_I_1_0_2 = n472_O_1_0_2; // @[Top.scala 820:12]
  assign n479_I_2_0_0 = n472_O_2_0_0; // @[Top.scala 820:12]
  assign n479_I_2_0_1 = n472_O_2_0_1; // @[Top.scala 820:12]
  assign n479_I_2_0_2 = n472_O_2_0_2; // @[Top.scala 820:12]
  assign n479_I_3_0_0 = n472_O_3_0_0; // @[Top.scala 820:12]
  assign n479_I_3_0_1 = n472_O_3_0_1; // @[Top.scala 820:12]
  assign n479_I_3_0_2 = n472_O_3_0_2; // @[Top.scala 820:12]
  assign n479_I_4_0_0 = n472_O_4_0_0; // @[Top.scala 820:12]
  assign n479_I_4_0_1 = n472_O_4_0_1; // @[Top.scala 820:12]
  assign n479_I_4_0_2 = n472_O_4_0_2; // @[Top.scala 820:12]
  assign n479_I_5_0_0 = n472_O_5_0_0; // @[Top.scala 820:12]
  assign n479_I_5_0_1 = n472_O_5_0_1; // @[Top.scala 820:12]
  assign n479_I_5_0_2 = n472_O_5_0_2; // @[Top.scala 820:12]
  assign n479_I_6_0_0 = n472_O_6_0_0; // @[Top.scala 820:12]
  assign n479_I_6_0_1 = n472_O_6_0_1; // @[Top.scala 820:12]
  assign n479_I_6_0_2 = n472_O_6_0_2; // @[Top.scala 820:12]
  assign n479_I_7_0_0 = n472_O_7_0_0; // @[Top.scala 820:12]
  assign n479_I_7_0_1 = n472_O_7_0_1; // @[Top.scala 820:12]
  assign n479_I_7_0_2 = n472_O_7_0_2; // @[Top.scala 820:12]
  assign n480_clock = clock;
  assign n480_valid_up = n452_valid_down; // @[Top.scala 824:19]
  assign n480_I_0 = n452_O_0; // @[Top.scala 823:12]
  assign n480_I_1 = n452_O_1; // @[Top.scala 823:12]
  assign n480_I_2 = n452_O_2; // @[Top.scala 823:12]
  assign n480_I_3 = n452_O_3; // @[Top.scala 823:12]
  assign n480_I_4 = n452_O_4; // @[Top.scala 823:12]
  assign n480_I_5 = n452_O_5; // @[Top.scala 823:12]
  assign n480_I_6 = n452_O_6; // @[Top.scala 823:12]
  assign n480_I_7 = n452_O_7; // @[Top.scala 823:12]
  assign n481_clock = clock;
  assign n481_valid_up = n480_valid_down; // @[Top.scala 827:19]
  assign n481_I_0 = n480_O_0; // @[Top.scala 826:12]
  assign n481_I_1 = n480_O_1; // @[Top.scala 826:12]
  assign n481_I_2 = n480_O_2; // @[Top.scala 826:12]
  assign n481_I_3 = n480_O_3; // @[Top.scala 826:12]
  assign n481_I_4 = n480_O_4; // @[Top.scala 826:12]
  assign n481_I_5 = n480_O_5; // @[Top.scala 826:12]
  assign n481_I_6 = n480_O_6; // @[Top.scala 826:12]
  assign n481_I_7 = n480_O_7; // @[Top.scala 826:12]
  assign n482_valid_up = n481_valid_down & n480_valid_down; // @[Top.scala 831:19]
  assign n482_I0_0 = n481_O_0; // @[Top.scala 829:13]
  assign n482_I0_1 = n481_O_1; // @[Top.scala 829:13]
  assign n482_I0_2 = n481_O_2; // @[Top.scala 829:13]
  assign n482_I0_3 = n481_O_3; // @[Top.scala 829:13]
  assign n482_I0_4 = n481_O_4; // @[Top.scala 829:13]
  assign n482_I0_5 = n481_O_5; // @[Top.scala 829:13]
  assign n482_I0_6 = n481_O_6; // @[Top.scala 829:13]
  assign n482_I0_7 = n481_O_7; // @[Top.scala 829:13]
  assign n482_I1_0 = n480_O_0; // @[Top.scala 830:13]
  assign n482_I1_1 = n480_O_1; // @[Top.scala 830:13]
  assign n482_I1_2 = n480_O_2; // @[Top.scala 830:13]
  assign n482_I1_3 = n480_O_3; // @[Top.scala 830:13]
  assign n482_I1_4 = n480_O_4; // @[Top.scala 830:13]
  assign n482_I1_5 = n480_O_5; // @[Top.scala 830:13]
  assign n482_I1_6 = n480_O_6; // @[Top.scala 830:13]
  assign n482_I1_7 = n480_O_7; // @[Top.scala 830:13]
  assign n489_valid_up = n482_valid_down & n452_valid_down; // @[Top.scala 835:19]
  assign n489_I0_0_0 = n482_O_0_0; // @[Top.scala 833:13]
  assign n489_I0_0_1 = n482_O_0_1; // @[Top.scala 833:13]
  assign n489_I0_1_0 = n482_O_1_0; // @[Top.scala 833:13]
  assign n489_I0_1_1 = n482_O_1_1; // @[Top.scala 833:13]
  assign n489_I0_2_0 = n482_O_2_0; // @[Top.scala 833:13]
  assign n489_I0_2_1 = n482_O_2_1; // @[Top.scala 833:13]
  assign n489_I0_3_0 = n482_O_3_0; // @[Top.scala 833:13]
  assign n489_I0_3_1 = n482_O_3_1; // @[Top.scala 833:13]
  assign n489_I0_4_0 = n482_O_4_0; // @[Top.scala 833:13]
  assign n489_I0_4_1 = n482_O_4_1; // @[Top.scala 833:13]
  assign n489_I0_5_0 = n482_O_5_0; // @[Top.scala 833:13]
  assign n489_I0_5_1 = n482_O_5_1; // @[Top.scala 833:13]
  assign n489_I0_6_0 = n482_O_6_0; // @[Top.scala 833:13]
  assign n489_I0_6_1 = n482_O_6_1; // @[Top.scala 833:13]
  assign n489_I0_7_0 = n482_O_7_0; // @[Top.scala 833:13]
  assign n489_I0_7_1 = n482_O_7_1; // @[Top.scala 833:13]
  assign n489_I1_0 = n452_O_0; // @[Top.scala 834:13]
  assign n489_I1_1 = n452_O_1; // @[Top.scala 834:13]
  assign n489_I1_2 = n452_O_2; // @[Top.scala 834:13]
  assign n489_I1_3 = n452_O_3; // @[Top.scala 834:13]
  assign n489_I1_4 = n452_O_4; // @[Top.scala 834:13]
  assign n489_I1_5 = n452_O_5; // @[Top.scala 834:13]
  assign n489_I1_6 = n452_O_6; // @[Top.scala 834:13]
  assign n489_I1_7 = n452_O_7; // @[Top.scala 834:13]
  assign n498_valid_up = n489_valid_down; // @[Top.scala 838:19]
  assign n498_I_0_0 = n489_O_0_0; // @[Top.scala 837:12]
  assign n498_I_0_1 = n489_O_0_1; // @[Top.scala 837:12]
  assign n498_I_0_2 = n489_O_0_2; // @[Top.scala 837:12]
  assign n498_I_1_0 = n489_O_1_0; // @[Top.scala 837:12]
  assign n498_I_1_1 = n489_O_1_1; // @[Top.scala 837:12]
  assign n498_I_1_2 = n489_O_1_2; // @[Top.scala 837:12]
  assign n498_I_2_0 = n489_O_2_0; // @[Top.scala 837:12]
  assign n498_I_2_1 = n489_O_2_1; // @[Top.scala 837:12]
  assign n498_I_2_2 = n489_O_2_2; // @[Top.scala 837:12]
  assign n498_I_3_0 = n489_O_3_0; // @[Top.scala 837:12]
  assign n498_I_3_1 = n489_O_3_1; // @[Top.scala 837:12]
  assign n498_I_3_2 = n489_O_3_2; // @[Top.scala 837:12]
  assign n498_I_4_0 = n489_O_4_0; // @[Top.scala 837:12]
  assign n498_I_4_1 = n489_O_4_1; // @[Top.scala 837:12]
  assign n498_I_4_2 = n489_O_4_2; // @[Top.scala 837:12]
  assign n498_I_5_0 = n489_O_5_0; // @[Top.scala 837:12]
  assign n498_I_5_1 = n489_O_5_1; // @[Top.scala 837:12]
  assign n498_I_5_2 = n489_O_5_2; // @[Top.scala 837:12]
  assign n498_I_6_0 = n489_O_6_0; // @[Top.scala 837:12]
  assign n498_I_6_1 = n489_O_6_1; // @[Top.scala 837:12]
  assign n498_I_6_2 = n489_O_6_2; // @[Top.scala 837:12]
  assign n498_I_7_0 = n489_O_7_0; // @[Top.scala 837:12]
  assign n498_I_7_1 = n489_O_7_1; // @[Top.scala 837:12]
  assign n498_I_7_2 = n489_O_7_2; // @[Top.scala 837:12]
  assign n505_valid_up = n498_valid_down; // @[Top.scala 841:19]
  assign n505_I_0_0_0 = n498_O_0_0_0; // @[Top.scala 840:12]
  assign n505_I_0_0_1 = n498_O_0_0_1; // @[Top.scala 840:12]
  assign n505_I_0_0_2 = n498_O_0_0_2; // @[Top.scala 840:12]
  assign n505_I_1_0_0 = n498_O_1_0_0; // @[Top.scala 840:12]
  assign n505_I_1_0_1 = n498_O_1_0_1; // @[Top.scala 840:12]
  assign n505_I_1_0_2 = n498_O_1_0_2; // @[Top.scala 840:12]
  assign n505_I_2_0_0 = n498_O_2_0_0; // @[Top.scala 840:12]
  assign n505_I_2_0_1 = n498_O_2_0_1; // @[Top.scala 840:12]
  assign n505_I_2_0_2 = n498_O_2_0_2; // @[Top.scala 840:12]
  assign n505_I_3_0_0 = n498_O_3_0_0; // @[Top.scala 840:12]
  assign n505_I_3_0_1 = n498_O_3_0_1; // @[Top.scala 840:12]
  assign n505_I_3_0_2 = n498_O_3_0_2; // @[Top.scala 840:12]
  assign n505_I_4_0_0 = n498_O_4_0_0; // @[Top.scala 840:12]
  assign n505_I_4_0_1 = n498_O_4_0_1; // @[Top.scala 840:12]
  assign n505_I_4_0_2 = n498_O_4_0_2; // @[Top.scala 840:12]
  assign n505_I_5_0_0 = n498_O_5_0_0; // @[Top.scala 840:12]
  assign n505_I_5_0_1 = n498_O_5_0_1; // @[Top.scala 840:12]
  assign n505_I_5_0_2 = n498_O_5_0_2; // @[Top.scala 840:12]
  assign n505_I_6_0_0 = n498_O_6_0_0; // @[Top.scala 840:12]
  assign n505_I_6_0_1 = n498_O_6_0_1; // @[Top.scala 840:12]
  assign n505_I_6_0_2 = n498_O_6_0_2; // @[Top.scala 840:12]
  assign n505_I_7_0_0 = n498_O_7_0_0; // @[Top.scala 840:12]
  assign n505_I_7_0_1 = n498_O_7_0_1; // @[Top.scala 840:12]
  assign n505_I_7_0_2 = n498_O_7_0_2; // @[Top.scala 840:12]
  assign n506_valid_up = n479_valid_down & n505_valid_down; // @[Top.scala 845:19]
  assign n506_I0_0_0 = n479_O_0_0; // @[Top.scala 843:13]
  assign n506_I0_0_1 = n479_O_0_1; // @[Top.scala 843:13]
  assign n506_I0_0_2 = n479_O_0_2; // @[Top.scala 843:13]
  assign n506_I0_1_0 = n479_O_1_0; // @[Top.scala 843:13]
  assign n506_I0_1_1 = n479_O_1_1; // @[Top.scala 843:13]
  assign n506_I0_1_2 = n479_O_1_2; // @[Top.scala 843:13]
  assign n506_I0_2_0 = n479_O_2_0; // @[Top.scala 843:13]
  assign n506_I0_2_1 = n479_O_2_1; // @[Top.scala 843:13]
  assign n506_I0_2_2 = n479_O_2_2; // @[Top.scala 843:13]
  assign n506_I0_3_0 = n479_O_3_0; // @[Top.scala 843:13]
  assign n506_I0_3_1 = n479_O_3_1; // @[Top.scala 843:13]
  assign n506_I0_3_2 = n479_O_3_2; // @[Top.scala 843:13]
  assign n506_I0_4_0 = n479_O_4_0; // @[Top.scala 843:13]
  assign n506_I0_4_1 = n479_O_4_1; // @[Top.scala 843:13]
  assign n506_I0_4_2 = n479_O_4_2; // @[Top.scala 843:13]
  assign n506_I0_5_0 = n479_O_5_0; // @[Top.scala 843:13]
  assign n506_I0_5_1 = n479_O_5_1; // @[Top.scala 843:13]
  assign n506_I0_5_2 = n479_O_5_2; // @[Top.scala 843:13]
  assign n506_I0_6_0 = n479_O_6_0; // @[Top.scala 843:13]
  assign n506_I0_6_1 = n479_O_6_1; // @[Top.scala 843:13]
  assign n506_I0_6_2 = n479_O_6_2; // @[Top.scala 843:13]
  assign n506_I0_7_0 = n479_O_7_0; // @[Top.scala 843:13]
  assign n506_I0_7_1 = n479_O_7_1; // @[Top.scala 843:13]
  assign n506_I0_7_2 = n479_O_7_2; // @[Top.scala 843:13]
  assign n506_I1_0_0 = n505_O_0_0; // @[Top.scala 844:13]
  assign n506_I1_0_1 = n505_O_0_1; // @[Top.scala 844:13]
  assign n506_I1_0_2 = n505_O_0_2; // @[Top.scala 844:13]
  assign n506_I1_1_0 = n505_O_1_0; // @[Top.scala 844:13]
  assign n506_I1_1_1 = n505_O_1_1; // @[Top.scala 844:13]
  assign n506_I1_1_2 = n505_O_1_2; // @[Top.scala 844:13]
  assign n506_I1_2_0 = n505_O_2_0; // @[Top.scala 844:13]
  assign n506_I1_2_1 = n505_O_2_1; // @[Top.scala 844:13]
  assign n506_I1_2_2 = n505_O_2_2; // @[Top.scala 844:13]
  assign n506_I1_3_0 = n505_O_3_0; // @[Top.scala 844:13]
  assign n506_I1_3_1 = n505_O_3_1; // @[Top.scala 844:13]
  assign n506_I1_3_2 = n505_O_3_2; // @[Top.scala 844:13]
  assign n506_I1_4_0 = n505_O_4_0; // @[Top.scala 844:13]
  assign n506_I1_4_1 = n505_O_4_1; // @[Top.scala 844:13]
  assign n506_I1_4_2 = n505_O_4_2; // @[Top.scala 844:13]
  assign n506_I1_5_0 = n505_O_5_0; // @[Top.scala 844:13]
  assign n506_I1_5_1 = n505_O_5_1; // @[Top.scala 844:13]
  assign n506_I1_5_2 = n505_O_5_2; // @[Top.scala 844:13]
  assign n506_I1_6_0 = n505_O_6_0; // @[Top.scala 844:13]
  assign n506_I1_6_1 = n505_O_6_1; // @[Top.scala 844:13]
  assign n506_I1_6_2 = n505_O_6_2; // @[Top.scala 844:13]
  assign n506_I1_7_0 = n505_O_7_0; // @[Top.scala 844:13]
  assign n506_I1_7_1 = n505_O_7_1; // @[Top.scala 844:13]
  assign n506_I1_7_2 = n505_O_7_2; // @[Top.scala 844:13]
  assign n513_clock = clock;
  assign n513_valid_up = n451_valid_down; // @[Top.scala 848:19]
  assign n513_I_0 = n451_O_0; // @[Top.scala 847:12]
  assign n513_I_1 = n451_O_1; // @[Top.scala 847:12]
  assign n513_I_2 = n451_O_2; // @[Top.scala 847:12]
  assign n513_I_3 = n451_O_3; // @[Top.scala 847:12]
  assign n513_I_4 = n451_O_4; // @[Top.scala 847:12]
  assign n513_I_5 = n451_O_5; // @[Top.scala 847:12]
  assign n513_I_6 = n451_O_6; // @[Top.scala 847:12]
  assign n513_I_7 = n451_O_7; // @[Top.scala 847:12]
  assign n514_clock = clock;
  assign n514_valid_up = n513_valid_down; // @[Top.scala 851:19]
  assign n514_I_0 = n513_O_0; // @[Top.scala 850:12]
  assign n514_I_1 = n513_O_1; // @[Top.scala 850:12]
  assign n514_I_2 = n513_O_2; // @[Top.scala 850:12]
  assign n514_I_3 = n513_O_3; // @[Top.scala 850:12]
  assign n514_I_4 = n513_O_4; // @[Top.scala 850:12]
  assign n514_I_5 = n513_O_5; // @[Top.scala 850:12]
  assign n514_I_6 = n513_O_6; // @[Top.scala 850:12]
  assign n514_I_7 = n513_O_7; // @[Top.scala 850:12]
  assign n515_valid_up = n514_valid_down & n513_valid_down; // @[Top.scala 855:19]
  assign n515_I0_0 = n514_O_0; // @[Top.scala 853:13]
  assign n515_I0_1 = n514_O_1; // @[Top.scala 853:13]
  assign n515_I0_2 = n514_O_2; // @[Top.scala 853:13]
  assign n515_I0_3 = n514_O_3; // @[Top.scala 853:13]
  assign n515_I0_4 = n514_O_4; // @[Top.scala 853:13]
  assign n515_I0_5 = n514_O_5; // @[Top.scala 853:13]
  assign n515_I0_6 = n514_O_6; // @[Top.scala 853:13]
  assign n515_I0_7 = n514_O_7; // @[Top.scala 853:13]
  assign n515_I1_0 = n513_O_0; // @[Top.scala 854:13]
  assign n515_I1_1 = n513_O_1; // @[Top.scala 854:13]
  assign n515_I1_2 = n513_O_2; // @[Top.scala 854:13]
  assign n515_I1_3 = n513_O_3; // @[Top.scala 854:13]
  assign n515_I1_4 = n513_O_4; // @[Top.scala 854:13]
  assign n515_I1_5 = n513_O_5; // @[Top.scala 854:13]
  assign n515_I1_6 = n513_O_6; // @[Top.scala 854:13]
  assign n515_I1_7 = n513_O_7; // @[Top.scala 854:13]
  assign n522_valid_up = n515_valid_down & n451_valid_down; // @[Top.scala 859:19]
  assign n522_I0_0_0 = n515_O_0_0; // @[Top.scala 857:13]
  assign n522_I0_0_1 = n515_O_0_1; // @[Top.scala 857:13]
  assign n522_I0_1_0 = n515_O_1_0; // @[Top.scala 857:13]
  assign n522_I0_1_1 = n515_O_1_1; // @[Top.scala 857:13]
  assign n522_I0_2_0 = n515_O_2_0; // @[Top.scala 857:13]
  assign n522_I0_2_1 = n515_O_2_1; // @[Top.scala 857:13]
  assign n522_I0_3_0 = n515_O_3_0; // @[Top.scala 857:13]
  assign n522_I0_3_1 = n515_O_3_1; // @[Top.scala 857:13]
  assign n522_I0_4_0 = n515_O_4_0; // @[Top.scala 857:13]
  assign n522_I0_4_1 = n515_O_4_1; // @[Top.scala 857:13]
  assign n522_I0_5_0 = n515_O_5_0; // @[Top.scala 857:13]
  assign n522_I0_5_1 = n515_O_5_1; // @[Top.scala 857:13]
  assign n522_I0_6_0 = n515_O_6_0; // @[Top.scala 857:13]
  assign n522_I0_6_1 = n515_O_6_1; // @[Top.scala 857:13]
  assign n522_I0_7_0 = n515_O_7_0; // @[Top.scala 857:13]
  assign n522_I0_7_1 = n515_O_7_1; // @[Top.scala 857:13]
  assign n522_I1_0 = n451_O_0; // @[Top.scala 858:13]
  assign n522_I1_1 = n451_O_1; // @[Top.scala 858:13]
  assign n522_I1_2 = n451_O_2; // @[Top.scala 858:13]
  assign n522_I1_3 = n451_O_3; // @[Top.scala 858:13]
  assign n522_I1_4 = n451_O_4; // @[Top.scala 858:13]
  assign n522_I1_5 = n451_O_5; // @[Top.scala 858:13]
  assign n522_I1_6 = n451_O_6; // @[Top.scala 858:13]
  assign n522_I1_7 = n451_O_7; // @[Top.scala 858:13]
  assign n531_valid_up = n522_valid_down; // @[Top.scala 862:19]
  assign n531_I_0_0 = n522_O_0_0; // @[Top.scala 861:12]
  assign n531_I_0_1 = n522_O_0_1; // @[Top.scala 861:12]
  assign n531_I_0_2 = n522_O_0_2; // @[Top.scala 861:12]
  assign n531_I_1_0 = n522_O_1_0; // @[Top.scala 861:12]
  assign n531_I_1_1 = n522_O_1_1; // @[Top.scala 861:12]
  assign n531_I_1_2 = n522_O_1_2; // @[Top.scala 861:12]
  assign n531_I_2_0 = n522_O_2_0; // @[Top.scala 861:12]
  assign n531_I_2_1 = n522_O_2_1; // @[Top.scala 861:12]
  assign n531_I_2_2 = n522_O_2_2; // @[Top.scala 861:12]
  assign n531_I_3_0 = n522_O_3_0; // @[Top.scala 861:12]
  assign n531_I_3_1 = n522_O_3_1; // @[Top.scala 861:12]
  assign n531_I_3_2 = n522_O_3_2; // @[Top.scala 861:12]
  assign n531_I_4_0 = n522_O_4_0; // @[Top.scala 861:12]
  assign n531_I_4_1 = n522_O_4_1; // @[Top.scala 861:12]
  assign n531_I_4_2 = n522_O_4_2; // @[Top.scala 861:12]
  assign n531_I_5_0 = n522_O_5_0; // @[Top.scala 861:12]
  assign n531_I_5_1 = n522_O_5_1; // @[Top.scala 861:12]
  assign n531_I_5_2 = n522_O_5_2; // @[Top.scala 861:12]
  assign n531_I_6_0 = n522_O_6_0; // @[Top.scala 861:12]
  assign n531_I_6_1 = n522_O_6_1; // @[Top.scala 861:12]
  assign n531_I_6_2 = n522_O_6_2; // @[Top.scala 861:12]
  assign n531_I_7_0 = n522_O_7_0; // @[Top.scala 861:12]
  assign n531_I_7_1 = n522_O_7_1; // @[Top.scala 861:12]
  assign n531_I_7_2 = n522_O_7_2; // @[Top.scala 861:12]
  assign n538_valid_up = n531_valid_down; // @[Top.scala 865:19]
  assign n538_I_0_0_0 = n531_O_0_0_0; // @[Top.scala 864:12]
  assign n538_I_0_0_1 = n531_O_0_0_1; // @[Top.scala 864:12]
  assign n538_I_0_0_2 = n531_O_0_0_2; // @[Top.scala 864:12]
  assign n538_I_1_0_0 = n531_O_1_0_0; // @[Top.scala 864:12]
  assign n538_I_1_0_1 = n531_O_1_0_1; // @[Top.scala 864:12]
  assign n538_I_1_0_2 = n531_O_1_0_2; // @[Top.scala 864:12]
  assign n538_I_2_0_0 = n531_O_2_0_0; // @[Top.scala 864:12]
  assign n538_I_2_0_1 = n531_O_2_0_1; // @[Top.scala 864:12]
  assign n538_I_2_0_2 = n531_O_2_0_2; // @[Top.scala 864:12]
  assign n538_I_3_0_0 = n531_O_3_0_0; // @[Top.scala 864:12]
  assign n538_I_3_0_1 = n531_O_3_0_1; // @[Top.scala 864:12]
  assign n538_I_3_0_2 = n531_O_3_0_2; // @[Top.scala 864:12]
  assign n538_I_4_0_0 = n531_O_4_0_0; // @[Top.scala 864:12]
  assign n538_I_4_0_1 = n531_O_4_0_1; // @[Top.scala 864:12]
  assign n538_I_4_0_2 = n531_O_4_0_2; // @[Top.scala 864:12]
  assign n538_I_5_0_0 = n531_O_5_0_0; // @[Top.scala 864:12]
  assign n538_I_5_0_1 = n531_O_5_0_1; // @[Top.scala 864:12]
  assign n538_I_5_0_2 = n531_O_5_0_2; // @[Top.scala 864:12]
  assign n538_I_6_0_0 = n531_O_6_0_0; // @[Top.scala 864:12]
  assign n538_I_6_0_1 = n531_O_6_0_1; // @[Top.scala 864:12]
  assign n538_I_6_0_2 = n531_O_6_0_2; // @[Top.scala 864:12]
  assign n538_I_7_0_0 = n531_O_7_0_0; // @[Top.scala 864:12]
  assign n538_I_7_0_1 = n531_O_7_0_1; // @[Top.scala 864:12]
  assign n538_I_7_0_2 = n531_O_7_0_2; // @[Top.scala 864:12]
  assign n539_valid_up = n506_valid_down & n538_valid_down; // @[Top.scala 869:19]
  assign n539_I0_0_0_0 = n506_O_0_0_0; // @[Top.scala 867:13]
  assign n539_I0_0_0_1 = n506_O_0_0_1; // @[Top.scala 867:13]
  assign n539_I0_0_0_2 = n506_O_0_0_2; // @[Top.scala 867:13]
  assign n539_I0_0_1_0 = n506_O_0_1_0; // @[Top.scala 867:13]
  assign n539_I0_0_1_1 = n506_O_0_1_1; // @[Top.scala 867:13]
  assign n539_I0_0_1_2 = n506_O_0_1_2; // @[Top.scala 867:13]
  assign n539_I0_1_0_0 = n506_O_1_0_0; // @[Top.scala 867:13]
  assign n539_I0_1_0_1 = n506_O_1_0_1; // @[Top.scala 867:13]
  assign n539_I0_1_0_2 = n506_O_1_0_2; // @[Top.scala 867:13]
  assign n539_I0_1_1_0 = n506_O_1_1_0; // @[Top.scala 867:13]
  assign n539_I0_1_1_1 = n506_O_1_1_1; // @[Top.scala 867:13]
  assign n539_I0_1_1_2 = n506_O_1_1_2; // @[Top.scala 867:13]
  assign n539_I0_2_0_0 = n506_O_2_0_0; // @[Top.scala 867:13]
  assign n539_I0_2_0_1 = n506_O_2_0_1; // @[Top.scala 867:13]
  assign n539_I0_2_0_2 = n506_O_2_0_2; // @[Top.scala 867:13]
  assign n539_I0_2_1_0 = n506_O_2_1_0; // @[Top.scala 867:13]
  assign n539_I0_2_1_1 = n506_O_2_1_1; // @[Top.scala 867:13]
  assign n539_I0_2_1_2 = n506_O_2_1_2; // @[Top.scala 867:13]
  assign n539_I0_3_0_0 = n506_O_3_0_0; // @[Top.scala 867:13]
  assign n539_I0_3_0_1 = n506_O_3_0_1; // @[Top.scala 867:13]
  assign n539_I0_3_0_2 = n506_O_3_0_2; // @[Top.scala 867:13]
  assign n539_I0_3_1_0 = n506_O_3_1_0; // @[Top.scala 867:13]
  assign n539_I0_3_1_1 = n506_O_3_1_1; // @[Top.scala 867:13]
  assign n539_I0_3_1_2 = n506_O_3_1_2; // @[Top.scala 867:13]
  assign n539_I0_4_0_0 = n506_O_4_0_0; // @[Top.scala 867:13]
  assign n539_I0_4_0_1 = n506_O_4_0_1; // @[Top.scala 867:13]
  assign n539_I0_4_0_2 = n506_O_4_0_2; // @[Top.scala 867:13]
  assign n539_I0_4_1_0 = n506_O_4_1_0; // @[Top.scala 867:13]
  assign n539_I0_4_1_1 = n506_O_4_1_1; // @[Top.scala 867:13]
  assign n539_I0_4_1_2 = n506_O_4_1_2; // @[Top.scala 867:13]
  assign n539_I0_5_0_0 = n506_O_5_0_0; // @[Top.scala 867:13]
  assign n539_I0_5_0_1 = n506_O_5_0_1; // @[Top.scala 867:13]
  assign n539_I0_5_0_2 = n506_O_5_0_2; // @[Top.scala 867:13]
  assign n539_I0_5_1_0 = n506_O_5_1_0; // @[Top.scala 867:13]
  assign n539_I0_5_1_1 = n506_O_5_1_1; // @[Top.scala 867:13]
  assign n539_I0_5_1_2 = n506_O_5_1_2; // @[Top.scala 867:13]
  assign n539_I0_6_0_0 = n506_O_6_0_0; // @[Top.scala 867:13]
  assign n539_I0_6_0_1 = n506_O_6_0_1; // @[Top.scala 867:13]
  assign n539_I0_6_0_2 = n506_O_6_0_2; // @[Top.scala 867:13]
  assign n539_I0_6_1_0 = n506_O_6_1_0; // @[Top.scala 867:13]
  assign n539_I0_6_1_1 = n506_O_6_1_1; // @[Top.scala 867:13]
  assign n539_I0_6_1_2 = n506_O_6_1_2; // @[Top.scala 867:13]
  assign n539_I0_7_0_0 = n506_O_7_0_0; // @[Top.scala 867:13]
  assign n539_I0_7_0_1 = n506_O_7_0_1; // @[Top.scala 867:13]
  assign n539_I0_7_0_2 = n506_O_7_0_2; // @[Top.scala 867:13]
  assign n539_I0_7_1_0 = n506_O_7_1_0; // @[Top.scala 867:13]
  assign n539_I0_7_1_1 = n506_O_7_1_1; // @[Top.scala 867:13]
  assign n539_I0_7_1_2 = n506_O_7_1_2; // @[Top.scala 867:13]
  assign n539_I1_0_0 = n538_O_0_0; // @[Top.scala 868:13]
  assign n539_I1_0_1 = n538_O_0_1; // @[Top.scala 868:13]
  assign n539_I1_0_2 = n538_O_0_2; // @[Top.scala 868:13]
  assign n539_I1_1_0 = n538_O_1_0; // @[Top.scala 868:13]
  assign n539_I1_1_1 = n538_O_1_1; // @[Top.scala 868:13]
  assign n539_I1_1_2 = n538_O_1_2; // @[Top.scala 868:13]
  assign n539_I1_2_0 = n538_O_2_0; // @[Top.scala 868:13]
  assign n539_I1_2_1 = n538_O_2_1; // @[Top.scala 868:13]
  assign n539_I1_2_2 = n538_O_2_2; // @[Top.scala 868:13]
  assign n539_I1_3_0 = n538_O_3_0; // @[Top.scala 868:13]
  assign n539_I1_3_1 = n538_O_3_1; // @[Top.scala 868:13]
  assign n539_I1_3_2 = n538_O_3_2; // @[Top.scala 868:13]
  assign n539_I1_4_0 = n538_O_4_0; // @[Top.scala 868:13]
  assign n539_I1_4_1 = n538_O_4_1; // @[Top.scala 868:13]
  assign n539_I1_4_2 = n538_O_4_2; // @[Top.scala 868:13]
  assign n539_I1_5_0 = n538_O_5_0; // @[Top.scala 868:13]
  assign n539_I1_5_1 = n538_O_5_1; // @[Top.scala 868:13]
  assign n539_I1_5_2 = n538_O_5_2; // @[Top.scala 868:13]
  assign n539_I1_6_0 = n538_O_6_0; // @[Top.scala 868:13]
  assign n539_I1_6_1 = n538_O_6_1; // @[Top.scala 868:13]
  assign n539_I1_6_2 = n538_O_6_2; // @[Top.scala 868:13]
  assign n539_I1_7_0 = n538_O_7_0; // @[Top.scala 868:13]
  assign n539_I1_7_1 = n538_O_7_1; // @[Top.scala 868:13]
  assign n539_I1_7_2 = n538_O_7_2; // @[Top.scala 868:13]
  assign n548_valid_up = n539_valid_down; // @[Top.scala 872:19]
  assign n548_I_0_0_0 = n539_O_0_0_0; // @[Top.scala 871:12]
  assign n548_I_0_0_1 = n539_O_0_0_1; // @[Top.scala 871:12]
  assign n548_I_0_0_2 = n539_O_0_0_2; // @[Top.scala 871:12]
  assign n548_I_0_1_0 = n539_O_0_1_0; // @[Top.scala 871:12]
  assign n548_I_0_1_1 = n539_O_0_1_1; // @[Top.scala 871:12]
  assign n548_I_0_1_2 = n539_O_0_1_2; // @[Top.scala 871:12]
  assign n548_I_0_2_0 = n539_O_0_2_0; // @[Top.scala 871:12]
  assign n548_I_0_2_1 = n539_O_0_2_1; // @[Top.scala 871:12]
  assign n548_I_0_2_2 = n539_O_0_2_2; // @[Top.scala 871:12]
  assign n548_I_1_0_0 = n539_O_1_0_0; // @[Top.scala 871:12]
  assign n548_I_1_0_1 = n539_O_1_0_1; // @[Top.scala 871:12]
  assign n548_I_1_0_2 = n539_O_1_0_2; // @[Top.scala 871:12]
  assign n548_I_1_1_0 = n539_O_1_1_0; // @[Top.scala 871:12]
  assign n548_I_1_1_1 = n539_O_1_1_1; // @[Top.scala 871:12]
  assign n548_I_1_1_2 = n539_O_1_1_2; // @[Top.scala 871:12]
  assign n548_I_1_2_0 = n539_O_1_2_0; // @[Top.scala 871:12]
  assign n548_I_1_2_1 = n539_O_1_2_1; // @[Top.scala 871:12]
  assign n548_I_1_2_2 = n539_O_1_2_2; // @[Top.scala 871:12]
  assign n548_I_2_0_0 = n539_O_2_0_0; // @[Top.scala 871:12]
  assign n548_I_2_0_1 = n539_O_2_0_1; // @[Top.scala 871:12]
  assign n548_I_2_0_2 = n539_O_2_0_2; // @[Top.scala 871:12]
  assign n548_I_2_1_0 = n539_O_2_1_0; // @[Top.scala 871:12]
  assign n548_I_2_1_1 = n539_O_2_1_1; // @[Top.scala 871:12]
  assign n548_I_2_1_2 = n539_O_2_1_2; // @[Top.scala 871:12]
  assign n548_I_2_2_0 = n539_O_2_2_0; // @[Top.scala 871:12]
  assign n548_I_2_2_1 = n539_O_2_2_1; // @[Top.scala 871:12]
  assign n548_I_2_2_2 = n539_O_2_2_2; // @[Top.scala 871:12]
  assign n548_I_3_0_0 = n539_O_3_0_0; // @[Top.scala 871:12]
  assign n548_I_3_0_1 = n539_O_3_0_1; // @[Top.scala 871:12]
  assign n548_I_3_0_2 = n539_O_3_0_2; // @[Top.scala 871:12]
  assign n548_I_3_1_0 = n539_O_3_1_0; // @[Top.scala 871:12]
  assign n548_I_3_1_1 = n539_O_3_1_1; // @[Top.scala 871:12]
  assign n548_I_3_1_2 = n539_O_3_1_2; // @[Top.scala 871:12]
  assign n548_I_3_2_0 = n539_O_3_2_0; // @[Top.scala 871:12]
  assign n548_I_3_2_1 = n539_O_3_2_1; // @[Top.scala 871:12]
  assign n548_I_3_2_2 = n539_O_3_2_2; // @[Top.scala 871:12]
  assign n548_I_4_0_0 = n539_O_4_0_0; // @[Top.scala 871:12]
  assign n548_I_4_0_1 = n539_O_4_0_1; // @[Top.scala 871:12]
  assign n548_I_4_0_2 = n539_O_4_0_2; // @[Top.scala 871:12]
  assign n548_I_4_1_0 = n539_O_4_1_0; // @[Top.scala 871:12]
  assign n548_I_4_1_1 = n539_O_4_1_1; // @[Top.scala 871:12]
  assign n548_I_4_1_2 = n539_O_4_1_2; // @[Top.scala 871:12]
  assign n548_I_4_2_0 = n539_O_4_2_0; // @[Top.scala 871:12]
  assign n548_I_4_2_1 = n539_O_4_2_1; // @[Top.scala 871:12]
  assign n548_I_4_2_2 = n539_O_4_2_2; // @[Top.scala 871:12]
  assign n548_I_5_0_0 = n539_O_5_0_0; // @[Top.scala 871:12]
  assign n548_I_5_0_1 = n539_O_5_0_1; // @[Top.scala 871:12]
  assign n548_I_5_0_2 = n539_O_5_0_2; // @[Top.scala 871:12]
  assign n548_I_5_1_0 = n539_O_5_1_0; // @[Top.scala 871:12]
  assign n548_I_5_1_1 = n539_O_5_1_1; // @[Top.scala 871:12]
  assign n548_I_5_1_2 = n539_O_5_1_2; // @[Top.scala 871:12]
  assign n548_I_5_2_0 = n539_O_5_2_0; // @[Top.scala 871:12]
  assign n548_I_5_2_1 = n539_O_5_2_1; // @[Top.scala 871:12]
  assign n548_I_5_2_2 = n539_O_5_2_2; // @[Top.scala 871:12]
  assign n548_I_6_0_0 = n539_O_6_0_0; // @[Top.scala 871:12]
  assign n548_I_6_0_1 = n539_O_6_0_1; // @[Top.scala 871:12]
  assign n548_I_6_0_2 = n539_O_6_0_2; // @[Top.scala 871:12]
  assign n548_I_6_1_0 = n539_O_6_1_0; // @[Top.scala 871:12]
  assign n548_I_6_1_1 = n539_O_6_1_1; // @[Top.scala 871:12]
  assign n548_I_6_1_2 = n539_O_6_1_2; // @[Top.scala 871:12]
  assign n548_I_6_2_0 = n539_O_6_2_0; // @[Top.scala 871:12]
  assign n548_I_6_2_1 = n539_O_6_2_1; // @[Top.scala 871:12]
  assign n548_I_6_2_2 = n539_O_6_2_2; // @[Top.scala 871:12]
  assign n548_I_7_0_0 = n539_O_7_0_0; // @[Top.scala 871:12]
  assign n548_I_7_0_1 = n539_O_7_0_1; // @[Top.scala 871:12]
  assign n548_I_7_0_2 = n539_O_7_0_2; // @[Top.scala 871:12]
  assign n548_I_7_1_0 = n539_O_7_1_0; // @[Top.scala 871:12]
  assign n548_I_7_1_1 = n539_O_7_1_1; // @[Top.scala 871:12]
  assign n548_I_7_1_2 = n539_O_7_1_2; // @[Top.scala 871:12]
  assign n548_I_7_2_0 = n539_O_7_2_0; // @[Top.scala 871:12]
  assign n548_I_7_2_1 = n539_O_7_2_1; // @[Top.scala 871:12]
  assign n548_I_7_2_2 = n539_O_7_2_2; // @[Top.scala 871:12]
  assign n555_valid_up = n548_valid_down; // @[Top.scala 875:19]
  assign n555_I_0_0_0_0 = n548_O_0_0_0_0; // @[Top.scala 874:12]
  assign n555_I_0_0_0_1 = n548_O_0_0_0_1; // @[Top.scala 874:12]
  assign n555_I_0_0_0_2 = n548_O_0_0_0_2; // @[Top.scala 874:12]
  assign n555_I_0_0_1_0 = n548_O_0_0_1_0; // @[Top.scala 874:12]
  assign n555_I_0_0_1_1 = n548_O_0_0_1_1; // @[Top.scala 874:12]
  assign n555_I_0_0_1_2 = n548_O_0_0_1_2; // @[Top.scala 874:12]
  assign n555_I_0_0_2_0 = n548_O_0_0_2_0; // @[Top.scala 874:12]
  assign n555_I_0_0_2_1 = n548_O_0_0_2_1; // @[Top.scala 874:12]
  assign n555_I_0_0_2_2 = n548_O_0_0_2_2; // @[Top.scala 874:12]
  assign n555_I_1_0_0_0 = n548_O_1_0_0_0; // @[Top.scala 874:12]
  assign n555_I_1_0_0_1 = n548_O_1_0_0_1; // @[Top.scala 874:12]
  assign n555_I_1_0_0_2 = n548_O_1_0_0_2; // @[Top.scala 874:12]
  assign n555_I_1_0_1_0 = n548_O_1_0_1_0; // @[Top.scala 874:12]
  assign n555_I_1_0_1_1 = n548_O_1_0_1_1; // @[Top.scala 874:12]
  assign n555_I_1_0_1_2 = n548_O_1_0_1_2; // @[Top.scala 874:12]
  assign n555_I_1_0_2_0 = n548_O_1_0_2_0; // @[Top.scala 874:12]
  assign n555_I_1_0_2_1 = n548_O_1_0_2_1; // @[Top.scala 874:12]
  assign n555_I_1_0_2_2 = n548_O_1_0_2_2; // @[Top.scala 874:12]
  assign n555_I_2_0_0_0 = n548_O_2_0_0_0; // @[Top.scala 874:12]
  assign n555_I_2_0_0_1 = n548_O_2_0_0_1; // @[Top.scala 874:12]
  assign n555_I_2_0_0_2 = n548_O_2_0_0_2; // @[Top.scala 874:12]
  assign n555_I_2_0_1_0 = n548_O_2_0_1_0; // @[Top.scala 874:12]
  assign n555_I_2_0_1_1 = n548_O_2_0_1_1; // @[Top.scala 874:12]
  assign n555_I_2_0_1_2 = n548_O_2_0_1_2; // @[Top.scala 874:12]
  assign n555_I_2_0_2_0 = n548_O_2_0_2_0; // @[Top.scala 874:12]
  assign n555_I_2_0_2_1 = n548_O_2_0_2_1; // @[Top.scala 874:12]
  assign n555_I_2_0_2_2 = n548_O_2_0_2_2; // @[Top.scala 874:12]
  assign n555_I_3_0_0_0 = n548_O_3_0_0_0; // @[Top.scala 874:12]
  assign n555_I_3_0_0_1 = n548_O_3_0_0_1; // @[Top.scala 874:12]
  assign n555_I_3_0_0_2 = n548_O_3_0_0_2; // @[Top.scala 874:12]
  assign n555_I_3_0_1_0 = n548_O_3_0_1_0; // @[Top.scala 874:12]
  assign n555_I_3_0_1_1 = n548_O_3_0_1_1; // @[Top.scala 874:12]
  assign n555_I_3_0_1_2 = n548_O_3_0_1_2; // @[Top.scala 874:12]
  assign n555_I_3_0_2_0 = n548_O_3_0_2_0; // @[Top.scala 874:12]
  assign n555_I_3_0_2_1 = n548_O_3_0_2_1; // @[Top.scala 874:12]
  assign n555_I_3_0_2_2 = n548_O_3_0_2_2; // @[Top.scala 874:12]
  assign n555_I_4_0_0_0 = n548_O_4_0_0_0; // @[Top.scala 874:12]
  assign n555_I_4_0_0_1 = n548_O_4_0_0_1; // @[Top.scala 874:12]
  assign n555_I_4_0_0_2 = n548_O_4_0_0_2; // @[Top.scala 874:12]
  assign n555_I_4_0_1_0 = n548_O_4_0_1_0; // @[Top.scala 874:12]
  assign n555_I_4_0_1_1 = n548_O_4_0_1_1; // @[Top.scala 874:12]
  assign n555_I_4_0_1_2 = n548_O_4_0_1_2; // @[Top.scala 874:12]
  assign n555_I_4_0_2_0 = n548_O_4_0_2_0; // @[Top.scala 874:12]
  assign n555_I_4_0_2_1 = n548_O_4_0_2_1; // @[Top.scala 874:12]
  assign n555_I_4_0_2_2 = n548_O_4_0_2_2; // @[Top.scala 874:12]
  assign n555_I_5_0_0_0 = n548_O_5_0_0_0; // @[Top.scala 874:12]
  assign n555_I_5_0_0_1 = n548_O_5_0_0_1; // @[Top.scala 874:12]
  assign n555_I_5_0_0_2 = n548_O_5_0_0_2; // @[Top.scala 874:12]
  assign n555_I_5_0_1_0 = n548_O_5_0_1_0; // @[Top.scala 874:12]
  assign n555_I_5_0_1_1 = n548_O_5_0_1_1; // @[Top.scala 874:12]
  assign n555_I_5_0_1_2 = n548_O_5_0_1_2; // @[Top.scala 874:12]
  assign n555_I_5_0_2_0 = n548_O_5_0_2_0; // @[Top.scala 874:12]
  assign n555_I_5_0_2_1 = n548_O_5_0_2_1; // @[Top.scala 874:12]
  assign n555_I_5_0_2_2 = n548_O_5_0_2_2; // @[Top.scala 874:12]
  assign n555_I_6_0_0_0 = n548_O_6_0_0_0; // @[Top.scala 874:12]
  assign n555_I_6_0_0_1 = n548_O_6_0_0_1; // @[Top.scala 874:12]
  assign n555_I_6_0_0_2 = n548_O_6_0_0_2; // @[Top.scala 874:12]
  assign n555_I_6_0_1_0 = n548_O_6_0_1_0; // @[Top.scala 874:12]
  assign n555_I_6_0_1_1 = n548_O_6_0_1_1; // @[Top.scala 874:12]
  assign n555_I_6_0_1_2 = n548_O_6_0_1_2; // @[Top.scala 874:12]
  assign n555_I_6_0_2_0 = n548_O_6_0_2_0; // @[Top.scala 874:12]
  assign n555_I_6_0_2_1 = n548_O_6_0_2_1; // @[Top.scala 874:12]
  assign n555_I_6_0_2_2 = n548_O_6_0_2_2; // @[Top.scala 874:12]
  assign n555_I_7_0_0_0 = n548_O_7_0_0_0; // @[Top.scala 874:12]
  assign n555_I_7_0_0_1 = n548_O_7_0_0_1; // @[Top.scala 874:12]
  assign n555_I_7_0_0_2 = n548_O_7_0_0_2; // @[Top.scala 874:12]
  assign n555_I_7_0_1_0 = n548_O_7_0_1_0; // @[Top.scala 874:12]
  assign n555_I_7_0_1_1 = n548_O_7_0_1_1; // @[Top.scala 874:12]
  assign n555_I_7_0_1_2 = n548_O_7_0_1_2; // @[Top.scala 874:12]
  assign n555_I_7_0_2_0 = n548_O_7_0_2_0; // @[Top.scala 874:12]
  assign n555_I_7_0_2_1 = n548_O_7_0_2_1; // @[Top.scala 874:12]
  assign n555_I_7_0_2_2 = n548_O_7_0_2_2; // @[Top.scala 874:12]
  assign n597_clock = clock;
  assign n597_reset = reset;
  assign n597_valid_up = n555_valid_down; // @[Top.scala 878:19]
  assign n597_I_0_0_0 = n555_O_0_0_0; // @[Top.scala 877:12]
  assign n597_I_0_0_1 = n555_O_0_0_1; // @[Top.scala 877:12]
  assign n597_I_0_0_2 = n555_O_0_0_2; // @[Top.scala 877:12]
  assign n597_I_0_1_0 = n555_O_0_1_0; // @[Top.scala 877:12]
  assign n597_I_0_1_1 = n555_O_0_1_1; // @[Top.scala 877:12]
  assign n597_I_0_1_2 = n555_O_0_1_2; // @[Top.scala 877:12]
  assign n597_I_0_2_0 = n555_O_0_2_0; // @[Top.scala 877:12]
  assign n597_I_0_2_1 = n555_O_0_2_1; // @[Top.scala 877:12]
  assign n597_I_0_2_2 = n555_O_0_2_2; // @[Top.scala 877:12]
  assign n597_I_1_0_0 = n555_O_1_0_0; // @[Top.scala 877:12]
  assign n597_I_1_0_1 = n555_O_1_0_1; // @[Top.scala 877:12]
  assign n597_I_1_0_2 = n555_O_1_0_2; // @[Top.scala 877:12]
  assign n597_I_1_1_0 = n555_O_1_1_0; // @[Top.scala 877:12]
  assign n597_I_1_1_1 = n555_O_1_1_1; // @[Top.scala 877:12]
  assign n597_I_1_1_2 = n555_O_1_1_2; // @[Top.scala 877:12]
  assign n597_I_1_2_0 = n555_O_1_2_0; // @[Top.scala 877:12]
  assign n597_I_1_2_1 = n555_O_1_2_1; // @[Top.scala 877:12]
  assign n597_I_1_2_2 = n555_O_1_2_2; // @[Top.scala 877:12]
  assign n597_I_2_0_0 = n555_O_2_0_0; // @[Top.scala 877:12]
  assign n597_I_2_0_1 = n555_O_2_0_1; // @[Top.scala 877:12]
  assign n597_I_2_0_2 = n555_O_2_0_2; // @[Top.scala 877:12]
  assign n597_I_2_1_0 = n555_O_2_1_0; // @[Top.scala 877:12]
  assign n597_I_2_1_1 = n555_O_2_1_1; // @[Top.scala 877:12]
  assign n597_I_2_1_2 = n555_O_2_1_2; // @[Top.scala 877:12]
  assign n597_I_2_2_0 = n555_O_2_2_0; // @[Top.scala 877:12]
  assign n597_I_2_2_1 = n555_O_2_2_1; // @[Top.scala 877:12]
  assign n597_I_2_2_2 = n555_O_2_2_2; // @[Top.scala 877:12]
  assign n597_I_3_0_0 = n555_O_3_0_0; // @[Top.scala 877:12]
  assign n597_I_3_0_1 = n555_O_3_0_1; // @[Top.scala 877:12]
  assign n597_I_3_0_2 = n555_O_3_0_2; // @[Top.scala 877:12]
  assign n597_I_3_1_0 = n555_O_3_1_0; // @[Top.scala 877:12]
  assign n597_I_3_1_1 = n555_O_3_1_1; // @[Top.scala 877:12]
  assign n597_I_3_1_2 = n555_O_3_1_2; // @[Top.scala 877:12]
  assign n597_I_3_2_0 = n555_O_3_2_0; // @[Top.scala 877:12]
  assign n597_I_3_2_1 = n555_O_3_2_1; // @[Top.scala 877:12]
  assign n597_I_3_2_2 = n555_O_3_2_2; // @[Top.scala 877:12]
  assign n597_I_4_0_0 = n555_O_4_0_0; // @[Top.scala 877:12]
  assign n597_I_4_0_1 = n555_O_4_0_1; // @[Top.scala 877:12]
  assign n597_I_4_0_2 = n555_O_4_0_2; // @[Top.scala 877:12]
  assign n597_I_4_1_0 = n555_O_4_1_0; // @[Top.scala 877:12]
  assign n597_I_4_1_1 = n555_O_4_1_1; // @[Top.scala 877:12]
  assign n597_I_4_1_2 = n555_O_4_1_2; // @[Top.scala 877:12]
  assign n597_I_4_2_0 = n555_O_4_2_0; // @[Top.scala 877:12]
  assign n597_I_4_2_1 = n555_O_4_2_1; // @[Top.scala 877:12]
  assign n597_I_4_2_2 = n555_O_4_2_2; // @[Top.scala 877:12]
  assign n597_I_5_0_0 = n555_O_5_0_0; // @[Top.scala 877:12]
  assign n597_I_5_0_1 = n555_O_5_0_1; // @[Top.scala 877:12]
  assign n597_I_5_0_2 = n555_O_5_0_2; // @[Top.scala 877:12]
  assign n597_I_5_1_0 = n555_O_5_1_0; // @[Top.scala 877:12]
  assign n597_I_5_1_1 = n555_O_5_1_1; // @[Top.scala 877:12]
  assign n597_I_5_1_2 = n555_O_5_1_2; // @[Top.scala 877:12]
  assign n597_I_5_2_0 = n555_O_5_2_0; // @[Top.scala 877:12]
  assign n597_I_5_2_1 = n555_O_5_2_1; // @[Top.scala 877:12]
  assign n597_I_5_2_2 = n555_O_5_2_2; // @[Top.scala 877:12]
  assign n597_I_6_0_0 = n555_O_6_0_0; // @[Top.scala 877:12]
  assign n597_I_6_0_1 = n555_O_6_0_1; // @[Top.scala 877:12]
  assign n597_I_6_0_2 = n555_O_6_0_2; // @[Top.scala 877:12]
  assign n597_I_6_1_0 = n555_O_6_1_0; // @[Top.scala 877:12]
  assign n597_I_6_1_1 = n555_O_6_1_1; // @[Top.scala 877:12]
  assign n597_I_6_1_2 = n555_O_6_1_2; // @[Top.scala 877:12]
  assign n597_I_6_2_0 = n555_O_6_2_0; // @[Top.scala 877:12]
  assign n597_I_6_2_1 = n555_O_6_2_1; // @[Top.scala 877:12]
  assign n597_I_6_2_2 = n555_O_6_2_2; // @[Top.scala 877:12]
  assign n597_I_7_0_0 = n555_O_7_0_0; // @[Top.scala 877:12]
  assign n597_I_7_0_1 = n555_O_7_0_1; // @[Top.scala 877:12]
  assign n597_I_7_0_2 = n555_O_7_0_2; // @[Top.scala 877:12]
  assign n597_I_7_1_0 = n555_O_7_1_0; // @[Top.scala 877:12]
  assign n597_I_7_1_1 = n555_O_7_1_1; // @[Top.scala 877:12]
  assign n597_I_7_1_2 = n555_O_7_1_2; // @[Top.scala 877:12]
  assign n597_I_7_2_0 = n555_O_7_2_0; // @[Top.scala 877:12]
  assign n597_I_7_2_1 = n555_O_7_2_1; // @[Top.scala 877:12]
  assign n597_I_7_2_2 = n555_O_7_2_2; // @[Top.scala 877:12]
  assign n598_valid_up = n597_valid_down; // @[Top.scala 881:19]
  assign n598_I_0_0_0 = n597_O_0_0_0; // @[Top.scala 880:12]
  assign n598_I_1_0_0 = n597_O_1_0_0; // @[Top.scala 880:12]
  assign n598_I_2_0_0 = n597_O_2_0_0; // @[Top.scala 880:12]
  assign n598_I_3_0_0 = n597_O_3_0_0; // @[Top.scala 880:12]
  assign n598_I_4_0_0 = n597_O_4_0_0; // @[Top.scala 880:12]
  assign n598_I_5_0_0 = n597_O_5_0_0; // @[Top.scala 880:12]
  assign n598_I_6_0_0 = n597_O_6_0_0; // @[Top.scala 880:12]
  assign n598_I_7_0_0 = n597_O_7_0_0; // @[Top.scala 880:12]
  assign n599_valid_up = n598_valid_down; // @[Top.scala 884:19]
  assign n599_I_0_0 = n598_O_0_0; // @[Top.scala 883:12]
  assign n599_I_1_0 = n598_O_1_0; // @[Top.scala 883:12]
  assign n599_I_2_0 = n598_O_2_0; // @[Top.scala 883:12]
  assign n599_I_3_0 = n598_O_3_0; // @[Top.scala 883:12]
  assign n599_I_4_0 = n598_O_4_0; // @[Top.scala 883:12]
  assign n599_I_5_0 = n598_O_5_0; // @[Top.scala 883:12]
  assign n599_I_6_0 = n598_O_6_0; // @[Top.scala 883:12]
  assign n599_I_7_0 = n598_O_7_0; // @[Top.scala 883:12]
  assign n600_clock = clock;
  assign n600_reset = reset;
  assign n600_valid_up = n451_valid_down; // @[Top.scala 887:19]
  assign n600_I_0 = n451_O_0; // @[Top.scala 886:12]
  assign n600_I_1 = n451_O_1; // @[Top.scala 886:12]
  assign n600_I_2 = n451_O_2; // @[Top.scala 886:12]
  assign n600_I_3 = n451_O_3; // @[Top.scala 886:12]
  assign n600_I_4 = n451_O_4; // @[Top.scala 886:12]
  assign n600_I_5 = n451_O_5; // @[Top.scala 886:12]
  assign n600_I_6 = n451_O_6; // @[Top.scala 886:12]
  assign n600_I_7 = n451_O_7; // @[Top.scala 886:12]
  assign n601_clock = clock;
  assign n601_reset = reset;
  assign n601_valid_up = n599_valid_down & n600_valid_down; // @[Top.scala 891:19]
  assign n601_I0_0 = n599_O_0; // @[Top.scala 889:13]
  assign n601_I0_1 = n599_O_1; // @[Top.scala 889:13]
  assign n601_I0_2 = n599_O_2; // @[Top.scala 889:13]
  assign n601_I0_3 = n599_O_3; // @[Top.scala 889:13]
  assign n601_I0_4 = n599_O_4; // @[Top.scala 889:13]
  assign n601_I0_5 = n599_O_5; // @[Top.scala 889:13]
  assign n601_I0_6 = n599_O_6; // @[Top.scala 889:13]
  assign n601_I0_7 = n599_O_7; // @[Top.scala 889:13]
  assign n601_I1_0 = n600_O_0; // @[Top.scala 890:13]
  assign n601_I1_1 = n600_O_1; // @[Top.scala 890:13]
  assign n601_I1_2 = n600_O_2; // @[Top.scala 890:13]
  assign n601_I1_3 = n600_O_3; // @[Top.scala 890:13]
  assign n601_I1_4 = n600_O_4; // @[Top.scala 890:13]
  assign n601_I1_5 = n600_O_5; // @[Top.scala 890:13]
  assign n601_I1_6 = n600_O_6; // @[Top.scala 890:13]
  assign n601_I1_7 = n600_O_7; // @[Top.scala 890:13]
  assign n637_valid_up = n446_valid_down; // @[Top.scala 894:19]
  assign n637_I_0_t1b_t0b = n446_O_0_t1b_t0b; // @[Top.scala 893:12]
  assign n637_I_0_t1b_t1b = n446_O_0_t1b_t1b; // @[Top.scala 893:12]
  assign n637_I_1_t1b_t0b = n446_O_1_t1b_t0b; // @[Top.scala 893:12]
  assign n637_I_1_t1b_t1b = n446_O_1_t1b_t1b; // @[Top.scala 893:12]
  assign n637_I_2_t1b_t0b = n446_O_2_t1b_t0b; // @[Top.scala 893:12]
  assign n637_I_2_t1b_t1b = n446_O_2_t1b_t1b; // @[Top.scala 893:12]
  assign n637_I_3_t1b_t0b = n446_O_3_t1b_t0b; // @[Top.scala 893:12]
  assign n637_I_3_t1b_t1b = n446_O_3_t1b_t1b; // @[Top.scala 893:12]
  assign n637_I_4_t1b_t0b = n446_O_4_t1b_t0b; // @[Top.scala 893:12]
  assign n637_I_4_t1b_t1b = n446_O_4_t1b_t1b; // @[Top.scala 893:12]
  assign n637_I_5_t1b_t0b = n446_O_5_t1b_t0b; // @[Top.scala 893:12]
  assign n637_I_5_t1b_t1b = n446_O_5_t1b_t1b; // @[Top.scala 893:12]
  assign n637_I_6_t1b_t0b = n446_O_6_t1b_t0b; // @[Top.scala 893:12]
  assign n637_I_6_t1b_t1b = n446_O_6_t1b_t1b; // @[Top.scala 893:12]
  assign n637_I_7_t1b_t0b = n446_O_7_t1b_t0b; // @[Top.scala 893:12]
  assign n637_I_7_t1b_t1b = n446_O_7_t1b_t1b; // @[Top.scala 893:12]
  assign n638_clock = clock;
  assign n638_reset = reset;
  assign n638_valid_up = n637_valid_down; // @[Top.scala 897:19]
  assign n638_I_0 = n637_O_0; // @[Top.scala 896:12]
  assign n638_I_1 = n637_O_1; // @[Top.scala 896:12]
  assign n638_I_2 = n637_O_2; // @[Top.scala 896:12]
  assign n638_I_3 = n637_O_3; // @[Top.scala 896:12]
  assign n638_I_4 = n637_O_4; // @[Top.scala 896:12]
  assign n638_I_5 = n637_O_5; // @[Top.scala 896:12]
  assign n638_I_6 = n637_O_6; // @[Top.scala 896:12]
  assign n638_I_7 = n637_O_7; // @[Top.scala 896:12]
  assign n639_clock = clock;
  assign n639_reset = reset;
  assign n639_valid_up = n638_valid_down; // @[Top.scala 900:19]
  assign n639_I_0 = n638_O_0; // @[Top.scala 899:12]
  assign n639_I_1 = n638_O_1; // @[Top.scala 899:12]
  assign n639_I_2 = n638_O_2; // @[Top.scala 899:12]
  assign n639_I_3 = n638_O_3; // @[Top.scala 899:12]
  assign n639_I_4 = n638_O_4; // @[Top.scala 899:12]
  assign n639_I_5 = n638_O_5; // @[Top.scala 899:12]
  assign n639_I_6 = n638_O_6; // @[Top.scala 899:12]
  assign n639_I_7 = n638_O_7; // @[Top.scala 899:12]
  assign n640_clock = clock;
  assign n640_valid_up = n639_valid_down; // @[Top.scala 903:19]
  assign n640_I_0 = n639_O_0; // @[Top.scala 902:12]
  assign n640_I_1 = n639_O_1; // @[Top.scala 902:12]
  assign n640_I_2 = n639_O_2; // @[Top.scala 902:12]
  assign n640_I_3 = n639_O_3; // @[Top.scala 902:12]
  assign n640_I_4 = n639_O_4; // @[Top.scala 902:12]
  assign n640_I_5 = n639_O_5; // @[Top.scala 902:12]
  assign n640_I_6 = n639_O_6; // @[Top.scala 902:12]
  assign n640_I_7 = n639_O_7; // @[Top.scala 902:12]
  assign n641_clock = clock;
  assign n641_valid_up = n640_valid_down; // @[Top.scala 906:19]
  assign n641_I_0 = n640_O_0; // @[Top.scala 905:12]
  assign n641_I_1 = n640_O_1; // @[Top.scala 905:12]
  assign n641_I_2 = n640_O_2; // @[Top.scala 905:12]
  assign n641_I_3 = n640_O_3; // @[Top.scala 905:12]
  assign n641_I_4 = n640_O_4; // @[Top.scala 905:12]
  assign n641_I_5 = n640_O_5; // @[Top.scala 905:12]
  assign n641_I_6 = n640_O_6; // @[Top.scala 905:12]
  assign n641_I_7 = n640_O_7; // @[Top.scala 905:12]
  assign n642_valid_up = n641_valid_down & n640_valid_down; // @[Top.scala 910:19]
  assign n642_I0_0 = n641_O_0; // @[Top.scala 908:13]
  assign n642_I0_1 = n641_O_1; // @[Top.scala 908:13]
  assign n642_I0_2 = n641_O_2; // @[Top.scala 908:13]
  assign n642_I0_3 = n641_O_3; // @[Top.scala 908:13]
  assign n642_I0_4 = n641_O_4; // @[Top.scala 908:13]
  assign n642_I0_5 = n641_O_5; // @[Top.scala 908:13]
  assign n642_I0_6 = n641_O_6; // @[Top.scala 908:13]
  assign n642_I0_7 = n641_O_7; // @[Top.scala 908:13]
  assign n642_I1_0 = n640_O_0; // @[Top.scala 909:13]
  assign n642_I1_1 = n640_O_1; // @[Top.scala 909:13]
  assign n642_I1_2 = n640_O_2; // @[Top.scala 909:13]
  assign n642_I1_3 = n640_O_3; // @[Top.scala 909:13]
  assign n642_I1_4 = n640_O_4; // @[Top.scala 909:13]
  assign n642_I1_5 = n640_O_5; // @[Top.scala 909:13]
  assign n642_I1_6 = n640_O_6; // @[Top.scala 909:13]
  assign n642_I1_7 = n640_O_7; // @[Top.scala 909:13]
  assign n649_valid_up = n642_valid_down & n639_valid_down; // @[Top.scala 914:19]
  assign n649_I0_0_0 = n642_O_0_0; // @[Top.scala 912:13]
  assign n649_I0_0_1 = n642_O_0_1; // @[Top.scala 912:13]
  assign n649_I0_1_0 = n642_O_1_0; // @[Top.scala 912:13]
  assign n649_I0_1_1 = n642_O_1_1; // @[Top.scala 912:13]
  assign n649_I0_2_0 = n642_O_2_0; // @[Top.scala 912:13]
  assign n649_I0_2_1 = n642_O_2_1; // @[Top.scala 912:13]
  assign n649_I0_3_0 = n642_O_3_0; // @[Top.scala 912:13]
  assign n649_I0_3_1 = n642_O_3_1; // @[Top.scala 912:13]
  assign n649_I0_4_0 = n642_O_4_0; // @[Top.scala 912:13]
  assign n649_I0_4_1 = n642_O_4_1; // @[Top.scala 912:13]
  assign n649_I0_5_0 = n642_O_5_0; // @[Top.scala 912:13]
  assign n649_I0_5_1 = n642_O_5_1; // @[Top.scala 912:13]
  assign n649_I0_6_0 = n642_O_6_0; // @[Top.scala 912:13]
  assign n649_I0_6_1 = n642_O_6_1; // @[Top.scala 912:13]
  assign n649_I0_7_0 = n642_O_7_0; // @[Top.scala 912:13]
  assign n649_I0_7_1 = n642_O_7_1; // @[Top.scala 912:13]
  assign n649_I1_0 = n639_O_0; // @[Top.scala 913:13]
  assign n649_I1_1 = n639_O_1; // @[Top.scala 913:13]
  assign n649_I1_2 = n639_O_2; // @[Top.scala 913:13]
  assign n649_I1_3 = n639_O_3; // @[Top.scala 913:13]
  assign n649_I1_4 = n639_O_4; // @[Top.scala 913:13]
  assign n649_I1_5 = n639_O_5; // @[Top.scala 913:13]
  assign n649_I1_6 = n639_O_6; // @[Top.scala 913:13]
  assign n649_I1_7 = n639_O_7; // @[Top.scala 913:13]
  assign n658_valid_up = n649_valid_down; // @[Top.scala 917:19]
  assign n658_I_0_0 = n649_O_0_0; // @[Top.scala 916:12]
  assign n658_I_0_1 = n649_O_0_1; // @[Top.scala 916:12]
  assign n658_I_0_2 = n649_O_0_2; // @[Top.scala 916:12]
  assign n658_I_1_0 = n649_O_1_0; // @[Top.scala 916:12]
  assign n658_I_1_1 = n649_O_1_1; // @[Top.scala 916:12]
  assign n658_I_1_2 = n649_O_1_2; // @[Top.scala 916:12]
  assign n658_I_2_0 = n649_O_2_0; // @[Top.scala 916:12]
  assign n658_I_2_1 = n649_O_2_1; // @[Top.scala 916:12]
  assign n658_I_2_2 = n649_O_2_2; // @[Top.scala 916:12]
  assign n658_I_3_0 = n649_O_3_0; // @[Top.scala 916:12]
  assign n658_I_3_1 = n649_O_3_1; // @[Top.scala 916:12]
  assign n658_I_3_2 = n649_O_3_2; // @[Top.scala 916:12]
  assign n658_I_4_0 = n649_O_4_0; // @[Top.scala 916:12]
  assign n658_I_4_1 = n649_O_4_1; // @[Top.scala 916:12]
  assign n658_I_4_2 = n649_O_4_2; // @[Top.scala 916:12]
  assign n658_I_5_0 = n649_O_5_0; // @[Top.scala 916:12]
  assign n658_I_5_1 = n649_O_5_1; // @[Top.scala 916:12]
  assign n658_I_5_2 = n649_O_5_2; // @[Top.scala 916:12]
  assign n658_I_6_0 = n649_O_6_0; // @[Top.scala 916:12]
  assign n658_I_6_1 = n649_O_6_1; // @[Top.scala 916:12]
  assign n658_I_6_2 = n649_O_6_2; // @[Top.scala 916:12]
  assign n658_I_7_0 = n649_O_7_0; // @[Top.scala 916:12]
  assign n658_I_7_1 = n649_O_7_1; // @[Top.scala 916:12]
  assign n658_I_7_2 = n649_O_7_2; // @[Top.scala 916:12]
  assign n665_valid_up = n658_valid_down; // @[Top.scala 920:19]
  assign n665_I_0_0_0 = n658_O_0_0_0; // @[Top.scala 919:12]
  assign n665_I_0_0_1 = n658_O_0_0_1; // @[Top.scala 919:12]
  assign n665_I_0_0_2 = n658_O_0_0_2; // @[Top.scala 919:12]
  assign n665_I_1_0_0 = n658_O_1_0_0; // @[Top.scala 919:12]
  assign n665_I_1_0_1 = n658_O_1_0_1; // @[Top.scala 919:12]
  assign n665_I_1_0_2 = n658_O_1_0_2; // @[Top.scala 919:12]
  assign n665_I_2_0_0 = n658_O_2_0_0; // @[Top.scala 919:12]
  assign n665_I_2_0_1 = n658_O_2_0_1; // @[Top.scala 919:12]
  assign n665_I_2_0_2 = n658_O_2_0_2; // @[Top.scala 919:12]
  assign n665_I_3_0_0 = n658_O_3_0_0; // @[Top.scala 919:12]
  assign n665_I_3_0_1 = n658_O_3_0_1; // @[Top.scala 919:12]
  assign n665_I_3_0_2 = n658_O_3_0_2; // @[Top.scala 919:12]
  assign n665_I_4_0_0 = n658_O_4_0_0; // @[Top.scala 919:12]
  assign n665_I_4_0_1 = n658_O_4_0_1; // @[Top.scala 919:12]
  assign n665_I_4_0_2 = n658_O_4_0_2; // @[Top.scala 919:12]
  assign n665_I_5_0_0 = n658_O_5_0_0; // @[Top.scala 919:12]
  assign n665_I_5_0_1 = n658_O_5_0_1; // @[Top.scala 919:12]
  assign n665_I_5_0_2 = n658_O_5_0_2; // @[Top.scala 919:12]
  assign n665_I_6_0_0 = n658_O_6_0_0; // @[Top.scala 919:12]
  assign n665_I_6_0_1 = n658_O_6_0_1; // @[Top.scala 919:12]
  assign n665_I_6_0_2 = n658_O_6_0_2; // @[Top.scala 919:12]
  assign n665_I_7_0_0 = n658_O_7_0_0; // @[Top.scala 919:12]
  assign n665_I_7_0_1 = n658_O_7_0_1; // @[Top.scala 919:12]
  assign n665_I_7_0_2 = n658_O_7_0_2; // @[Top.scala 919:12]
  assign n666_clock = clock;
  assign n666_valid_up = n638_valid_down; // @[Top.scala 923:19]
  assign n666_I_0 = n638_O_0; // @[Top.scala 922:12]
  assign n666_I_1 = n638_O_1; // @[Top.scala 922:12]
  assign n666_I_2 = n638_O_2; // @[Top.scala 922:12]
  assign n666_I_3 = n638_O_3; // @[Top.scala 922:12]
  assign n666_I_4 = n638_O_4; // @[Top.scala 922:12]
  assign n666_I_5 = n638_O_5; // @[Top.scala 922:12]
  assign n666_I_6 = n638_O_6; // @[Top.scala 922:12]
  assign n666_I_7 = n638_O_7; // @[Top.scala 922:12]
  assign n667_clock = clock;
  assign n667_valid_up = n666_valid_down; // @[Top.scala 926:19]
  assign n667_I_0 = n666_O_0; // @[Top.scala 925:12]
  assign n667_I_1 = n666_O_1; // @[Top.scala 925:12]
  assign n667_I_2 = n666_O_2; // @[Top.scala 925:12]
  assign n667_I_3 = n666_O_3; // @[Top.scala 925:12]
  assign n667_I_4 = n666_O_4; // @[Top.scala 925:12]
  assign n667_I_5 = n666_O_5; // @[Top.scala 925:12]
  assign n667_I_6 = n666_O_6; // @[Top.scala 925:12]
  assign n667_I_7 = n666_O_7; // @[Top.scala 925:12]
  assign n668_valid_up = n667_valid_down & n666_valid_down; // @[Top.scala 930:19]
  assign n668_I0_0 = n667_O_0; // @[Top.scala 928:13]
  assign n668_I0_1 = n667_O_1; // @[Top.scala 928:13]
  assign n668_I0_2 = n667_O_2; // @[Top.scala 928:13]
  assign n668_I0_3 = n667_O_3; // @[Top.scala 928:13]
  assign n668_I0_4 = n667_O_4; // @[Top.scala 928:13]
  assign n668_I0_5 = n667_O_5; // @[Top.scala 928:13]
  assign n668_I0_6 = n667_O_6; // @[Top.scala 928:13]
  assign n668_I0_7 = n667_O_7; // @[Top.scala 928:13]
  assign n668_I1_0 = n666_O_0; // @[Top.scala 929:13]
  assign n668_I1_1 = n666_O_1; // @[Top.scala 929:13]
  assign n668_I1_2 = n666_O_2; // @[Top.scala 929:13]
  assign n668_I1_3 = n666_O_3; // @[Top.scala 929:13]
  assign n668_I1_4 = n666_O_4; // @[Top.scala 929:13]
  assign n668_I1_5 = n666_O_5; // @[Top.scala 929:13]
  assign n668_I1_6 = n666_O_6; // @[Top.scala 929:13]
  assign n668_I1_7 = n666_O_7; // @[Top.scala 929:13]
  assign n675_valid_up = n668_valid_down & n638_valid_down; // @[Top.scala 934:19]
  assign n675_I0_0_0 = n668_O_0_0; // @[Top.scala 932:13]
  assign n675_I0_0_1 = n668_O_0_1; // @[Top.scala 932:13]
  assign n675_I0_1_0 = n668_O_1_0; // @[Top.scala 932:13]
  assign n675_I0_1_1 = n668_O_1_1; // @[Top.scala 932:13]
  assign n675_I0_2_0 = n668_O_2_0; // @[Top.scala 932:13]
  assign n675_I0_2_1 = n668_O_2_1; // @[Top.scala 932:13]
  assign n675_I0_3_0 = n668_O_3_0; // @[Top.scala 932:13]
  assign n675_I0_3_1 = n668_O_3_1; // @[Top.scala 932:13]
  assign n675_I0_4_0 = n668_O_4_0; // @[Top.scala 932:13]
  assign n675_I0_4_1 = n668_O_4_1; // @[Top.scala 932:13]
  assign n675_I0_5_0 = n668_O_5_0; // @[Top.scala 932:13]
  assign n675_I0_5_1 = n668_O_5_1; // @[Top.scala 932:13]
  assign n675_I0_6_0 = n668_O_6_0; // @[Top.scala 932:13]
  assign n675_I0_6_1 = n668_O_6_1; // @[Top.scala 932:13]
  assign n675_I0_7_0 = n668_O_7_0; // @[Top.scala 932:13]
  assign n675_I0_7_1 = n668_O_7_1; // @[Top.scala 932:13]
  assign n675_I1_0 = n638_O_0; // @[Top.scala 933:13]
  assign n675_I1_1 = n638_O_1; // @[Top.scala 933:13]
  assign n675_I1_2 = n638_O_2; // @[Top.scala 933:13]
  assign n675_I1_3 = n638_O_3; // @[Top.scala 933:13]
  assign n675_I1_4 = n638_O_4; // @[Top.scala 933:13]
  assign n675_I1_5 = n638_O_5; // @[Top.scala 933:13]
  assign n675_I1_6 = n638_O_6; // @[Top.scala 933:13]
  assign n675_I1_7 = n638_O_7; // @[Top.scala 933:13]
  assign n684_valid_up = n675_valid_down; // @[Top.scala 937:19]
  assign n684_I_0_0 = n675_O_0_0; // @[Top.scala 936:12]
  assign n684_I_0_1 = n675_O_0_1; // @[Top.scala 936:12]
  assign n684_I_0_2 = n675_O_0_2; // @[Top.scala 936:12]
  assign n684_I_1_0 = n675_O_1_0; // @[Top.scala 936:12]
  assign n684_I_1_1 = n675_O_1_1; // @[Top.scala 936:12]
  assign n684_I_1_2 = n675_O_1_2; // @[Top.scala 936:12]
  assign n684_I_2_0 = n675_O_2_0; // @[Top.scala 936:12]
  assign n684_I_2_1 = n675_O_2_1; // @[Top.scala 936:12]
  assign n684_I_2_2 = n675_O_2_2; // @[Top.scala 936:12]
  assign n684_I_3_0 = n675_O_3_0; // @[Top.scala 936:12]
  assign n684_I_3_1 = n675_O_3_1; // @[Top.scala 936:12]
  assign n684_I_3_2 = n675_O_3_2; // @[Top.scala 936:12]
  assign n684_I_4_0 = n675_O_4_0; // @[Top.scala 936:12]
  assign n684_I_4_1 = n675_O_4_1; // @[Top.scala 936:12]
  assign n684_I_4_2 = n675_O_4_2; // @[Top.scala 936:12]
  assign n684_I_5_0 = n675_O_5_0; // @[Top.scala 936:12]
  assign n684_I_5_1 = n675_O_5_1; // @[Top.scala 936:12]
  assign n684_I_5_2 = n675_O_5_2; // @[Top.scala 936:12]
  assign n684_I_6_0 = n675_O_6_0; // @[Top.scala 936:12]
  assign n684_I_6_1 = n675_O_6_1; // @[Top.scala 936:12]
  assign n684_I_6_2 = n675_O_6_2; // @[Top.scala 936:12]
  assign n684_I_7_0 = n675_O_7_0; // @[Top.scala 936:12]
  assign n684_I_7_1 = n675_O_7_1; // @[Top.scala 936:12]
  assign n684_I_7_2 = n675_O_7_2; // @[Top.scala 936:12]
  assign n691_valid_up = n684_valid_down; // @[Top.scala 940:19]
  assign n691_I_0_0_0 = n684_O_0_0_0; // @[Top.scala 939:12]
  assign n691_I_0_0_1 = n684_O_0_0_1; // @[Top.scala 939:12]
  assign n691_I_0_0_2 = n684_O_0_0_2; // @[Top.scala 939:12]
  assign n691_I_1_0_0 = n684_O_1_0_0; // @[Top.scala 939:12]
  assign n691_I_1_0_1 = n684_O_1_0_1; // @[Top.scala 939:12]
  assign n691_I_1_0_2 = n684_O_1_0_2; // @[Top.scala 939:12]
  assign n691_I_2_0_0 = n684_O_2_0_0; // @[Top.scala 939:12]
  assign n691_I_2_0_1 = n684_O_2_0_1; // @[Top.scala 939:12]
  assign n691_I_2_0_2 = n684_O_2_0_2; // @[Top.scala 939:12]
  assign n691_I_3_0_0 = n684_O_3_0_0; // @[Top.scala 939:12]
  assign n691_I_3_0_1 = n684_O_3_0_1; // @[Top.scala 939:12]
  assign n691_I_3_0_2 = n684_O_3_0_2; // @[Top.scala 939:12]
  assign n691_I_4_0_0 = n684_O_4_0_0; // @[Top.scala 939:12]
  assign n691_I_4_0_1 = n684_O_4_0_1; // @[Top.scala 939:12]
  assign n691_I_4_0_2 = n684_O_4_0_2; // @[Top.scala 939:12]
  assign n691_I_5_0_0 = n684_O_5_0_0; // @[Top.scala 939:12]
  assign n691_I_5_0_1 = n684_O_5_0_1; // @[Top.scala 939:12]
  assign n691_I_5_0_2 = n684_O_5_0_2; // @[Top.scala 939:12]
  assign n691_I_6_0_0 = n684_O_6_0_0; // @[Top.scala 939:12]
  assign n691_I_6_0_1 = n684_O_6_0_1; // @[Top.scala 939:12]
  assign n691_I_6_0_2 = n684_O_6_0_2; // @[Top.scala 939:12]
  assign n691_I_7_0_0 = n684_O_7_0_0; // @[Top.scala 939:12]
  assign n691_I_7_0_1 = n684_O_7_0_1; // @[Top.scala 939:12]
  assign n691_I_7_0_2 = n684_O_7_0_2; // @[Top.scala 939:12]
  assign n692_valid_up = n665_valid_down & n691_valid_down; // @[Top.scala 944:19]
  assign n692_I0_0_0 = n665_O_0_0; // @[Top.scala 942:13]
  assign n692_I0_0_1 = n665_O_0_1; // @[Top.scala 942:13]
  assign n692_I0_0_2 = n665_O_0_2; // @[Top.scala 942:13]
  assign n692_I0_1_0 = n665_O_1_0; // @[Top.scala 942:13]
  assign n692_I0_1_1 = n665_O_1_1; // @[Top.scala 942:13]
  assign n692_I0_1_2 = n665_O_1_2; // @[Top.scala 942:13]
  assign n692_I0_2_0 = n665_O_2_0; // @[Top.scala 942:13]
  assign n692_I0_2_1 = n665_O_2_1; // @[Top.scala 942:13]
  assign n692_I0_2_2 = n665_O_2_2; // @[Top.scala 942:13]
  assign n692_I0_3_0 = n665_O_3_0; // @[Top.scala 942:13]
  assign n692_I0_3_1 = n665_O_3_1; // @[Top.scala 942:13]
  assign n692_I0_3_2 = n665_O_3_2; // @[Top.scala 942:13]
  assign n692_I0_4_0 = n665_O_4_0; // @[Top.scala 942:13]
  assign n692_I0_4_1 = n665_O_4_1; // @[Top.scala 942:13]
  assign n692_I0_4_2 = n665_O_4_2; // @[Top.scala 942:13]
  assign n692_I0_5_0 = n665_O_5_0; // @[Top.scala 942:13]
  assign n692_I0_5_1 = n665_O_5_1; // @[Top.scala 942:13]
  assign n692_I0_5_2 = n665_O_5_2; // @[Top.scala 942:13]
  assign n692_I0_6_0 = n665_O_6_0; // @[Top.scala 942:13]
  assign n692_I0_6_1 = n665_O_6_1; // @[Top.scala 942:13]
  assign n692_I0_6_2 = n665_O_6_2; // @[Top.scala 942:13]
  assign n692_I0_7_0 = n665_O_7_0; // @[Top.scala 942:13]
  assign n692_I0_7_1 = n665_O_7_1; // @[Top.scala 942:13]
  assign n692_I0_7_2 = n665_O_7_2; // @[Top.scala 942:13]
  assign n692_I1_0_0 = n691_O_0_0; // @[Top.scala 943:13]
  assign n692_I1_0_1 = n691_O_0_1; // @[Top.scala 943:13]
  assign n692_I1_0_2 = n691_O_0_2; // @[Top.scala 943:13]
  assign n692_I1_1_0 = n691_O_1_0; // @[Top.scala 943:13]
  assign n692_I1_1_1 = n691_O_1_1; // @[Top.scala 943:13]
  assign n692_I1_1_2 = n691_O_1_2; // @[Top.scala 943:13]
  assign n692_I1_2_0 = n691_O_2_0; // @[Top.scala 943:13]
  assign n692_I1_2_1 = n691_O_2_1; // @[Top.scala 943:13]
  assign n692_I1_2_2 = n691_O_2_2; // @[Top.scala 943:13]
  assign n692_I1_3_0 = n691_O_3_0; // @[Top.scala 943:13]
  assign n692_I1_3_1 = n691_O_3_1; // @[Top.scala 943:13]
  assign n692_I1_3_2 = n691_O_3_2; // @[Top.scala 943:13]
  assign n692_I1_4_0 = n691_O_4_0; // @[Top.scala 943:13]
  assign n692_I1_4_1 = n691_O_4_1; // @[Top.scala 943:13]
  assign n692_I1_4_2 = n691_O_4_2; // @[Top.scala 943:13]
  assign n692_I1_5_0 = n691_O_5_0; // @[Top.scala 943:13]
  assign n692_I1_5_1 = n691_O_5_1; // @[Top.scala 943:13]
  assign n692_I1_5_2 = n691_O_5_2; // @[Top.scala 943:13]
  assign n692_I1_6_0 = n691_O_6_0; // @[Top.scala 943:13]
  assign n692_I1_6_1 = n691_O_6_1; // @[Top.scala 943:13]
  assign n692_I1_6_2 = n691_O_6_2; // @[Top.scala 943:13]
  assign n692_I1_7_0 = n691_O_7_0; // @[Top.scala 943:13]
  assign n692_I1_7_1 = n691_O_7_1; // @[Top.scala 943:13]
  assign n692_I1_7_2 = n691_O_7_2; // @[Top.scala 943:13]
  assign n699_clock = clock;
  assign n699_valid_up = n637_valid_down; // @[Top.scala 947:19]
  assign n699_I_0 = n637_O_0; // @[Top.scala 946:12]
  assign n699_I_1 = n637_O_1; // @[Top.scala 946:12]
  assign n699_I_2 = n637_O_2; // @[Top.scala 946:12]
  assign n699_I_3 = n637_O_3; // @[Top.scala 946:12]
  assign n699_I_4 = n637_O_4; // @[Top.scala 946:12]
  assign n699_I_5 = n637_O_5; // @[Top.scala 946:12]
  assign n699_I_6 = n637_O_6; // @[Top.scala 946:12]
  assign n699_I_7 = n637_O_7; // @[Top.scala 946:12]
  assign n700_clock = clock;
  assign n700_valid_up = n699_valid_down; // @[Top.scala 950:19]
  assign n700_I_0 = n699_O_0; // @[Top.scala 949:12]
  assign n700_I_1 = n699_O_1; // @[Top.scala 949:12]
  assign n700_I_2 = n699_O_2; // @[Top.scala 949:12]
  assign n700_I_3 = n699_O_3; // @[Top.scala 949:12]
  assign n700_I_4 = n699_O_4; // @[Top.scala 949:12]
  assign n700_I_5 = n699_O_5; // @[Top.scala 949:12]
  assign n700_I_6 = n699_O_6; // @[Top.scala 949:12]
  assign n700_I_7 = n699_O_7; // @[Top.scala 949:12]
  assign n701_valid_up = n700_valid_down & n699_valid_down; // @[Top.scala 954:19]
  assign n701_I0_0 = n700_O_0; // @[Top.scala 952:13]
  assign n701_I0_1 = n700_O_1; // @[Top.scala 952:13]
  assign n701_I0_2 = n700_O_2; // @[Top.scala 952:13]
  assign n701_I0_3 = n700_O_3; // @[Top.scala 952:13]
  assign n701_I0_4 = n700_O_4; // @[Top.scala 952:13]
  assign n701_I0_5 = n700_O_5; // @[Top.scala 952:13]
  assign n701_I0_6 = n700_O_6; // @[Top.scala 952:13]
  assign n701_I0_7 = n700_O_7; // @[Top.scala 952:13]
  assign n701_I1_0 = n699_O_0; // @[Top.scala 953:13]
  assign n701_I1_1 = n699_O_1; // @[Top.scala 953:13]
  assign n701_I1_2 = n699_O_2; // @[Top.scala 953:13]
  assign n701_I1_3 = n699_O_3; // @[Top.scala 953:13]
  assign n701_I1_4 = n699_O_4; // @[Top.scala 953:13]
  assign n701_I1_5 = n699_O_5; // @[Top.scala 953:13]
  assign n701_I1_6 = n699_O_6; // @[Top.scala 953:13]
  assign n701_I1_7 = n699_O_7; // @[Top.scala 953:13]
  assign n708_valid_up = n701_valid_down & n637_valid_down; // @[Top.scala 958:19]
  assign n708_I0_0_0 = n701_O_0_0; // @[Top.scala 956:13]
  assign n708_I0_0_1 = n701_O_0_1; // @[Top.scala 956:13]
  assign n708_I0_1_0 = n701_O_1_0; // @[Top.scala 956:13]
  assign n708_I0_1_1 = n701_O_1_1; // @[Top.scala 956:13]
  assign n708_I0_2_0 = n701_O_2_0; // @[Top.scala 956:13]
  assign n708_I0_2_1 = n701_O_2_1; // @[Top.scala 956:13]
  assign n708_I0_3_0 = n701_O_3_0; // @[Top.scala 956:13]
  assign n708_I0_3_1 = n701_O_3_1; // @[Top.scala 956:13]
  assign n708_I0_4_0 = n701_O_4_0; // @[Top.scala 956:13]
  assign n708_I0_4_1 = n701_O_4_1; // @[Top.scala 956:13]
  assign n708_I0_5_0 = n701_O_5_0; // @[Top.scala 956:13]
  assign n708_I0_5_1 = n701_O_5_1; // @[Top.scala 956:13]
  assign n708_I0_6_0 = n701_O_6_0; // @[Top.scala 956:13]
  assign n708_I0_6_1 = n701_O_6_1; // @[Top.scala 956:13]
  assign n708_I0_7_0 = n701_O_7_0; // @[Top.scala 956:13]
  assign n708_I0_7_1 = n701_O_7_1; // @[Top.scala 956:13]
  assign n708_I1_0 = n637_O_0; // @[Top.scala 957:13]
  assign n708_I1_1 = n637_O_1; // @[Top.scala 957:13]
  assign n708_I1_2 = n637_O_2; // @[Top.scala 957:13]
  assign n708_I1_3 = n637_O_3; // @[Top.scala 957:13]
  assign n708_I1_4 = n637_O_4; // @[Top.scala 957:13]
  assign n708_I1_5 = n637_O_5; // @[Top.scala 957:13]
  assign n708_I1_6 = n637_O_6; // @[Top.scala 957:13]
  assign n708_I1_7 = n637_O_7; // @[Top.scala 957:13]
  assign n717_valid_up = n708_valid_down; // @[Top.scala 961:19]
  assign n717_I_0_0 = n708_O_0_0; // @[Top.scala 960:12]
  assign n717_I_0_1 = n708_O_0_1; // @[Top.scala 960:12]
  assign n717_I_0_2 = n708_O_0_2; // @[Top.scala 960:12]
  assign n717_I_1_0 = n708_O_1_0; // @[Top.scala 960:12]
  assign n717_I_1_1 = n708_O_1_1; // @[Top.scala 960:12]
  assign n717_I_1_2 = n708_O_1_2; // @[Top.scala 960:12]
  assign n717_I_2_0 = n708_O_2_0; // @[Top.scala 960:12]
  assign n717_I_2_1 = n708_O_2_1; // @[Top.scala 960:12]
  assign n717_I_2_2 = n708_O_2_2; // @[Top.scala 960:12]
  assign n717_I_3_0 = n708_O_3_0; // @[Top.scala 960:12]
  assign n717_I_3_1 = n708_O_3_1; // @[Top.scala 960:12]
  assign n717_I_3_2 = n708_O_3_2; // @[Top.scala 960:12]
  assign n717_I_4_0 = n708_O_4_0; // @[Top.scala 960:12]
  assign n717_I_4_1 = n708_O_4_1; // @[Top.scala 960:12]
  assign n717_I_4_2 = n708_O_4_2; // @[Top.scala 960:12]
  assign n717_I_5_0 = n708_O_5_0; // @[Top.scala 960:12]
  assign n717_I_5_1 = n708_O_5_1; // @[Top.scala 960:12]
  assign n717_I_5_2 = n708_O_5_2; // @[Top.scala 960:12]
  assign n717_I_6_0 = n708_O_6_0; // @[Top.scala 960:12]
  assign n717_I_6_1 = n708_O_6_1; // @[Top.scala 960:12]
  assign n717_I_6_2 = n708_O_6_2; // @[Top.scala 960:12]
  assign n717_I_7_0 = n708_O_7_0; // @[Top.scala 960:12]
  assign n717_I_7_1 = n708_O_7_1; // @[Top.scala 960:12]
  assign n717_I_7_2 = n708_O_7_2; // @[Top.scala 960:12]
  assign n724_valid_up = n717_valid_down; // @[Top.scala 964:19]
  assign n724_I_0_0_0 = n717_O_0_0_0; // @[Top.scala 963:12]
  assign n724_I_0_0_1 = n717_O_0_0_1; // @[Top.scala 963:12]
  assign n724_I_0_0_2 = n717_O_0_0_2; // @[Top.scala 963:12]
  assign n724_I_1_0_0 = n717_O_1_0_0; // @[Top.scala 963:12]
  assign n724_I_1_0_1 = n717_O_1_0_1; // @[Top.scala 963:12]
  assign n724_I_1_0_2 = n717_O_1_0_2; // @[Top.scala 963:12]
  assign n724_I_2_0_0 = n717_O_2_0_0; // @[Top.scala 963:12]
  assign n724_I_2_0_1 = n717_O_2_0_1; // @[Top.scala 963:12]
  assign n724_I_2_0_2 = n717_O_2_0_2; // @[Top.scala 963:12]
  assign n724_I_3_0_0 = n717_O_3_0_0; // @[Top.scala 963:12]
  assign n724_I_3_0_1 = n717_O_3_0_1; // @[Top.scala 963:12]
  assign n724_I_3_0_2 = n717_O_3_0_2; // @[Top.scala 963:12]
  assign n724_I_4_0_0 = n717_O_4_0_0; // @[Top.scala 963:12]
  assign n724_I_4_0_1 = n717_O_4_0_1; // @[Top.scala 963:12]
  assign n724_I_4_0_2 = n717_O_4_0_2; // @[Top.scala 963:12]
  assign n724_I_5_0_0 = n717_O_5_0_0; // @[Top.scala 963:12]
  assign n724_I_5_0_1 = n717_O_5_0_1; // @[Top.scala 963:12]
  assign n724_I_5_0_2 = n717_O_5_0_2; // @[Top.scala 963:12]
  assign n724_I_6_0_0 = n717_O_6_0_0; // @[Top.scala 963:12]
  assign n724_I_6_0_1 = n717_O_6_0_1; // @[Top.scala 963:12]
  assign n724_I_6_0_2 = n717_O_6_0_2; // @[Top.scala 963:12]
  assign n724_I_7_0_0 = n717_O_7_0_0; // @[Top.scala 963:12]
  assign n724_I_7_0_1 = n717_O_7_0_1; // @[Top.scala 963:12]
  assign n724_I_7_0_2 = n717_O_7_0_2; // @[Top.scala 963:12]
  assign n725_valid_up = n692_valid_down & n724_valid_down; // @[Top.scala 968:19]
  assign n725_I0_0_0_0 = n692_O_0_0_0; // @[Top.scala 966:13]
  assign n725_I0_0_0_1 = n692_O_0_0_1; // @[Top.scala 966:13]
  assign n725_I0_0_0_2 = n692_O_0_0_2; // @[Top.scala 966:13]
  assign n725_I0_0_1_0 = n692_O_0_1_0; // @[Top.scala 966:13]
  assign n725_I0_0_1_1 = n692_O_0_1_1; // @[Top.scala 966:13]
  assign n725_I0_0_1_2 = n692_O_0_1_2; // @[Top.scala 966:13]
  assign n725_I0_1_0_0 = n692_O_1_0_0; // @[Top.scala 966:13]
  assign n725_I0_1_0_1 = n692_O_1_0_1; // @[Top.scala 966:13]
  assign n725_I0_1_0_2 = n692_O_1_0_2; // @[Top.scala 966:13]
  assign n725_I0_1_1_0 = n692_O_1_1_0; // @[Top.scala 966:13]
  assign n725_I0_1_1_1 = n692_O_1_1_1; // @[Top.scala 966:13]
  assign n725_I0_1_1_2 = n692_O_1_1_2; // @[Top.scala 966:13]
  assign n725_I0_2_0_0 = n692_O_2_0_0; // @[Top.scala 966:13]
  assign n725_I0_2_0_1 = n692_O_2_0_1; // @[Top.scala 966:13]
  assign n725_I0_2_0_2 = n692_O_2_0_2; // @[Top.scala 966:13]
  assign n725_I0_2_1_0 = n692_O_2_1_0; // @[Top.scala 966:13]
  assign n725_I0_2_1_1 = n692_O_2_1_1; // @[Top.scala 966:13]
  assign n725_I0_2_1_2 = n692_O_2_1_2; // @[Top.scala 966:13]
  assign n725_I0_3_0_0 = n692_O_3_0_0; // @[Top.scala 966:13]
  assign n725_I0_3_0_1 = n692_O_3_0_1; // @[Top.scala 966:13]
  assign n725_I0_3_0_2 = n692_O_3_0_2; // @[Top.scala 966:13]
  assign n725_I0_3_1_0 = n692_O_3_1_0; // @[Top.scala 966:13]
  assign n725_I0_3_1_1 = n692_O_3_1_1; // @[Top.scala 966:13]
  assign n725_I0_3_1_2 = n692_O_3_1_2; // @[Top.scala 966:13]
  assign n725_I0_4_0_0 = n692_O_4_0_0; // @[Top.scala 966:13]
  assign n725_I0_4_0_1 = n692_O_4_0_1; // @[Top.scala 966:13]
  assign n725_I0_4_0_2 = n692_O_4_0_2; // @[Top.scala 966:13]
  assign n725_I0_4_1_0 = n692_O_4_1_0; // @[Top.scala 966:13]
  assign n725_I0_4_1_1 = n692_O_4_1_1; // @[Top.scala 966:13]
  assign n725_I0_4_1_2 = n692_O_4_1_2; // @[Top.scala 966:13]
  assign n725_I0_5_0_0 = n692_O_5_0_0; // @[Top.scala 966:13]
  assign n725_I0_5_0_1 = n692_O_5_0_1; // @[Top.scala 966:13]
  assign n725_I0_5_0_2 = n692_O_5_0_2; // @[Top.scala 966:13]
  assign n725_I0_5_1_0 = n692_O_5_1_0; // @[Top.scala 966:13]
  assign n725_I0_5_1_1 = n692_O_5_1_1; // @[Top.scala 966:13]
  assign n725_I0_5_1_2 = n692_O_5_1_2; // @[Top.scala 966:13]
  assign n725_I0_6_0_0 = n692_O_6_0_0; // @[Top.scala 966:13]
  assign n725_I0_6_0_1 = n692_O_6_0_1; // @[Top.scala 966:13]
  assign n725_I0_6_0_2 = n692_O_6_0_2; // @[Top.scala 966:13]
  assign n725_I0_6_1_0 = n692_O_6_1_0; // @[Top.scala 966:13]
  assign n725_I0_6_1_1 = n692_O_6_1_1; // @[Top.scala 966:13]
  assign n725_I0_6_1_2 = n692_O_6_1_2; // @[Top.scala 966:13]
  assign n725_I0_7_0_0 = n692_O_7_0_0; // @[Top.scala 966:13]
  assign n725_I0_7_0_1 = n692_O_7_0_1; // @[Top.scala 966:13]
  assign n725_I0_7_0_2 = n692_O_7_0_2; // @[Top.scala 966:13]
  assign n725_I0_7_1_0 = n692_O_7_1_0; // @[Top.scala 966:13]
  assign n725_I0_7_1_1 = n692_O_7_1_1; // @[Top.scala 966:13]
  assign n725_I0_7_1_2 = n692_O_7_1_2; // @[Top.scala 966:13]
  assign n725_I1_0_0 = n724_O_0_0; // @[Top.scala 967:13]
  assign n725_I1_0_1 = n724_O_0_1; // @[Top.scala 967:13]
  assign n725_I1_0_2 = n724_O_0_2; // @[Top.scala 967:13]
  assign n725_I1_1_0 = n724_O_1_0; // @[Top.scala 967:13]
  assign n725_I1_1_1 = n724_O_1_1; // @[Top.scala 967:13]
  assign n725_I1_1_2 = n724_O_1_2; // @[Top.scala 967:13]
  assign n725_I1_2_0 = n724_O_2_0; // @[Top.scala 967:13]
  assign n725_I1_2_1 = n724_O_2_1; // @[Top.scala 967:13]
  assign n725_I1_2_2 = n724_O_2_2; // @[Top.scala 967:13]
  assign n725_I1_3_0 = n724_O_3_0; // @[Top.scala 967:13]
  assign n725_I1_3_1 = n724_O_3_1; // @[Top.scala 967:13]
  assign n725_I1_3_2 = n724_O_3_2; // @[Top.scala 967:13]
  assign n725_I1_4_0 = n724_O_4_0; // @[Top.scala 967:13]
  assign n725_I1_4_1 = n724_O_4_1; // @[Top.scala 967:13]
  assign n725_I1_4_2 = n724_O_4_2; // @[Top.scala 967:13]
  assign n725_I1_5_0 = n724_O_5_0; // @[Top.scala 967:13]
  assign n725_I1_5_1 = n724_O_5_1; // @[Top.scala 967:13]
  assign n725_I1_5_2 = n724_O_5_2; // @[Top.scala 967:13]
  assign n725_I1_6_0 = n724_O_6_0; // @[Top.scala 967:13]
  assign n725_I1_6_1 = n724_O_6_1; // @[Top.scala 967:13]
  assign n725_I1_6_2 = n724_O_6_2; // @[Top.scala 967:13]
  assign n725_I1_7_0 = n724_O_7_0; // @[Top.scala 967:13]
  assign n725_I1_7_1 = n724_O_7_1; // @[Top.scala 967:13]
  assign n725_I1_7_2 = n724_O_7_2; // @[Top.scala 967:13]
  assign n734_valid_up = n725_valid_down; // @[Top.scala 971:19]
  assign n734_I_0_0_0 = n725_O_0_0_0; // @[Top.scala 970:12]
  assign n734_I_0_0_1 = n725_O_0_0_1; // @[Top.scala 970:12]
  assign n734_I_0_0_2 = n725_O_0_0_2; // @[Top.scala 970:12]
  assign n734_I_0_1_0 = n725_O_0_1_0; // @[Top.scala 970:12]
  assign n734_I_0_1_1 = n725_O_0_1_1; // @[Top.scala 970:12]
  assign n734_I_0_1_2 = n725_O_0_1_2; // @[Top.scala 970:12]
  assign n734_I_0_2_0 = n725_O_0_2_0; // @[Top.scala 970:12]
  assign n734_I_0_2_1 = n725_O_0_2_1; // @[Top.scala 970:12]
  assign n734_I_0_2_2 = n725_O_0_2_2; // @[Top.scala 970:12]
  assign n734_I_1_0_0 = n725_O_1_0_0; // @[Top.scala 970:12]
  assign n734_I_1_0_1 = n725_O_1_0_1; // @[Top.scala 970:12]
  assign n734_I_1_0_2 = n725_O_1_0_2; // @[Top.scala 970:12]
  assign n734_I_1_1_0 = n725_O_1_1_0; // @[Top.scala 970:12]
  assign n734_I_1_1_1 = n725_O_1_1_1; // @[Top.scala 970:12]
  assign n734_I_1_1_2 = n725_O_1_1_2; // @[Top.scala 970:12]
  assign n734_I_1_2_0 = n725_O_1_2_0; // @[Top.scala 970:12]
  assign n734_I_1_2_1 = n725_O_1_2_1; // @[Top.scala 970:12]
  assign n734_I_1_2_2 = n725_O_1_2_2; // @[Top.scala 970:12]
  assign n734_I_2_0_0 = n725_O_2_0_0; // @[Top.scala 970:12]
  assign n734_I_2_0_1 = n725_O_2_0_1; // @[Top.scala 970:12]
  assign n734_I_2_0_2 = n725_O_2_0_2; // @[Top.scala 970:12]
  assign n734_I_2_1_0 = n725_O_2_1_0; // @[Top.scala 970:12]
  assign n734_I_2_1_1 = n725_O_2_1_1; // @[Top.scala 970:12]
  assign n734_I_2_1_2 = n725_O_2_1_2; // @[Top.scala 970:12]
  assign n734_I_2_2_0 = n725_O_2_2_0; // @[Top.scala 970:12]
  assign n734_I_2_2_1 = n725_O_2_2_1; // @[Top.scala 970:12]
  assign n734_I_2_2_2 = n725_O_2_2_2; // @[Top.scala 970:12]
  assign n734_I_3_0_0 = n725_O_3_0_0; // @[Top.scala 970:12]
  assign n734_I_3_0_1 = n725_O_3_0_1; // @[Top.scala 970:12]
  assign n734_I_3_0_2 = n725_O_3_0_2; // @[Top.scala 970:12]
  assign n734_I_3_1_0 = n725_O_3_1_0; // @[Top.scala 970:12]
  assign n734_I_3_1_1 = n725_O_3_1_1; // @[Top.scala 970:12]
  assign n734_I_3_1_2 = n725_O_3_1_2; // @[Top.scala 970:12]
  assign n734_I_3_2_0 = n725_O_3_2_0; // @[Top.scala 970:12]
  assign n734_I_3_2_1 = n725_O_3_2_1; // @[Top.scala 970:12]
  assign n734_I_3_2_2 = n725_O_3_2_2; // @[Top.scala 970:12]
  assign n734_I_4_0_0 = n725_O_4_0_0; // @[Top.scala 970:12]
  assign n734_I_4_0_1 = n725_O_4_0_1; // @[Top.scala 970:12]
  assign n734_I_4_0_2 = n725_O_4_0_2; // @[Top.scala 970:12]
  assign n734_I_4_1_0 = n725_O_4_1_0; // @[Top.scala 970:12]
  assign n734_I_4_1_1 = n725_O_4_1_1; // @[Top.scala 970:12]
  assign n734_I_4_1_2 = n725_O_4_1_2; // @[Top.scala 970:12]
  assign n734_I_4_2_0 = n725_O_4_2_0; // @[Top.scala 970:12]
  assign n734_I_4_2_1 = n725_O_4_2_1; // @[Top.scala 970:12]
  assign n734_I_4_2_2 = n725_O_4_2_2; // @[Top.scala 970:12]
  assign n734_I_5_0_0 = n725_O_5_0_0; // @[Top.scala 970:12]
  assign n734_I_5_0_1 = n725_O_5_0_1; // @[Top.scala 970:12]
  assign n734_I_5_0_2 = n725_O_5_0_2; // @[Top.scala 970:12]
  assign n734_I_5_1_0 = n725_O_5_1_0; // @[Top.scala 970:12]
  assign n734_I_5_1_1 = n725_O_5_1_1; // @[Top.scala 970:12]
  assign n734_I_5_1_2 = n725_O_5_1_2; // @[Top.scala 970:12]
  assign n734_I_5_2_0 = n725_O_5_2_0; // @[Top.scala 970:12]
  assign n734_I_5_2_1 = n725_O_5_2_1; // @[Top.scala 970:12]
  assign n734_I_5_2_2 = n725_O_5_2_2; // @[Top.scala 970:12]
  assign n734_I_6_0_0 = n725_O_6_0_0; // @[Top.scala 970:12]
  assign n734_I_6_0_1 = n725_O_6_0_1; // @[Top.scala 970:12]
  assign n734_I_6_0_2 = n725_O_6_0_2; // @[Top.scala 970:12]
  assign n734_I_6_1_0 = n725_O_6_1_0; // @[Top.scala 970:12]
  assign n734_I_6_1_1 = n725_O_6_1_1; // @[Top.scala 970:12]
  assign n734_I_6_1_2 = n725_O_6_1_2; // @[Top.scala 970:12]
  assign n734_I_6_2_0 = n725_O_6_2_0; // @[Top.scala 970:12]
  assign n734_I_6_2_1 = n725_O_6_2_1; // @[Top.scala 970:12]
  assign n734_I_6_2_2 = n725_O_6_2_2; // @[Top.scala 970:12]
  assign n734_I_7_0_0 = n725_O_7_0_0; // @[Top.scala 970:12]
  assign n734_I_7_0_1 = n725_O_7_0_1; // @[Top.scala 970:12]
  assign n734_I_7_0_2 = n725_O_7_0_2; // @[Top.scala 970:12]
  assign n734_I_7_1_0 = n725_O_7_1_0; // @[Top.scala 970:12]
  assign n734_I_7_1_1 = n725_O_7_1_1; // @[Top.scala 970:12]
  assign n734_I_7_1_2 = n725_O_7_1_2; // @[Top.scala 970:12]
  assign n734_I_7_2_0 = n725_O_7_2_0; // @[Top.scala 970:12]
  assign n734_I_7_2_1 = n725_O_7_2_1; // @[Top.scala 970:12]
  assign n734_I_7_2_2 = n725_O_7_2_2; // @[Top.scala 970:12]
  assign n741_valid_up = n734_valid_down; // @[Top.scala 974:19]
  assign n741_I_0_0_0_0 = n734_O_0_0_0_0; // @[Top.scala 973:12]
  assign n741_I_0_0_0_1 = n734_O_0_0_0_1; // @[Top.scala 973:12]
  assign n741_I_0_0_0_2 = n734_O_0_0_0_2; // @[Top.scala 973:12]
  assign n741_I_0_0_1_0 = n734_O_0_0_1_0; // @[Top.scala 973:12]
  assign n741_I_0_0_1_1 = n734_O_0_0_1_1; // @[Top.scala 973:12]
  assign n741_I_0_0_1_2 = n734_O_0_0_1_2; // @[Top.scala 973:12]
  assign n741_I_0_0_2_0 = n734_O_0_0_2_0; // @[Top.scala 973:12]
  assign n741_I_0_0_2_1 = n734_O_0_0_2_1; // @[Top.scala 973:12]
  assign n741_I_0_0_2_2 = n734_O_0_0_2_2; // @[Top.scala 973:12]
  assign n741_I_1_0_0_0 = n734_O_1_0_0_0; // @[Top.scala 973:12]
  assign n741_I_1_0_0_1 = n734_O_1_0_0_1; // @[Top.scala 973:12]
  assign n741_I_1_0_0_2 = n734_O_1_0_0_2; // @[Top.scala 973:12]
  assign n741_I_1_0_1_0 = n734_O_1_0_1_0; // @[Top.scala 973:12]
  assign n741_I_1_0_1_1 = n734_O_1_0_1_1; // @[Top.scala 973:12]
  assign n741_I_1_0_1_2 = n734_O_1_0_1_2; // @[Top.scala 973:12]
  assign n741_I_1_0_2_0 = n734_O_1_0_2_0; // @[Top.scala 973:12]
  assign n741_I_1_0_2_1 = n734_O_1_0_2_1; // @[Top.scala 973:12]
  assign n741_I_1_0_2_2 = n734_O_1_0_2_2; // @[Top.scala 973:12]
  assign n741_I_2_0_0_0 = n734_O_2_0_0_0; // @[Top.scala 973:12]
  assign n741_I_2_0_0_1 = n734_O_2_0_0_1; // @[Top.scala 973:12]
  assign n741_I_2_0_0_2 = n734_O_2_0_0_2; // @[Top.scala 973:12]
  assign n741_I_2_0_1_0 = n734_O_2_0_1_0; // @[Top.scala 973:12]
  assign n741_I_2_0_1_1 = n734_O_2_0_1_1; // @[Top.scala 973:12]
  assign n741_I_2_0_1_2 = n734_O_2_0_1_2; // @[Top.scala 973:12]
  assign n741_I_2_0_2_0 = n734_O_2_0_2_0; // @[Top.scala 973:12]
  assign n741_I_2_0_2_1 = n734_O_2_0_2_1; // @[Top.scala 973:12]
  assign n741_I_2_0_2_2 = n734_O_2_0_2_2; // @[Top.scala 973:12]
  assign n741_I_3_0_0_0 = n734_O_3_0_0_0; // @[Top.scala 973:12]
  assign n741_I_3_0_0_1 = n734_O_3_0_0_1; // @[Top.scala 973:12]
  assign n741_I_3_0_0_2 = n734_O_3_0_0_2; // @[Top.scala 973:12]
  assign n741_I_3_0_1_0 = n734_O_3_0_1_0; // @[Top.scala 973:12]
  assign n741_I_3_0_1_1 = n734_O_3_0_1_1; // @[Top.scala 973:12]
  assign n741_I_3_0_1_2 = n734_O_3_0_1_2; // @[Top.scala 973:12]
  assign n741_I_3_0_2_0 = n734_O_3_0_2_0; // @[Top.scala 973:12]
  assign n741_I_3_0_2_1 = n734_O_3_0_2_1; // @[Top.scala 973:12]
  assign n741_I_3_0_2_2 = n734_O_3_0_2_2; // @[Top.scala 973:12]
  assign n741_I_4_0_0_0 = n734_O_4_0_0_0; // @[Top.scala 973:12]
  assign n741_I_4_0_0_1 = n734_O_4_0_0_1; // @[Top.scala 973:12]
  assign n741_I_4_0_0_2 = n734_O_4_0_0_2; // @[Top.scala 973:12]
  assign n741_I_4_0_1_0 = n734_O_4_0_1_0; // @[Top.scala 973:12]
  assign n741_I_4_0_1_1 = n734_O_4_0_1_1; // @[Top.scala 973:12]
  assign n741_I_4_0_1_2 = n734_O_4_0_1_2; // @[Top.scala 973:12]
  assign n741_I_4_0_2_0 = n734_O_4_0_2_0; // @[Top.scala 973:12]
  assign n741_I_4_0_2_1 = n734_O_4_0_2_1; // @[Top.scala 973:12]
  assign n741_I_4_0_2_2 = n734_O_4_0_2_2; // @[Top.scala 973:12]
  assign n741_I_5_0_0_0 = n734_O_5_0_0_0; // @[Top.scala 973:12]
  assign n741_I_5_0_0_1 = n734_O_5_0_0_1; // @[Top.scala 973:12]
  assign n741_I_5_0_0_2 = n734_O_5_0_0_2; // @[Top.scala 973:12]
  assign n741_I_5_0_1_0 = n734_O_5_0_1_0; // @[Top.scala 973:12]
  assign n741_I_5_0_1_1 = n734_O_5_0_1_1; // @[Top.scala 973:12]
  assign n741_I_5_0_1_2 = n734_O_5_0_1_2; // @[Top.scala 973:12]
  assign n741_I_5_0_2_0 = n734_O_5_0_2_0; // @[Top.scala 973:12]
  assign n741_I_5_0_2_1 = n734_O_5_0_2_1; // @[Top.scala 973:12]
  assign n741_I_5_0_2_2 = n734_O_5_0_2_2; // @[Top.scala 973:12]
  assign n741_I_6_0_0_0 = n734_O_6_0_0_0; // @[Top.scala 973:12]
  assign n741_I_6_0_0_1 = n734_O_6_0_0_1; // @[Top.scala 973:12]
  assign n741_I_6_0_0_2 = n734_O_6_0_0_2; // @[Top.scala 973:12]
  assign n741_I_6_0_1_0 = n734_O_6_0_1_0; // @[Top.scala 973:12]
  assign n741_I_6_0_1_1 = n734_O_6_0_1_1; // @[Top.scala 973:12]
  assign n741_I_6_0_1_2 = n734_O_6_0_1_2; // @[Top.scala 973:12]
  assign n741_I_6_0_2_0 = n734_O_6_0_2_0; // @[Top.scala 973:12]
  assign n741_I_6_0_2_1 = n734_O_6_0_2_1; // @[Top.scala 973:12]
  assign n741_I_6_0_2_2 = n734_O_6_0_2_2; // @[Top.scala 973:12]
  assign n741_I_7_0_0_0 = n734_O_7_0_0_0; // @[Top.scala 973:12]
  assign n741_I_7_0_0_1 = n734_O_7_0_0_1; // @[Top.scala 973:12]
  assign n741_I_7_0_0_2 = n734_O_7_0_0_2; // @[Top.scala 973:12]
  assign n741_I_7_0_1_0 = n734_O_7_0_1_0; // @[Top.scala 973:12]
  assign n741_I_7_0_1_1 = n734_O_7_0_1_1; // @[Top.scala 973:12]
  assign n741_I_7_0_1_2 = n734_O_7_0_1_2; // @[Top.scala 973:12]
  assign n741_I_7_0_2_0 = n734_O_7_0_2_0; // @[Top.scala 973:12]
  assign n741_I_7_0_2_1 = n734_O_7_0_2_1; // @[Top.scala 973:12]
  assign n741_I_7_0_2_2 = n734_O_7_0_2_2; // @[Top.scala 973:12]
  assign n783_clock = clock;
  assign n783_reset = reset;
  assign n783_valid_up = n741_valid_down; // @[Top.scala 977:19]
  assign n783_I_0_0_0 = n741_O_0_0_0; // @[Top.scala 976:12]
  assign n783_I_0_0_1 = n741_O_0_0_1; // @[Top.scala 976:12]
  assign n783_I_0_0_2 = n741_O_0_0_2; // @[Top.scala 976:12]
  assign n783_I_0_1_0 = n741_O_0_1_0; // @[Top.scala 976:12]
  assign n783_I_0_1_1 = n741_O_0_1_1; // @[Top.scala 976:12]
  assign n783_I_0_1_2 = n741_O_0_1_2; // @[Top.scala 976:12]
  assign n783_I_0_2_0 = n741_O_0_2_0; // @[Top.scala 976:12]
  assign n783_I_0_2_1 = n741_O_0_2_1; // @[Top.scala 976:12]
  assign n783_I_0_2_2 = n741_O_0_2_2; // @[Top.scala 976:12]
  assign n783_I_1_0_0 = n741_O_1_0_0; // @[Top.scala 976:12]
  assign n783_I_1_0_1 = n741_O_1_0_1; // @[Top.scala 976:12]
  assign n783_I_1_0_2 = n741_O_1_0_2; // @[Top.scala 976:12]
  assign n783_I_1_1_0 = n741_O_1_1_0; // @[Top.scala 976:12]
  assign n783_I_1_1_1 = n741_O_1_1_1; // @[Top.scala 976:12]
  assign n783_I_1_1_2 = n741_O_1_1_2; // @[Top.scala 976:12]
  assign n783_I_1_2_0 = n741_O_1_2_0; // @[Top.scala 976:12]
  assign n783_I_1_2_1 = n741_O_1_2_1; // @[Top.scala 976:12]
  assign n783_I_1_2_2 = n741_O_1_2_2; // @[Top.scala 976:12]
  assign n783_I_2_0_0 = n741_O_2_0_0; // @[Top.scala 976:12]
  assign n783_I_2_0_1 = n741_O_2_0_1; // @[Top.scala 976:12]
  assign n783_I_2_0_2 = n741_O_2_0_2; // @[Top.scala 976:12]
  assign n783_I_2_1_0 = n741_O_2_1_0; // @[Top.scala 976:12]
  assign n783_I_2_1_1 = n741_O_2_1_1; // @[Top.scala 976:12]
  assign n783_I_2_1_2 = n741_O_2_1_2; // @[Top.scala 976:12]
  assign n783_I_2_2_0 = n741_O_2_2_0; // @[Top.scala 976:12]
  assign n783_I_2_2_1 = n741_O_2_2_1; // @[Top.scala 976:12]
  assign n783_I_2_2_2 = n741_O_2_2_2; // @[Top.scala 976:12]
  assign n783_I_3_0_0 = n741_O_3_0_0; // @[Top.scala 976:12]
  assign n783_I_3_0_1 = n741_O_3_0_1; // @[Top.scala 976:12]
  assign n783_I_3_0_2 = n741_O_3_0_2; // @[Top.scala 976:12]
  assign n783_I_3_1_0 = n741_O_3_1_0; // @[Top.scala 976:12]
  assign n783_I_3_1_1 = n741_O_3_1_1; // @[Top.scala 976:12]
  assign n783_I_3_1_2 = n741_O_3_1_2; // @[Top.scala 976:12]
  assign n783_I_3_2_0 = n741_O_3_2_0; // @[Top.scala 976:12]
  assign n783_I_3_2_1 = n741_O_3_2_1; // @[Top.scala 976:12]
  assign n783_I_3_2_2 = n741_O_3_2_2; // @[Top.scala 976:12]
  assign n783_I_4_0_0 = n741_O_4_0_0; // @[Top.scala 976:12]
  assign n783_I_4_0_1 = n741_O_4_0_1; // @[Top.scala 976:12]
  assign n783_I_4_0_2 = n741_O_4_0_2; // @[Top.scala 976:12]
  assign n783_I_4_1_0 = n741_O_4_1_0; // @[Top.scala 976:12]
  assign n783_I_4_1_1 = n741_O_4_1_1; // @[Top.scala 976:12]
  assign n783_I_4_1_2 = n741_O_4_1_2; // @[Top.scala 976:12]
  assign n783_I_4_2_0 = n741_O_4_2_0; // @[Top.scala 976:12]
  assign n783_I_4_2_1 = n741_O_4_2_1; // @[Top.scala 976:12]
  assign n783_I_4_2_2 = n741_O_4_2_2; // @[Top.scala 976:12]
  assign n783_I_5_0_0 = n741_O_5_0_0; // @[Top.scala 976:12]
  assign n783_I_5_0_1 = n741_O_5_0_1; // @[Top.scala 976:12]
  assign n783_I_5_0_2 = n741_O_5_0_2; // @[Top.scala 976:12]
  assign n783_I_5_1_0 = n741_O_5_1_0; // @[Top.scala 976:12]
  assign n783_I_5_1_1 = n741_O_5_1_1; // @[Top.scala 976:12]
  assign n783_I_5_1_2 = n741_O_5_1_2; // @[Top.scala 976:12]
  assign n783_I_5_2_0 = n741_O_5_2_0; // @[Top.scala 976:12]
  assign n783_I_5_2_1 = n741_O_5_2_1; // @[Top.scala 976:12]
  assign n783_I_5_2_2 = n741_O_5_2_2; // @[Top.scala 976:12]
  assign n783_I_6_0_0 = n741_O_6_0_0; // @[Top.scala 976:12]
  assign n783_I_6_0_1 = n741_O_6_0_1; // @[Top.scala 976:12]
  assign n783_I_6_0_2 = n741_O_6_0_2; // @[Top.scala 976:12]
  assign n783_I_6_1_0 = n741_O_6_1_0; // @[Top.scala 976:12]
  assign n783_I_6_1_1 = n741_O_6_1_1; // @[Top.scala 976:12]
  assign n783_I_6_1_2 = n741_O_6_1_2; // @[Top.scala 976:12]
  assign n783_I_6_2_0 = n741_O_6_2_0; // @[Top.scala 976:12]
  assign n783_I_6_2_1 = n741_O_6_2_1; // @[Top.scala 976:12]
  assign n783_I_6_2_2 = n741_O_6_2_2; // @[Top.scala 976:12]
  assign n783_I_7_0_0 = n741_O_7_0_0; // @[Top.scala 976:12]
  assign n783_I_7_0_1 = n741_O_7_0_1; // @[Top.scala 976:12]
  assign n783_I_7_0_2 = n741_O_7_0_2; // @[Top.scala 976:12]
  assign n783_I_7_1_0 = n741_O_7_1_0; // @[Top.scala 976:12]
  assign n783_I_7_1_1 = n741_O_7_1_1; // @[Top.scala 976:12]
  assign n783_I_7_1_2 = n741_O_7_1_2; // @[Top.scala 976:12]
  assign n783_I_7_2_0 = n741_O_7_2_0; // @[Top.scala 976:12]
  assign n783_I_7_2_1 = n741_O_7_2_1; // @[Top.scala 976:12]
  assign n783_I_7_2_2 = n741_O_7_2_2; // @[Top.scala 976:12]
  assign n784_valid_up = n783_valid_down; // @[Top.scala 980:19]
  assign n784_I_0_0_0 = n783_O_0_0_0; // @[Top.scala 979:12]
  assign n784_I_1_0_0 = n783_O_1_0_0; // @[Top.scala 979:12]
  assign n784_I_2_0_0 = n783_O_2_0_0; // @[Top.scala 979:12]
  assign n784_I_3_0_0 = n783_O_3_0_0; // @[Top.scala 979:12]
  assign n784_I_4_0_0 = n783_O_4_0_0; // @[Top.scala 979:12]
  assign n784_I_5_0_0 = n783_O_5_0_0; // @[Top.scala 979:12]
  assign n784_I_6_0_0 = n783_O_6_0_0; // @[Top.scala 979:12]
  assign n784_I_7_0_0 = n783_O_7_0_0; // @[Top.scala 979:12]
  assign n785_valid_up = n784_valid_down; // @[Top.scala 983:19]
  assign n785_I_0_0 = n784_O_0_0; // @[Top.scala 982:12]
  assign n785_I_1_0 = n784_O_1_0; // @[Top.scala 982:12]
  assign n785_I_2_0 = n784_O_2_0; // @[Top.scala 982:12]
  assign n785_I_3_0 = n784_O_3_0; // @[Top.scala 982:12]
  assign n785_I_4_0 = n784_O_4_0; // @[Top.scala 982:12]
  assign n785_I_5_0 = n784_O_5_0; // @[Top.scala 982:12]
  assign n785_I_6_0 = n784_O_6_0; // @[Top.scala 982:12]
  assign n785_I_7_0 = n784_O_7_0; // @[Top.scala 982:12]
  assign n786_clock = clock;
  assign n786_reset = reset;
  assign n786_valid_up = n637_valid_down; // @[Top.scala 986:19]
  assign n786_I_0 = n637_O_0; // @[Top.scala 985:12]
  assign n786_I_1 = n637_O_1; // @[Top.scala 985:12]
  assign n786_I_2 = n637_O_2; // @[Top.scala 985:12]
  assign n786_I_3 = n637_O_3; // @[Top.scala 985:12]
  assign n786_I_4 = n637_O_4; // @[Top.scala 985:12]
  assign n786_I_5 = n637_O_5; // @[Top.scala 985:12]
  assign n786_I_6 = n637_O_6; // @[Top.scala 985:12]
  assign n786_I_7 = n637_O_7; // @[Top.scala 985:12]
  assign n787_clock = clock;
  assign n787_reset = reset;
  assign n787_valid_up = n785_valid_down & n786_valid_down; // @[Top.scala 990:19]
  assign n787_I0_0 = n785_O_0; // @[Top.scala 988:13]
  assign n787_I0_1 = n785_O_1; // @[Top.scala 988:13]
  assign n787_I0_2 = n785_O_2; // @[Top.scala 988:13]
  assign n787_I0_3 = n785_O_3; // @[Top.scala 988:13]
  assign n787_I0_4 = n785_O_4; // @[Top.scala 988:13]
  assign n787_I0_5 = n785_O_5; // @[Top.scala 988:13]
  assign n787_I0_6 = n785_O_6; // @[Top.scala 988:13]
  assign n787_I0_7 = n785_O_7; // @[Top.scala 988:13]
  assign n787_I1_0 = n786_O_0; // @[Top.scala 989:13]
  assign n787_I1_1 = n786_O_1; // @[Top.scala 989:13]
  assign n787_I1_2 = n786_O_2; // @[Top.scala 989:13]
  assign n787_I1_3 = n786_O_3; // @[Top.scala 989:13]
  assign n787_I1_4 = n786_O_4; // @[Top.scala 989:13]
  assign n787_I1_5 = n786_O_5; // @[Top.scala 989:13]
  assign n787_I1_6 = n786_O_6; // @[Top.scala 989:13]
  assign n787_I1_7 = n786_O_7; // @[Top.scala 989:13]
  assign n823_valid_up = n446_valid_down; // @[Top.scala 993:19]
  assign n823_I_0_t1b_t0b = n446_O_0_t1b_t0b; // @[Top.scala 992:12]
  assign n823_I_0_t1b_t1b = n446_O_0_t1b_t1b; // @[Top.scala 992:12]
  assign n823_I_1_t1b_t0b = n446_O_1_t1b_t0b; // @[Top.scala 992:12]
  assign n823_I_1_t1b_t1b = n446_O_1_t1b_t1b; // @[Top.scala 992:12]
  assign n823_I_2_t1b_t0b = n446_O_2_t1b_t0b; // @[Top.scala 992:12]
  assign n823_I_2_t1b_t1b = n446_O_2_t1b_t1b; // @[Top.scala 992:12]
  assign n823_I_3_t1b_t0b = n446_O_3_t1b_t0b; // @[Top.scala 992:12]
  assign n823_I_3_t1b_t1b = n446_O_3_t1b_t1b; // @[Top.scala 992:12]
  assign n823_I_4_t1b_t0b = n446_O_4_t1b_t0b; // @[Top.scala 992:12]
  assign n823_I_4_t1b_t1b = n446_O_4_t1b_t1b; // @[Top.scala 992:12]
  assign n823_I_5_t1b_t0b = n446_O_5_t1b_t0b; // @[Top.scala 992:12]
  assign n823_I_5_t1b_t1b = n446_O_5_t1b_t1b; // @[Top.scala 992:12]
  assign n823_I_6_t1b_t0b = n446_O_6_t1b_t0b; // @[Top.scala 992:12]
  assign n823_I_6_t1b_t1b = n446_O_6_t1b_t1b; // @[Top.scala 992:12]
  assign n823_I_7_t1b_t0b = n446_O_7_t1b_t0b; // @[Top.scala 992:12]
  assign n823_I_7_t1b_t1b = n446_O_7_t1b_t1b; // @[Top.scala 992:12]
  assign n824_clock = clock;
  assign n824_reset = reset;
  assign n824_valid_up = n823_valid_down; // @[Top.scala 996:19]
  assign n824_I_0 = n823_O_0; // @[Top.scala 995:12]
  assign n824_I_1 = n823_O_1; // @[Top.scala 995:12]
  assign n824_I_2 = n823_O_2; // @[Top.scala 995:12]
  assign n824_I_3 = n823_O_3; // @[Top.scala 995:12]
  assign n824_I_4 = n823_O_4; // @[Top.scala 995:12]
  assign n824_I_5 = n823_O_5; // @[Top.scala 995:12]
  assign n824_I_6 = n823_O_6; // @[Top.scala 995:12]
  assign n824_I_7 = n823_O_7; // @[Top.scala 995:12]
  assign n825_clock = clock;
  assign n825_reset = reset;
  assign n825_valid_up = n824_valid_down; // @[Top.scala 999:19]
  assign n825_I_0 = n824_O_0; // @[Top.scala 998:12]
  assign n825_I_1 = n824_O_1; // @[Top.scala 998:12]
  assign n825_I_2 = n824_O_2; // @[Top.scala 998:12]
  assign n825_I_3 = n824_O_3; // @[Top.scala 998:12]
  assign n825_I_4 = n824_O_4; // @[Top.scala 998:12]
  assign n825_I_5 = n824_O_5; // @[Top.scala 998:12]
  assign n825_I_6 = n824_O_6; // @[Top.scala 998:12]
  assign n825_I_7 = n824_O_7; // @[Top.scala 998:12]
  assign n826_clock = clock;
  assign n826_valid_up = n825_valid_down; // @[Top.scala 1002:19]
  assign n826_I_0 = n825_O_0; // @[Top.scala 1001:12]
  assign n826_I_1 = n825_O_1; // @[Top.scala 1001:12]
  assign n826_I_2 = n825_O_2; // @[Top.scala 1001:12]
  assign n826_I_3 = n825_O_3; // @[Top.scala 1001:12]
  assign n826_I_4 = n825_O_4; // @[Top.scala 1001:12]
  assign n826_I_5 = n825_O_5; // @[Top.scala 1001:12]
  assign n826_I_6 = n825_O_6; // @[Top.scala 1001:12]
  assign n826_I_7 = n825_O_7; // @[Top.scala 1001:12]
  assign n827_clock = clock;
  assign n827_valid_up = n826_valid_down; // @[Top.scala 1005:19]
  assign n827_I_0 = n826_O_0; // @[Top.scala 1004:12]
  assign n827_I_1 = n826_O_1; // @[Top.scala 1004:12]
  assign n827_I_2 = n826_O_2; // @[Top.scala 1004:12]
  assign n827_I_3 = n826_O_3; // @[Top.scala 1004:12]
  assign n827_I_4 = n826_O_4; // @[Top.scala 1004:12]
  assign n827_I_5 = n826_O_5; // @[Top.scala 1004:12]
  assign n827_I_6 = n826_O_6; // @[Top.scala 1004:12]
  assign n827_I_7 = n826_O_7; // @[Top.scala 1004:12]
  assign n828_valid_up = n827_valid_down & n826_valid_down; // @[Top.scala 1009:19]
  assign n828_I0_0 = n827_O_0; // @[Top.scala 1007:13]
  assign n828_I0_1 = n827_O_1; // @[Top.scala 1007:13]
  assign n828_I0_2 = n827_O_2; // @[Top.scala 1007:13]
  assign n828_I0_3 = n827_O_3; // @[Top.scala 1007:13]
  assign n828_I0_4 = n827_O_4; // @[Top.scala 1007:13]
  assign n828_I0_5 = n827_O_5; // @[Top.scala 1007:13]
  assign n828_I0_6 = n827_O_6; // @[Top.scala 1007:13]
  assign n828_I0_7 = n827_O_7; // @[Top.scala 1007:13]
  assign n828_I1_0 = n826_O_0; // @[Top.scala 1008:13]
  assign n828_I1_1 = n826_O_1; // @[Top.scala 1008:13]
  assign n828_I1_2 = n826_O_2; // @[Top.scala 1008:13]
  assign n828_I1_3 = n826_O_3; // @[Top.scala 1008:13]
  assign n828_I1_4 = n826_O_4; // @[Top.scala 1008:13]
  assign n828_I1_5 = n826_O_5; // @[Top.scala 1008:13]
  assign n828_I1_6 = n826_O_6; // @[Top.scala 1008:13]
  assign n828_I1_7 = n826_O_7; // @[Top.scala 1008:13]
  assign n835_valid_up = n828_valid_down & n825_valid_down; // @[Top.scala 1013:19]
  assign n835_I0_0_0 = n828_O_0_0; // @[Top.scala 1011:13]
  assign n835_I0_0_1 = n828_O_0_1; // @[Top.scala 1011:13]
  assign n835_I0_1_0 = n828_O_1_0; // @[Top.scala 1011:13]
  assign n835_I0_1_1 = n828_O_1_1; // @[Top.scala 1011:13]
  assign n835_I0_2_0 = n828_O_2_0; // @[Top.scala 1011:13]
  assign n835_I0_2_1 = n828_O_2_1; // @[Top.scala 1011:13]
  assign n835_I0_3_0 = n828_O_3_0; // @[Top.scala 1011:13]
  assign n835_I0_3_1 = n828_O_3_1; // @[Top.scala 1011:13]
  assign n835_I0_4_0 = n828_O_4_0; // @[Top.scala 1011:13]
  assign n835_I0_4_1 = n828_O_4_1; // @[Top.scala 1011:13]
  assign n835_I0_5_0 = n828_O_5_0; // @[Top.scala 1011:13]
  assign n835_I0_5_1 = n828_O_5_1; // @[Top.scala 1011:13]
  assign n835_I0_6_0 = n828_O_6_0; // @[Top.scala 1011:13]
  assign n835_I0_6_1 = n828_O_6_1; // @[Top.scala 1011:13]
  assign n835_I0_7_0 = n828_O_7_0; // @[Top.scala 1011:13]
  assign n835_I0_7_1 = n828_O_7_1; // @[Top.scala 1011:13]
  assign n835_I1_0 = n825_O_0; // @[Top.scala 1012:13]
  assign n835_I1_1 = n825_O_1; // @[Top.scala 1012:13]
  assign n835_I1_2 = n825_O_2; // @[Top.scala 1012:13]
  assign n835_I1_3 = n825_O_3; // @[Top.scala 1012:13]
  assign n835_I1_4 = n825_O_4; // @[Top.scala 1012:13]
  assign n835_I1_5 = n825_O_5; // @[Top.scala 1012:13]
  assign n835_I1_6 = n825_O_6; // @[Top.scala 1012:13]
  assign n835_I1_7 = n825_O_7; // @[Top.scala 1012:13]
  assign n844_valid_up = n835_valid_down; // @[Top.scala 1016:19]
  assign n844_I_0_0 = n835_O_0_0; // @[Top.scala 1015:12]
  assign n844_I_0_1 = n835_O_0_1; // @[Top.scala 1015:12]
  assign n844_I_0_2 = n835_O_0_2; // @[Top.scala 1015:12]
  assign n844_I_1_0 = n835_O_1_0; // @[Top.scala 1015:12]
  assign n844_I_1_1 = n835_O_1_1; // @[Top.scala 1015:12]
  assign n844_I_1_2 = n835_O_1_2; // @[Top.scala 1015:12]
  assign n844_I_2_0 = n835_O_2_0; // @[Top.scala 1015:12]
  assign n844_I_2_1 = n835_O_2_1; // @[Top.scala 1015:12]
  assign n844_I_2_2 = n835_O_2_2; // @[Top.scala 1015:12]
  assign n844_I_3_0 = n835_O_3_0; // @[Top.scala 1015:12]
  assign n844_I_3_1 = n835_O_3_1; // @[Top.scala 1015:12]
  assign n844_I_3_2 = n835_O_3_2; // @[Top.scala 1015:12]
  assign n844_I_4_0 = n835_O_4_0; // @[Top.scala 1015:12]
  assign n844_I_4_1 = n835_O_4_1; // @[Top.scala 1015:12]
  assign n844_I_4_2 = n835_O_4_2; // @[Top.scala 1015:12]
  assign n844_I_5_0 = n835_O_5_0; // @[Top.scala 1015:12]
  assign n844_I_5_1 = n835_O_5_1; // @[Top.scala 1015:12]
  assign n844_I_5_2 = n835_O_5_2; // @[Top.scala 1015:12]
  assign n844_I_6_0 = n835_O_6_0; // @[Top.scala 1015:12]
  assign n844_I_6_1 = n835_O_6_1; // @[Top.scala 1015:12]
  assign n844_I_6_2 = n835_O_6_2; // @[Top.scala 1015:12]
  assign n844_I_7_0 = n835_O_7_0; // @[Top.scala 1015:12]
  assign n844_I_7_1 = n835_O_7_1; // @[Top.scala 1015:12]
  assign n844_I_7_2 = n835_O_7_2; // @[Top.scala 1015:12]
  assign n851_valid_up = n844_valid_down; // @[Top.scala 1019:19]
  assign n851_I_0_0_0 = n844_O_0_0_0; // @[Top.scala 1018:12]
  assign n851_I_0_0_1 = n844_O_0_0_1; // @[Top.scala 1018:12]
  assign n851_I_0_0_2 = n844_O_0_0_2; // @[Top.scala 1018:12]
  assign n851_I_1_0_0 = n844_O_1_0_0; // @[Top.scala 1018:12]
  assign n851_I_1_0_1 = n844_O_1_0_1; // @[Top.scala 1018:12]
  assign n851_I_1_0_2 = n844_O_1_0_2; // @[Top.scala 1018:12]
  assign n851_I_2_0_0 = n844_O_2_0_0; // @[Top.scala 1018:12]
  assign n851_I_2_0_1 = n844_O_2_0_1; // @[Top.scala 1018:12]
  assign n851_I_2_0_2 = n844_O_2_0_2; // @[Top.scala 1018:12]
  assign n851_I_3_0_0 = n844_O_3_0_0; // @[Top.scala 1018:12]
  assign n851_I_3_0_1 = n844_O_3_0_1; // @[Top.scala 1018:12]
  assign n851_I_3_0_2 = n844_O_3_0_2; // @[Top.scala 1018:12]
  assign n851_I_4_0_0 = n844_O_4_0_0; // @[Top.scala 1018:12]
  assign n851_I_4_0_1 = n844_O_4_0_1; // @[Top.scala 1018:12]
  assign n851_I_4_0_2 = n844_O_4_0_2; // @[Top.scala 1018:12]
  assign n851_I_5_0_0 = n844_O_5_0_0; // @[Top.scala 1018:12]
  assign n851_I_5_0_1 = n844_O_5_0_1; // @[Top.scala 1018:12]
  assign n851_I_5_0_2 = n844_O_5_0_2; // @[Top.scala 1018:12]
  assign n851_I_6_0_0 = n844_O_6_0_0; // @[Top.scala 1018:12]
  assign n851_I_6_0_1 = n844_O_6_0_1; // @[Top.scala 1018:12]
  assign n851_I_6_0_2 = n844_O_6_0_2; // @[Top.scala 1018:12]
  assign n851_I_7_0_0 = n844_O_7_0_0; // @[Top.scala 1018:12]
  assign n851_I_7_0_1 = n844_O_7_0_1; // @[Top.scala 1018:12]
  assign n851_I_7_0_2 = n844_O_7_0_2; // @[Top.scala 1018:12]
  assign n852_clock = clock;
  assign n852_valid_up = n824_valid_down; // @[Top.scala 1022:19]
  assign n852_I_0 = n824_O_0; // @[Top.scala 1021:12]
  assign n852_I_1 = n824_O_1; // @[Top.scala 1021:12]
  assign n852_I_2 = n824_O_2; // @[Top.scala 1021:12]
  assign n852_I_3 = n824_O_3; // @[Top.scala 1021:12]
  assign n852_I_4 = n824_O_4; // @[Top.scala 1021:12]
  assign n852_I_5 = n824_O_5; // @[Top.scala 1021:12]
  assign n852_I_6 = n824_O_6; // @[Top.scala 1021:12]
  assign n852_I_7 = n824_O_7; // @[Top.scala 1021:12]
  assign n853_clock = clock;
  assign n853_valid_up = n852_valid_down; // @[Top.scala 1025:19]
  assign n853_I_0 = n852_O_0; // @[Top.scala 1024:12]
  assign n853_I_1 = n852_O_1; // @[Top.scala 1024:12]
  assign n853_I_2 = n852_O_2; // @[Top.scala 1024:12]
  assign n853_I_3 = n852_O_3; // @[Top.scala 1024:12]
  assign n853_I_4 = n852_O_4; // @[Top.scala 1024:12]
  assign n853_I_5 = n852_O_5; // @[Top.scala 1024:12]
  assign n853_I_6 = n852_O_6; // @[Top.scala 1024:12]
  assign n853_I_7 = n852_O_7; // @[Top.scala 1024:12]
  assign n854_valid_up = n853_valid_down & n852_valid_down; // @[Top.scala 1029:19]
  assign n854_I0_0 = n853_O_0; // @[Top.scala 1027:13]
  assign n854_I0_1 = n853_O_1; // @[Top.scala 1027:13]
  assign n854_I0_2 = n853_O_2; // @[Top.scala 1027:13]
  assign n854_I0_3 = n853_O_3; // @[Top.scala 1027:13]
  assign n854_I0_4 = n853_O_4; // @[Top.scala 1027:13]
  assign n854_I0_5 = n853_O_5; // @[Top.scala 1027:13]
  assign n854_I0_6 = n853_O_6; // @[Top.scala 1027:13]
  assign n854_I0_7 = n853_O_7; // @[Top.scala 1027:13]
  assign n854_I1_0 = n852_O_0; // @[Top.scala 1028:13]
  assign n854_I1_1 = n852_O_1; // @[Top.scala 1028:13]
  assign n854_I1_2 = n852_O_2; // @[Top.scala 1028:13]
  assign n854_I1_3 = n852_O_3; // @[Top.scala 1028:13]
  assign n854_I1_4 = n852_O_4; // @[Top.scala 1028:13]
  assign n854_I1_5 = n852_O_5; // @[Top.scala 1028:13]
  assign n854_I1_6 = n852_O_6; // @[Top.scala 1028:13]
  assign n854_I1_7 = n852_O_7; // @[Top.scala 1028:13]
  assign n861_valid_up = n854_valid_down & n824_valid_down; // @[Top.scala 1033:19]
  assign n861_I0_0_0 = n854_O_0_0; // @[Top.scala 1031:13]
  assign n861_I0_0_1 = n854_O_0_1; // @[Top.scala 1031:13]
  assign n861_I0_1_0 = n854_O_1_0; // @[Top.scala 1031:13]
  assign n861_I0_1_1 = n854_O_1_1; // @[Top.scala 1031:13]
  assign n861_I0_2_0 = n854_O_2_0; // @[Top.scala 1031:13]
  assign n861_I0_2_1 = n854_O_2_1; // @[Top.scala 1031:13]
  assign n861_I0_3_0 = n854_O_3_0; // @[Top.scala 1031:13]
  assign n861_I0_3_1 = n854_O_3_1; // @[Top.scala 1031:13]
  assign n861_I0_4_0 = n854_O_4_0; // @[Top.scala 1031:13]
  assign n861_I0_4_1 = n854_O_4_1; // @[Top.scala 1031:13]
  assign n861_I0_5_0 = n854_O_5_0; // @[Top.scala 1031:13]
  assign n861_I0_5_1 = n854_O_5_1; // @[Top.scala 1031:13]
  assign n861_I0_6_0 = n854_O_6_0; // @[Top.scala 1031:13]
  assign n861_I0_6_1 = n854_O_6_1; // @[Top.scala 1031:13]
  assign n861_I0_7_0 = n854_O_7_0; // @[Top.scala 1031:13]
  assign n861_I0_7_1 = n854_O_7_1; // @[Top.scala 1031:13]
  assign n861_I1_0 = n824_O_0; // @[Top.scala 1032:13]
  assign n861_I1_1 = n824_O_1; // @[Top.scala 1032:13]
  assign n861_I1_2 = n824_O_2; // @[Top.scala 1032:13]
  assign n861_I1_3 = n824_O_3; // @[Top.scala 1032:13]
  assign n861_I1_4 = n824_O_4; // @[Top.scala 1032:13]
  assign n861_I1_5 = n824_O_5; // @[Top.scala 1032:13]
  assign n861_I1_6 = n824_O_6; // @[Top.scala 1032:13]
  assign n861_I1_7 = n824_O_7; // @[Top.scala 1032:13]
  assign n870_valid_up = n861_valid_down; // @[Top.scala 1036:19]
  assign n870_I_0_0 = n861_O_0_0; // @[Top.scala 1035:12]
  assign n870_I_0_1 = n861_O_0_1; // @[Top.scala 1035:12]
  assign n870_I_0_2 = n861_O_0_2; // @[Top.scala 1035:12]
  assign n870_I_1_0 = n861_O_1_0; // @[Top.scala 1035:12]
  assign n870_I_1_1 = n861_O_1_1; // @[Top.scala 1035:12]
  assign n870_I_1_2 = n861_O_1_2; // @[Top.scala 1035:12]
  assign n870_I_2_0 = n861_O_2_0; // @[Top.scala 1035:12]
  assign n870_I_2_1 = n861_O_2_1; // @[Top.scala 1035:12]
  assign n870_I_2_2 = n861_O_2_2; // @[Top.scala 1035:12]
  assign n870_I_3_0 = n861_O_3_0; // @[Top.scala 1035:12]
  assign n870_I_3_1 = n861_O_3_1; // @[Top.scala 1035:12]
  assign n870_I_3_2 = n861_O_3_2; // @[Top.scala 1035:12]
  assign n870_I_4_0 = n861_O_4_0; // @[Top.scala 1035:12]
  assign n870_I_4_1 = n861_O_4_1; // @[Top.scala 1035:12]
  assign n870_I_4_2 = n861_O_4_2; // @[Top.scala 1035:12]
  assign n870_I_5_0 = n861_O_5_0; // @[Top.scala 1035:12]
  assign n870_I_5_1 = n861_O_5_1; // @[Top.scala 1035:12]
  assign n870_I_5_2 = n861_O_5_2; // @[Top.scala 1035:12]
  assign n870_I_6_0 = n861_O_6_0; // @[Top.scala 1035:12]
  assign n870_I_6_1 = n861_O_6_1; // @[Top.scala 1035:12]
  assign n870_I_6_2 = n861_O_6_2; // @[Top.scala 1035:12]
  assign n870_I_7_0 = n861_O_7_0; // @[Top.scala 1035:12]
  assign n870_I_7_1 = n861_O_7_1; // @[Top.scala 1035:12]
  assign n870_I_7_2 = n861_O_7_2; // @[Top.scala 1035:12]
  assign n877_valid_up = n870_valid_down; // @[Top.scala 1039:19]
  assign n877_I_0_0_0 = n870_O_0_0_0; // @[Top.scala 1038:12]
  assign n877_I_0_0_1 = n870_O_0_0_1; // @[Top.scala 1038:12]
  assign n877_I_0_0_2 = n870_O_0_0_2; // @[Top.scala 1038:12]
  assign n877_I_1_0_0 = n870_O_1_0_0; // @[Top.scala 1038:12]
  assign n877_I_1_0_1 = n870_O_1_0_1; // @[Top.scala 1038:12]
  assign n877_I_1_0_2 = n870_O_1_0_2; // @[Top.scala 1038:12]
  assign n877_I_2_0_0 = n870_O_2_0_0; // @[Top.scala 1038:12]
  assign n877_I_2_0_1 = n870_O_2_0_1; // @[Top.scala 1038:12]
  assign n877_I_2_0_2 = n870_O_2_0_2; // @[Top.scala 1038:12]
  assign n877_I_3_0_0 = n870_O_3_0_0; // @[Top.scala 1038:12]
  assign n877_I_3_0_1 = n870_O_3_0_1; // @[Top.scala 1038:12]
  assign n877_I_3_0_2 = n870_O_3_0_2; // @[Top.scala 1038:12]
  assign n877_I_4_0_0 = n870_O_4_0_0; // @[Top.scala 1038:12]
  assign n877_I_4_0_1 = n870_O_4_0_1; // @[Top.scala 1038:12]
  assign n877_I_4_0_2 = n870_O_4_0_2; // @[Top.scala 1038:12]
  assign n877_I_5_0_0 = n870_O_5_0_0; // @[Top.scala 1038:12]
  assign n877_I_5_0_1 = n870_O_5_0_1; // @[Top.scala 1038:12]
  assign n877_I_5_0_2 = n870_O_5_0_2; // @[Top.scala 1038:12]
  assign n877_I_6_0_0 = n870_O_6_0_0; // @[Top.scala 1038:12]
  assign n877_I_6_0_1 = n870_O_6_0_1; // @[Top.scala 1038:12]
  assign n877_I_6_0_2 = n870_O_6_0_2; // @[Top.scala 1038:12]
  assign n877_I_7_0_0 = n870_O_7_0_0; // @[Top.scala 1038:12]
  assign n877_I_7_0_1 = n870_O_7_0_1; // @[Top.scala 1038:12]
  assign n877_I_7_0_2 = n870_O_7_0_2; // @[Top.scala 1038:12]
  assign n878_valid_up = n851_valid_down & n877_valid_down; // @[Top.scala 1043:19]
  assign n878_I0_0_0 = n851_O_0_0; // @[Top.scala 1041:13]
  assign n878_I0_0_1 = n851_O_0_1; // @[Top.scala 1041:13]
  assign n878_I0_0_2 = n851_O_0_2; // @[Top.scala 1041:13]
  assign n878_I0_1_0 = n851_O_1_0; // @[Top.scala 1041:13]
  assign n878_I0_1_1 = n851_O_1_1; // @[Top.scala 1041:13]
  assign n878_I0_1_2 = n851_O_1_2; // @[Top.scala 1041:13]
  assign n878_I0_2_0 = n851_O_2_0; // @[Top.scala 1041:13]
  assign n878_I0_2_1 = n851_O_2_1; // @[Top.scala 1041:13]
  assign n878_I0_2_2 = n851_O_2_2; // @[Top.scala 1041:13]
  assign n878_I0_3_0 = n851_O_3_0; // @[Top.scala 1041:13]
  assign n878_I0_3_1 = n851_O_3_1; // @[Top.scala 1041:13]
  assign n878_I0_3_2 = n851_O_3_2; // @[Top.scala 1041:13]
  assign n878_I0_4_0 = n851_O_4_0; // @[Top.scala 1041:13]
  assign n878_I0_4_1 = n851_O_4_1; // @[Top.scala 1041:13]
  assign n878_I0_4_2 = n851_O_4_2; // @[Top.scala 1041:13]
  assign n878_I0_5_0 = n851_O_5_0; // @[Top.scala 1041:13]
  assign n878_I0_5_1 = n851_O_5_1; // @[Top.scala 1041:13]
  assign n878_I0_5_2 = n851_O_5_2; // @[Top.scala 1041:13]
  assign n878_I0_6_0 = n851_O_6_0; // @[Top.scala 1041:13]
  assign n878_I0_6_1 = n851_O_6_1; // @[Top.scala 1041:13]
  assign n878_I0_6_2 = n851_O_6_2; // @[Top.scala 1041:13]
  assign n878_I0_7_0 = n851_O_7_0; // @[Top.scala 1041:13]
  assign n878_I0_7_1 = n851_O_7_1; // @[Top.scala 1041:13]
  assign n878_I0_7_2 = n851_O_7_2; // @[Top.scala 1041:13]
  assign n878_I1_0_0 = n877_O_0_0; // @[Top.scala 1042:13]
  assign n878_I1_0_1 = n877_O_0_1; // @[Top.scala 1042:13]
  assign n878_I1_0_2 = n877_O_0_2; // @[Top.scala 1042:13]
  assign n878_I1_1_0 = n877_O_1_0; // @[Top.scala 1042:13]
  assign n878_I1_1_1 = n877_O_1_1; // @[Top.scala 1042:13]
  assign n878_I1_1_2 = n877_O_1_2; // @[Top.scala 1042:13]
  assign n878_I1_2_0 = n877_O_2_0; // @[Top.scala 1042:13]
  assign n878_I1_2_1 = n877_O_2_1; // @[Top.scala 1042:13]
  assign n878_I1_2_2 = n877_O_2_2; // @[Top.scala 1042:13]
  assign n878_I1_3_0 = n877_O_3_0; // @[Top.scala 1042:13]
  assign n878_I1_3_1 = n877_O_3_1; // @[Top.scala 1042:13]
  assign n878_I1_3_2 = n877_O_3_2; // @[Top.scala 1042:13]
  assign n878_I1_4_0 = n877_O_4_0; // @[Top.scala 1042:13]
  assign n878_I1_4_1 = n877_O_4_1; // @[Top.scala 1042:13]
  assign n878_I1_4_2 = n877_O_4_2; // @[Top.scala 1042:13]
  assign n878_I1_5_0 = n877_O_5_0; // @[Top.scala 1042:13]
  assign n878_I1_5_1 = n877_O_5_1; // @[Top.scala 1042:13]
  assign n878_I1_5_2 = n877_O_5_2; // @[Top.scala 1042:13]
  assign n878_I1_6_0 = n877_O_6_0; // @[Top.scala 1042:13]
  assign n878_I1_6_1 = n877_O_6_1; // @[Top.scala 1042:13]
  assign n878_I1_6_2 = n877_O_6_2; // @[Top.scala 1042:13]
  assign n878_I1_7_0 = n877_O_7_0; // @[Top.scala 1042:13]
  assign n878_I1_7_1 = n877_O_7_1; // @[Top.scala 1042:13]
  assign n878_I1_7_2 = n877_O_7_2; // @[Top.scala 1042:13]
  assign n885_clock = clock;
  assign n885_valid_up = n823_valid_down; // @[Top.scala 1046:19]
  assign n885_I_0 = n823_O_0; // @[Top.scala 1045:12]
  assign n885_I_1 = n823_O_1; // @[Top.scala 1045:12]
  assign n885_I_2 = n823_O_2; // @[Top.scala 1045:12]
  assign n885_I_3 = n823_O_3; // @[Top.scala 1045:12]
  assign n885_I_4 = n823_O_4; // @[Top.scala 1045:12]
  assign n885_I_5 = n823_O_5; // @[Top.scala 1045:12]
  assign n885_I_6 = n823_O_6; // @[Top.scala 1045:12]
  assign n885_I_7 = n823_O_7; // @[Top.scala 1045:12]
  assign n886_clock = clock;
  assign n886_valid_up = n885_valid_down; // @[Top.scala 1049:19]
  assign n886_I_0 = n885_O_0; // @[Top.scala 1048:12]
  assign n886_I_1 = n885_O_1; // @[Top.scala 1048:12]
  assign n886_I_2 = n885_O_2; // @[Top.scala 1048:12]
  assign n886_I_3 = n885_O_3; // @[Top.scala 1048:12]
  assign n886_I_4 = n885_O_4; // @[Top.scala 1048:12]
  assign n886_I_5 = n885_O_5; // @[Top.scala 1048:12]
  assign n886_I_6 = n885_O_6; // @[Top.scala 1048:12]
  assign n886_I_7 = n885_O_7; // @[Top.scala 1048:12]
  assign n887_valid_up = n886_valid_down & n885_valid_down; // @[Top.scala 1053:19]
  assign n887_I0_0 = n886_O_0; // @[Top.scala 1051:13]
  assign n887_I0_1 = n886_O_1; // @[Top.scala 1051:13]
  assign n887_I0_2 = n886_O_2; // @[Top.scala 1051:13]
  assign n887_I0_3 = n886_O_3; // @[Top.scala 1051:13]
  assign n887_I0_4 = n886_O_4; // @[Top.scala 1051:13]
  assign n887_I0_5 = n886_O_5; // @[Top.scala 1051:13]
  assign n887_I0_6 = n886_O_6; // @[Top.scala 1051:13]
  assign n887_I0_7 = n886_O_7; // @[Top.scala 1051:13]
  assign n887_I1_0 = n885_O_0; // @[Top.scala 1052:13]
  assign n887_I1_1 = n885_O_1; // @[Top.scala 1052:13]
  assign n887_I1_2 = n885_O_2; // @[Top.scala 1052:13]
  assign n887_I1_3 = n885_O_3; // @[Top.scala 1052:13]
  assign n887_I1_4 = n885_O_4; // @[Top.scala 1052:13]
  assign n887_I1_5 = n885_O_5; // @[Top.scala 1052:13]
  assign n887_I1_6 = n885_O_6; // @[Top.scala 1052:13]
  assign n887_I1_7 = n885_O_7; // @[Top.scala 1052:13]
  assign n894_valid_up = n887_valid_down & n823_valid_down; // @[Top.scala 1057:19]
  assign n894_I0_0_0 = n887_O_0_0; // @[Top.scala 1055:13]
  assign n894_I0_0_1 = n887_O_0_1; // @[Top.scala 1055:13]
  assign n894_I0_1_0 = n887_O_1_0; // @[Top.scala 1055:13]
  assign n894_I0_1_1 = n887_O_1_1; // @[Top.scala 1055:13]
  assign n894_I0_2_0 = n887_O_2_0; // @[Top.scala 1055:13]
  assign n894_I0_2_1 = n887_O_2_1; // @[Top.scala 1055:13]
  assign n894_I0_3_0 = n887_O_3_0; // @[Top.scala 1055:13]
  assign n894_I0_3_1 = n887_O_3_1; // @[Top.scala 1055:13]
  assign n894_I0_4_0 = n887_O_4_0; // @[Top.scala 1055:13]
  assign n894_I0_4_1 = n887_O_4_1; // @[Top.scala 1055:13]
  assign n894_I0_5_0 = n887_O_5_0; // @[Top.scala 1055:13]
  assign n894_I0_5_1 = n887_O_5_1; // @[Top.scala 1055:13]
  assign n894_I0_6_0 = n887_O_6_0; // @[Top.scala 1055:13]
  assign n894_I0_6_1 = n887_O_6_1; // @[Top.scala 1055:13]
  assign n894_I0_7_0 = n887_O_7_0; // @[Top.scala 1055:13]
  assign n894_I0_7_1 = n887_O_7_1; // @[Top.scala 1055:13]
  assign n894_I1_0 = n823_O_0; // @[Top.scala 1056:13]
  assign n894_I1_1 = n823_O_1; // @[Top.scala 1056:13]
  assign n894_I1_2 = n823_O_2; // @[Top.scala 1056:13]
  assign n894_I1_3 = n823_O_3; // @[Top.scala 1056:13]
  assign n894_I1_4 = n823_O_4; // @[Top.scala 1056:13]
  assign n894_I1_5 = n823_O_5; // @[Top.scala 1056:13]
  assign n894_I1_6 = n823_O_6; // @[Top.scala 1056:13]
  assign n894_I1_7 = n823_O_7; // @[Top.scala 1056:13]
  assign n903_valid_up = n894_valid_down; // @[Top.scala 1060:19]
  assign n903_I_0_0 = n894_O_0_0; // @[Top.scala 1059:12]
  assign n903_I_0_1 = n894_O_0_1; // @[Top.scala 1059:12]
  assign n903_I_0_2 = n894_O_0_2; // @[Top.scala 1059:12]
  assign n903_I_1_0 = n894_O_1_0; // @[Top.scala 1059:12]
  assign n903_I_1_1 = n894_O_1_1; // @[Top.scala 1059:12]
  assign n903_I_1_2 = n894_O_1_2; // @[Top.scala 1059:12]
  assign n903_I_2_0 = n894_O_2_0; // @[Top.scala 1059:12]
  assign n903_I_2_1 = n894_O_2_1; // @[Top.scala 1059:12]
  assign n903_I_2_2 = n894_O_2_2; // @[Top.scala 1059:12]
  assign n903_I_3_0 = n894_O_3_0; // @[Top.scala 1059:12]
  assign n903_I_3_1 = n894_O_3_1; // @[Top.scala 1059:12]
  assign n903_I_3_2 = n894_O_3_2; // @[Top.scala 1059:12]
  assign n903_I_4_0 = n894_O_4_0; // @[Top.scala 1059:12]
  assign n903_I_4_1 = n894_O_4_1; // @[Top.scala 1059:12]
  assign n903_I_4_2 = n894_O_4_2; // @[Top.scala 1059:12]
  assign n903_I_5_0 = n894_O_5_0; // @[Top.scala 1059:12]
  assign n903_I_5_1 = n894_O_5_1; // @[Top.scala 1059:12]
  assign n903_I_5_2 = n894_O_5_2; // @[Top.scala 1059:12]
  assign n903_I_6_0 = n894_O_6_0; // @[Top.scala 1059:12]
  assign n903_I_6_1 = n894_O_6_1; // @[Top.scala 1059:12]
  assign n903_I_6_2 = n894_O_6_2; // @[Top.scala 1059:12]
  assign n903_I_7_0 = n894_O_7_0; // @[Top.scala 1059:12]
  assign n903_I_7_1 = n894_O_7_1; // @[Top.scala 1059:12]
  assign n903_I_7_2 = n894_O_7_2; // @[Top.scala 1059:12]
  assign n910_valid_up = n903_valid_down; // @[Top.scala 1063:19]
  assign n910_I_0_0_0 = n903_O_0_0_0; // @[Top.scala 1062:12]
  assign n910_I_0_0_1 = n903_O_0_0_1; // @[Top.scala 1062:12]
  assign n910_I_0_0_2 = n903_O_0_0_2; // @[Top.scala 1062:12]
  assign n910_I_1_0_0 = n903_O_1_0_0; // @[Top.scala 1062:12]
  assign n910_I_1_0_1 = n903_O_1_0_1; // @[Top.scala 1062:12]
  assign n910_I_1_0_2 = n903_O_1_0_2; // @[Top.scala 1062:12]
  assign n910_I_2_0_0 = n903_O_2_0_0; // @[Top.scala 1062:12]
  assign n910_I_2_0_1 = n903_O_2_0_1; // @[Top.scala 1062:12]
  assign n910_I_2_0_2 = n903_O_2_0_2; // @[Top.scala 1062:12]
  assign n910_I_3_0_0 = n903_O_3_0_0; // @[Top.scala 1062:12]
  assign n910_I_3_0_1 = n903_O_3_0_1; // @[Top.scala 1062:12]
  assign n910_I_3_0_2 = n903_O_3_0_2; // @[Top.scala 1062:12]
  assign n910_I_4_0_0 = n903_O_4_0_0; // @[Top.scala 1062:12]
  assign n910_I_4_0_1 = n903_O_4_0_1; // @[Top.scala 1062:12]
  assign n910_I_4_0_2 = n903_O_4_0_2; // @[Top.scala 1062:12]
  assign n910_I_5_0_0 = n903_O_5_0_0; // @[Top.scala 1062:12]
  assign n910_I_5_0_1 = n903_O_5_0_1; // @[Top.scala 1062:12]
  assign n910_I_5_0_2 = n903_O_5_0_2; // @[Top.scala 1062:12]
  assign n910_I_6_0_0 = n903_O_6_0_0; // @[Top.scala 1062:12]
  assign n910_I_6_0_1 = n903_O_6_0_1; // @[Top.scala 1062:12]
  assign n910_I_6_0_2 = n903_O_6_0_2; // @[Top.scala 1062:12]
  assign n910_I_7_0_0 = n903_O_7_0_0; // @[Top.scala 1062:12]
  assign n910_I_7_0_1 = n903_O_7_0_1; // @[Top.scala 1062:12]
  assign n910_I_7_0_2 = n903_O_7_0_2; // @[Top.scala 1062:12]
  assign n911_valid_up = n878_valid_down & n910_valid_down; // @[Top.scala 1067:19]
  assign n911_I0_0_0_0 = n878_O_0_0_0; // @[Top.scala 1065:13]
  assign n911_I0_0_0_1 = n878_O_0_0_1; // @[Top.scala 1065:13]
  assign n911_I0_0_0_2 = n878_O_0_0_2; // @[Top.scala 1065:13]
  assign n911_I0_0_1_0 = n878_O_0_1_0; // @[Top.scala 1065:13]
  assign n911_I0_0_1_1 = n878_O_0_1_1; // @[Top.scala 1065:13]
  assign n911_I0_0_1_2 = n878_O_0_1_2; // @[Top.scala 1065:13]
  assign n911_I0_1_0_0 = n878_O_1_0_0; // @[Top.scala 1065:13]
  assign n911_I0_1_0_1 = n878_O_1_0_1; // @[Top.scala 1065:13]
  assign n911_I0_1_0_2 = n878_O_1_0_2; // @[Top.scala 1065:13]
  assign n911_I0_1_1_0 = n878_O_1_1_0; // @[Top.scala 1065:13]
  assign n911_I0_1_1_1 = n878_O_1_1_1; // @[Top.scala 1065:13]
  assign n911_I0_1_1_2 = n878_O_1_1_2; // @[Top.scala 1065:13]
  assign n911_I0_2_0_0 = n878_O_2_0_0; // @[Top.scala 1065:13]
  assign n911_I0_2_0_1 = n878_O_2_0_1; // @[Top.scala 1065:13]
  assign n911_I0_2_0_2 = n878_O_2_0_2; // @[Top.scala 1065:13]
  assign n911_I0_2_1_0 = n878_O_2_1_0; // @[Top.scala 1065:13]
  assign n911_I0_2_1_1 = n878_O_2_1_1; // @[Top.scala 1065:13]
  assign n911_I0_2_1_2 = n878_O_2_1_2; // @[Top.scala 1065:13]
  assign n911_I0_3_0_0 = n878_O_3_0_0; // @[Top.scala 1065:13]
  assign n911_I0_3_0_1 = n878_O_3_0_1; // @[Top.scala 1065:13]
  assign n911_I0_3_0_2 = n878_O_3_0_2; // @[Top.scala 1065:13]
  assign n911_I0_3_1_0 = n878_O_3_1_0; // @[Top.scala 1065:13]
  assign n911_I0_3_1_1 = n878_O_3_1_1; // @[Top.scala 1065:13]
  assign n911_I0_3_1_2 = n878_O_3_1_2; // @[Top.scala 1065:13]
  assign n911_I0_4_0_0 = n878_O_4_0_0; // @[Top.scala 1065:13]
  assign n911_I0_4_0_1 = n878_O_4_0_1; // @[Top.scala 1065:13]
  assign n911_I0_4_0_2 = n878_O_4_0_2; // @[Top.scala 1065:13]
  assign n911_I0_4_1_0 = n878_O_4_1_0; // @[Top.scala 1065:13]
  assign n911_I0_4_1_1 = n878_O_4_1_1; // @[Top.scala 1065:13]
  assign n911_I0_4_1_2 = n878_O_4_1_2; // @[Top.scala 1065:13]
  assign n911_I0_5_0_0 = n878_O_5_0_0; // @[Top.scala 1065:13]
  assign n911_I0_5_0_1 = n878_O_5_0_1; // @[Top.scala 1065:13]
  assign n911_I0_5_0_2 = n878_O_5_0_2; // @[Top.scala 1065:13]
  assign n911_I0_5_1_0 = n878_O_5_1_0; // @[Top.scala 1065:13]
  assign n911_I0_5_1_1 = n878_O_5_1_1; // @[Top.scala 1065:13]
  assign n911_I0_5_1_2 = n878_O_5_1_2; // @[Top.scala 1065:13]
  assign n911_I0_6_0_0 = n878_O_6_0_0; // @[Top.scala 1065:13]
  assign n911_I0_6_0_1 = n878_O_6_0_1; // @[Top.scala 1065:13]
  assign n911_I0_6_0_2 = n878_O_6_0_2; // @[Top.scala 1065:13]
  assign n911_I0_6_1_0 = n878_O_6_1_0; // @[Top.scala 1065:13]
  assign n911_I0_6_1_1 = n878_O_6_1_1; // @[Top.scala 1065:13]
  assign n911_I0_6_1_2 = n878_O_6_1_2; // @[Top.scala 1065:13]
  assign n911_I0_7_0_0 = n878_O_7_0_0; // @[Top.scala 1065:13]
  assign n911_I0_7_0_1 = n878_O_7_0_1; // @[Top.scala 1065:13]
  assign n911_I0_7_0_2 = n878_O_7_0_2; // @[Top.scala 1065:13]
  assign n911_I0_7_1_0 = n878_O_7_1_0; // @[Top.scala 1065:13]
  assign n911_I0_7_1_1 = n878_O_7_1_1; // @[Top.scala 1065:13]
  assign n911_I0_7_1_2 = n878_O_7_1_2; // @[Top.scala 1065:13]
  assign n911_I1_0_0 = n910_O_0_0; // @[Top.scala 1066:13]
  assign n911_I1_0_1 = n910_O_0_1; // @[Top.scala 1066:13]
  assign n911_I1_0_2 = n910_O_0_2; // @[Top.scala 1066:13]
  assign n911_I1_1_0 = n910_O_1_0; // @[Top.scala 1066:13]
  assign n911_I1_1_1 = n910_O_1_1; // @[Top.scala 1066:13]
  assign n911_I1_1_2 = n910_O_1_2; // @[Top.scala 1066:13]
  assign n911_I1_2_0 = n910_O_2_0; // @[Top.scala 1066:13]
  assign n911_I1_2_1 = n910_O_2_1; // @[Top.scala 1066:13]
  assign n911_I1_2_2 = n910_O_2_2; // @[Top.scala 1066:13]
  assign n911_I1_3_0 = n910_O_3_0; // @[Top.scala 1066:13]
  assign n911_I1_3_1 = n910_O_3_1; // @[Top.scala 1066:13]
  assign n911_I1_3_2 = n910_O_3_2; // @[Top.scala 1066:13]
  assign n911_I1_4_0 = n910_O_4_0; // @[Top.scala 1066:13]
  assign n911_I1_4_1 = n910_O_4_1; // @[Top.scala 1066:13]
  assign n911_I1_4_2 = n910_O_4_2; // @[Top.scala 1066:13]
  assign n911_I1_5_0 = n910_O_5_0; // @[Top.scala 1066:13]
  assign n911_I1_5_1 = n910_O_5_1; // @[Top.scala 1066:13]
  assign n911_I1_5_2 = n910_O_5_2; // @[Top.scala 1066:13]
  assign n911_I1_6_0 = n910_O_6_0; // @[Top.scala 1066:13]
  assign n911_I1_6_1 = n910_O_6_1; // @[Top.scala 1066:13]
  assign n911_I1_6_2 = n910_O_6_2; // @[Top.scala 1066:13]
  assign n911_I1_7_0 = n910_O_7_0; // @[Top.scala 1066:13]
  assign n911_I1_7_1 = n910_O_7_1; // @[Top.scala 1066:13]
  assign n911_I1_7_2 = n910_O_7_2; // @[Top.scala 1066:13]
  assign n920_valid_up = n911_valid_down; // @[Top.scala 1070:19]
  assign n920_I_0_0_0 = n911_O_0_0_0; // @[Top.scala 1069:12]
  assign n920_I_0_0_1 = n911_O_0_0_1; // @[Top.scala 1069:12]
  assign n920_I_0_0_2 = n911_O_0_0_2; // @[Top.scala 1069:12]
  assign n920_I_0_1_0 = n911_O_0_1_0; // @[Top.scala 1069:12]
  assign n920_I_0_1_1 = n911_O_0_1_1; // @[Top.scala 1069:12]
  assign n920_I_0_1_2 = n911_O_0_1_2; // @[Top.scala 1069:12]
  assign n920_I_0_2_0 = n911_O_0_2_0; // @[Top.scala 1069:12]
  assign n920_I_0_2_1 = n911_O_0_2_1; // @[Top.scala 1069:12]
  assign n920_I_0_2_2 = n911_O_0_2_2; // @[Top.scala 1069:12]
  assign n920_I_1_0_0 = n911_O_1_0_0; // @[Top.scala 1069:12]
  assign n920_I_1_0_1 = n911_O_1_0_1; // @[Top.scala 1069:12]
  assign n920_I_1_0_2 = n911_O_1_0_2; // @[Top.scala 1069:12]
  assign n920_I_1_1_0 = n911_O_1_1_0; // @[Top.scala 1069:12]
  assign n920_I_1_1_1 = n911_O_1_1_1; // @[Top.scala 1069:12]
  assign n920_I_1_1_2 = n911_O_1_1_2; // @[Top.scala 1069:12]
  assign n920_I_1_2_0 = n911_O_1_2_0; // @[Top.scala 1069:12]
  assign n920_I_1_2_1 = n911_O_1_2_1; // @[Top.scala 1069:12]
  assign n920_I_1_2_2 = n911_O_1_2_2; // @[Top.scala 1069:12]
  assign n920_I_2_0_0 = n911_O_2_0_0; // @[Top.scala 1069:12]
  assign n920_I_2_0_1 = n911_O_2_0_1; // @[Top.scala 1069:12]
  assign n920_I_2_0_2 = n911_O_2_0_2; // @[Top.scala 1069:12]
  assign n920_I_2_1_0 = n911_O_2_1_0; // @[Top.scala 1069:12]
  assign n920_I_2_1_1 = n911_O_2_1_1; // @[Top.scala 1069:12]
  assign n920_I_2_1_2 = n911_O_2_1_2; // @[Top.scala 1069:12]
  assign n920_I_2_2_0 = n911_O_2_2_0; // @[Top.scala 1069:12]
  assign n920_I_2_2_1 = n911_O_2_2_1; // @[Top.scala 1069:12]
  assign n920_I_2_2_2 = n911_O_2_2_2; // @[Top.scala 1069:12]
  assign n920_I_3_0_0 = n911_O_3_0_0; // @[Top.scala 1069:12]
  assign n920_I_3_0_1 = n911_O_3_0_1; // @[Top.scala 1069:12]
  assign n920_I_3_0_2 = n911_O_3_0_2; // @[Top.scala 1069:12]
  assign n920_I_3_1_0 = n911_O_3_1_0; // @[Top.scala 1069:12]
  assign n920_I_3_1_1 = n911_O_3_1_1; // @[Top.scala 1069:12]
  assign n920_I_3_1_2 = n911_O_3_1_2; // @[Top.scala 1069:12]
  assign n920_I_3_2_0 = n911_O_3_2_0; // @[Top.scala 1069:12]
  assign n920_I_3_2_1 = n911_O_3_2_1; // @[Top.scala 1069:12]
  assign n920_I_3_2_2 = n911_O_3_2_2; // @[Top.scala 1069:12]
  assign n920_I_4_0_0 = n911_O_4_0_0; // @[Top.scala 1069:12]
  assign n920_I_4_0_1 = n911_O_4_0_1; // @[Top.scala 1069:12]
  assign n920_I_4_0_2 = n911_O_4_0_2; // @[Top.scala 1069:12]
  assign n920_I_4_1_0 = n911_O_4_1_0; // @[Top.scala 1069:12]
  assign n920_I_4_1_1 = n911_O_4_1_1; // @[Top.scala 1069:12]
  assign n920_I_4_1_2 = n911_O_4_1_2; // @[Top.scala 1069:12]
  assign n920_I_4_2_0 = n911_O_4_2_0; // @[Top.scala 1069:12]
  assign n920_I_4_2_1 = n911_O_4_2_1; // @[Top.scala 1069:12]
  assign n920_I_4_2_2 = n911_O_4_2_2; // @[Top.scala 1069:12]
  assign n920_I_5_0_0 = n911_O_5_0_0; // @[Top.scala 1069:12]
  assign n920_I_5_0_1 = n911_O_5_0_1; // @[Top.scala 1069:12]
  assign n920_I_5_0_2 = n911_O_5_0_2; // @[Top.scala 1069:12]
  assign n920_I_5_1_0 = n911_O_5_1_0; // @[Top.scala 1069:12]
  assign n920_I_5_1_1 = n911_O_5_1_1; // @[Top.scala 1069:12]
  assign n920_I_5_1_2 = n911_O_5_1_2; // @[Top.scala 1069:12]
  assign n920_I_5_2_0 = n911_O_5_2_0; // @[Top.scala 1069:12]
  assign n920_I_5_2_1 = n911_O_5_2_1; // @[Top.scala 1069:12]
  assign n920_I_5_2_2 = n911_O_5_2_2; // @[Top.scala 1069:12]
  assign n920_I_6_0_0 = n911_O_6_0_0; // @[Top.scala 1069:12]
  assign n920_I_6_0_1 = n911_O_6_0_1; // @[Top.scala 1069:12]
  assign n920_I_6_0_2 = n911_O_6_0_2; // @[Top.scala 1069:12]
  assign n920_I_6_1_0 = n911_O_6_1_0; // @[Top.scala 1069:12]
  assign n920_I_6_1_1 = n911_O_6_1_1; // @[Top.scala 1069:12]
  assign n920_I_6_1_2 = n911_O_6_1_2; // @[Top.scala 1069:12]
  assign n920_I_6_2_0 = n911_O_6_2_0; // @[Top.scala 1069:12]
  assign n920_I_6_2_1 = n911_O_6_2_1; // @[Top.scala 1069:12]
  assign n920_I_6_2_2 = n911_O_6_2_2; // @[Top.scala 1069:12]
  assign n920_I_7_0_0 = n911_O_7_0_0; // @[Top.scala 1069:12]
  assign n920_I_7_0_1 = n911_O_7_0_1; // @[Top.scala 1069:12]
  assign n920_I_7_0_2 = n911_O_7_0_2; // @[Top.scala 1069:12]
  assign n920_I_7_1_0 = n911_O_7_1_0; // @[Top.scala 1069:12]
  assign n920_I_7_1_1 = n911_O_7_1_1; // @[Top.scala 1069:12]
  assign n920_I_7_1_2 = n911_O_7_1_2; // @[Top.scala 1069:12]
  assign n920_I_7_2_0 = n911_O_7_2_0; // @[Top.scala 1069:12]
  assign n920_I_7_2_1 = n911_O_7_2_1; // @[Top.scala 1069:12]
  assign n920_I_7_2_2 = n911_O_7_2_2; // @[Top.scala 1069:12]
  assign n927_valid_up = n920_valid_down; // @[Top.scala 1073:19]
  assign n927_I_0_0_0_0 = n920_O_0_0_0_0; // @[Top.scala 1072:12]
  assign n927_I_0_0_0_1 = n920_O_0_0_0_1; // @[Top.scala 1072:12]
  assign n927_I_0_0_0_2 = n920_O_0_0_0_2; // @[Top.scala 1072:12]
  assign n927_I_0_0_1_0 = n920_O_0_0_1_0; // @[Top.scala 1072:12]
  assign n927_I_0_0_1_1 = n920_O_0_0_1_1; // @[Top.scala 1072:12]
  assign n927_I_0_0_1_2 = n920_O_0_0_1_2; // @[Top.scala 1072:12]
  assign n927_I_0_0_2_0 = n920_O_0_0_2_0; // @[Top.scala 1072:12]
  assign n927_I_0_0_2_1 = n920_O_0_0_2_1; // @[Top.scala 1072:12]
  assign n927_I_0_0_2_2 = n920_O_0_0_2_2; // @[Top.scala 1072:12]
  assign n927_I_1_0_0_0 = n920_O_1_0_0_0; // @[Top.scala 1072:12]
  assign n927_I_1_0_0_1 = n920_O_1_0_0_1; // @[Top.scala 1072:12]
  assign n927_I_1_0_0_2 = n920_O_1_0_0_2; // @[Top.scala 1072:12]
  assign n927_I_1_0_1_0 = n920_O_1_0_1_0; // @[Top.scala 1072:12]
  assign n927_I_1_0_1_1 = n920_O_1_0_1_1; // @[Top.scala 1072:12]
  assign n927_I_1_0_1_2 = n920_O_1_0_1_2; // @[Top.scala 1072:12]
  assign n927_I_1_0_2_0 = n920_O_1_0_2_0; // @[Top.scala 1072:12]
  assign n927_I_1_0_2_1 = n920_O_1_0_2_1; // @[Top.scala 1072:12]
  assign n927_I_1_0_2_2 = n920_O_1_0_2_2; // @[Top.scala 1072:12]
  assign n927_I_2_0_0_0 = n920_O_2_0_0_0; // @[Top.scala 1072:12]
  assign n927_I_2_0_0_1 = n920_O_2_0_0_1; // @[Top.scala 1072:12]
  assign n927_I_2_0_0_2 = n920_O_2_0_0_2; // @[Top.scala 1072:12]
  assign n927_I_2_0_1_0 = n920_O_2_0_1_0; // @[Top.scala 1072:12]
  assign n927_I_2_0_1_1 = n920_O_2_0_1_1; // @[Top.scala 1072:12]
  assign n927_I_2_0_1_2 = n920_O_2_0_1_2; // @[Top.scala 1072:12]
  assign n927_I_2_0_2_0 = n920_O_2_0_2_0; // @[Top.scala 1072:12]
  assign n927_I_2_0_2_1 = n920_O_2_0_2_1; // @[Top.scala 1072:12]
  assign n927_I_2_0_2_2 = n920_O_2_0_2_2; // @[Top.scala 1072:12]
  assign n927_I_3_0_0_0 = n920_O_3_0_0_0; // @[Top.scala 1072:12]
  assign n927_I_3_0_0_1 = n920_O_3_0_0_1; // @[Top.scala 1072:12]
  assign n927_I_3_0_0_2 = n920_O_3_0_0_2; // @[Top.scala 1072:12]
  assign n927_I_3_0_1_0 = n920_O_3_0_1_0; // @[Top.scala 1072:12]
  assign n927_I_3_0_1_1 = n920_O_3_0_1_1; // @[Top.scala 1072:12]
  assign n927_I_3_0_1_2 = n920_O_3_0_1_2; // @[Top.scala 1072:12]
  assign n927_I_3_0_2_0 = n920_O_3_0_2_0; // @[Top.scala 1072:12]
  assign n927_I_3_0_2_1 = n920_O_3_0_2_1; // @[Top.scala 1072:12]
  assign n927_I_3_0_2_2 = n920_O_3_0_2_2; // @[Top.scala 1072:12]
  assign n927_I_4_0_0_0 = n920_O_4_0_0_0; // @[Top.scala 1072:12]
  assign n927_I_4_0_0_1 = n920_O_4_0_0_1; // @[Top.scala 1072:12]
  assign n927_I_4_0_0_2 = n920_O_4_0_0_2; // @[Top.scala 1072:12]
  assign n927_I_4_0_1_0 = n920_O_4_0_1_0; // @[Top.scala 1072:12]
  assign n927_I_4_0_1_1 = n920_O_4_0_1_1; // @[Top.scala 1072:12]
  assign n927_I_4_0_1_2 = n920_O_4_0_1_2; // @[Top.scala 1072:12]
  assign n927_I_4_0_2_0 = n920_O_4_0_2_0; // @[Top.scala 1072:12]
  assign n927_I_4_0_2_1 = n920_O_4_0_2_1; // @[Top.scala 1072:12]
  assign n927_I_4_0_2_2 = n920_O_4_0_2_2; // @[Top.scala 1072:12]
  assign n927_I_5_0_0_0 = n920_O_5_0_0_0; // @[Top.scala 1072:12]
  assign n927_I_5_0_0_1 = n920_O_5_0_0_1; // @[Top.scala 1072:12]
  assign n927_I_5_0_0_2 = n920_O_5_0_0_2; // @[Top.scala 1072:12]
  assign n927_I_5_0_1_0 = n920_O_5_0_1_0; // @[Top.scala 1072:12]
  assign n927_I_5_0_1_1 = n920_O_5_0_1_1; // @[Top.scala 1072:12]
  assign n927_I_5_0_1_2 = n920_O_5_0_1_2; // @[Top.scala 1072:12]
  assign n927_I_5_0_2_0 = n920_O_5_0_2_0; // @[Top.scala 1072:12]
  assign n927_I_5_0_2_1 = n920_O_5_0_2_1; // @[Top.scala 1072:12]
  assign n927_I_5_0_2_2 = n920_O_5_0_2_2; // @[Top.scala 1072:12]
  assign n927_I_6_0_0_0 = n920_O_6_0_0_0; // @[Top.scala 1072:12]
  assign n927_I_6_0_0_1 = n920_O_6_0_0_1; // @[Top.scala 1072:12]
  assign n927_I_6_0_0_2 = n920_O_6_0_0_2; // @[Top.scala 1072:12]
  assign n927_I_6_0_1_0 = n920_O_6_0_1_0; // @[Top.scala 1072:12]
  assign n927_I_6_0_1_1 = n920_O_6_0_1_1; // @[Top.scala 1072:12]
  assign n927_I_6_0_1_2 = n920_O_6_0_1_2; // @[Top.scala 1072:12]
  assign n927_I_6_0_2_0 = n920_O_6_0_2_0; // @[Top.scala 1072:12]
  assign n927_I_6_0_2_1 = n920_O_6_0_2_1; // @[Top.scala 1072:12]
  assign n927_I_6_0_2_2 = n920_O_6_0_2_2; // @[Top.scala 1072:12]
  assign n927_I_7_0_0_0 = n920_O_7_0_0_0; // @[Top.scala 1072:12]
  assign n927_I_7_0_0_1 = n920_O_7_0_0_1; // @[Top.scala 1072:12]
  assign n927_I_7_0_0_2 = n920_O_7_0_0_2; // @[Top.scala 1072:12]
  assign n927_I_7_0_1_0 = n920_O_7_0_1_0; // @[Top.scala 1072:12]
  assign n927_I_7_0_1_1 = n920_O_7_0_1_1; // @[Top.scala 1072:12]
  assign n927_I_7_0_1_2 = n920_O_7_0_1_2; // @[Top.scala 1072:12]
  assign n927_I_7_0_2_0 = n920_O_7_0_2_0; // @[Top.scala 1072:12]
  assign n927_I_7_0_2_1 = n920_O_7_0_2_1; // @[Top.scala 1072:12]
  assign n927_I_7_0_2_2 = n920_O_7_0_2_2; // @[Top.scala 1072:12]
  assign n969_clock = clock;
  assign n969_reset = reset;
  assign n969_valid_up = n927_valid_down; // @[Top.scala 1076:19]
  assign n969_I_0_0_0 = n927_O_0_0_0; // @[Top.scala 1075:12]
  assign n969_I_0_0_1 = n927_O_0_0_1; // @[Top.scala 1075:12]
  assign n969_I_0_0_2 = n927_O_0_0_2; // @[Top.scala 1075:12]
  assign n969_I_0_1_0 = n927_O_0_1_0; // @[Top.scala 1075:12]
  assign n969_I_0_1_1 = n927_O_0_1_1; // @[Top.scala 1075:12]
  assign n969_I_0_1_2 = n927_O_0_1_2; // @[Top.scala 1075:12]
  assign n969_I_0_2_0 = n927_O_0_2_0; // @[Top.scala 1075:12]
  assign n969_I_0_2_1 = n927_O_0_2_1; // @[Top.scala 1075:12]
  assign n969_I_0_2_2 = n927_O_0_2_2; // @[Top.scala 1075:12]
  assign n969_I_1_0_0 = n927_O_1_0_0; // @[Top.scala 1075:12]
  assign n969_I_1_0_1 = n927_O_1_0_1; // @[Top.scala 1075:12]
  assign n969_I_1_0_2 = n927_O_1_0_2; // @[Top.scala 1075:12]
  assign n969_I_1_1_0 = n927_O_1_1_0; // @[Top.scala 1075:12]
  assign n969_I_1_1_1 = n927_O_1_1_1; // @[Top.scala 1075:12]
  assign n969_I_1_1_2 = n927_O_1_1_2; // @[Top.scala 1075:12]
  assign n969_I_1_2_0 = n927_O_1_2_0; // @[Top.scala 1075:12]
  assign n969_I_1_2_1 = n927_O_1_2_1; // @[Top.scala 1075:12]
  assign n969_I_1_2_2 = n927_O_1_2_2; // @[Top.scala 1075:12]
  assign n969_I_2_0_0 = n927_O_2_0_0; // @[Top.scala 1075:12]
  assign n969_I_2_0_1 = n927_O_2_0_1; // @[Top.scala 1075:12]
  assign n969_I_2_0_2 = n927_O_2_0_2; // @[Top.scala 1075:12]
  assign n969_I_2_1_0 = n927_O_2_1_0; // @[Top.scala 1075:12]
  assign n969_I_2_1_1 = n927_O_2_1_1; // @[Top.scala 1075:12]
  assign n969_I_2_1_2 = n927_O_2_1_2; // @[Top.scala 1075:12]
  assign n969_I_2_2_0 = n927_O_2_2_0; // @[Top.scala 1075:12]
  assign n969_I_2_2_1 = n927_O_2_2_1; // @[Top.scala 1075:12]
  assign n969_I_2_2_2 = n927_O_2_2_2; // @[Top.scala 1075:12]
  assign n969_I_3_0_0 = n927_O_3_0_0; // @[Top.scala 1075:12]
  assign n969_I_3_0_1 = n927_O_3_0_1; // @[Top.scala 1075:12]
  assign n969_I_3_0_2 = n927_O_3_0_2; // @[Top.scala 1075:12]
  assign n969_I_3_1_0 = n927_O_3_1_0; // @[Top.scala 1075:12]
  assign n969_I_3_1_1 = n927_O_3_1_1; // @[Top.scala 1075:12]
  assign n969_I_3_1_2 = n927_O_3_1_2; // @[Top.scala 1075:12]
  assign n969_I_3_2_0 = n927_O_3_2_0; // @[Top.scala 1075:12]
  assign n969_I_3_2_1 = n927_O_3_2_1; // @[Top.scala 1075:12]
  assign n969_I_3_2_2 = n927_O_3_2_2; // @[Top.scala 1075:12]
  assign n969_I_4_0_0 = n927_O_4_0_0; // @[Top.scala 1075:12]
  assign n969_I_4_0_1 = n927_O_4_0_1; // @[Top.scala 1075:12]
  assign n969_I_4_0_2 = n927_O_4_0_2; // @[Top.scala 1075:12]
  assign n969_I_4_1_0 = n927_O_4_1_0; // @[Top.scala 1075:12]
  assign n969_I_4_1_1 = n927_O_4_1_1; // @[Top.scala 1075:12]
  assign n969_I_4_1_2 = n927_O_4_1_2; // @[Top.scala 1075:12]
  assign n969_I_4_2_0 = n927_O_4_2_0; // @[Top.scala 1075:12]
  assign n969_I_4_2_1 = n927_O_4_2_1; // @[Top.scala 1075:12]
  assign n969_I_4_2_2 = n927_O_4_2_2; // @[Top.scala 1075:12]
  assign n969_I_5_0_0 = n927_O_5_0_0; // @[Top.scala 1075:12]
  assign n969_I_5_0_1 = n927_O_5_0_1; // @[Top.scala 1075:12]
  assign n969_I_5_0_2 = n927_O_5_0_2; // @[Top.scala 1075:12]
  assign n969_I_5_1_0 = n927_O_5_1_0; // @[Top.scala 1075:12]
  assign n969_I_5_1_1 = n927_O_5_1_1; // @[Top.scala 1075:12]
  assign n969_I_5_1_2 = n927_O_5_1_2; // @[Top.scala 1075:12]
  assign n969_I_5_2_0 = n927_O_5_2_0; // @[Top.scala 1075:12]
  assign n969_I_5_2_1 = n927_O_5_2_1; // @[Top.scala 1075:12]
  assign n969_I_5_2_2 = n927_O_5_2_2; // @[Top.scala 1075:12]
  assign n969_I_6_0_0 = n927_O_6_0_0; // @[Top.scala 1075:12]
  assign n969_I_6_0_1 = n927_O_6_0_1; // @[Top.scala 1075:12]
  assign n969_I_6_0_2 = n927_O_6_0_2; // @[Top.scala 1075:12]
  assign n969_I_6_1_0 = n927_O_6_1_0; // @[Top.scala 1075:12]
  assign n969_I_6_1_1 = n927_O_6_1_1; // @[Top.scala 1075:12]
  assign n969_I_6_1_2 = n927_O_6_1_2; // @[Top.scala 1075:12]
  assign n969_I_6_2_0 = n927_O_6_2_0; // @[Top.scala 1075:12]
  assign n969_I_6_2_1 = n927_O_6_2_1; // @[Top.scala 1075:12]
  assign n969_I_6_2_2 = n927_O_6_2_2; // @[Top.scala 1075:12]
  assign n969_I_7_0_0 = n927_O_7_0_0; // @[Top.scala 1075:12]
  assign n969_I_7_0_1 = n927_O_7_0_1; // @[Top.scala 1075:12]
  assign n969_I_7_0_2 = n927_O_7_0_2; // @[Top.scala 1075:12]
  assign n969_I_7_1_0 = n927_O_7_1_0; // @[Top.scala 1075:12]
  assign n969_I_7_1_1 = n927_O_7_1_1; // @[Top.scala 1075:12]
  assign n969_I_7_1_2 = n927_O_7_1_2; // @[Top.scala 1075:12]
  assign n969_I_7_2_0 = n927_O_7_2_0; // @[Top.scala 1075:12]
  assign n969_I_7_2_1 = n927_O_7_2_1; // @[Top.scala 1075:12]
  assign n969_I_7_2_2 = n927_O_7_2_2; // @[Top.scala 1075:12]
  assign n970_valid_up = n969_valid_down; // @[Top.scala 1079:19]
  assign n970_I_0_0_0 = n969_O_0_0_0; // @[Top.scala 1078:12]
  assign n970_I_1_0_0 = n969_O_1_0_0; // @[Top.scala 1078:12]
  assign n970_I_2_0_0 = n969_O_2_0_0; // @[Top.scala 1078:12]
  assign n970_I_3_0_0 = n969_O_3_0_0; // @[Top.scala 1078:12]
  assign n970_I_4_0_0 = n969_O_4_0_0; // @[Top.scala 1078:12]
  assign n970_I_5_0_0 = n969_O_5_0_0; // @[Top.scala 1078:12]
  assign n970_I_6_0_0 = n969_O_6_0_0; // @[Top.scala 1078:12]
  assign n970_I_7_0_0 = n969_O_7_0_0; // @[Top.scala 1078:12]
  assign n971_valid_up = n970_valid_down; // @[Top.scala 1082:19]
  assign n971_I_0_0 = n970_O_0_0; // @[Top.scala 1081:12]
  assign n971_I_1_0 = n970_O_1_0; // @[Top.scala 1081:12]
  assign n971_I_2_0 = n970_O_2_0; // @[Top.scala 1081:12]
  assign n971_I_3_0 = n970_O_3_0; // @[Top.scala 1081:12]
  assign n971_I_4_0 = n970_O_4_0; // @[Top.scala 1081:12]
  assign n971_I_5_0 = n970_O_5_0; // @[Top.scala 1081:12]
  assign n971_I_6_0 = n970_O_6_0; // @[Top.scala 1081:12]
  assign n971_I_7_0 = n970_O_7_0; // @[Top.scala 1081:12]
  assign n972_clock = clock;
  assign n972_reset = reset;
  assign n972_valid_up = n823_valid_down; // @[Top.scala 1085:19]
  assign n972_I_0 = n823_O_0; // @[Top.scala 1084:12]
  assign n972_I_1 = n823_O_1; // @[Top.scala 1084:12]
  assign n972_I_2 = n823_O_2; // @[Top.scala 1084:12]
  assign n972_I_3 = n823_O_3; // @[Top.scala 1084:12]
  assign n972_I_4 = n823_O_4; // @[Top.scala 1084:12]
  assign n972_I_5 = n823_O_5; // @[Top.scala 1084:12]
  assign n972_I_6 = n823_O_6; // @[Top.scala 1084:12]
  assign n972_I_7 = n823_O_7; // @[Top.scala 1084:12]
  assign n973_clock = clock;
  assign n973_reset = reset;
  assign n973_valid_up = n971_valid_down & n972_valid_down; // @[Top.scala 1089:19]
  assign n973_I0_0 = n971_O_0; // @[Top.scala 1087:13]
  assign n973_I0_1 = n971_O_1; // @[Top.scala 1087:13]
  assign n973_I0_2 = n971_O_2; // @[Top.scala 1087:13]
  assign n973_I0_3 = n971_O_3; // @[Top.scala 1087:13]
  assign n973_I0_4 = n971_O_4; // @[Top.scala 1087:13]
  assign n973_I0_5 = n971_O_5; // @[Top.scala 1087:13]
  assign n973_I0_6 = n971_O_6; // @[Top.scala 1087:13]
  assign n973_I0_7 = n971_O_7; // @[Top.scala 1087:13]
  assign n973_I1_0 = n972_O_0; // @[Top.scala 1088:13]
  assign n973_I1_1 = n972_O_1; // @[Top.scala 1088:13]
  assign n973_I1_2 = n972_O_2; // @[Top.scala 1088:13]
  assign n973_I1_3 = n972_O_3; // @[Top.scala 1088:13]
  assign n973_I1_4 = n972_O_4; // @[Top.scala 1088:13]
  assign n973_I1_5 = n972_O_5; // @[Top.scala 1088:13]
  assign n973_I1_6 = n972_O_6; // @[Top.scala 1088:13]
  assign n973_I1_7 = n972_O_7; // @[Top.scala 1088:13]
  assign n1004_valid_up = n787_valid_down & n973_valid_down; // @[Top.scala 1093:20]
  assign n1004_I0_0 = n787_O_0; // @[Top.scala 1091:14]
  assign n1004_I0_1 = n787_O_1; // @[Top.scala 1091:14]
  assign n1004_I0_2 = n787_O_2; // @[Top.scala 1091:14]
  assign n1004_I0_3 = n787_O_3; // @[Top.scala 1091:14]
  assign n1004_I0_4 = n787_O_4; // @[Top.scala 1091:14]
  assign n1004_I0_5 = n787_O_5; // @[Top.scala 1091:14]
  assign n1004_I0_6 = n787_O_6; // @[Top.scala 1091:14]
  assign n1004_I0_7 = n787_O_7; // @[Top.scala 1091:14]
  assign n1004_I1_0 = n973_O_0; // @[Top.scala 1092:14]
  assign n1004_I1_1 = n973_O_1; // @[Top.scala 1092:14]
  assign n1004_I1_2 = n973_O_2; // @[Top.scala 1092:14]
  assign n1004_I1_3 = n973_O_3; // @[Top.scala 1092:14]
  assign n1004_I1_4 = n973_O_4; // @[Top.scala 1092:14]
  assign n1004_I1_5 = n973_O_5; // @[Top.scala 1092:14]
  assign n1004_I1_6 = n973_O_6; // @[Top.scala 1092:14]
  assign n1004_I1_7 = n973_O_7; // @[Top.scala 1092:14]
  assign n1011_valid_up = n601_valid_down & n1004_valid_down; // @[Top.scala 1097:20]
  assign n1011_I0_0 = n601_O_0; // @[Top.scala 1095:14]
  assign n1011_I0_1 = n601_O_1; // @[Top.scala 1095:14]
  assign n1011_I0_2 = n601_O_2; // @[Top.scala 1095:14]
  assign n1011_I0_3 = n601_O_3; // @[Top.scala 1095:14]
  assign n1011_I0_4 = n601_O_4; // @[Top.scala 1095:14]
  assign n1011_I0_5 = n601_O_5; // @[Top.scala 1095:14]
  assign n1011_I0_6 = n601_O_6; // @[Top.scala 1095:14]
  assign n1011_I0_7 = n601_O_7; // @[Top.scala 1095:14]
  assign n1011_I1_0_t0b = n1004_O_0_t0b; // @[Top.scala 1096:14]
  assign n1011_I1_0_t1b = n1004_O_0_t1b; // @[Top.scala 1096:14]
  assign n1011_I1_1_t0b = n1004_O_1_t0b; // @[Top.scala 1096:14]
  assign n1011_I1_1_t1b = n1004_O_1_t1b; // @[Top.scala 1096:14]
  assign n1011_I1_2_t0b = n1004_O_2_t0b; // @[Top.scala 1096:14]
  assign n1011_I1_2_t1b = n1004_O_2_t1b; // @[Top.scala 1096:14]
  assign n1011_I1_3_t0b = n1004_O_3_t0b; // @[Top.scala 1096:14]
  assign n1011_I1_3_t1b = n1004_O_3_t1b; // @[Top.scala 1096:14]
  assign n1011_I1_4_t0b = n1004_O_4_t0b; // @[Top.scala 1096:14]
  assign n1011_I1_4_t1b = n1004_O_4_t1b; // @[Top.scala 1096:14]
  assign n1011_I1_5_t0b = n1004_O_5_t0b; // @[Top.scala 1096:14]
  assign n1011_I1_5_t1b = n1004_O_5_t1b; // @[Top.scala 1096:14]
  assign n1011_I1_6_t0b = n1004_O_6_t0b; // @[Top.scala 1096:14]
  assign n1011_I1_6_t1b = n1004_O_6_t1b; // @[Top.scala 1096:14]
  assign n1011_I1_7_t0b = n1004_O_7_t0b; // @[Top.scala 1096:14]
  assign n1011_I1_7_t1b = n1004_O_7_t1b; // @[Top.scala 1096:14]
  assign n1018_clock = clock;
  assign n1018_reset = reset;
  assign n1018_valid_up = n1011_valid_down; // @[Top.scala 1100:20]
  assign n1018_I_0_t0b = n1011_O_0_t0b; // @[Top.scala 1099:13]
  assign n1018_I_0_t1b_t0b = n1011_O_0_t1b_t0b; // @[Top.scala 1099:13]
  assign n1018_I_0_t1b_t1b = n1011_O_0_t1b_t1b; // @[Top.scala 1099:13]
  assign n1018_I_1_t0b = n1011_O_1_t0b; // @[Top.scala 1099:13]
  assign n1018_I_1_t1b_t0b = n1011_O_1_t1b_t0b; // @[Top.scala 1099:13]
  assign n1018_I_1_t1b_t1b = n1011_O_1_t1b_t1b; // @[Top.scala 1099:13]
  assign n1018_I_2_t0b = n1011_O_2_t0b; // @[Top.scala 1099:13]
  assign n1018_I_2_t1b_t0b = n1011_O_2_t1b_t0b; // @[Top.scala 1099:13]
  assign n1018_I_2_t1b_t1b = n1011_O_2_t1b_t1b; // @[Top.scala 1099:13]
  assign n1018_I_3_t0b = n1011_O_3_t0b; // @[Top.scala 1099:13]
  assign n1018_I_3_t1b_t0b = n1011_O_3_t1b_t0b; // @[Top.scala 1099:13]
  assign n1018_I_3_t1b_t1b = n1011_O_3_t1b_t1b; // @[Top.scala 1099:13]
  assign n1018_I_4_t0b = n1011_O_4_t0b; // @[Top.scala 1099:13]
  assign n1018_I_4_t1b_t0b = n1011_O_4_t1b_t0b; // @[Top.scala 1099:13]
  assign n1018_I_4_t1b_t1b = n1011_O_4_t1b_t1b; // @[Top.scala 1099:13]
  assign n1018_I_5_t0b = n1011_O_5_t0b; // @[Top.scala 1099:13]
  assign n1018_I_5_t1b_t0b = n1011_O_5_t1b_t0b; // @[Top.scala 1099:13]
  assign n1018_I_5_t1b_t1b = n1011_O_5_t1b_t1b; // @[Top.scala 1099:13]
  assign n1018_I_6_t0b = n1011_O_6_t0b; // @[Top.scala 1099:13]
  assign n1018_I_6_t1b_t0b = n1011_O_6_t1b_t0b; // @[Top.scala 1099:13]
  assign n1018_I_6_t1b_t1b = n1011_O_6_t1b_t1b; // @[Top.scala 1099:13]
  assign n1018_I_7_t0b = n1011_O_7_t0b; // @[Top.scala 1099:13]
  assign n1018_I_7_t1b_t0b = n1011_O_7_t1b_t0b; // @[Top.scala 1099:13]
  assign n1018_I_7_t1b_t1b = n1011_O_7_t1b_t1b; // @[Top.scala 1099:13]
  assign n1019_clock = clock;
  assign n1019_reset = reset;
  assign n1019_valid_up = n1018_valid_down; // @[Top.scala 1103:20]
  assign n1019_I_0_t0b = n1018_O_0_t0b; // @[Top.scala 1102:13]
  assign n1019_I_0_t1b_t0b = n1018_O_0_t1b_t0b; // @[Top.scala 1102:13]
  assign n1019_I_0_t1b_t1b = n1018_O_0_t1b_t1b; // @[Top.scala 1102:13]
  assign n1019_I_1_t0b = n1018_O_1_t0b; // @[Top.scala 1102:13]
  assign n1019_I_1_t1b_t0b = n1018_O_1_t1b_t0b; // @[Top.scala 1102:13]
  assign n1019_I_1_t1b_t1b = n1018_O_1_t1b_t1b; // @[Top.scala 1102:13]
  assign n1019_I_2_t0b = n1018_O_2_t0b; // @[Top.scala 1102:13]
  assign n1019_I_2_t1b_t0b = n1018_O_2_t1b_t0b; // @[Top.scala 1102:13]
  assign n1019_I_2_t1b_t1b = n1018_O_2_t1b_t1b; // @[Top.scala 1102:13]
  assign n1019_I_3_t0b = n1018_O_3_t0b; // @[Top.scala 1102:13]
  assign n1019_I_3_t1b_t0b = n1018_O_3_t1b_t0b; // @[Top.scala 1102:13]
  assign n1019_I_3_t1b_t1b = n1018_O_3_t1b_t1b; // @[Top.scala 1102:13]
  assign n1019_I_4_t0b = n1018_O_4_t0b; // @[Top.scala 1102:13]
  assign n1019_I_4_t1b_t0b = n1018_O_4_t1b_t0b; // @[Top.scala 1102:13]
  assign n1019_I_4_t1b_t1b = n1018_O_4_t1b_t1b; // @[Top.scala 1102:13]
  assign n1019_I_5_t0b = n1018_O_5_t0b; // @[Top.scala 1102:13]
  assign n1019_I_5_t1b_t0b = n1018_O_5_t1b_t0b; // @[Top.scala 1102:13]
  assign n1019_I_5_t1b_t1b = n1018_O_5_t1b_t1b; // @[Top.scala 1102:13]
  assign n1019_I_6_t0b = n1018_O_6_t0b; // @[Top.scala 1102:13]
  assign n1019_I_6_t1b_t0b = n1018_O_6_t1b_t0b; // @[Top.scala 1102:13]
  assign n1019_I_6_t1b_t1b = n1018_O_6_t1b_t1b; // @[Top.scala 1102:13]
  assign n1019_I_7_t0b = n1018_O_7_t0b; // @[Top.scala 1102:13]
  assign n1019_I_7_t1b_t0b = n1018_O_7_t1b_t0b; // @[Top.scala 1102:13]
  assign n1019_I_7_t1b_t1b = n1018_O_7_t1b_t1b; // @[Top.scala 1102:13]
  assign n1020_clock = clock;
  assign n1020_reset = reset;
  assign n1020_valid_up = n1019_valid_down; // @[Top.scala 1106:20]
  assign n1020_I_0_t0b = n1019_O_0_t0b; // @[Top.scala 1105:13]
  assign n1020_I_0_t1b_t0b = n1019_O_0_t1b_t0b; // @[Top.scala 1105:13]
  assign n1020_I_0_t1b_t1b = n1019_O_0_t1b_t1b; // @[Top.scala 1105:13]
  assign n1020_I_1_t0b = n1019_O_1_t0b; // @[Top.scala 1105:13]
  assign n1020_I_1_t1b_t0b = n1019_O_1_t1b_t0b; // @[Top.scala 1105:13]
  assign n1020_I_1_t1b_t1b = n1019_O_1_t1b_t1b; // @[Top.scala 1105:13]
  assign n1020_I_2_t0b = n1019_O_2_t0b; // @[Top.scala 1105:13]
  assign n1020_I_2_t1b_t0b = n1019_O_2_t1b_t0b; // @[Top.scala 1105:13]
  assign n1020_I_2_t1b_t1b = n1019_O_2_t1b_t1b; // @[Top.scala 1105:13]
  assign n1020_I_3_t0b = n1019_O_3_t0b; // @[Top.scala 1105:13]
  assign n1020_I_3_t1b_t0b = n1019_O_3_t1b_t0b; // @[Top.scala 1105:13]
  assign n1020_I_3_t1b_t1b = n1019_O_3_t1b_t1b; // @[Top.scala 1105:13]
  assign n1020_I_4_t0b = n1019_O_4_t0b; // @[Top.scala 1105:13]
  assign n1020_I_4_t1b_t0b = n1019_O_4_t1b_t0b; // @[Top.scala 1105:13]
  assign n1020_I_4_t1b_t1b = n1019_O_4_t1b_t1b; // @[Top.scala 1105:13]
  assign n1020_I_5_t0b = n1019_O_5_t0b; // @[Top.scala 1105:13]
  assign n1020_I_5_t1b_t0b = n1019_O_5_t1b_t0b; // @[Top.scala 1105:13]
  assign n1020_I_5_t1b_t1b = n1019_O_5_t1b_t1b; // @[Top.scala 1105:13]
  assign n1020_I_6_t0b = n1019_O_6_t0b; // @[Top.scala 1105:13]
  assign n1020_I_6_t1b_t0b = n1019_O_6_t1b_t0b; // @[Top.scala 1105:13]
  assign n1020_I_6_t1b_t1b = n1019_O_6_t1b_t1b; // @[Top.scala 1105:13]
  assign n1020_I_7_t0b = n1019_O_7_t0b; // @[Top.scala 1105:13]
  assign n1020_I_7_t1b_t0b = n1019_O_7_t1b_t0b; // @[Top.scala 1105:13]
  assign n1020_I_7_t1b_t1b = n1019_O_7_t1b_t1b; // @[Top.scala 1105:13]
endmodule
