// Latency = 4
module top(
  input CLK/*verilator public*/, 
  input [7:0] I_0_0_0/*verilator public*/, 
  output [7:0] O_0_0_0/*verilator public*/, 
  input [7:0] I_1_0_0/*verilator public*/, 
  output [7:0] O_1_0_0/*verilator public*/, 
  input [7:0] I_2_0_0/*verilator public*/, 
  output [7:0] O_2_0_0/*verilator public*/, 
  input [7:0] I_3_0_0/*verilator public*/, 
  output [7:0] O_3_0_0/*verilator public*/, 
  output valid_down/*verilator public*/, 
  input valid_up/*verilator public*/
);
  wire dontcare;
  wire [31:0] io_output_counts_1;
  wire [31:0] io_output_counts_0;

  x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1 sampler_box ( // @[m_x55_ctr_0.scala 26:17:@1721.4]
    .clock(CLK), // @[:@1296.4]
    .reset('b0), // @[:@1297.4]
    .io_in_x316_TREADY(dontcare), // @[:@1298.4]
    .io_in_x316_TDATA({I_0_0_0,I_1_0_0,I_2_0_0,I_3_0_0}), // @[:@1298.4]
    .io_in_x316_TID(8'h0),
    .io_in_x316_TDEST(8'h0),
    .io_in_x317_TVALID(valid_down), // @[:@1298.4]
    .io_in_x317_TDATA({O_0_0_0,O_1_0_0,O_2_0_0,O_3_0_0}), // @[:@1298.4]
    .io_in_x317_TREADY(1'b1), // @[:@1298.4]
    .io_sigsIn_datapathEn(valid_up), // @[:@1298.4]
    .io_sigsIn_backpressure(1'b1), // @[:@20563.4]
    .io_sigsIn_break(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_1(io_output_counts_1), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_0(io_output_counts_0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_0(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_1(1'b0), // @[:@20563.4]
    .io_rr('b1) // @[:@1298.4]
  );

  wire dontcare2;

  wire io_output_oobs_0;
  wire io_output_oobs_1;
  x324_ctrchain cchain ( // @[:@2879.2]
    .clock(CLK), // @[:@2880.4]
    .reset(1'b0), // @[:@2881.4]
    .io_input_reset(1'b0), // @[:@2882.4]
    .io_input_enable(valid_up), // @[:@2882.4]
    .io_output_counts_1(io_output_counts_1), // @[:@2882.4]
    .io_output_counts_0(io_output_counts_0), // @[:@2882.4]
    .io_output_oobs_0(io_output_oobs_0), // @[:@2882.4]
    .io_output_oobs_1(io_output_oobs_1), // @[:@2882.4]
    .io_output_done(dontcare2) // @[:@2882.4]
  );

endmodule

module RetimeShiftRegister
#(
    parameter WIDTH = 1,
    parameter STAGES = 1)
(
    input clock,
    input reset,
    input flow,
    input [WIDTH-1:0] init,
    input [WIDTH-1:0] in,
    output reg [WIDTH-1:0] out
);
  integer i;
  reg [WIDTH-1:0] sr[STAGES:0]; // Create 'STAGES' number of register, each 'WIDTH' bits wide

   /* synopsys dc_tcl_script_begin
    set_ungroup [current_design] true
    set_flatten true -effort high -phase true -design [current_design]
    set_dont_retime [current_design] false
    set_optimize_registers true -design [current_design]
    */
  always @(posedge clock) begin
    if (reset) begin
      for(i=0; i<STAGES; i=i+1) begin
        sr[i] <= init;
      end
    end else begin
      if (flow) begin 
        sr[0] <= in;
        for(i=1; i<STAGES; i=i+1) begin
          sr[i] <= sr[i-1];
        end
      end
    end
  end

  always @(*) begin
    out = sr[STAGES-1];
  end
endmodule
module FF( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  output [31:0] io_rPort_0_output_0, // @[:@6.4]
  input  [31:0] io_wPort_0_data_0, // @[:@6.4]
  input         io_wPort_0_reset, // @[:@6.4]
  input         io_wPort_0_en_0 // @[:@6.4]
);
  reg [31:0] ff; // @[MemPrimitives.scala 173:19:@21.4]
  reg [31:0] _RAND_0;
  wire [31:0] _T_68; // @[MemPrimitives.scala 177:32:@23.4]
  wire [31:0] _T_69; // @[MemPrimitives.scala 177:12:@24.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 177:32:@23.4]
  assign _T_69 = io_wPort_0_reset ? 32'h0 : _T_68; // @[MemPrimitives.scala 177:12:@24.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 178:34:@26.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 32'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 32'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SRFF( // @[:@28.2]
  input   clock, // @[:@29.4]
  input   reset, // @[:@30.4]
  input   io_input_set, // @[:@31.4]
  input   io_input_reset, // @[:@31.4]
  input   io_input_asyn_reset, // @[:@31.4]
  output  io_output // @[:@31.4]
);
  reg  _T_15; // @[SRFF.scala 20:21:@33.4]
  reg [31:0] _RAND_0;
  wire  _T_19; // @[SRFF.scala 21:74:@34.4]
  wire  _T_20; // @[SRFF.scala 21:48:@35.4]
  wire  _T_21; // @[SRFF.scala 21:14:@36.4]
  assign _T_19 = io_input_reset ? 1'h0 : _T_15; // @[SRFF.scala 21:74:@34.4]
  assign _T_20 = io_input_set ? 1'h1 : _T_19; // @[SRFF.scala 21:48:@35.4]
  assign _T_21 = io_input_asyn_reset ? 1'h0 : _T_20; // @[SRFF.scala 21:14:@36.4]
  assign io_output = io_input_asyn_reset ? 1'h0 : _T_15; // @[SRFF.scala 22:15:@39.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_15 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_15 <= 1'h0;
    end else begin
      if (io_input_asyn_reset) begin
        _T_15 <= 1'h0;
      end else begin
        if (io_input_set) begin
          _T_15 <= 1'h1;
        end else begin
          if (io_input_reset) begin
            _T_15 <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module SingleCounter( // @[:@41.2]
  input   clock, // @[:@42.4]
  input   reset, // @[:@43.4]
  input   io_input_reset, // @[:@44.4]
  output  io_output_done // @[:@44.4]
);
  wire  bases_0_clock; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_reset; // @[Counter.scala 253:53:@57.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 253:53:@57.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 253:53:@57.4]
  wire  SRFF_clock; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_set; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_output; // @[Counter.scala 255:22:@73.4]
  wire [31:0] _T_48; // @[Counter.scala 279:52:@101.4]
  wire [32:0] _T_50; // @[Counter.scala 283:33:@102.4]
  wire [31:0] _T_51; // @[Counter.scala 283:33:@103.4]
  wire [31:0] _T_52; // @[Counter.scala 283:33:@104.4]
  wire  _T_57; // @[Counter.scala 285:18:@106.4]
  wire [31:0] _T_68; // @[Counter.scala 291:115:@114.4]
  wire [31:0] _T_71; // @[Counter.scala 291:152:@117.4]
  wire [31:0] _T_72; // @[Counter.scala 291:74:@118.4]
  FF bases_0 ( // @[Counter.scala 253:53:@57.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 255:22:@73.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 279:52:@101.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@102.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@103.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 283:33:@104.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'shf); // @[Counter.scala 285:18:@106.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 291:115:@114.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 291:152:@117.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 291:74:@118.4]
  assign io_output_done = $signed(_T_52) >= $signed(32'shf); // @[Counter.scala 325:20:@127.4]
  assign bases_0_clock = clock; // @[:@58.4]
  assign bases_0_reset = reset; // @[:@59.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 291:31:@120.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 273:27:@99.4]
  assign bases_0_io_wPort_0_en_0 = 1'h1; // @[Counter.scala 276:29:@100.4]
  assign SRFF_clock = clock; // @[:@74.4]
  assign SRFF_reset = reset; // @[:@75.4]
  assign SRFF_io_input_set = io_input_reset == 1'h0; // @[Counter.scala 256:23:@78.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 257:25:@80.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 258:30:@81.4]
endmodule
module RetimeWrapper( // @[:@144.2]
  input   clock, // @[:@145.4]
  input   reset, // @[:@146.4]
  input   io_flow, // @[:@147.4]
  input   io_in, // @[:@147.4]
  output  io_out // @[:@147.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@149.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@149.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@162.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@161.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@160.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@159.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@158.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@156.4]
endmodule
module RootController_sm( // @[:@312.2]
  input   clock, // @[:@313.4]
  input   reset, // @[:@314.4]
  input   io_enable, // @[:@315.4]
  output  io_done, // @[:@315.4]
  input   io_rst, // @[:@315.4]
  input   io_ctrDone, // @[:@315.4]
  output  io_ctrInc, // @[:@315.4]
  input   io_doneIn_0, // @[:@315.4]
  output  io_enableOut_0, // @[:@315.4]
  output  io_childAck_0 // @[:@315.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@318.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@321.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@338.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@433.4]
  wire  finished; // @[Controllers.scala 81:26:@324.4]
  wire  synchronize; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  wire  _T_122; // @[Controllers.scala 128:33:@371.4]
  wire  _T_124; // @[Controllers.scala 128:54:@372.4]
  wire  _T_125; // @[Controllers.scala 128:52:@373.4]
  wire  _T_126; // @[Controllers.scala 128:66:@374.4]
  wire  _T_128; // @[Controllers.scala 128:98:@376.4]
  wire  _T_129; // @[Controllers.scala 128:96:@377.4]
  wire  _T_131; // @[Controllers.scala 128:123:@378.4]
  wire  _T_133; // @[Controllers.scala 129:48:@381.4]
  wire  _T_138; // @[Controllers.scala 130:52:@386.4]
  wire  _T_139; // @[Controllers.scala 130:50:@387.4]
  wire  _T_147; // @[Controllers.scala 130:129:@393.4]
  wire  _T_150; // @[Controllers.scala 131:45:@396.4]
  wire  _T_154; // @[Controllers.scala 213:68:@402.4]
  wire  _T_156; // @[Controllers.scala 213:90:@404.4]
  wire  _T_158; // @[Controllers.scala 213:132:@406.4]
  wire  _T_159; // @[Controllers.scala 213:130:@407.4]
  wire  _T_160; // @[Controllers.scala 213:156:@408.4]
  reg  _T_166; // @[package.scala 48:56:@412.4]
  reg [31:0] _RAND_0;
  reg  _T_180; // @[package.scala 48:56:@430.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@318.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@321.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@338.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@357.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@416.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@433.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  assign finished = done_0_io_output | io_done; // @[Controllers.scala 81:26:@324.4]
  assign synchronize = RetimeWrapper_io_out; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  assign _T_122 = done_0_io_output == 1'h0; // @[Controllers.scala 128:33:@371.4]
  assign _T_124 = io_ctrDone == 1'h0; // @[Controllers.scala 128:54:@372.4]
  assign _T_125 = _T_122 & _T_124; // @[Controllers.scala 128:52:@373.4]
  assign _T_126 = _T_125 & io_enable; // @[Controllers.scala 128:66:@374.4]
  assign _T_128 = ~ iterDone_0_io_output; // @[Controllers.scala 128:98:@376.4]
  assign _T_129 = _T_126 & _T_128; // @[Controllers.scala 128:96:@377.4]
  assign _T_131 = io_doneIn_0 == 1'h0; // @[Controllers.scala 128:123:@378.4]
  assign _T_133 = io_doneIn_0 | io_rst; // @[Controllers.scala 129:48:@381.4]
  assign _T_138 = synchronize == 1'h0; // @[Controllers.scala 130:52:@386.4]
  assign _T_139 = io_doneIn_0 & _T_138; // @[Controllers.scala 130:50:@387.4]
  assign _T_147 = finished == 1'h0; // @[Controllers.scala 130:129:@393.4]
  assign _T_150 = io_rst == 1'h0; // @[Controllers.scala 131:45:@396.4]
  assign _T_154 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@402.4]
  assign _T_156 = _T_154 & _T_128; // @[Controllers.scala 213:90:@404.4]
  assign _T_158 = ~ done_0_io_output; // @[Controllers.scala 213:132:@406.4]
  assign _T_159 = _T_156 & _T_158; // @[Controllers.scala 213:130:@407.4]
  assign _T_160 = ~ io_ctrDone; // @[Controllers.scala 213:156:@408.4]
  assign io_done = RetimeWrapper_2_io_out; // @[Controllers.scala 245:13:@440.4]
  assign io_ctrInc = io_doneIn_0; // @[Controllers.scala 122:17:@356.4]
  assign io_enableOut_0 = _T_159 & _T_160; // @[Controllers.scala 213:55:@410.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@401.4]
  assign active_0_clock = clock; // @[:@319.4]
  assign active_0_reset = reset; // @[:@320.4]
  assign active_0_io_input_set = _T_129 & _T_131; // @[Controllers.scala 128:30:@380.4]
  assign active_0_io_input_reset = _T_133 | done_0_io_output; // @[Controllers.scala 129:32:@385.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@326.4]
  assign done_0_clock = clock; // @[:@322.4]
  assign done_0_reset = reset; // @[:@323.4]
  assign done_0_io_input_set = io_ctrDone & _T_150; // @[Controllers.scala 131:28:@399.4]
  assign done_0_io_input_reset = io_rst | done_0_io_output; // @[Controllers.scala 86:33:@336.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@327.4]
  assign iterDone_0_clock = clock; // @[:@339.4]
  assign iterDone_0_reset = reset; // @[:@340.4]
  assign iterDone_0_io_input_set = _T_139 & _T_147; // @[Controllers.scala 130:32:@395.4]
  assign iterDone_0_io_input_reset = synchronize | io_rst; // @[Controllers.scala 92:37:@350.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@341.4]
  assign RetimeWrapper_clock = clock; // @[:@358.4]
  assign RetimeWrapper_reset = reset; // @[:@359.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@361.4]
  assign RetimeWrapper_io_in = io_doneIn_0; // @[package.scala 94:16:@360.4]
  assign RetimeWrapper_1_clock = clock; // @[:@417.4]
  assign RetimeWrapper_1_reset = reset; // @[:@418.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@420.4]
  assign RetimeWrapper_1_io_in = done_0_io_output & _T_166; // @[package.scala 94:16:@419.4]
  assign RetimeWrapper_2_clock = clock; // @[:@434.4]
  assign RetimeWrapper_2_reset = reset; // @[:@435.4]
  assign RetimeWrapper_2_io_flow = io_enable; // @[package.scala 95:18:@437.4]
  assign RetimeWrapper_2_io_in = done_0_io_output & _T_180; // @[package.scala 94:16:@436.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_166 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_180 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_166 <= 1'h0;
    end else begin
      _T_166 <= _T_122;
    end
    if (reset) begin
      _T_180 <= 1'h0;
    end else begin
      _T_180 <= _T_122;
    end
  end
endmodule
module x593_outr_UnitPipe_sm( // @[:@2389.2]
  input   clock, // @[:@2390.4]
  input   reset, // @[:@2391.4]
  input   io_enable, // @[:@2392.4]
  output  io_done, // @[:@2392.4]
  input   io_parentAck, // @[:@2392.4]
  input   io_doneIn_0, // @[:@2392.4]
  output  io_enableOut_0, // @[:@2392.4]
  output  io_childAck_0, // @[:@2392.4]
  input   io_ctrCopyDone_0 // @[:@2392.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@2395.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@2395.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@2395.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@2395.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@2395.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@2395.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@2398.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@2398.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@2398.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@2398.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@2398.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@2398.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@2415.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@2415.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@2415.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@2415.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@2415.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@2415.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@2446.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@2446.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@2446.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@2446.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@2446.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@2460.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@2460.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@2460.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@2460.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@2460.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@2478.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@2478.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@2478.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@2478.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@2478.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@2515.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@2515.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@2515.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@2515.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@2515.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@2532.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@2532.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@2532.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@2532.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@2532.4]
  wire  _T_105; // @[Controllers.scala 165:35:@2430.4]
  wire  _T_107; // @[Controllers.scala 165:60:@2431.4]
  wire  _T_108; // @[Controllers.scala 165:58:@2432.4]
  wire  _T_110; // @[Controllers.scala 165:76:@2433.4]
  wire  _T_111; // @[Controllers.scala 165:74:@2434.4]
  wire  _T_115; // @[Controllers.scala 165:109:@2437.4]
  wire  _T_118; // @[Controllers.scala 165:141:@2439.4]
  wire  _T_126; // @[package.scala 96:25:@2451.4 package.scala 96:25:@2452.4]
  wire  _T_130; // @[Controllers.scala 167:54:@2454.4]
  wire  _T_131; // @[Controllers.scala 167:52:@2455.4]
  wire  _T_138; // @[package.scala 96:25:@2465.4 package.scala 96:25:@2466.4]
  wire  _T_156; // @[package.scala 96:25:@2483.4 package.scala 96:25:@2484.4]
  wire  _T_160; // @[Controllers.scala 169:67:@2486.4]
  wire  _T_161; // @[Controllers.scala 169:86:@2487.4]
  wire  _T_174; // @[Controllers.scala 213:68:@2501.4]
  wire  _T_176; // @[Controllers.scala 213:90:@2503.4]
  wire  _T_178; // @[Controllers.scala 213:132:@2505.4]
  reg  _T_186; // @[package.scala 48:56:@2511.4]
  reg [31:0] _RAND_0;
  wire  _T_187; // @[package.scala 100:41:@2513.4]
  reg  _T_200; // @[package.scala 48:56:@2529.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@2395.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@2398.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@2415.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@2446.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@2460.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@2478.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@2515.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@2532.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_105 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@2430.4]
  assign _T_107 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@2431.4]
  assign _T_108 = _T_105 & _T_107; // @[Controllers.scala 165:58:@2432.4]
  assign _T_110 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@2433.4]
  assign _T_111 = _T_108 & _T_110; // @[Controllers.scala 165:74:@2434.4]
  assign _T_115 = _T_111 & io_enable; // @[Controllers.scala 165:109:@2437.4]
  assign _T_118 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@2439.4]
  assign _T_126 = RetimeWrapper_io_out; // @[package.scala 96:25:@2451.4 package.scala 96:25:@2452.4]
  assign _T_130 = _T_126 == 1'h0; // @[Controllers.scala 167:54:@2454.4]
  assign _T_131 = io_doneIn_0 | _T_130; // @[Controllers.scala 167:52:@2455.4]
  assign _T_138 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@2465.4 package.scala 96:25:@2466.4]
  assign _T_156 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@2483.4 package.scala 96:25:@2484.4]
  assign _T_160 = _T_156 == 1'h0; // @[Controllers.scala 169:67:@2486.4]
  assign _T_161 = _T_160 & io_enable; // @[Controllers.scala 169:86:@2487.4]
  assign _T_174 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@2501.4]
  assign _T_176 = _T_174 & _T_105; // @[Controllers.scala 213:90:@2503.4]
  assign _T_178 = ~ done_0_io_output; // @[Controllers.scala 213:132:@2505.4]
  assign _T_187 = done_0_io_output & _T_186; // @[package.scala 100:41:@2513.4]
  assign io_done = RetimeWrapper_4_io_out; // @[Controllers.scala 245:13:@2539.4]
  assign io_enableOut_0 = _T_176 & _T_178; // @[Controllers.scala 213:55:@2509.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@2500.4]
  assign active_0_clock = clock; // @[:@2396.4]
  assign active_0_reset = reset; // @[:@2397.4]
  assign active_0_io_input_set = _T_115 & _T_118; // @[Controllers.scala 165:32:@2441.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@2445.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@2403.4]
  assign done_0_clock = clock; // @[:@2399.4]
  assign done_0_reset = reset; // @[:@2400.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_161; // @[Controllers.scala 169:30:@2491.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@2413.4 Controllers.scala 170:32:@2498.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@2404.4]
  assign iterDone_0_clock = clock; // @[:@2416.4]
  assign iterDone_0_reset = reset; // @[:@2417.4]
  assign iterDone_0_io_input_set = _T_131 & io_enable; // @[Controllers.scala 167:34:@2459.4]
  assign iterDone_0_io_input_reset = _T_138 | io_parentAck; // @[Controllers.scala 92:37:@2427.4 Controllers.scala 168:36:@2475.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@2418.4]
  assign RetimeWrapper_clock = clock; // @[:@2447.4]
  assign RetimeWrapper_reset = reset; // @[:@2448.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@2450.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@2449.4]
  assign RetimeWrapper_1_clock = clock; // @[:@2461.4]
  assign RetimeWrapper_1_reset = reset; // @[:@2462.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@2464.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@2463.4]
  assign RetimeWrapper_2_clock = clock; // @[:@2479.4]
  assign RetimeWrapper_2_reset = reset; // @[:@2480.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@2482.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@2481.4]
  assign RetimeWrapper_3_clock = clock; // @[:@2516.4]
  assign RetimeWrapper_3_reset = reset; // @[:@2517.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@2519.4]
  assign RetimeWrapper_3_io_in = _T_187 | io_parentAck; // @[package.scala 94:16:@2518.4]
  assign RetimeWrapper_4_clock = clock; // @[:@2533.4]
  assign RetimeWrapper_4_reset = reset; // @[:@2534.4]
  assign RetimeWrapper_4_io_flow = io_enable; // @[package.scala 95:18:@2536.4]
  assign RetimeWrapper_4_io_in = done_0_io_output & _T_200; // @[package.scala 94:16:@2535.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_186 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_200 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_186 <= 1'h0;
    end else begin
      _T_186 <= _T_110;
    end
    if (reset) begin
      _T_200 <= 1'h0;
    end else begin
      _T_200 <= _T_110;
    end
  end
endmodule
module SingleCounter_1( // @[:@2659.2]
  input         clock, // @[:@2660.4]
  input         reset, // @[:@2661.4]
  input         io_input_reset, // @[:@2662.4]
  input         io_input_enable, // @[:@2662.4]
  output [31:0] io_output_count_0, // @[:@2662.4]
  output        io_output_oobs_0, // @[:@2662.4]
  output        io_output_done, // @[:@2662.4]
  output        io_output_saturated // @[:@2662.4]
);
  wire  bases_0_clock; // @[Counter.scala 253:53:@2675.4]
  wire  bases_0_reset; // @[Counter.scala 253:53:@2675.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 253:53:@2675.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 253:53:@2675.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 253:53:@2675.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 253:53:@2675.4]
  wire  SRFF_clock; // @[Counter.scala 255:22:@2691.4]
  wire  SRFF_reset; // @[Counter.scala 255:22:@2691.4]
  wire  SRFF_io_input_set; // @[Counter.scala 255:22:@2691.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 255:22:@2691.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 255:22:@2691.4]
  wire  SRFF_io_output; // @[Counter.scala 255:22:@2691.4]
  wire  _T_36; // @[Counter.scala 256:45:@2694.4]
  wire [31:0] _T_48; // @[Counter.scala 279:52:@2719.4]
  wire [32:0] _T_50; // @[Counter.scala 283:33:@2720.4]
  wire [31:0] _T_51; // @[Counter.scala 283:33:@2721.4]
  wire [31:0] _T_52; // @[Counter.scala 283:33:@2722.4]
  wire  _T_57; // @[Counter.scala 285:18:@2724.4]
  wire [31:0] _T_68; // @[Counter.scala 291:115:@2732.4]
  wire [31:0] _T_71; // @[Counter.scala 291:152:@2735.4]
  wire [31:0] _T_72; // @[Counter.scala 291:74:@2736.4]
  wire  _T_75; // @[Counter.scala 314:102:@2740.4]
  wire  _T_77; // @[Counter.scala 314:130:@2741.4]
  FF bases_0 ( // @[Counter.scala 253:53:@2675.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 255:22:@2691.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 256:45:@2694.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 279:52:@2719.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@2720.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@2721.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 283:33:@2722.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh4); // @[Counter.scala 285:18:@2724.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 291:115:@2732.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 291:152:@2735.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 291:74:@2736.4]
  assign _T_75 = $signed(_T_48) < $signed(32'sh0); // @[Counter.scala 314:102:@2740.4]
  assign _T_77 = $signed(_T_48) >= $signed(32'sh4); // @[Counter.scala 314:130:@2741.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 296:28:@2739.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 314:60:@2743.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 325:20:@2745.4]
  assign io_output_saturated = $signed(_T_52) >= $signed(32'sh4); // @[Counter.scala 332:25:@2748.4]
  assign bases_0_clock = clock; // @[:@2676.4]
  assign bases_0_reset = reset; // @[:@2677.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 291:31:@2738.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 273:27:@2717.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 276:29:@2718.4]
  assign SRFF_clock = clock; // @[:@2692.4]
  assign SRFF_reset = reset; // @[:@2693.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 256:23:@2696.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 257:25:@2698.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 258:30:@2699.4]
endmodule
module SingleCounter_2( // @[:@2788.2]
  input         clock, // @[:@2789.4]
  input         reset, // @[:@2790.4]
  input         io_setup_saturate, // @[:@2791.4]
  input         io_input_reset, // @[:@2791.4]
  input         io_input_enable, // @[:@2791.4]
  output [31:0] io_output_count_0, // @[:@2791.4]
  output        io_output_oobs_0, // @[:@2791.4]
  output        io_output_done // @[:@2791.4]
);
  wire  bases_0_clock; // @[Counter.scala 253:53:@2804.4]
  wire  bases_0_reset; // @[Counter.scala 253:53:@2804.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 253:53:@2804.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 253:53:@2804.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 253:53:@2804.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 253:53:@2804.4]
  wire  SRFF_clock; // @[Counter.scala 255:22:@2820.4]
  wire  SRFF_reset; // @[Counter.scala 255:22:@2820.4]
  wire  SRFF_io_input_set; // @[Counter.scala 255:22:@2820.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 255:22:@2820.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 255:22:@2820.4]
  wire  SRFF_io_output; // @[Counter.scala 255:22:@2820.4]
  wire  _T_36; // @[Counter.scala 256:45:@2823.4]
  wire [31:0] _T_48; // @[Counter.scala 279:52:@2848.4]
  wire [32:0] _T_50; // @[Counter.scala 283:33:@2849.4]
  wire [31:0] _T_51; // @[Counter.scala 283:33:@2850.4]
  wire [31:0] _T_52; // @[Counter.scala 283:33:@2851.4]
  wire  _T_57; // @[Counter.scala 285:18:@2853.4]
  wire [31:0] _T_68; // @[Counter.scala 291:115:@2861.4]
  wire [31:0] _T_70; // @[Counter.scala 291:85:@2863.4]
  wire [31:0] _T_71; // @[Counter.scala 291:152:@2864.4]
  wire [31:0] _T_72; // @[Counter.scala 291:74:@2865.4]
  wire  _T_75; // @[Counter.scala 314:102:@2869.4]
  wire  _T_77; // @[Counter.scala 314:130:@2870.4]
  FF bases_0 ( // @[Counter.scala 253:53:@2804.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 255:22:@2820.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 256:45:@2823.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 279:52:@2848.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh4); // @[Counter.scala 283:33:@2849.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh4); // @[Counter.scala 283:33:@2850.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 283:33:@2851.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh4); // @[Counter.scala 285:18:@2853.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 291:115:@2861.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 32'h0; // @[Counter.scala 291:85:@2863.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 291:152:@2864.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 291:74:@2865.4]
  assign _T_75 = $signed(_T_48) < $signed(32'sh0); // @[Counter.scala 314:102:@2869.4]
  assign _T_77 = $signed(_T_48) >= $signed(32'sh4); // @[Counter.scala 314:130:@2870.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 296:28:@2868.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 314:60:@2872.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 325:20:@2874.4]
  assign bases_0_clock = clock; // @[:@2805.4]
  assign bases_0_reset = reset; // @[:@2806.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 291:31:@2867.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 273:27:@2846.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 276:29:@2847.4]
  assign SRFF_clock = clock; // @[:@2821.4]
  assign SRFF_reset = reset; // @[:@2822.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 256:23:@2825.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 257:25:@2827.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 258:30:@2828.4]
endmodule
module x324_ctrchain( // @[:@2879.2]
  input         clock, // @[:@2880.4]
  input         reset, // @[:@2881.4]
  input         io_input_reset, // @[:@2882.4]
  input         io_input_enable, // @[:@2882.4]
  output [31:0] io_output_counts_1, // @[:@2882.4]
  output [31:0] io_output_counts_0, // @[:@2882.4]
  output        io_output_oobs_0, // @[:@2882.4]
  output        io_output_oobs_1, // @[:@2882.4]
  output        io_output_done // @[:@2882.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_reset; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 505:46:@2884.4]
  wire [31:0] ctrs_0_io_output_count_0; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_io_output_saturated; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_1_clock; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_reset; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_io_setup_saturate; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_io_input_reset; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_io_input_enable; // @[Counter.scala 505:46:@2887.4]
  wire [31:0] ctrs_1_io_output_count_0; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_io_output_oobs_0; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_io_output_done; // @[Counter.scala 505:46:@2887.4]
  wire  isDone; // @[Counter.scala 533:51:@2904.4]
  reg  wasDone; // @[Counter.scala 534:24:@2905.4]
  reg [31:0] _RAND_0;
  wire  _T_64; // @[Counter.scala 538:69:@2913.4]
  wire  _T_66; // @[Counter.scala 538:80:@2914.4]
  reg  doneLatch; // @[Counter.scala 542:26:@2919.4]
  reg [31:0] _RAND_1;
  wire  _T_73; // @[Counter.scala 543:48:@2920.4]
  wire  _T_74; // @[Counter.scala 543:19:@2921.4]
  SingleCounter_1 ctrs_0 ( // @[Counter.scala 505:46:@2884.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done),
    .io_output_saturated(ctrs_0_io_output_saturated)
  );
  SingleCounter_2 ctrs_1 ( // @[Counter.scala 505:46:@2887.4]
    .clock(ctrs_1_clock),
    .reset(ctrs_1_reset),
    .io_setup_saturate(ctrs_1_io_setup_saturate),
    .io_input_reset(ctrs_1_io_input_reset),
    .io_input_enable(ctrs_1_io_input_enable),
    .io_output_count_0(ctrs_1_io_output_count_0),
    .io_output_oobs_0(ctrs_1_io_output_oobs_0),
    .io_output_done(ctrs_1_io_output_done)
  );
  assign isDone = ctrs_0_io_output_done & ctrs_1_io_output_done; // @[Counter.scala 533:51:@2904.4]
  assign _T_64 = io_input_enable & isDone; // @[Counter.scala 538:69:@2913.4]
  assign _T_66 = wasDone == 1'h0; // @[Counter.scala 538:80:@2914.4]
  assign _T_73 = isDone ? 1'h1 : doneLatch; // @[Counter.scala 543:48:@2920.4]
  assign _T_74 = io_input_reset ? 1'h0 : _T_73; // @[Counter.scala 543:19:@2921.4]
  assign io_output_counts_1 = ctrs_1_io_output_count_0; // @[Counter.scala 549:32:@2926.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 549:32:@2923.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 550:30:@2925.4]
  assign io_output_oobs_1 = ctrs_1_io_output_oobs_0 | doneLatch; // @[Counter.scala 550:30:@2928.4]
  assign io_output_done = _T_64 & _T_66; // @[Counter.scala 538:18:@2916.4]
  assign ctrs_0_clock = clock; // @[:@2885.4]
  assign ctrs_0_reset = reset; // @[:@2886.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 512:24:@2893.4]
  assign ctrs_0_io_input_enable = ctrs_1_io_output_done & io_input_enable; // @[Counter.scala 518:29:@2900.4]
  assign ctrs_1_clock = clock; // @[:@2888.4]
  assign ctrs_1_reset = reset; // @[:@2889.4]
  assign ctrs_1_io_setup_saturate = ctrs_0_io_output_saturated; // @[Counter.scala 524:31:@2903.4]
  assign ctrs_1_io_input_reset = io_input_reset; // @[Counter.scala 512:24:@2897.4]
  assign ctrs_1_io_input_enable = io_input_enable; // @[Counter.scala 516:33:@2898.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= isDone;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (isDone) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module RetimeWrapper_12( // @[:@2968.2]
  input   clock, // @[:@2969.4]
  input   reset, // @[:@2970.4]
  input   io_flow, // @[:@2971.4]
  input   io_in, // @[:@2971.4]
  output  io_out // @[:@2971.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(15)) sr ( // @[RetimeShiftRegister.scala 15:20:@2973.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@2986.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@2985.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@2984.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@2983.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@2982.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@2980.4]
endmodule
module RetimeWrapper_16( // @[:@3096.2]
  input   clock, // @[:@3097.4]
  input   reset, // @[:@3098.4]
  input   io_flow, // @[:@3099.4]
  input   io_in, // @[:@3099.4]
  output  io_out // @[:@3099.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(14)) sr ( // @[RetimeShiftRegister.scala 15:20:@3101.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3114.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3113.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3112.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3111.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3110.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3108.4]
endmodule
module x592_inr_Foreach_SAMPLER_BOX_sm( // @[:@3116.2]
  input   clock, // @[:@3117.4]
  input   reset, // @[:@3118.4]
  input   io_enable, // @[:@3119.4]
  output  io_done, // @[:@3119.4]
  output  io_doneLatch, // @[:@3119.4]
  input   io_ctrDone, // @[:@3119.4]
  output  io_datapathEn, // @[:@3119.4]
  output  io_ctrInc, // @[:@3119.4]
  output  io_ctrRst, // @[:@3119.4]
  input   io_parentAck, // @[:@3119.4]
  input   io_backpressure, // @[:@3119.4]
  input   io_break // @[:@3119.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@3121.4]
  wire  active_reset; // @[Controllers.scala 261:22:@3121.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@3121.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@3121.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@3121.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@3121.4]
  wire  done_clock; // @[Controllers.scala 262:20:@3124.4]
  wire  done_reset; // @[Controllers.scala 262:20:@3124.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@3124.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@3124.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@3124.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@3124.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3158.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3158.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3158.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@3158.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@3158.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@3180.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@3180.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@3180.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@3180.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@3180.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@3192.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@3192.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@3192.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@3192.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@3192.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@3200.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@3200.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@3200.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@3200.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@3200.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@3216.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@3216.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@3216.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@3216.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@3216.4]
  wire  _T_80; // @[Controllers.scala 264:48:@3129.4]
  wire  _T_81; // @[Controllers.scala 264:46:@3130.4]
  wire  _T_82; // @[Controllers.scala 264:62:@3131.4]
  wire  _T_83; // @[Controllers.scala 264:60:@3132.4]
  wire  _T_100; // @[package.scala 100:49:@3149.4]
  reg  _T_103; // @[package.scala 48:56:@3150.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@3163.4 package.scala 96:25:@3164.4]
  wire  _T_110; // @[package.scala 100:49:@3165.4]
  reg  _T_113; // @[package.scala 48:56:@3166.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@3168.4]
  wire  _T_118; // @[Controllers.scala 283:41:@3173.4]
  wire  _T_119; // @[Controllers.scala 283:59:@3174.4]
  wire  _T_121; // @[Controllers.scala 284:37:@3177.4]
  wire  _T_124; // @[package.scala 96:25:@3185.4 package.scala 96:25:@3186.4]
  wire  _T_126; // @[package.scala 100:49:@3187.4]
  reg  _T_129; // @[package.scala 48:56:@3188.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@3210.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@3212.4]
  reg  _T_153; // @[package.scala 48:56:@3213.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@3221.4 package.scala 96:25:@3222.4]
  wire  _T_158; // @[Controllers.scala 292:61:@3223.4]
  wire  _T_159; // @[Controllers.scala 292:24:@3224.4]
  SRFF active ( // @[Controllers.scala 261:22:@3121.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@3124.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_12 RetimeWrapper ( // @[package.scala 93:22:@3158.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_12 RetimeWrapper_1 ( // @[package.scala 93:22:@3180.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@3192.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@3200.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_16 RetimeWrapper_4 ( // @[package.scala 93:22:@3216.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@3129.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@3130.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@3131.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@3132.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@3149.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@3163.4 package.scala 96:25:@3164.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@3165.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@3168.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@3173.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@3174.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@3177.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@3185.4 package.scala 96:25:@3186.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@3187.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@3212.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@3221.4 package.scala 96:25:@3222.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@3223.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@3224.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@3191.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@3226.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@3176.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@3179.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@3171.4]
  assign active_clock = clock; // @[:@3122.4]
  assign active_reset = reset; // @[:@3123.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@3134.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@3138.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@3139.4]
  assign done_clock = clock; // @[:@3125.4]
  assign done_reset = reset; // @[:@3126.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@3154.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@3147.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@3148.4]
  assign RetimeWrapper_clock = clock; // @[:@3159.4]
  assign RetimeWrapper_reset = reset; // @[:@3160.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@3162.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@3161.4]
  assign RetimeWrapper_1_clock = clock; // @[:@3181.4]
  assign RetimeWrapper_1_reset = reset; // @[:@3182.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@3184.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@3183.4]
  assign RetimeWrapper_2_clock = clock; // @[:@3193.4]
  assign RetimeWrapper_2_reset = reset; // @[:@3194.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@3196.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@3195.4]
  assign RetimeWrapper_3_clock = clock; // @[:@3201.4]
  assign RetimeWrapper_3_reset = reset; // @[:@3202.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@3204.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@3203.4]
  assign RetimeWrapper_4_clock = clock; // @[:@3217.4]
  assign RetimeWrapper_4_reset = reset; // @[:@3218.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@3220.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@3219.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module SimBlackBoxesfix2fixBox( // @[:@3332.2]
  input  [31:0] io_a, // @[:@3335.4]
  output [31:0] io_b // @[:@3335.4]
);
  assign io_b = io_a; // @[SimBlackBoxes.scala 99:40:@3345.4]
endmodule
module _( // @[:@3347.2]
  input  [31:0] io_b, // @[:@3350.4]
  output [31:0] io_result // @[:@3350.4]
);
  wire [31:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@3355.4]
  wire [31:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@3355.4]
  SimBlackBoxesfix2fixBox SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@3355.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@3368.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@3363.4]
endmodule
module RetimeWrapper_21( // @[:@3452.2]
  input        clock, // @[:@3453.4]
  input        reset, // @[:@3454.4]
  input        io_flow, // @[:@3455.4]
  input  [7:0] io_in, // @[:@3455.4]
  output [7:0] io_out // @[:@3455.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@3457.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3470.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3469.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@3468.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3467.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3466.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3464.4]
endmodule
module Mem1D_4( // @[:@3472.2]
  input        clock, // @[:@3473.4]
  input        reset, // @[:@3474.4]
  input        io_r_ofs_0, // @[:@3475.4]
  input        io_r_backpressure, // @[:@3475.4]
  input        io_w_ofs_0, // @[:@3475.4]
  input  [7:0] io_w_data_0, // @[:@3475.4]
  input        io_w_en_0, // @[:@3475.4]
  output [7:0] io_output // @[:@3475.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3485.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3485.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3485.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@3485.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@3485.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@3494.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@3494.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@3494.4]
  wire [7:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@3494.4]
  wire [7:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@3494.4]
  reg [7:0] _T_127; // @[MemPrimitives.scala 560:26:@3479.4]
  reg [31:0] _RAND_0;
  wire  _T_130; // @[MemPrimitives.scala 561:61:@3481.4]
  wire  _T_131; // @[MemPrimitives.scala 561:44:@3482.4]
  wire [7:0] _T_132; // @[MemPrimitives.scala 561:19:@3483.4]
  wire  _T_135; // @[package.scala 96:25:@3490.4 package.scala 96:25:@3491.4]
  wire  _T_137; // @[Mux.scala 46:19:@3492.4]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@3485.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_1 ( // @[package.scala 93:22:@3494.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign _T_130 = io_w_ofs_0 == 1'h0; // @[MemPrimitives.scala 561:61:@3481.4]
  assign _T_131 = io_w_en_0 & _T_130; // @[MemPrimitives.scala 561:44:@3482.4]
  assign _T_132 = _T_131 ? io_w_data_0 : _T_127; // @[MemPrimitives.scala 561:19:@3483.4]
  assign _T_135 = RetimeWrapper_io_out; // @[package.scala 96:25:@3490.4 package.scala 96:25:@3491.4]
  assign _T_137 = 1'h0 == _T_135; // @[Mux.scala 46:19:@3492.4]
  assign io_output = RetimeWrapper_1_io_out; // @[MemPrimitives.scala 565:17:@3501.4]
  assign RetimeWrapper_clock = clock; // @[:@3486.4]
  assign RetimeWrapper_reset = reset; // @[:@3487.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@3489.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@3488.4]
  assign RetimeWrapper_1_clock = clock; // @[:@3495.4]
  assign RetimeWrapper_1_reset = reset; // @[:@3496.4]
  assign RetimeWrapper_1_io_flow = io_r_backpressure; // @[package.scala 95:18:@3498.4]
  assign RetimeWrapper_1_io_in = _T_137 ? _T_127 : 8'h0; // @[package.scala 94:16:@3497.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_127 = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_127 <= 8'h0;
    end else begin
      if (_T_131) begin
        _T_127 <= io_w_data_0;
      end
    end
  end
endmodule
module StickySelects( // @[:@4928.2]
  input   clock, // @[:@4929.4]
  input   reset, // @[:@4930.4]
  input   io_ins_0, // @[:@4931.4]
  input   io_ins_1, // @[:@4931.4]
  input   io_ins_2, // @[:@4931.4]
  output  io_outs_0, // @[:@4931.4]
  output  io_outs_1, // @[:@4931.4]
  output  io_outs_2 // @[:@4931.4]
);
  reg  _T_19; // @[StickySelects.scala 21:22:@4933.4]
  reg [31:0] _RAND_0;
  wire  _T_20; // @[StickySelects.scala 22:54:@4934.4]
  wire  _T_22; // @[StickySelects.scala 24:52:@4935.4]
  wire  _T_23; // @[StickySelects.scala 24:21:@4936.4]
  reg  _T_26; // @[StickySelects.scala 21:22:@4938.4]
  reg [31:0] _RAND_1;
  wire  _T_27; // @[StickySelects.scala 22:54:@4939.4]
  wire  _T_29; // @[StickySelects.scala 24:52:@4940.4]
  wire  _T_30; // @[StickySelects.scala 24:21:@4941.4]
  reg  _T_33; // @[StickySelects.scala 21:22:@4943.4]
  reg [31:0] _RAND_2;
  wire  _T_34; // @[StickySelects.scala 22:54:@4944.4]
  wire  _T_36; // @[StickySelects.scala 24:52:@4945.4]
  wire  _T_37; // @[StickySelects.scala 24:21:@4946.4]
  assign _T_20 = io_ins_1 | io_ins_2; // @[StickySelects.scala 22:54:@4934.4]
  assign _T_22 = io_ins_0 | _T_19; // @[StickySelects.scala 24:52:@4935.4]
  assign _T_23 = _T_20 ? 1'h0 : _T_22; // @[StickySelects.scala 24:21:@4936.4]
  assign _T_27 = io_ins_0 | io_ins_2; // @[StickySelects.scala 22:54:@4939.4]
  assign _T_29 = io_ins_1 | _T_26; // @[StickySelects.scala 24:52:@4940.4]
  assign _T_30 = _T_27 ? 1'h0 : _T_29; // @[StickySelects.scala 24:21:@4941.4]
  assign _T_34 = io_ins_0 | io_ins_1; // @[StickySelects.scala 22:54:@4944.4]
  assign _T_36 = io_ins_2 | _T_33; // @[StickySelects.scala 24:52:@4945.4]
  assign _T_37 = _T_34 ? 1'h0 : _T_36; // @[StickySelects.scala 24:21:@4946.4]
  assign io_outs_0 = _T_20 ? 1'h0 : _T_22; // @[StickySelects.scala 28:52:@4948.4]
  assign io_outs_1 = _T_27 ? 1'h0 : _T_29; // @[StickySelects.scala 28:52:@4949.4]
  assign io_outs_2 = _T_34 ? 1'h0 : _T_36; // @[StickySelects.scala 28:52:@4950.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_26 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_33 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (_T_20) begin
        _T_19 <= 1'h0;
      end else begin
        _T_19 <= _T_22;
      end
    end
    if (reset) begin
      _T_26 <= 1'h0;
    end else begin
      if (_T_27) begin
        _T_26 <= 1'h0;
      end else begin
        _T_26 <= _T_29;
      end
    end
    if (reset) begin
      _T_33 <= 1'h0;
    end else begin
      if (_T_34) begin
        _T_33 <= 1'h0;
      end else begin
        _T_33 <= _T_36;
      end
    end
  end
endmodule
module StickySelects_2( // @[:@4976.2]
  input   clock, // @[:@4977.4]
  input   reset, // @[:@4978.4]
  input   io_ins_0, // @[:@4979.4]
  input   io_ins_1, // @[:@4979.4]
  input   io_ins_2, // @[:@4979.4]
  input   io_ins_3, // @[:@4979.4]
  input   io_ins_4, // @[:@4979.4]
  input   io_ins_5, // @[:@4979.4]
  output  io_outs_0, // @[:@4979.4]
  output  io_outs_1, // @[:@4979.4]
  output  io_outs_2, // @[:@4979.4]
  output  io_outs_3, // @[:@4979.4]
  output  io_outs_4, // @[:@4979.4]
  output  io_outs_5 // @[:@4979.4]
);
  reg  _T_19; // @[StickySelects.scala 21:22:@4981.4]
  reg [31:0] _RAND_0;
  wire  _T_20; // @[StickySelects.scala 22:54:@4982.4]
  wire  _T_21; // @[StickySelects.scala 22:54:@4983.4]
  wire  _T_22; // @[StickySelects.scala 22:54:@4984.4]
  wire  _T_23; // @[StickySelects.scala 22:54:@4985.4]
  wire  _T_25; // @[StickySelects.scala 24:52:@4986.4]
  wire  _T_26; // @[StickySelects.scala 24:21:@4987.4]
  reg  _T_29; // @[StickySelects.scala 21:22:@4989.4]
  reg [31:0] _RAND_1;
  wire  _T_30; // @[StickySelects.scala 22:54:@4990.4]
  wire  _T_31; // @[StickySelects.scala 22:54:@4991.4]
  wire  _T_32; // @[StickySelects.scala 22:54:@4992.4]
  wire  _T_33; // @[StickySelects.scala 22:54:@4993.4]
  wire  _T_35; // @[StickySelects.scala 24:52:@4994.4]
  wire  _T_36; // @[StickySelects.scala 24:21:@4995.4]
  reg  _T_39; // @[StickySelects.scala 21:22:@4997.4]
  reg [31:0] _RAND_2;
  wire  _T_40; // @[StickySelects.scala 22:54:@4998.4]
  wire  _T_41; // @[StickySelects.scala 22:54:@4999.4]
  wire  _T_42; // @[StickySelects.scala 22:54:@5000.4]
  wire  _T_43; // @[StickySelects.scala 22:54:@5001.4]
  wire  _T_45; // @[StickySelects.scala 24:52:@5002.4]
  wire  _T_46; // @[StickySelects.scala 24:21:@5003.4]
  reg  _T_49; // @[StickySelects.scala 21:22:@5005.4]
  reg [31:0] _RAND_3;
  wire  _T_51; // @[StickySelects.scala 22:54:@5007.4]
  wire  _T_52; // @[StickySelects.scala 22:54:@5008.4]
  wire  _T_53; // @[StickySelects.scala 22:54:@5009.4]
  wire  _T_55; // @[StickySelects.scala 24:52:@5010.4]
  wire  _T_56; // @[StickySelects.scala 24:21:@5011.4]
  reg  _T_59; // @[StickySelects.scala 21:22:@5013.4]
  reg [31:0] _RAND_4;
  wire  _T_62; // @[StickySelects.scala 22:54:@5016.4]
  wire  _T_63; // @[StickySelects.scala 22:54:@5017.4]
  wire  _T_65; // @[StickySelects.scala 24:52:@5018.4]
  wire  _T_66; // @[StickySelects.scala 24:21:@5019.4]
  reg  _T_69; // @[StickySelects.scala 21:22:@5021.4]
  reg [31:0] _RAND_5;
  wire  _T_73; // @[StickySelects.scala 22:54:@5025.4]
  wire  _T_75; // @[StickySelects.scala 24:52:@5026.4]
  wire  _T_76; // @[StickySelects.scala 24:21:@5027.4]
  assign _T_20 = io_ins_1 | io_ins_2; // @[StickySelects.scala 22:54:@4982.4]
  assign _T_21 = _T_20 | io_ins_3; // @[StickySelects.scala 22:54:@4983.4]
  assign _T_22 = _T_21 | io_ins_4; // @[StickySelects.scala 22:54:@4984.4]
  assign _T_23 = _T_22 | io_ins_5; // @[StickySelects.scala 22:54:@4985.4]
  assign _T_25 = io_ins_0 | _T_19; // @[StickySelects.scala 24:52:@4986.4]
  assign _T_26 = _T_23 ? 1'h0 : _T_25; // @[StickySelects.scala 24:21:@4987.4]
  assign _T_30 = io_ins_0 | io_ins_2; // @[StickySelects.scala 22:54:@4990.4]
  assign _T_31 = _T_30 | io_ins_3; // @[StickySelects.scala 22:54:@4991.4]
  assign _T_32 = _T_31 | io_ins_4; // @[StickySelects.scala 22:54:@4992.4]
  assign _T_33 = _T_32 | io_ins_5; // @[StickySelects.scala 22:54:@4993.4]
  assign _T_35 = io_ins_1 | _T_29; // @[StickySelects.scala 24:52:@4994.4]
  assign _T_36 = _T_33 ? 1'h0 : _T_35; // @[StickySelects.scala 24:21:@4995.4]
  assign _T_40 = io_ins_0 | io_ins_1; // @[StickySelects.scala 22:54:@4998.4]
  assign _T_41 = _T_40 | io_ins_3; // @[StickySelects.scala 22:54:@4999.4]
  assign _T_42 = _T_41 | io_ins_4; // @[StickySelects.scala 22:54:@5000.4]
  assign _T_43 = _T_42 | io_ins_5; // @[StickySelects.scala 22:54:@5001.4]
  assign _T_45 = io_ins_2 | _T_39; // @[StickySelects.scala 24:52:@5002.4]
  assign _T_46 = _T_43 ? 1'h0 : _T_45; // @[StickySelects.scala 24:21:@5003.4]
  assign _T_51 = _T_40 | io_ins_2; // @[StickySelects.scala 22:54:@5007.4]
  assign _T_52 = _T_51 | io_ins_4; // @[StickySelects.scala 22:54:@5008.4]
  assign _T_53 = _T_52 | io_ins_5; // @[StickySelects.scala 22:54:@5009.4]
  assign _T_55 = io_ins_3 | _T_49; // @[StickySelects.scala 24:52:@5010.4]
  assign _T_56 = _T_53 ? 1'h0 : _T_55; // @[StickySelects.scala 24:21:@5011.4]
  assign _T_62 = _T_51 | io_ins_3; // @[StickySelects.scala 22:54:@5016.4]
  assign _T_63 = _T_62 | io_ins_5; // @[StickySelects.scala 22:54:@5017.4]
  assign _T_65 = io_ins_4 | _T_59; // @[StickySelects.scala 24:52:@5018.4]
  assign _T_66 = _T_63 ? 1'h0 : _T_65; // @[StickySelects.scala 24:21:@5019.4]
  assign _T_73 = _T_62 | io_ins_4; // @[StickySelects.scala 22:54:@5025.4]
  assign _T_75 = io_ins_5 | _T_69; // @[StickySelects.scala 24:52:@5026.4]
  assign _T_76 = _T_73 ? 1'h0 : _T_75; // @[StickySelects.scala 24:21:@5027.4]
  assign io_outs_0 = _T_23 ? 1'h0 : _T_25; // @[StickySelects.scala 28:52:@5029.4]
  assign io_outs_1 = _T_33 ? 1'h0 : _T_35; // @[StickySelects.scala 28:52:@5030.4]
  assign io_outs_2 = _T_43 ? 1'h0 : _T_45; // @[StickySelects.scala 28:52:@5031.4]
  assign io_outs_3 = _T_53 ? 1'h0 : _T_55; // @[StickySelects.scala 28:52:@5032.4]
  assign io_outs_4 = _T_63 ? 1'h0 : _T_65; // @[StickySelects.scala 28:52:@5033.4]
  assign io_outs_5 = _T_73 ? 1'h0 : _T_75; // @[StickySelects.scala 28:52:@5034.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_29 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_39 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_49 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_59 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_69 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (_T_23) begin
        _T_19 <= 1'h0;
      end else begin
        _T_19 <= _T_25;
      end
    end
    if (reset) begin
      _T_29 <= 1'h0;
    end else begin
      if (_T_33) begin
        _T_29 <= 1'h0;
      end else begin
        _T_29 <= _T_35;
      end
    end
    if (reset) begin
      _T_39 <= 1'h0;
    end else begin
      if (_T_43) begin
        _T_39 <= 1'h0;
      end else begin
        _T_39 <= _T_45;
      end
    end
    if (reset) begin
      _T_49 <= 1'h0;
    end else begin
      if (_T_53) begin
        _T_49 <= 1'h0;
      end else begin
        _T_49 <= _T_55;
      end
    end
    if (reset) begin
      _T_59 <= 1'h0;
    end else begin
      if (_T_63) begin
        _T_59 <= 1'h0;
      end else begin
        _T_59 <= _T_65;
      end
    end
    if (reset) begin
      _T_69 <= 1'h0;
    end else begin
      if (_T_73) begin
        _T_69 <= 1'h0;
      end else begin
        _T_69 <= _T_75;
      end
    end
  end
endmodule
module RetimeWrapper_52( // @[:@5612.2]
  input   clock, // @[:@5613.4]
  input   reset, // @[:@5614.4]
  input   io_flow, // @[:@5615.4]
  input   io_in, // @[:@5615.4]
  output  io_out // @[:@5615.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@5617.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@5617.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@5617.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@5617.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@5617.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@5617.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@5617.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@5630.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@5629.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@5628.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@5627.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@5626.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@5624.4]
endmodule
module x329_lb_0( // @[:@7904.2]
  input        clock, // @[:@7905.4]
  input        reset, // @[:@7906.4]
  input  [2:0] io_rPort_17_banks_0, // @[:@7907.4]
  input        io_rPort_17_ofs_0, // @[:@7907.4]
  input        io_rPort_17_en_0, // @[:@7907.4]
  input        io_rPort_17_backpressure, // @[:@7907.4]
  output [7:0] io_rPort_17_output_0, // @[:@7907.4]
  input  [2:0] io_rPort_16_banks_0, // @[:@7907.4]
  input        io_rPort_16_ofs_0, // @[:@7907.4]
  input        io_rPort_16_en_0, // @[:@7907.4]
  input        io_rPort_16_backpressure, // @[:@7907.4]
  output [7:0] io_rPort_16_output_0, // @[:@7907.4]
  input  [2:0] io_rPort_15_banks_0, // @[:@7907.4]
  input        io_rPort_15_ofs_0, // @[:@7907.4]
  input        io_rPort_15_en_0, // @[:@7907.4]
  input        io_rPort_15_backpressure, // @[:@7907.4]
  output [7:0] io_rPort_15_output_0, // @[:@7907.4]
  input  [2:0] io_rPort_14_banks_0, // @[:@7907.4]
  input        io_rPort_14_ofs_0, // @[:@7907.4]
  input        io_rPort_14_en_0, // @[:@7907.4]
  input        io_rPort_14_backpressure, // @[:@7907.4]
  output [7:0] io_rPort_14_output_0, // @[:@7907.4]
  input  [2:0] io_rPort_13_banks_0, // @[:@7907.4]
  input        io_rPort_13_ofs_0, // @[:@7907.4]
  input        io_rPort_13_en_0, // @[:@7907.4]
  input        io_rPort_13_backpressure, // @[:@7907.4]
  output [7:0] io_rPort_13_output_0, // @[:@7907.4]
  input  [2:0] io_rPort_12_banks_0, // @[:@7907.4]
  input        io_rPort_12_ofs_0, // @[:@7907.4]
  input        io_rPort_12_en_0, // @[:@7907.4]
  input        io_rPort_12_backpressure, // @[:@7907.4]
  output [7:0] io_rPort_12_output_0, // @[:@7907.4]
  input  [2:0] io_rPort_11_banks_0, // @[:@7907.4]
  input        io_rPort_11_ofs_0, // @[:@7907.4]
  input        io_rPort_11_en_0, // @[:@7907.4]
  input        io_rPort_11_backpressure, // @[:@7907.4]
  output [7:0] io_rPort_11_output_0, // @[:@7907.4]
  input  [2:0] io_rPort_10_banks_0, // @[:@7907.4]
  input        io_rPort_10_ofs_0, // @[:@7907.4]
  input        io_rPort_10_en_0, // @[:@7907.4]
  input        io_rPort_10_backpressure, // @[:@7907.4]
  output [7:0] io_rPort_10_output_0, // @[:@7907.4]
  input  [2:0] io_rPort_9_banks_0, // @[:@7907.4]
  input        io_rPort_9_ofs_0, // @[:@7907.4]
  input        io_rPort_9_en_0, // @[:@7907.4]
  input        io_rPort_9_backpressure, // @[:@7907.4]
  output [7:0] io_rPort_9_output_0, // @[:@7907.4]
  input  [2:0] io_rPort_8_banks_0, // @[:@7907.4]
  input        io_rPort_8_ofs_0, // @[:@7907.4]
  input        io_rPort_8_en_0, // @[:@7907.4]
  input        io_rPort_8_backpressure, // @[:@7907.4]
  output [7:0] io_rPort_8_output_0, // @[:@7907.4]
  input  [2:0] io_rPort_7_banks_0, // @[:@7907.4]
  input        io_rPort_7_ofs_0, // @[:@7907.4]
  input        io_rPort_7_en_0, // @[:@7907.4]
  input        io_rPort_7_backpressure, // @[:@7907.4]
  output [7:0] io_rPort_7_output_0, // @[:@7907.4]
  input  [2:0] io_rPort_6_banks_0, // @[:@7907.4]
  input        io_rPort_6_ofs_0, // @[:@7907.4]
  input        io_rPort_6_en_0, // @[:@7907.4]
  input        io_rPort_6_backpressure, // @[:@7907.4]
  output [7:0] io_rPort_6_output_0, // @[:@7907.4]
  input  [2:0] io_rPort_5_banks_0, // @[:@7907.4]
  input        io_rPort_5_ofs_0, // @[:@7907.4]
  input        io_rPort_5_en_0, // @[:@7907.4]
  input        io_rPort_5_backpressure, // @[:@7907.4]
  output [7:0] io_rPort_5_output_0, // @[:@7907.4]
  input  [2:0] io_rPort_4_banks_0, // @[:@7907.4]
  input        io_rPort_4_ofs_0, // @[:@7907.4]
  input        io_rPort_4_en_0, // @[:@7907.4]
  input        io_rPort_4_backpressure, // @[:@7907.4]
  output [7:0] io_rPort_4_output_0, // @[:@7907.4]
  input  [2:0] io_rPort_3_banks_0, // @[:@7907.4]
  input        io_rPort_3_ofs_0, // @[:@7907.4]
  input        io_rPort_3_en_0, // @[:@7907.4]
  input        io_rPort_3_backpressure, // @[:@7907.4]
  output [7:0] io_rPort_3_output_0, // @[:@7907.4]
  input  [2:0] io_rPort_2_banks_0, // @[:@7907.4]
  input        io_rPort_2_ofs_0, // @[:@7907.4]
  input        io_rPort_2_en_0, // @[:@7907.4]
  input        io_rPort_2_backpressure, // @[:@7907.4]
  output [7:0] io_rPort_2_output_0, // @[:@7907.4]
  input  [2:0] io_rPort_1_banks_0, // @[:@7907.4]
  input        io_rPort_1_ofs_0, // @[:@7907.4]
  input        io_rPort_1_en_0, // @[:@7907.4]
  input        io_rPort_1_backpressure, // @[:@7907.4]
  output [7:0] io_rPort_1_output_0, // @[:@7907.4]
  input  [2:0] io_rPort_0_banks_0, // @[:@7907.4]
  input        io_rPort_0_ofs_0, // @[:@7907.4]
  input        io_rPort_0_en_0, // @[:@7907.4]
  input        io_rPort_0_backpressure, // @[:@7907.4]
  output [7:0] io_rPort_0_output_0, // @[:@7907.4]
  input  [2:0] io_wPort_3_banks_0, // @[:@7907.4]
  input        io_wPort_3_ofs_0, // @[:@7907.4]
  input  [7:0] io_wPort_3_data_0, // @[:@7907.4]
  input        io_wPort_3_en_0, // @[:@7907.4]
  input  [2:0] io_wPort_2_banks_0, // @[:@7907.4]
  input        io_wPort_2_ofs_0, // @[:@7907.4]
  input  [7:0] io_wPort_2_data_0, // @[:@7907.4]
  input        io_wPort_2_en_0, // @[:@7907.4]
  input  [2:0] io_wPort_1_banks_0, // @[:@7907.4]
  input        io_wPort_1_ofs_0, // @[:@7907.4]
  input  [7:0] io_wPort_1_data_0, // @[:@7907.4]
  input        io_wPort_1_en_0, // @[:@7907.4]
  input  [2:0] io_wPort_0_banks_0, // @[:@7907.4]
  input        io_wPort_0_ofs_0, // @[:@7907.4]
  input  [7:0] io_wPort_0_data_0, // @[:@7907.4]
  input        io_wPort_0_en_0 // @[:@7907.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@8050.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@8050.4]
  wire  Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@8050.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@8050.4]
  wire  Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@8050.4]
  wire [7:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@8050.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@8050.4]
  wire [7:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@8050.4]
  wire  Mem1D_1_clock; // @[MemPrimitives.scala 64:21:@8066.4]
  wire  Mem1D_1_reset; // @[MemPrimitives.scala 64:21:@8066.4]
  wire  Mem1D_1_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@8066.4]
  wire  Mem1D_1_io_r_backpressure; // @[MemPrimitives.scala 64:21:@8066.4]
  wire  Mem1D_1_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@8066.4]
  wire [7:0] Mem1D_1_io_w_data_0; // @[MemPrimitives.scala 64:21:@8066.4]
  wire  Mem1D_1_io_w_en_0; // @[MemPrimitives.scala 64:21:@8066.4]
  wire [7:0] Mem1D_1_io_output; // @[MemPrimitives.scala 64:21:@8066.4]
  wire  Mem1D_2_clock; // @[MemPrimitives.scala 64:21:@8082.4]
  wire  Mem1D_2_reset; // @[MemPrimitives.scala 64:21:@8082.4]
  wire  Mem1D_2_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@8082.4]
  wire  Mem1D_2_io_r_backpressure; // @[MemPrimitives.scala 64:21:@8082.4]
  wire  Mem1D_2_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@8082.4]
  wire [7:0] Mem1D_2_io_w_data_0; // @[MemPrimitives.scala 64:21:@8082.4]
  wire  Mem1D_2_io_w_en_0; // @[MemPrimitives.scala 64:21:@8082.4]
  wire [7:0] Mem1D_2_io_output; // @[MemPrimitives.scala 64:21:@8082.4]
  wire  Mem1D_3_clock; // @[MemPrimitives.scala 64:21:@8098.4]
  wire  Mem1D_3_reset; // @[MemPrimitives.scala 64:21:@8098.4]
  wire  Mem1D_3_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@8098.4]
  wire  Mem1D_3_io_r_backpressure; // @[MemPrimitives.scala 64:21:@8098.4]
  wire  Mem1D_3_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@8098.4]
  wire [7:0] Mem1D_3_io_w_data_0; // @[MemPrimitives.scala 64:21:@8098.4]
  wire  Mem1D_3_io_w_en_0; // @[MemPrimitives.scala 64:21:@8098.4]
  wire [7:0] Mem1D_3_io_output; // @[MemPrimitives.scala 64:21:@8098.4]
  wire  Mem1D_4_clock; // @[MemPrimitives.scala 64:21:@8114.4]
  wire  Mem1D_4_reset; // @[MemPrimitives.scala 64:21:@8114.4]
  wire  Mem1D_4_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@8114.4]
  wire  Mem1D_4_io_r_backpressure; // @[MemPrimitives.scala 64:21:@8114.4]
  wire  Mem1D_4_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@8114.4]
  wire [7:0] Mem1D_4_io_w_data_0; // @[MemPrimitives.scala 64:21:@8114.4]
  wire  Mem1D_4_io_w_en_0; // @[MemPrimitives.scala 64:21:@8114.4]
  wire [7:0] Mem1D_4_io_output; // @[MemPrimitives.scala 64:21:@8114.4]
  wire  Mem1D_5_clock; // @[MemPrimitives.scala 64:21:@8130.4]
  wire  Mem1D_5_reset; // @[MemPrimitives.scala 64:21:@8130.4]
  wire  Mem1D_5_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@8130.4]
  wire  Mem1D_5_io_r_backpressure; // @[MemPrimitives.scala 64:21:@8130.4]
  wire  Mem1D_5_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@8130.4]
  wire [7:0] Mem1D_5_io_w_data_0; // @[MemPrimitives.scala 64:21:@8130.4]
  wire  Mem1D_5_io_w_en_0; // @[MemPrimitives.scala 64:21:@8130.4]
  wire [7:0] Mem1D_5_io_output; // @[MemPrimitives.scala 64:21:@8130.4]
  wire  Mem1D_6_clock; // @[MemPrimitives.scala 64:21:@8146.4]
  wire  Mem1D_6_reset; // @[MemPrimitives.scala 64:21:@8146.4]
  wire  Mem1D_6_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@8146.4]
  wire  Mem1D_6_io_r_backpressure; // @[MemPrimitives.scala 64:21:@8146.4]
  wire  Mem1D_6_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@8146.4]
  wire [7:0] Mem1D_6_io_w_data_0; // @[MemPrimitives.scala 64:21:@8146.4]
  wire  Mem1D_6_io_w_en_0; // @[MemPrimitives.scala 64:21:@8146.4]
  wire [7:0] Mem1D_6_io_output; // @[MemPrimitives.scala 64:21:@8146.4]
  wire  Mem1D_7_clock; // @[MemPrimitives.scala 64:21:@8162.4]
  wire  Mem1D_7_reset; // @[MemPrimitives.scala 64:21:@8162.4]
  wire  Mem1D_7_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@8162.4]
  wire  Mem1D_7_io_r_backpressure; // @[MemPrimitives.scala 64:21:@8162.4]
  wire  Mem1D_7_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@8162.4]
  wire [7:0] Mem1D_7_io_w_data_0; // @[MemPrimitives.scala 64:21:@8162.4]
  wire  Mem1D_7_io_w_en_0; // @[MemPrimitives.scala 64:21:@8162.4]
  wire [7:0] Mem1D_7_io_output; // @[MemPrimitives.scala 64:21:@8162.4]
  wire  Mem1D_8_clock; // @[MemPrimitives.scala 64:21:@8178.4]
  wire  Mem1D_8_reset; // @[MemPrimitives.scala 64:21:@8178.4]
  wire  Mem1D_8_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@8178.4]
  wire  Mem1D_8_io_r_backpressure; // @[MemPrimitives.scala 64:21:@8178.4]
  wire  Mem1D_8_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@8178.4]
  wire [7:0] Mem1D_8_io_w_data_0; // @[MemPrimitives.scala 64:21:@8178.4]
  wire  Mem1D_8_io_w_en_0; // @[MemPrimitives.scala 64:21:@8178.4]
  wire [7:0] Mem1D_8_io_output; // @[MemPrimitives.scala 64:21:@8178.4]
  wire  Mem1D_9_clock; // @[MemPrimitives.scala 64:21:@8194.4]
  wire  Mem1D_9_reset; // @[MemPrimitives.scala 64:21:@8194.4]
  wire  Mem1D_9_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@8194.4]
  wire  Mem1D_9_io_r_backpressure; // @[MemPrimitives.scala 64:21:@8194.4]
  wire  Mem1D_9_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@8194.4]
  wire [7:0] Mem1D_9_io_w_data_0; // @[MemPrimitives.scala 64:21:@8194.4]
  wire  Mem1D_9_io_w_en_0; // @[MemPrimitives.scala 64:21:@8194.4]
  wire [7:0] Mem1D_9_io_output; // @[MemPrimitives.scala 64:21:@8194.4]
  wire  Mem1D_10_clock; // @[MemPrimitives.scala 64:21:@8210.4]
  wire  Mem1D_10_reset; // @[MemPrimitives.scala 64:21:@8210.4]
  wire  Mem1D_10_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@8210.4]
  wire  Mem1D_10_io_r_backpressure; // @[MemPrimitives.scala 64:21:@8210.4]
  wire  Mem1D_10_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@8210.4]
  wire [7:0] Mem1D_10_io_w_data_0; // @[MemPrimitives.scala 64:21:@8210.4]
  wire  Mem1D_10_io_w_en_0; // @[MemPrimitives.scala 64:21:@8210.4]
  wire [7:0] Mem1D_10_io_output; // @[MemPrimitives.scala 64:21:@8210.4]
  wire  Mem1D_11_clock; // @[MemPrimitives.scala 64:21:@8226.4]
  wire  Mem1D_11_reset; // @[MemPrimitives.scala 64:21:@8226.4]
  wire  Mem1D_11_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@8226.4]
  wire  Mem1D_11_io_r_backpressure; // @[MemPrimitives.scala 64:21:@8226.4]
  wire  Mem1D_11_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@8226.4]
  wire [7:0] Mem1D_11_io_w_data_0; // @[MemPrimitives.scala 64:21:@8226.4]
  wire  Mem1D_11_io_w_en_0; // @[MemPrimitives.scala 64:21:@8226.4]
  wire [7:0] Mem1D_11_io_output; // @[MemPrimitives.scala 64:21:@8226.4]
  wire  Mem1D_12_clock; // @[MemPrimitives.scala 64:21:@8242.4]
  wire  Mem1D_12_reset; // @[MemPrimitives.scala 64:21:@8242.4]
  wire  Mem1D_12_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@8242.4]
  wire  Mem1D_12_io_r_backpressure; // @[MemPrimitives.scala 64:21:@8242.4]
  wire  Mem1D_12_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@8242.4]
  wire [7:0] Mem1D_12_io_w_data_0; // @[MemPrimitives.scala 64:21:@8242.4]
  wire  Mem1D_12_io_w_en_0; // @[MemPrimitives.scala 64:21:@8242.4]
  wire [7:0] Mem1D_12_io_output; // @[MemPrimitives.scala 64:21:@8242.4]
  wire  Mem1D_13_clock; // @[MemPrimitives.scala 64:21:@8258.4]
  wire  Mem1D_13_reset; // @[MemPrimitives.scala 64:21:@8258.4]
  wire  Mem1D_13_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@8258.4]
  wire  Mem1D_13_io_r_backpressure; // @[MemPrimitives.scala 64:21:@8258.4]
  wire  Mem1D_13_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@8258.4]
  wire [7:0] Mem1D_13_io_w_data_0; // @[MemPrimitives.scala 64:21:@8258.4]
  wire  Mem1D_13_io_w_en_0; // @[MemPrimitives.scala 64:21:@8258.4]
  wire [7:0] Mem1D_13_io_output; // @[MemPrimitives.scala 64:21:@8258.4]
  wire  Mem1D_14_clock; // @[MemPrimitives.scala 64:21:@8274.4]
  wire  Mem1D_14_reset; // @[MemPrimitives.scala 64:21:@8274.4]
  wire  Mem1D_14_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@8274.4]
  wire  Mem1D_14_io_r_backpressure; // @[MemPrimitives.scala 64:21:@8274.4]
  wire  Mem1D_14_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@8274.4]
  wire [7:0] Mem1D_14_io_w_data_0; // @[MemPrimitives.scala 64:21:@8274.4]
  wire  Mem1D_14_io_w_en_0; // @[MemPrimitives.scala 64:21:@8274.4]
  wire [7:0] Mem1D_14_io_output; // @[MemPrimitives.scala 64:21:@8274.4]
  wire  Mem1D_15_clock; // @[MemPrimitives.scala 64:21:@8290.4]
  wire  Mem1D_15_reset; // @[MemPrimitives.scala 64:21:@8290.4]
  wire  Mem1D_15_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@8290.4]
  wire  Mem1D_15_io_r_backpressure; // @[MemPrimitives.scala 64:21:@8290.4]
  wire  Mem1D_15_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@8290.4]
  wire [7:0] Mem1D_15_io_w_data_0; // @[MemPrimitives.scala 64:21:@8290.4]
  wire  Mem1D_15_io_w_en_0; // @[MemPrimitives.scala 64:21:@8290.4]
  wire [7:0] Mem1D_15_io_output; // @[MemPrimitives.scala 64:21:@8290.4]
  wire  StickySelects_clock; // @[MemPrimitives.scala 121:29:@8491.4]
  wire  StickySelects_reset; // @[MemPrimitives.scala 121:29:@8491.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 121:29:@8491.4]
  wire  StickySelects_io_ins_1; // @[MemPrimitives.scala 121:29:@8491.4]
  wire  StickySelects_io_ins_2; // @[MemPrimitives.scala 121:29:@8491.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 121:29:@8491.4]
  wire  StickySelects_io_outs_1; // @[MemPrimitives.scala 121:29:@8491.4]
  wire  StickySelects_io_outs_2; // @[MemPrimitives.scala 121:29:@8491.4]
  wire  StickySelects_1_clock; // @[MemPrimitives.scala 121:29:@8523.4]
  wire  StickySelects_1_reset; // @[MemPrimitives.scala 121:29:@8523.4]
  wire  StickySelects_1_io_ins_0; // @[MemPrimitives.scala 121:29:@8523.4]
  wire  StickySelects_1_io_ins_1; // @[MemPrimitives.scala 121:29:@8523.4]
  wire  StickySelects_1_io_ins_2; // @[MemPrimitives.scala 121:29:@8523.4]
  wire  StickySelects_1_io_outs_0; // @[MemPrimitives.scala 121:29:@8523.4]
  wire  StickySelects_1_io_outs_1; // @[MemPrimitives.scala 121:29:@8523.4]
  wire  StickySelects_1_io_outs_2; // @[MemPrimitives.scala 121:29:@8523.4]
  wire  StickySelects_2_clock; // @[MemPrimitives.scala 121:29:@8564.4]
  wire  StickySelects_2_reset; // @[MemPrimitives.scala 121:29:@8564.4]
  wire  StickySelects_2_io_ins_0; // @[MemPrimitives.scala 121:29:@8564.4]
  wire  StickySelects_2_io_ins_1; // @[MemPrimitives.scala 121:29:@8564.4]
  wire  StickySelects_2_io_ins_2; // @[MemPrimitives.scala 121:29:@8564.4]
  wire  StickySelects_2_io_ins_3; // @[MemPrimitives.scala 121:29:@8564.4]
  wire  StickySelects_2_io_ins_4; // @[MemPrimitives.scala 121:29:@8564.4]
  wire  StickySelects_2_io_ins_5; // @[MemPrimitives.scala 121:29:@8564.4]
  wire  StickySelects_2_io_outs_0; // @[MemPrimitives.scala 121:29:@8564.4]
  wire  StickySelects_2_io_outs_1; // @[MemPrimitives.scala 121:29:@8564.4]
  wire  StickySelects_2_io_outs_2; // @[MemPrimitives.scala 121:29:@8564.4]
  wire  StickySelects_2_io_outs_3; // @[MemPrimitives.scala 121:29:@8564.4]
  wire  StickySelects_2_io_outs_4; // @[MemPrimitives.scala 121:29:@8564.4]
  wire  StickySelects_2_io_outs_5; // @[MemPrimitives.scala 121:29:@8564.4]
  wire  StickySelects_3_clock; // @[MemPrimitives.scala 121:29:@8620.4]
  wire  StickySelects_3_reset; // @[MemPrimitives.scala 121:29:@8620.4]
  wire  StickySelects_3_io_ins_0; // @[MemPrimitives.scala 121:29:@8620.4]
  wire  StickySelects_3_io_ins_1; // @[MemPrimitives.scala 121:29:@8620.4]
  wire  StickySelects_3_io_ins_2; // @[MemPrimitives.scala 121:29:@8620.4]
  wire  StickySelects_3_io_ins_3; // @[MemPrimitives.scala 121:29:@8620.4]
  wire  StickySelects_3_io_ins_4; // @[MemPrimitives.scala 121:29:@8620.4]
  wire  StickySelects_3_io_ins_5; // @[MemPrimitives.scala 121:29:@8620.4]
  wire  StickySelects_3_io_outs_0; // @[MemPrimitives.scala 121:29:@8620.4]
  wire  StickySelects_3_io_outs_1; // @[MemPrimitives.scala 121:29:@8620.4]
  wire  StickySelects_3_io_outs_2; // @[MemPrimitives.scala 121:29:@8620.4]
  wire  StickySelects_3_io_outs_3; // @[MemPrimitives.scala 121:29:@8620.4]
  wire  StickySelects_3_io_outs_4; // @[MemPrimitives.scala 121:29:@8620.4]
  wire  StickySelects_3_io_outs_5; // @[MemPrimitives.scala 121:29:@8620.4]
  wire  StickySelects_4_clock; // @[MemPrimitives.scala 121:29:@8667.4]
  wire  StickySelects_4_reset; // @[MemPrimitives.scala 121:29:@8667.4]
  wire  StickySelects_4_io_ins_0; // @[MemPrimitives.scala 121:29:@8667.4]
  wire  StickySelects_4_io_ins_1; // @[MemPrimitives.scala 121:29:@8667.4]
  wire  StickySelects_4_io_ins_2; // @[MemPrimitives.scala 121:29:@8667.4]
  wire  StickySelects_4_io_outs_0; // @[MemPrimitives.scala 121:29:@8667.4]
  wire  StickySelects_4_io_outs_1; // @[MemPrimitives.scala 121:29:@8667.4]
  wire  StickySelects_4_io_outs_2; // @[MemPrimitives.scala 121:29:@8667.4]
  wire  StickySelects_5_clock; // @[MemPrimitives.scala 121:29:@8699.4]
  wire  StickySelects_5_reset; // @[MemPrimitives.scala 121:29:@8699.4]
  wire  StickySelects_5_io_ins_0; // @[MemPrimitives.scala 121:29:@8699.4]
  wire  StickySelects_5_io_ins_1; // @[MemPrimitives.scala 121:29:@8699.4]
  wire  StickySelects_5_io_ins_2; // @[MemPrimitives.scala 121:29:@8699.4]
  wire  StickySelects_5_io_outs_0; // @[MemPrimitives.scala 121:29:@8699.4]
  wire  StickySelects_5_io_outs_1; // @[MemPrimitives.scala 121:29:@8699.4]
  wire  StickySelects_5_io_outs_2; // @[MemPrimitives.scala 121:29:@8699.4]
  wire  StickySelects_6_clock; // @[MemPrimitives.scala 121:29:@8740.4]
  wire  StickySelects_6_reset; // @[MemPrimitives.scala 121:29:@8740.4]
  wire  StickySelects_6_io_ins_0; // @[MemPrimitives.scala 121:29:@8740.4]
  wire  StickySelects_6_io_ins_1; // @[MemPrimitives.scala 121:29:@8740.4]
  wire  StickySelects_6_io_ins_2; // @[MemPrimitives.scala 121:29:@8740.4]
  wire  StickySelects_6_io_ins_3; // @[MemPrimitives.scala 121:29:@8740.4]
  wire  StickySelects_6_io_ins_4; // @[MemPrimitives.scala 121:29:@8740.4]
  wire  StickySelects_6_io_ins_5; // @[MemPrimitives.scala 121:29:@8740.4]
  wire  StickySelects_6_io_outs_0; // @[MemPrimitives.scala 121:29:@8740.4]
  wire  StickySelects_6_io_outs_1; // @[MemPrimitives.scala 121:29:@8740.4]
  wire  StickySelects_6_io_outs_2; // @[MemPrimitives.scala 121:29:@8740.4]
  wire  StickySelects_6_io_outs_3; // @[MemPrimitives.scala 121:29:@8740.4]
  wire  StickySelects_6_io_outs_4; // @[MemPrimitives.scala 121:29:@8740.4]
  wire  StickySelects_6_io_outs_5; // @[MemPrimitives.scala 121:29:@8740.4]
  wire  StickySelects_7_clock; // @[MemPrimitives.scala 121:29:@8796.4]
  wire  StickySelects_7_reset; // @[MemPrimitives.scala 121:29:@8796.4]
  wire  StickySelects_7_io_ins_0; // @[MemPrimitives.scala 121:29:@8796.4]
  wire  StickySelects_7_io_ins_1; // @[MemPrimitives.scala 121:29:@8796.4]
  wire  StickySelects_7_io_ins_2; // @[MemPrimitives.scala 121:29:@8796.4]
  wire  StickySelects_7_io_ins_3; // @[MemPrimitives.scala 121:29:@8796.4]
  wire  StickySelects_7_io_ins_4; // @[MemPrimitives.scala 121:29:@8796.4]
  wire  StickySelects_7_io_ins_5; // @[MemPrimitives.scala 121:29:@8796.4]
  wire  StickySelects_7_io_outs_0; // @[MemPrimitives.scala 121:29:@8796.4]
  wire  StickySelects_7_io_outs_1; // @[MemPrimitives.scala 121:29:@8796.4]
  wire  StickySelects_7_io_outs_2; // @[MemPrimitives.scala 121:29:@8796.4]
  wire  StickySelects_7_io_outs_3; // @[MemPrimitives.scala 121:29:@8796.4]
  wire  StickySelects_7_io_outs_4; // @[MemPrimitives.scala 121:29:@8796.4]
  wire  StickySelects_7_io_outs_5; // @[MemPrimitives.scala 121:29:@8796.4]
  wire  StickySelects_8_clock; // @[MemPrimitives.scala 121:29:@8843.4]
  wire  StickySelects_8_reset; // @[MemPrimitives.scala 121:29:@8843.4]
  wire  StickySelects_8_io_ins_0; // @[MemPrimitives.scala 121:29:@8843.4]
  wire  StickySelects_8_io_ins_1; // @[MemPrimitives.scala 121:29:@8843.4]
  wire  StickySelects_8_io_ins_2; // @[MemPrimitives.scala 121:29:@8843.4]
  wire  StickySelects_8_io_outs_0; // @[MemPrimitives.scala 121:29:@8843.4]
  wire  StickySelects_8_io_outs_1; // @[MemPrimitives.scala 121:29:@8843.4]
  wire  StickySelects_8_io_outs_2; // @[MemPrimitives.scala 121:29:@8843.4]
  wire  StickySelects_9_clock; // @[MemPrimitives.scala 121:29:@8875.4]
  wire  StickySelects_9_reset; // @[MemPrimitives.scala 121:29:@8875.4]
  wire  StickySelects_9_io_ins_0; // @[MemPrimitives.scala 121:29:@8875.4]
  wire  StickySelects_9_io_ins_1; // @[MemPrimitives.scala 121:29:@8875.4]
  wire  StickySelects_9_io_ins_2; // @[MemPrimitives.scala 121:29:@8875.4]
  wire  StickySelects_9_io_outs_0; // @[MemPrimitives.scala 121:29:@8875.4]
  wire  StickySelects_9_io_outs_1; // @[MemPrimitives.scala 121:29:@8875.4]
  wire  StickySelects_9_io_outs_2; // @[MemPrimitives.scala 121:29:@8875.4]
  wire  StickySelects_10_clock; // @[MemPrimitives.scala 121:29:@8916.4]
  wire  StickySelects_10_reset; // @[MemPrimitives.scala 121:29:@8916.4]
  wire  StickySelects_10_io_ins_0; // @[MemPrimitives.scala 121:29:@8916.4]
  wire  StickySelects_10_io_ins_1; // @[MemPrimitives.scala 121:29:@8916.4]
  wire  StickySelects_10_io_ins_2; // @[MemPrimitives.scala 121:29:@8916.4]
  wire  StickySelects_10_io_ins_3; // @[MemPrimitives.scala 121:29:@8916.4]
  wire  StickySelects_10_io_ins_4; // @[MemPrimitives.scala 121:29:@8916.4]
  wire  StickySelects_10_io_ins_5; // @[MemPrimitives.scala 121:29:@8916.4]
  wire  StickySelects_10_io_outs_0; // @[MemPrimitives.scala 121:29:@8916.4]
  wire  StickySelects_10_io_outs_1; // @[MemPrimitives.scala 121:29:@8916.4]
  wire  StickySelects_10_io_outs_2; // @[MemPrimitives.scala 121:29:@8916.4]
  wire  StickySelects_10_io_outs_3; // @[MemPrimitives.scala 121:29:@8916.4]
  wire  StickySelects_10_io_outs_4; // @[MemPrimitives.scala 121:29:@8916.4]
  wire  StickySelects_10_io_outs_5; // @[MemPrimitives.scala 121:29:@8916.4]
  wire  StickySelects_11_clock; // @[MemPrimitives.scala 121:29:@8972.4]
  wire  StickySelects_11_reset; // @[MemPrimitives.scala 121:29:@8972.4]
  wire  StickySelects_11_io_ins_0; // @[MemPrimitives.scala 121:29:@8972.4]
  wire  StickySelects_11_io_ins_1; // @[MemPrimitives.scala 121:29:@8972.4]
  wire  StickySelects_11_io_ins_2; // @[MemPrimitives.scala 121:29:@8972.4]
  wire  StickySelects_11_io_ins_3; // @[MemPrimitives.scala 121:29:@8972.4]
  wire  StickySelects_11_io_ins_4; // @[MemPrimitives.scala 121:29:@8972.4]
  wire  StickySelects_11_io_ins_5; // @[MemPrimitives.scala 121:29:@8972.4]
  wire  StickySelects_11_io_outs_0; // @[MemPrimitives.scala 121:29:@8972.4]
  wire  StickySelects_11_io_outs_1; // @[MemPrimitives.scala 121:29:@8972.4]
  wire  StickySelects_11_io_outs_2; // @[MemPrimitives.scala 121:29:@8972.4]
  wire  StickySelects_11_io_outs_3; // @[MemPrimitives.scala 121:29:@8972.4]
  wire  StickySelects_11_io_outs_4; // @[MemPrimitives.scala 121:29:@8972.4]
  wire  StickySelects_11_io_outs_5; // @[MemPrimitives.scala 121:29:@8972.4]
  wire  StickySelects_12_clock; // @[MemPrimitives.scala 121:29:@9019.4]
  wire  StickySelects_12_reset; // @[MemPrimitives.scala 121:29:@9019.4]
  wire  StickySelects_12_io_ins_0; // @[MemPrimitives.scala 121:29:@9019.4]
  wire  StickySelects_12_io_ins_1; // @[MemPrimitives.scala 121:29:@9019.4]
  wire  StickySelects_12_io_ins_2; // @[MemPrimitives.scala 121:29:@9019.4]
  wire  StickySelects_12_io_outs_0; // @[MemPrimitives.scala 121:29:@9019.4]
  wire  StickySelects_12_io_outs_1; // @[MemPrimitives.scala 121:29:@9019.4]
  wire  StickySelects_12_io_outs_2; // @[MemPrimitives.scala 121:29:@9019.4]
  wire  StickySelects_13_clock; // @[MemPrimitives.scala 121:29:@9051.4]
  wire  StickySelects_13_reset; // @[MemPrimitives.scala 121:29:@9051.4]
  wire  StickySelects_13_io_ins_0; // @[MemPrimitives.scala 121:29:@9051.4]
  wire  StickySelects_13_io_ins_1; // @[MemPrimitives.scala 121:29:@9051.4]
  wire  StickySelects_13_io_ins_2; // @[MemPrimitives.scala 121:29:@9051.4]
  wire  StickySelects_13_io_outs_0; // @[MemPrimitives.scala 121:29:@9051.4]
  wire  StickySelects_13_io_outs_1; // @[MemPrimitives.scala 121:29:@9051.4]
  wire  StickySelects_13_io_outs_2; // @[MemPrimitives.scala 121:29:@9051.4]
  wire  StickySelects_14_clock; // @[MemPrimitives.scala 121:29:@9092.4]
  wire  StickySelects_14_reset; // @[MemPrimitives.scala 121:29:@9092.4]
  wire  StickySelects_14_io_ins_0; // @[MemPrimitives.scala 121:29:@9092.4]
  wire  StickySelects_14_io_ins_1; // @[MemPrimitives.scala 121:29:@9092.4]
  wire  StickySelects_14_io_ins_2; // @[MemPrimitives.scala 121:29:@9092.4]
  wire  StickySelects_14_io_ins_3; // @[MemPrimitives.scala 121:29:@9092.4]
  wire  StickySelects_14_io_ins_4; // @[MemPrimitives.scala 121:29:@9092.4]
  wire  StickySelects_14_io_ins_5; // @[MemPrimitives.scala 121:29:@9092.4]
  wire  StickySelects_14_io_outs_0; // @[MemPrimitives.scala 121:29:@9092.4]
  wire  StickySelects_14_io_outs_1; // @[MemPrimitives.scala 121:29:@9092.4]
  wire  StickySelects_14_io_outs_2; // @[MemPrimitives.scala 121:29:@9092.4]
  wire  StickySelects_14_io_outs_3; // @[MemPrimitives.scala 121:29:@9092.4]
  wire  StickySelects_14_io_outs_4; // @[MemPrimitives.scala 121:29:@9092.4]
  wire  StickySelects_14_io_outs_5; // @[MemPrimitives.scala 121:29:@9092.4]
  wire  StickySelects_15_clock; // @[MemPrimitives.scala 121:29:@9148.4]
  wire  StickySelects_15_reset; // @[MemPrimitives.scala 121:29:@9148.4]
  wire  StickySelects_15_io_ins_0; // @[MemPrimitives.scala 121:29:@9148.4]
  wire  StickySelects_15_io_ins_1; // @[MemPrimitives.scala 121:29:@9148.4]
  wire  StickySelects_15_io_ins_2; // @[MemPrimitives.scala 121:29:@9148.4]
  wire  StickySelects_15_io_ins_3; // @[MemPrimitives.scala 121:29:@9148.4]
  wire  StickySelects_15_io_ins_4; // @[MemPrimitives.scala 121:29:@9148.4]
  wire  StickySelects_15_io_ins_5; // @[MemPrimitives.scala 121:29:@9148.4]
  wire  StickySelects_15_io_outs_0; // @[MemPrimitives.scala 121:29:@9148.4]
  wire  StickySelects_15_io_outs_1; // @[MemPrimitives.scala 121:29:@9148.4]
  wire  StickySelects_15_io_outs_2; // @[MemPrimitives.scala 121:29:@9148.4]
  wire  StickySelects_15_io_outs_3; // @[MemPrimitives.scala 121:29:@9148.4]
  wire  StickySelects_15_io_outs_4; // @[MemPrimitives.scala 121:29:@9148.4]
  wire  StickySelects_15_io_outs_5; // @[MemPrimitives.scala 121:29:@9148.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@9199.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@9199.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@9199.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@9199.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@9199.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@9207.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@9207.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@9207.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@9207.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@9207.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@9215.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@9215.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@9215.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@9215.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@9215.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@9223.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@9223.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@9223.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@9223.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@9223.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@9247.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@9247.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@9247.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@9247.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@9247.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@9255.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@9255.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@9255.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@9255.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@9255.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@9263.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@9263.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@9263.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@9263.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@9263.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@9271.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@9271.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@9271.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@9271.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@9271.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@9295.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@9295.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@9295.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@9295.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@9295.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@9303.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@9303.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@9303.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@9303.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@9303.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@9311.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@9311.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@9311.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@9311.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@9311.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@9319.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@9319.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@9319.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@9319.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@9319.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@9343.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@9343.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@9343.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@9343.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@9343.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@9351.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@9351.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@9351.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@9351.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@9351.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@9359.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@9359.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@9359.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@9359.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@9359.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@9367.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@9367.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@9367.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@9367.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@9367.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@9391.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@9391.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@9391.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@9391.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@9391.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@9399.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@9399.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@9399.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@9399.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@9399.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@9407.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@9407.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@9407.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@9407.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@9407.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@9415.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@9415.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@9415.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@9415.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@9415.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@9439.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@9439.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@9439.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@9439.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@9439.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@9447.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@9447.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@9447.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@9447.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@9447.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@9455.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@9455.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@9455.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@9455.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@9455.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@9463.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@9463.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@9463.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@9463.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@9463.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@9487.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@9487.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@9487.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@9487.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@9487.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@9495.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@9495.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@9495.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@9495.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@9495.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@9503.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@9503.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@9503.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@9503.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@9503.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@9511.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@9511.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@9511.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@9511.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@9511.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@9535.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@9535.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@9535.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@9535.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@9535.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@9543.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@9543.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@9543.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@9543.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@9543.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@9551.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@9551.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@9551.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@9551.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@9551.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@9559.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@9559.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@9559.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@9559.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@9559.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@9583.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@9583.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@9583.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@9583.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@9583.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@9591.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@9591.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@9591.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@9591.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@9591.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@9599.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@9599.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@9599.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@9599.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@9599.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@9607.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@9607.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@9607.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@9607.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@9607.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@9631.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@9631.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@9631.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@9631.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@9631.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@9639.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@9639.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@9639.4]
  wire  RetimeWrapper_37_io_in; // @[package.scala 93:22:@9639.4]
  wire  RetimeWrapper_37_io_out; // @[package.scala 93:22:@9639.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@9647.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@9647.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@9647.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@9647.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@9647.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@9655.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@9655.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@9655.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@9655.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@9655.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@9679.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@9679.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@9679.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@9679.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@9679.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@9687.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@9687.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@9687.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@9687.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@9687.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@9695.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@9695.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@9695.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@9695.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@9695.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@9703.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@9703.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@9703.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@9703.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@9703.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@9727.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@9727.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@9727.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@9727.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@9727.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@9735.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@9735.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@9735.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@9735.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@9735.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@9743.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@9743.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@9743.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@9743.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@9743.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@9751.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@9751.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@9751.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@9751.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@9751.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@9775.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@9775.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@9775.4]
  wire  RetimeWrapper_48_io_in; // @[package.scala 93:22:@9775.4]
  wire  RetimeWrapper_48_io_out; // @[package.scala 93:22:@9775.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@9783.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@9783.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@9783.4]
  wire  RetimeWrapper_49_io_in; // @[package.scala 93:22:@9783.4]
  wire  RetimeWrapper_49_io_out; // @[package.scala 93:22:@9783.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@9791.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@9791.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@9791.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@9791.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@9791.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@9799.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@9799.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@9799.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@9799.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@9799.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@9823.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@9823.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@9823.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@9823.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@9823.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@9831.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@9831.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@9831.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@9831.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@9831.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@9839.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@9839.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@9839.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@9839.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@9839.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@9847.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@9847.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@9847.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@9847.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@9847.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@9871.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@9871.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@9871.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@9871.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@9871.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@9879.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@9879.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@9879.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@9879.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@9879.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@9887.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@9887.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@9887.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@9887.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@9887.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@9895.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@9895.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@9895.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@9895.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@9895.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@9919.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@9919.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@9919.4]
  wire  RetimeWrapper_60_io_in; // @[package.scala 93:22:@9919.4]
  wire  RetimeWrapper_60_io_out; // @[package.scala 93:22:@9919.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@9927.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@9927.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@9927.4]
  wire  RetimeWrapper_61_io_in; // @[package.scala 93:22:@9927.4]
  wire  RetimeWrapper_61_io_out; // @[package.scala 93:22:@9927.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@9935.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@9935.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@9935.4]
  wire  RetimeWrapper_62_io_in; // @[package.scala 93:22:@9935.4]
  wire  RetimeWrapper_62_io_out; // @[package.scala 93:22:@9935.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@9943.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@9943.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@9943.4]
  wire  RetimeWrapper_63_io_in; // @[package.scala 93:22:@9943.4]
  wire  RetimeWrapper_63_io_out; // @[package.scala 93:22:@9943.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@9967.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@9967.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@9967.4]
  wire  RetimeWrapper_64_io_in; // @[package.scala 93:22:@9967.4]
  wire  RetimeWrapper_64_io_out; // @[package.scala 93:22:@9967.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@9975.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@9975.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@9975.4]
  wire  RetimeWrapper_65_io_in; // @[package.scala 93:22:@9975.4]
  wire  RetimeWrapper_65_io_out; // @[package.scala 93:22:@9975.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@9983.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@9983.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@9983.4]
  wire  RetimeWrapper_66_io_in; // @[package.scala 93:22:@9983.4]
  wire  RetimeWrapper_66_io_out; // @[package.scala 93:22:@9983.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@9991.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@9991.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@9991.4]
  wire  RetimeWrapper_67_io_in; // @[package.scala 93:22:@9991.4]
  wire  RetimeWrapper_67_io_out; // @[package.scala 93:22:@9991.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@10015.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@10015.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@10015.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@10015.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@10015.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@10023.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@10023.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@10023.4]
  wire  RetimeWrapper_69_io_in; // @[package.scala 93:22:@10023.4]
  wire  RetimeWrapper_69_io_out; // @[package.scala 93:22:@10023.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@10031.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@10031.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@10031.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@10031.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@10031.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@10039.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@10039.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@10039.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@10039.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@10039.4]
  wire  _T_700; // @[MemPrimitives.scala 82:210:@8306.4]
  wire  _T_703; // @[MemPrimitives.scala 83:102:@8308.4]
  wire [9:0] _T_705; // @[Cat.scala 30:58:@8310.4]
  wire  _T_710; // @[MemPrimitives.scala 82:210:@8317.4]
  wire  _T_713; // @[MemPrimitives.scala 83:102:@8319.4]
  wire [9:0] _T_715; // @[Cat.scala 30:58:@8321.4]
  wire  _T_720; // @[MemPrimitives.scala 82:210:@8328.4]
  wire  _T_723; // @[MemPrimitives.scala 83:102:@8330.4]
  wire [9:0] _T_725; // @[Cat.scala 30:58:@8332.4]
  wire  _T_730; // @[MemPrimitives.scala 82:210:@8339.4]
  wire  _T_733; // @[MemPrimitives.scala 83:102:@8341.4]
  wire [9:0] _T_735; // @[Cat.scala 30:58:@8343.4]
  wire  _T_740; // @[MemPrimitives.scala 82:210:@8350.4]
  wire  _T_743; // @[MemPrimitives.scala 83:102:@8352.4]
  wire [9:0] _T_745; // @[Cat.scala 30:58:@8354.4]
  wire  _T_750; // @[MemPrimitives.scala 82:210:@8361.4]
  wire  _T_753; // @[MemPrimitives.scala 83:102:@8363.4]
  wire [9:0] _T_755; // @[Cat.scala 30:58:@8365.4]
  wire  _T_760; // @[MemPrimitives.scala 82:210:@8372.4]
  wire  _T_763; // @[MemPrimitives.scala 83:102:@8374.4]
  wire [9:0] _T_765; // @[Cat.scala 30:58:@8376.4]
  wire  _T_770; // @[MemPrimitives.scala 82:210:@8383.4]
  wire  _T_773; // @[MemPrimitives.scala 83:102:@8385.4]
  wire [9:0] _T_775; // @[Cat.scala 30:58:@8387.4]
  wire  _T_780; // @[MemPrimitives.scala 82:210:@8394.4]
  wire  _T_783; // @[MemPrimitives.scala 83:102:@8396.4]
  wire [9:0] _T_785; // @[Cat.scala 30:58:@8398.4]
  wire  _T_790; // @[MemPrimitives.scala 82:210:@8405.4]
  wire  _T_793; // @[MemPrimitives.scala 83:102:@8407.4]
  wire [9:0] _T_795; // @[Cat.scala 30:58:@8409.4]
  wire  _T_800; // @[MemPrimitives.scala 82:210:@8416.4]
  wire  _T_803; // @[MemPrimitives.scala 83:102:@8418.4]
  wire [9:0] _T_805; // @[Cat.scala 30:58:@8420.4]
  wire  _T_810; // @[MemPrimitives.scala 82:210:@8427.4]
  wire  _T_813; // @[MemPrimitives.scala 83:102:@8429.4]
  wire [9:0] _T_815; // @[Cat.scala 30:58:@8431.4]
  wire  _T_820; // @[MemPrimitives.scala 82:210:@8438.4]
  wire  _T_823; // @[MemPrimitives.scala 83:102:@8440.4]
  wire [9:0] _T_825; // @[Cat.scala 30:58:@8442.4]
  wire  _T_830; // @[MemPrimitives.scala 82:210:@8449.4]
  wire  _T_833; // @[MemPrimitives.scala 83:102:@8451.4]
  wire [9:0] _T_835; // @[Cat.scala 30:58:@8453.4]
  wire  _T_840; // @[MemPrimitives.scala 82:210:@8460.4]
  wire  _T_843; // @[MemPrimitives.scala 83:102:@8462.4]
  wire [9:0] _T_845; // @[Cat.scala 30:58:@8464.4]
  wire  _T_850; // @[MemPrimitives.scala 82:210:@8471.4]
  wire  _T_853; // @[MemPrimitives.scala 83:102:@8473.4]
  wire [9:0] _T_855; // @[Cat.scala 30:58:@8475.4]
  wire  _T_860; // @[MemPrimitives.scala 110:210:@8482.4]
  wire  _T_865; // @[MemPrimitives.scala 110:210:@8485.4]
  wire  _T_870; // @[MemPrimitives.scala 110:210:@8488.4]
  wire  _T_874; // @[MemPrimitives.scala 123:41:@8497.4]
  wire  _T_875; // @[MemPrimitives.scala 123:41:@8498.4]
  wire  _T_876; // @[MemPrimitives.scala 123:41:@8499.4]
  wire [2:0] _T_878; // @[Cat.scala 30:58:@8501.4]
  wire [2:0] _T_880; // @[Cat.scala 30:58:@8503.4]
  wire [2:0] _T_882; // @[Cat.scala 30:58:@8505.4]
  wire [2:0] _T_883; // @[Mux.scala 31:69:@8506.4]
  wire [2:0] _T_884; // @[Mux.scala 31:69:@8507.4]
  wire  _T_889; // @[MemPrimitives.scala 110:210:@8514.4]
  wire  _T_894; // @[MemPrimitives.scala 110:210:@8517.4]
  wire  _T_899; // @[MemPrimitives.scala 110:210:@8520.4]
  wire  _T_903; // @[MemPrimitives.scala 123:41:@8529.4]
  wire  _T_904; // @[MemPrimitives.scala 123:41:@8530.4]
  wire  _T_905; // @[MemPrimitives.scala 123:41:@8531.4]
  wire [2:0] _T_907; // @[Cat.scala 30:58:@8533.4]
  wire [2:0] _T_909; // @[Cat.scala 30:58:@8535.4]
  wire [2:0] _T_911; // @[Cat.scala 30:58:@8537.4]
  wire [2:0] _T_912; // @[Mux.scala 31:69:@8538.4]
  wire [2:0] _T_913; // @[Mux.scala 31:69:@8539.4]
  wire  _T_918; // @[MemPrimitives.scala 110:210:@8546.4]
  wire  _T_923; // @[MemPrimitives.scala 110:210:@8549.4]
  wire  _T_928; // @[MemPrimitives.scala 110:210:@8552.4]
  wire  _T_933; // @[MemPrimitives.scala 110:210:@8555.4]
  wire  _T_938; // @[MemPrimitives.scala 110:210:@8558.4]
  wire  _T_943; // @[MemPrimitives.scala 110:210:@8561.4]
  wire  _T_947; // @[MemPrimitives.scala 123:41:@8573.4]
  wire  _T_948; // @[MemPrimitives.scala 123:41:@8574.4]
  wire  _T_949; // @[MemPrimitives.scala 123:41:@8575.4]
  wire  _T_950; // @[MemPrimitives.scala 123:41:@8576.4]
  wire  _T_951; // @[MemPrimitives.scala 123:41:@8577.4]
  wire  _T_952; // @[MemPrimitives.scala 123:41:@8578.4]
  wire [2:0] _T_954; // @[Cat.scala 30:58:@8580.4]
  wire [2:0] _T_956; // @[Cat.scala 30:58:@8582.4]
  wire [2:0] _T_958; // @[Cat.scala 30:58:@8584.4]
  wire [2:0] _T_960; // @[Cat.scala 30:58:@8586.4]
  wire [2:0] _T_962; // @[Cat.scala 30:58:@8588.4]
  wire [2:0] _T_964; // @[Cat.scala 30:58:@8590.4]
  wire [2:0] _T_965; // @[Mux.scala 31:69:@8591.4]
  wire [2:0] _T_966; // @[Mux.scala 31:69:@8592.4]
  wire [2:0] _T_967; // @[Mux.scala 31:69:@8593.4]
  wire [2:0] _T_968; // @[Mux.scala 31:69:@8594.4]
  wire [2:0] _T_969; // @[Mux.scala 31:69:@8595.4]
  wire  _T_974; // @[MemPrimitives.scala 110:210:@8602.4]
  wire  _T_979; // @[MemPrimitives.scala 110:210:@8605.4]
  wire  _T_984; // @[MemPrimitives.scala 110:210:@8608.4]
  wire  _T_989; // @[MemPrimitives.scala 110:210:@8611.4]
  wire  _T_994; // @[MemPrimitives.scala 110:210:@8614.4]
  wire  _T_999; // @[MemPrimitives.scala 110:210:@8617.4]
  wire  _T_1003; // @[MemPrimitives.scala 123:41:@8629.4]
  wire  _T_1004; // @[MemPrimitives.scala 123:41:@8630.4]
  wire  _T_1005; // @[MemPrimitives.scala 123:41:@8631.4]
  wire  _T_1006; // @[MemPrimitives.scala 123:41:@8632.4]
  wire  _T_1007; // @[MemPrimitives.scala 123:41:@8633.4]
  wire  _T_1008; // @[MemPrimitives.scala 123:41:@8634.4]
  wire [2:0] _T_1010; // @[Cat.scala 30:58:@8636.4]
  wire [2:0] _T_1012; // @[Cat.scala 30:58:@8638.4]
  wire [2:0] _T_1014; // @[Cat.scala 30:58:@8640.4]
  wire [2:0] _T_1016; // @[Cat.scala 30:58:@8642.4]
  wire [2:0] _T_1018; // @[Cat.scala 30:58:@8644.4]
  wire [2:0] _T_1020; // @[Cat.scala 30:58:@8646.4]
  wire [2:0] _T_1021; // @[Mux.scala 31:69:@8647.4]
  wire [2:0] _T_1022; // @[Mux.scala 31:69:@8648.4]
  wire [2:0] _T_1023; // @[Mux.scala 31:69:@8649.4]
  wire [2:0] _T_1024; // @[Mux.scala 31:69:@8650.4]
  wire [2:0] _T_1025; // @[Mux.scala 31:69:@8651.4]
  wire  _T_1030; // @[MemPrimitives.scala 110:210:@8658.4]
  wire  _T_1035; // @[MemPrimitives.scala 110:210:@8661.4]
  wire  _T_1040; // @[MemPrimitives.scala 110:210:@8664.4]
  wire  _T_1044; // @[MemPrimitives.scala 123:41:@8673.4]
  wire  _T_1045; // @[MemPrimitives.scala 123:41:@8674.4]
  wire  _T_1046; // @[MemPrimitives.scala 123:41:@8675.4]
  wire [2:0] _T_1048; // @[Cat.scala 30:58:@8677.4]
  wire [2:0] _T_1050; // @[Cat.scala 30:58:@8679.4]
  wire [2:0] _T_1052; // @[Cat.scala 30:58:@8681.4]
  wire [2:0] _T_1053; // @[Mux.scala 31:69:@8682.4]
  wire [2:0] _T_1054; // @[Mux.scala 31:69:@8683.4]
  wire  _T_1059; // @[MemPrimitives.scala 110:210:@8690.4]
  wire  _T_1064; // @[MemPrimitives.scala 110:210:@8693.4]
  wire  _T_1069; // @[MemPrimitives.scala 110:210:@8696.4]
  wire  _T_1073; // @[MemPrimitives.scala 123:41:@8705.4]
  wire  _T_1074; // @[MemPrimitives.scala 123:41:@8706.4]
  wire  _T_1075; // @[MemPrimitives.scala 123:41:@8707.4]
  wire [2:0] _T_1077; // @[Cat.scala 30:58:@8709.4]
  wire [2:0] _T_1079; // @[Cat.scala 30:58:@8711.4]
  wire [2:0] _T_1081; // @[Cat.scala 30:58:@8713.4]
  wire [2:0] _T_1082; // @[Mux.scala 31:69:@8714.4]
  wire [2:0] _T_1083; // @[Mux.scala 31:69:@8715.4]
  wire  _T_1088; // @[MemPrimitives.scala 110:210:@8722.4]
  wire  _T_1093; // @[MemPrimitives.scala 110:210:@8725.4]
  wire  _T_1098; // @[MemPrimitives.scala 110:210:@8728.4]
  wire  _T_1103; // @[MemPrimitives.scala 110:210:@8731.4]
  wire  _T_1108; // @[MemPrimitives.scala 110:210:@8734.4]
  wire  _T_1113; // @[MemPrimitives.scala 110:210:@8737.4]
  wire  _T_1117; // @[MemPrimitives.scala 123:41:@8749.4]
  wire  _T_1118; // @[MemPrimitives.scala 123:41:@8750.4]
  wire  _T_1119; // @[MemPrimitives.scala 123:41:@8751.4]
  wire  _T_1120; // @[MemPrimitives.scala 123:41:@8752.4]
  wire  _T_1121; // @[MemPrimitives.scala 123:41:@8753.4]
  wire  _T_1122; // @[MemPrimitives.scala 123:41:@8754.4]
  wire [2:0] _T_1124; // @[Cat.scala 30:58:@8756.4]
  wire [2:0] _T_1126; // @[Cat.scala 30:58:@8758.4]
  wire [2:0] _T_1128; // @[Cat.scala 30:58:@8760.4]
  wire [2:0] _T_1130; // @[Cat.scala 30:58:@8762.4]
  wire [2:0] _T_1132; // @[Cat.scala 30:58:@8764.4]
  wire [2:0] _T_1134; // @[Cat.scala 30:58:@8766.4]
  wire [2:0] _T_1135; // @[Mux.scala 31:69:@8767.4]
  wire [2:0] _T_1136; // @[Mux.scala 31:69:@8768.4]
  wire [2:0] _T_1137; // @[Mux.scala 31:69:@8769.4]
  wire [2:0] _T_1138; // @[Mux.scala 31:69:@8770.4]
  wire [2:0] _T_1139; // @[Mux.scala 31:69:@8771.4]
  wire  _T_1144; // @[MemPrimitives.scala 110:210:@8778.4]
  wire  _T_1149; // @[MemPrimitives.scala 110:210:@8781.4]
  wire  _T_1154; // @[MemPrimitives.scala 110:210:@8784.4]
  wire  _T_1159; // @[MemPrimitives.scala 110:210:@8787.4]
  wire  _T_1164; // @[MemPrimitives.scala 110:210:@8790.4]
  wire  _T_1169; // @[MemPrimitives.scala 110:210:@8793.4]
  wire  _T_1173; // @[MemPrimitives.scala 123:41:@8805.4]
  wire  _T_1174; // @[MemPrimitives.scala 123:41:@8806.4]
  wire  _T_1175; // @[MemPrimitives.scala 123:41:@8807.4]
  wire  _T_1176; // @[MemPrimitives.scala 123:41:@8808.4]
  wire  _T_1177; // @[MemPrimitives.scala 123:41:@8809.4]
  wire  _T_1178; // @[MemPrimitives.scala 123:41:@8810.4]
  wire [2:0] _T_1180; // @[Cat.scala 30:58:@8812.4]
  wire [2:0] _T_1182; // @[Cat.scala 30:58:@8814.4]
  wire [2:0] _T_1184; // @[Cat.scala 30:58:@8816.4]
  wire [2:0] _T_1186; // @[Cat.scala 30:58:@8818.4]
  wire [2:0] _T_1188; // @[Cat.scala 30:58:@8820.4]
  wire [2:0] _T_1190; // @[Cat.scala 30:58:@8822.4]
  wire [2:0] _T_1191; // @[Mux.scala 31:69:@8823.4]
  wire [2:0] _T_1192; // @[Mux.scala 31:69:@8824.4]
  wire [2:0] _T_1193; // @[Mux.scala 31:69:@8825.4]
  wire [2:0] _T_1194; // @[Mux.scala 31:69:@8826.4]
  wire [2:0] _T_1195; // @[Mux.scala 31:69:@8827.4]
  wire  _T_1200; // @[MemPrimitives.scala 110:210:@8834.4]
  wire  _T_1205; // @[MemPrimitives.scala 110:210:@8837.4]
  wire  _T_1210; // @[MemPrimitives.scala 110:210:@8840.4]
  wire  _T_1214; // @[MemPrimitives.scala 123:41:@8849.4]
  wire  _T_1215; // @[MemPrimitives.scala 123:41:@8850.4]
  wire  _T_1216; // @[MemPrimitives.scala 123:41:@8851.4]
  wire [2:0] _T_1218; // @[Cat.scala 30:58:@8853.4]
  wire [2:0] _T_1220; // @[Cat.scala 30:58:@8855.4]
  wire [2:0] _T_1222; // @[Cat.scala 30:58:@8857.4]
  wire [2:0] _T_1223; // @[Mux.scala 31:69:@8858.4]
  wire [2:0] _T_1224; // @[Mux.scala 31:69:@8859.4]
  wire  _T_1229; // @[MemPrimitives.scala 110:210:@8866.4]
  wire  _T_1234; // @[MemPrimitives.scala 110:210:@8869.4]
  wire  _T_1239; // @[MemPrimitives.scala 110:210:@8872.4]
  wire  _T_1243; // @[MemPrimitives.scala 123:41:@8881.4]
  wire  _T_1244; // @[MemPrimitives.scala 123:41:@8882.4]
  wire  _T_1245; // @[MemPrimitives.scala 123:41:@8883.4]
  wire [2:0] _T_1247; // @[Cat.scala 30:58:@8885.4]
  wire [2:0] _T_1249; // @[Cat.scala 30:58:@8887.4]
  wire [2:0] _T_1251; // @[Cat.scala 30:58:@8889.4]
  wire [2:0] _T_1252; // @[Mux.scala 31:69:@8890.4]
  wire [2:0] _T_1253; // @[Mux.scala 31:69:@8891.4]
  wire  _T_1258; // @[MemPrimitives.scala 110:210:@8898.4]
  wire  _T_1263; // @[MemPrimitives.scala 110:210:@8901.4]
  wire  _T_1268; // @[MemPrimitives.scala 110:210:@8904.4]
  wire  _T_1273; // @[MemPrimitives.scala 110:210:@8907.4]
  wire  _T_1278; // @[MemPrimitives.scala 110:210:@8910.4]
  wire  _T_1283; // @[MemPrimitives.scala 110:210:@8913.4]
  wire  _T_1287; // @[MemPrimitives.scala 123:41:@8925.4]
  wire  _T_1288; // @[MemPrimitives.scala 123:41:@8926.4]
  wire  _T_1289; // @[MemPrimitives.scala 123:41:@8927.4]
  wire  _T_1290; // @[MemPrimitives.scala 123:41:@8928.4]
  wire  _T_1291; // @[MemPrimitives.scala 123:41:@8929.4]
  wire  _T_1292; // @[MemPrimitives.scala 123:41:@8930.4]
  wire [2:0] _T_1294; // @[Cat.scala 30:58:@8932.4]
  wire [2:0] _T_1296; // @[Cat.scala 30:58:@8934.4]
  wire [2:0] _T_1298; // @[Cat.scala 30:58:@8936.4]
  wire [2:0] _T_1300; // @[Cat.scala 30:58:@8938.4]
  wire [2:0] _T_1302; // @[Cat.scala 30:58:@8940.4]
  wire [2:0] _T_1304; // @[Cat.scala 30:58:@8942.4]
  wire [2:0] _T_1305; // @[Mux.scala 31:69:@8943.4]
  wire [2:0] _T_1306; // @[Mux.scala 31:69:@8944.4]
  wire [2:0] _T_1307; // @[Mux.scala 31:69:@8945.4]
  wire [2:0] _T_1308; // @[Mux.scala 31:69:@8946.4]
  wire [2:0] _T_1309; // @[Mux.scala 31:69:@8947.4]
  wire  _T_1314; // @[MemPrimitives.scala 110:210:@8954.4]
  wire  _T_1319; // @[MemPrimitives.scala 110:210:@8957.4]
  wire  _T_1324; // @[MemPrimitives.scala 110:210:@8960.4]
  wire  _T_1329; // @[MemPrimitives.scala 110:210:@8963.4]
  wire  _T_1334; // @[MemPrimitives.scala 110:210:@8966.4]
  wire  _T_1339; // @[MemPrimitives.scala 110:210:@8969.4]
  wire  _T_1343; // @[MemPrimitives.scala 123:41:@8981.4]
  wire  _T_1344; // @[MemPrimitives.scala 123:41:@8982.4]
  wire  _T_1345; // @[MemPrimitives.scala 123:41:@8983.4]
  wire  _T_1346; // @[MemPrimitives.scala 123:41:@8984.4]
  wire  _T_1347; // @[MemPrimitives.scala 123:41:@8985.4]
  wire  _T_1348; // @[MemPrimitives.scala 123:41:@8986.4]
  wire [2:0] _T_1350; // @[Cat.scala 30:58:@8988.4]
  wire [2:0] _T_1352; // @[Cat.scala 30:58:@8990.4]
  wire [2:0] _T_1354; // @[Cat.scala 30:58:@8992.4]
  wire [2:0] _T_1356; // @[Cat.scala 30:58:@8994.4]
  wire [2:0] _T_1358; // @[Cat.scala 30:58:@8996.4]
  wire [2:0] _T_1360; // @[Cat.scala 30:58:@8998.4]
  wire [2:0] _T_1361; // @[Mux.scala 31:69:@8999.4]
  wire [2:0] _T_1362; // @[Mux.scala 31:69:@9000.4]
  wire [2:0] _T_1363; // @[Mux.scala 31:69:@9001.4]
  wire [2:0] _T_1364; // @[Mux.scala 31:69:@9002.4]
  wire [2:0] _T_1365; // @[Mux.scala 31:69:@9003.4]
  wire  _T_1370; // @[MemPrimitives.scala 110:210:@9010.4]
  wire  _T_1375; // @[MemPrimitives.scala 110:210:@9013.4]
  wire  _T_1380; // @[MemPrimitives.scala 110:210:@9016.4]
  wire  _T_1384; // @[MemPrimitives.scala 123:41:@9025.4]
  wire  _T_1385; // @[MemPrimitives.scala 123:41:@9026.4]
  wire  _T_1386; // @[MemPrimitives.scala 123:41:@9027.4]
  wire [2:0] _T_1388; // @[Cat.scala 30:58:@9029.4]
  wire [2:0] _T_1390; // @[Cat.scala 30:58:@9031.4]
  wire [2:0] _T_1392; // @[Cat.scala 30:58:@9033.4]
  wire [2:0] _T_1393; // @[Mux.scala 31:69:@9034.4]
  wire [2:0] _T_1394; // @[Mux.scala 31:69:@9035.4]
  wire  _T_1399; // @[MemPrimitives.scala 110:210:@9042.4]
  wire  _T_1404; // @[MemPrimitives.scala 110:210:@9045.4]
  wire  _T_1409; // @[MemPrimitives.scala 110:210:@9048.4]
  wire  _T_1413; // @[MemPrimitives.scala 123:41:@9057.4]
  wire  _T_1414; // @[MemPrimitives.scala 123:41:@9058.4]
  wire  _T_1415; // @[MemPrimitives.scala 123:41:@9059.4]
  wire [2:0] _T_1417; // @[Cat.scala 30:58:@9061.4]
  wire [2:0] _T_1419; // @[Cat.scala 30:58:@9063.4]
  wire [2:0] _T_1421; // @[Cat.scala 30:58:@9065.4]
  wire [2:0] _T_1422; // @[Mux.scala 31:69:@9066.4]
  wire [2:0] _T_1423; // @[Mux.scala 31:69:@9067.4]
  wire  _T_1428; // @[MemPrimitives.scala 110:210:@9074.4]
  wire  _T_1433; // @[MemPrimitives.scala 110:210:@9077.4]
  wire  _T_1438; // @[MemPrimitives.scala 110:210:@9080.4]
  wire  _T_1443; // @[MemPrimitives.scala 110:210:@9083.4]
  wire  _T_1448; // @[MemPrimitives.scala 110:210:@9086.4]
  wire  _T_1453; // @[MemPrimitives.scala 110:210:@9089.4]
  wire  _T_1457; // @[MemPrimitives.scala 123:41:@9101.4]
  wire  _T_1458; // @[MemPrimitives.scala 123:41:@9102.4]
  wire  _T_1459; // @[MemPrimitives.scala 123:41:@9103.4]
  wire  _T_1460; // @[MemPrimitives.scala 123:41:@9104.4]
  wire  _T_1461; // @[MemPrimitives.scala 123:41:@9105.4]
  wire  _T_1462; // @[MemPrimitives.scala 123:41:@9106.4]
  wire [2:0] _T_1464; // @[Cat.scala 30:58:@9108.4]
  wire [2:0] _T_1466; // @[Cat.scala 30:58:@9110.4]
  wire [2:0] _T_1468; // @[Cat.scala 30:58:@9112.4]
  wire [2:0] _T_1470; // @[Cat.scala 30:58:@9114.4]
  wire [2:0] _T_1472; // @[Cat.scala 30:58:@9116.4]
  wire [2:0] _T_1474; // @[Cat.scala 30:58:@9118.4]
  wire [2:0] _T_1475; // @[Mux.scala 31:69:@9119.4]
  wire [2:0] _T_1476; // @[Mux.scala 31:69:@9120.4]
  wire [2:0] _T_1477; // @[Mux.scala 31:69:@9121.4]
  wire [2:0] _T_1478; // @[Mux.scala 31:69:@9122.4]
  wire [2:0] _T_1479; // @[Mux.scala 31:69:@9123.4]
  wire  _T_1484; // @[MemPrimitives.scala 110:210:@9130.4]
  wire  _T_1489; // @[MemPrimitives.scala 110:210:@9133.4]
  wire  _T_1494; // @[MemPrimitives.scala 110:210:@9136.4]
  wire  _T_1499; // @[MemPrimitives.scala 110:210:@9139.4]
  wire  _T_1504; // @[MemPrimitives.scala 110:210:@9142.4]
  wire  _T_1509; // @[MemPrimitives.scala 110:210:@9145.4]
  wire  _T_1513; // @[MemPrimitives.scala 123:41:@9157.4]
  wire  _T_1514; // @[MemPrimitives.scala 123:41:@9158.4]
  wire  _T_1515; // @[MemPrimitives.scala 123:41:@9159.4]
  wire  _T_1516; // @[MemPrimitives.scala 123:41:@9160.4]
  wire  _T_1517; // @[MemPrimitives.scala 123:41:@9161.4]
  wire  _T_1518; // @[MemPrimitives.scala 123:41:@9162.4]
  wire [2:0] _T_1520; // @[Cat.scala 30:58:@9164.4]
  wire [2:0] _T_1522; // @[Cat.scala 30:58:@9166.4]
  wire [2:0] _T_1524; // @[Cat.scala 30:58:@9168.4]
  wire [2:0] _T_1526; // @[Cat.scala 30:58:@9170.4]
  wire [2:0] _T_1528; // @[Cat.scala 30:58:@9172.4]
  wire [2:0] _T_1530; // @[Cat.scala 30:58:@9174.4]
  wire [2:0] _T_1531; // @[Mux.scala 31:69:@9175.4]
  wire [2:0] _T_1532; // @[Mux.scala 31:69:@9176.4]
  wire [2:0] _T_1533; // @[Mux.scala 31:69:@9177.4]
  wire [2:0] _T_1534; // @[Mux.scala 31:69:@9178.4]
  wire [2:0] _T_1535; // @[Mux.scala 31:69:@9179.4]
  wire  _T_1567; // @[package.scala 96:25:@9220.4 package.scala 96:25:@9221.4]
  wire [7:0] _T_1571; // @[Mux.scala 31:69:@9230.4]
  wire  _T_1564; // @[package.scala 96:25:@9212.4 package.scala 96:25:@9213.4]
  wire [7:0] _T_1572; // @[Mux.scala 31:69:@9231.4]
  wire  _T_1561; // @[package.scala 96:25:@9204.4 package.scala 96:25:@9205.4]
  wire  _T_1602; // @[package.scala 96:25:@9268.4 package.scala 96:25:@9269.4]
  wire [7:0] _T_1606; // @[Mux.scala 31:69:@9278.4]
  wire  _T_1599; // @[package.scala 96:25:@9260.4 package.scala 96:25:@9261.4]
  wire [7:0] _T_1607; // @[Mux.scala 31:69:@9279.4]
  wire  _T_1596; // @[package.scala 96:25:@9252.4 package.scala 96:25:@9253.4]
  wire  _T_1637; // @[package.scala 96:25:@9316.4 package.scala 96:25:@9317.4]
  wire [7:0] _T_1641; // @[Mux.scala 31:69:@9326.4]
  wire  _T_1634; // @[package.scala 96:25:@9308.4 package.scala 96:25:@9309.4]
  wire [7:0] _T_1642; // @[Mux.scala 31:69:@9327.4]
  wire  _T_1631; // @[package.scala 96:25:@9300.4 package.scala 96:25:@9301.4]
  wire  _T_1672; // @[package.scala 96:25:@9364.4 package.scala 96:25:@9365.4]
  wire [7:0] _T_1676; // @[Mux.scala 31:69:@9374.4]
  wire  _T_1669; // @[package.scala 96:25:@9356.4 package.scala 96:25:@9357.4]
  wire [7:0] _T_1677; // @[Mux.scala 31:69:@9375.4]
  wire  _T_1666; // @[package.scala 96:25:@9348.4 package.scala 96:25:@9349.4]
  wire  _T_1707; // @[package.scala 96:25:@9412.4 package.scala 96:25:@9413.4]
  wire [7:0] _T_1711; // @[Mux.scala 31:69:@9422.4]
  wire  _T_1704; // @[package.scala 96:25:@9404.4 package.scala 96:25:@9405.4]
  wire [7:0] _T_1712; // @[Mux.scala 31:69:@9423.4]
  wire  _T_1701; // @[package.scala 96:25:@9396.4 package.scala 96:25:@9397.4]
  wire  _T_1742; // @[package.scala 96:25:@9460.4 package.scala 96:25:@9461.4]
  wire [7:0] _T_1746; // @[Mux.scala 31:69:@9470.4]
  wire  _T_1739; // @[package.scala 96:25:@9452.4 package.scala 96:25:@9453.4]
  wire [7:0] _T_1747; // @[Mux.scala 31:69:@9471.4]
  wire  _T_1736; // @[package.scala 96:25:@9444.4 package.scala 96:25:@9445.4]
  wire  _T_1777; // @[package.scala 96:25:@9508.4 package.scala 96:25:@9509.4]
  wire [7:0] _T_1781; // @[Mux.scala 31:69:@9518.4]
  wire  _T_1774; // @[package.scala 96:25:@9500.4 package.scala 96:25:@9501.4]
  wire [7:0] _T_1782; // @[Mux.scala 31:69:@9519.4]
  wire  _T_1771; // @[package.scala 96:25:@9492.4 package.scala 96:25:@9493.4]
  wire  _T_1812; // @[package.scala 96:25:@9556.4 package.scala 96:25:@9557.4]
  wire [7:0] _T_1816; // @[Mux.scala 31:69:@9566.4]
  wire  _T_1809; // @[package.scala 96:25:@9548.4 package.scala 96:25:@9549.4]
  wire [7:0] _T_1817; // @[Mux.scala 31:69:@9567.4]
  wire  _T_1806; // @[package.scala 96:25:@9540.4 package.scala 96:25:@9541.4]
  wire  _T_1847; // @[package.scala 96:25:@9604.4 package.scala 96:25:@9605.4]
  wire [7:0] _T_1851; // @[Mux.scala 31:69:@9614.4]
  wire  _T_1844; // @[package.scala 96:25:@9596.4 package.scala 96:25:@9597.4]
  wire [7:0] _T_1852; // @[Mux.scala 31:69:@9615.4]
  wire  _T_1841; // @[package.scala 96:25:@9588.4 package.scala 96:25:@9589.4]
  wire  _T_1882; // @[package.scala 96:25:@9652.4 package.scala 96:25:@9653.4]
  wire [7:0] _T_1886; // @[Mux.scala 31:69:@9662.4]
  wire  _T_1879; // @[package.scala 96:25:@9644.4 package.scala 96:25:@9645.4]
  wire [7:0] _T_1887; // @[Mux.scala 31:69:@9663.4]
  wire  _T_1876; // @[package.scala 96:25:@9636.4 package.scala 96:25:@9637.4]
  wire  _T_1917; // @[package.scala 96:25:@9700.4 package.scala 96:25:@9701.4]
  wire [7:0] _T_1921; // @[Mux.scala 31:69:@9710.4]
  wire  _T_1914; // @[package.scala 96:25:@9692.4 package.scala 96:25:@9693.4]
  wire [7:0] _T_1922; // @[Mux.scala 31:69:@9711.4]
  wire  _T_1911; // @[package.scala 96:25:@9684.4 package.scala 96:25:@9685.4]
  wire  _T_1952; // @[package.scala 96:25:@9748.4 package.scala 96:25:@9749.4]
  wire [7:0] _T_1956; // @[Mux.scala 31:69:@9758.4]
  wire  _T_1949; // @[package.scala 96:25:@9740.4 package.scala 96:25:@9741.4]
  wire [7:0] _T_1957; // @[Mux.scala 31:69:@9759.4]
  wire  _T_1946; // @[package.scala 96:25:@9732.4 package.scala 96:25:@9733.4]
  wire  _T_1987; // @[package.scala 96:25:@9796.4 package.scala 96:25:@9797.4]
  wire [7:0] _T_1991; // @[Mux.scala 31:69:@9806.4]
  wire  _T_1984; // @[package.scala 96:25:@9788.4 package.scala 96:25:@9789.4]
  wire [7:0] _T_1992; // @[Mux.scala 31:69:@9807.4]
  wire  _T_1981; // @[package.scala 96:25:@9780.4 package.scala 96:25:@9781.4]
  wire  _T_2022; // @[package.scala 96:25:@9844.4 package.scala 96:25:@9845.4]
  wire [7:0] _T_2026; // @[Mux.scala 31:69:@9854.4]
  wire  _T_2019; // @[package.scala 96:25:@9836.4 package.scala 96:25:@9837.4]
  wire [7:0] _T_2027; // @[Mux.scala 31:69:@9855.4]
  wire  _T_2016; // @[package.scala 96:25:@9828.4 package.scala 96:25:@9829.4]
  wire  _T_2057; // @[package.scala 96:25:@9892.4 package.scala 96:25:@9893.4]
  wire [7:0] _T_2061; // @[Mux.scala 31:69:@9902.4]
  wire  _T_2054; // @[package.scala 96:25:@9884.4 package.scala 96:25:@9885.4]
  wire [7:0] _T_2062; // @[Mux.scala 31:69:@9903.4]
  wire  _T_2051; // @[package.scala 96:25:@9876.4 package.scala 96:25:@9877.4]
  wire  _T_2092; // @[package.scala 96:25:@9940.4 package.scala 96:25:@9941.4]
  wire [7:0] _T_2096; // @[Mux.scala 31:69:@9950.4]
  wire  _T_2089; // @[package.scala 96:25:@9932.4 package.scala 96:25:@9933.4]
  wire [7:0] _T_2097; // @[Mux.scala 31:69:@9951.4]
  wire  _T_2086; // @[package.scala 96:25:@9924.4 package.scala 96:25:@9925.4]
  wire  _T_2127; // @[package.scala 96:25:@9988.4 package.scala 96:25:@9989.4]
  wire [7:0] _T_2131; // @[Mux.scala 31:69:@9998.4]
  wire  _T_2124; // @[package.scala 96:25:@9980.4 package.scala 96:25:@9981.4]
  wire [7:0] _T_2132; // @[Mux.scala 31:69:@9999.4]
  wire  _T_2121; // @[package.scala 96:25:@9972.4 package.scala 96:25:@9973.4]
  wire  _T_2162; // @[package.scala 96:25:@10036.4 package.scala 96:25:@10037.4]
  wire [7:0] _T_2166; // @[Mux.scala 31:69:@10046.4]
  wire  _T_2159; // @[package.scala 96:25:@10028.4 package.scala 96:25:@10029.4]
  wire [7:0] _T_2167; // @[Mux.scala 31:69:@10047.4]
  wire  _T_2156; // @[package.scala 96:25:@10020.4 package.scala 96:25:@10021.4]
  Mem1D_4 Mem1D ( // @[MemPrimitives.scala 64:21:@8050.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  Mem1D_4 Mem1D_1 ( // @[MemPrimitives.scala 64:21:@8066.4]
    .clock(Mem1D_1_clock),
    .reset(Mem1D_1_reset),
    .io_r_ofs_0(Mem1D_1_io_r_ofs_0),
    .io_r_backpressure(Mem1D_1_io_r_backpressure),
    .io_w_ofs_0(Mem1D_1_io_w_ofs_0),
    .io_w_data_0(Mem1D_1_io_w_data_0),
    .io_w_en_0(Mem1D_1_io_w_en_0),
    .io_output(Mem1D_1_io_output)
  );
  Mem1D_4 Mem1D_2 ( // @[MemPrimitives.scala 64:21:@8082.4]
    .clock(Mem1D_2_clock),
    .reset(Mem1D_2_reset),
    .io_r_ofs_0(Mem1D_2_io_r_ofs_0),
    .io_r_backpressure(Mem1D_2_io_r_backpressure),
    .io_w_ofs_0(Mem1D_2_io_w_ofs_0),
    .io_w_data_0(Mem1D_2_io_w_data_0),
    .io_w_en_0(Mem1D_2_io_w_en_0),
    .io_output(Mem1D_2_io_output)
  );
  Mem1D_4 Mem1D_3 ( // @[MemPrimitives.scala 64:21:@8098.4]
    .clock(Mem1D_3_clock),
    .reset(Mem1D_3_reset),
    .io_r_ofs_0(Mem1D_3_io_r_ofs_0),
    .io_r_backpressure(Mem1D_3_io_r_backpressure),
    .io_w_ofs_0(Mem1D_3_io_w_ofs_0),
    .io_w_data_0(Mem1D_3_io_w_data_0),
    .io_w_en_0(Mem1D_3_io_w_en_0),
    .io_output(Mem1D_3_io_output)
  );
  Mem1D_4 Mem1D_4 ( // @[MemPrimitives.scala 64:21:@8114.4]
    .clock(Mem1D_4_clock),
    .reset(Mem1D_4_reset),
    .io_r_ofs_0(Mem1D_4_io_r_ofs_0),
    .io_r_backpressure(Mem1D_4_io_r_backpressure),
    .io_w_ofs_0(Mem1D_4_io_w_ofs_0),
    .io_w_data_0(Mem1D_4_io_w_data_0),
    .io_w_en_0(Mem1D_4_io_w_en_0),
    .io_output(Mem1D_4_io_output)
  );
  Mem1D_4 Mem1D_5 ( // @[MemPrimitives.scala 64:21:@8130.4]
    .clock(Mem1D_5_clock),
    .reset(Mem1D_5_reset),
    .io_r_ofs_0(Mem1D_5_io_r_ofs_0),
    .io_r_backpressure(Mem1D_5_io_r_backpressure),
    .io_w_ofs_0(Mem1D_5_io_w_ofs_0),
    .io_w_data_0(Mem1D_5_io_w_data_0),
    .io_w_en_0(Mem1D_5_io_w_en_0),
    .io_output(Mem1D_5_io_output)
  );
  Mem1D_4 Mem1D_6 ( // @[MemPrimitives.scala 64:21:@8146.4]
    .clock(Mem1D_6_clock),
    .reset(Mem1D_6_reset),
    .io_r_ofs_0(Mem1D_6_io_r_ofs_0),
    .io_r_backpressure(Mem1D_6_io_r_backpressure),
    .io_w_ofs_0(Mem1D_6_io_w_ofs_0),
    .io_w_data_0(Mem1D_6_io_w_data_0),
    .io_w_en_0(Mem1D_6_io_w_en_0),
    .io_output(Mem1D_6_io_output)
  );
  Mem1D_4 Mem1D_7 ( // @[MemPrimitives.scala 64:21:@8162.4]
    .clock(Mem1D_7_clock),
    .reset(Mem1D_7_reset),
    .io_r_ofs_0(Mem1D_7_io_r_ofs_0),
    .io_r_backpressure(Mem1D_7_io_r_backpressure),
    .io_w_ofs_0(Mem1D_7_io_w_ofs_0),
    .io_w_data_0(Mem1D_7_io_w_data_0),
    .io_w_en_0(Mem1D_7_io_w_en_0),
    .io_output(Mem1D_7_io_output)
  );
  Mem1D_4 Mem1D_8 ( // @[MemPrimitives.scala 64:21:@8178.4]
    .clock(Mem1D_8_clock),
    .reset(Mem1D_8_reset),
    .io_r_ofs_0(Mem1D_8_io_r_ofs_0),
    .io_r_backpressure(Mem1D_8_io_r_backpressure),
    .io_w_ofs_0(Mem1D_8_io_w_ofs_0),
    .io_w_data_0(Mem1D_8_io_w_data_0),
    .io_w_en_0(Mem1D_8_io_w_en_0),
    .io_output(Mem1D_8_io_output)
  );
  Mem1D_4 Mem1D_9 ( // @[MemPrimitives.scala 64:21:@8194.4]
    .clock(Mem1D_9_clock),
    .reset(Mem1D_9_reset),
    .io_r_ofs_0(Mem1D_9_io_r_ofs_0),
    .io_r_backpressure(Mem1D_9_io_r_backpressure),
    .io_w_ofs_0(Mem1D_9_io_w_ofs_0),
    .io_w_data_0(Mem1D_9_io_w_data_0),
    .io_w_en_0(Mem1D_9_io_w_en_0),
    .io_output(Mem1D_9_io_output)
  );
  Mem1D_4 Mem1D_10 ( // @[MemPrimitives.scala 64:21:@8210.4]
    .clock(Mem1D_10_clock),
    .reset(Mem1D_10_reset),
    .io_r_ofs_0(Mem1D_10_io_r_ofs_0),
    .io_r_backpressure(Mem1D_10_io_r_backpressure),
    .io_w_ofs_0(Mem1D_10_io_w_ofs_0),
    .io_w_data_0(Mem1D_10_io_w_data_0),
    .io_w_en_0(Mem1D_10_io_w_en_0),
    .io_output(Mem1D_10_io_output)
  );
  Mem1D_4 Mem1D_11 ( // @[MemPrimitives.scala 64:21:@8226.4]
    .clock(Mem1D_11_clock),
    .reset(Mem1D_11_reset),
    .io_r_ofs_0(Mem1D_11_io_r_ofs_0),
    .io_r_backpressure(Mem1D_11_io_r_backpressure),
    .io_w_ofs_0(Mem1D_11_io_w_ofs_0),
    .io_w_data_0(Mem1D_11_io_w_data_0),
    .io_w_en_0(Mem1D_11_io_w_en_0),
    .io_output(Mem1D_11_io_output)
  );
  Mem1D_4 Mem1D_12 ( // @[MemPrimitives.scala 64:21:@8242.4]
    .clock(Mem1D_12_clock),
    .reset(Mem1D_12_reset),
    .io_r_ofs_0(Mem1D_12_io_r_ofs_0),
    .io_r_backpressure(Mem1D_12_io_r_backpressure),
    .io_w_ofs_0(Mem1D_12_io_w_ofs_0),
    .io_w_data_0(Mem1D_12_io_w_data_0),
    .io_w_en_0(Mem1D_12_io_w_en_0),
    .io_output(Mem1D_12_io_output)
  );
  Mem1D_4 Mem1D_13 ( // @[MemPrimitives.scala 64:21:@8258.4]
    .clock(Mem1D_13_clock),
    .reset(Mem1D_13_reset),
    .io_r_ofs_0(Mem1D_13_io_r_ofs_0),
    .io_r_backpressure(Mem1D_13_io_r_backpressure),
    .io_w_ofs_0(Mem1D_13_io_w_ofs_0),
    .io_w_data_0(Mem1D_13_io_w_data_0),
    .io_w_en_0(Mem1D_13_io_w_en_0),
    .io_output(Mem1D_13_io_output)
  );
  Mem1D_4 Mem1D_14 ( // @[MemPrimitives.scala 64:21:@8274.4]
    .clock(Mem1D_14_clock),
    .reset(Mem1D_14_reset),
    .io_r_ofs_0(Mem1D_14_io_r_ofs_0),
    .io_r_backpressure(Mem1D_14_io_r_backpressure),
    .io_w_ofs_0(Mem1D_14_io_w_ofs_0),
    .io_w_data_0(Mem1D_14_io_w_data_0),
    .io_w_en_0(Mem1D_14_io_w_en_0),
    .io_output(Mem1D_14_io_output)
  );
  Mem1D_4 Mem1D_15 ( // @[MemPrimitives.scala 64:21:@8290.4]
    .clock(Mem1D_15_clock),
    .reset(Mem1D_15_reset),
    .io_r_ofs_0(Mem1D_15_io_r_ofs_0),
    .io_r_backpressure(Mem1D_15_io_r_backpressure),
    .io_w_ofs_0(Mem1D_15_io_w_ofs_0),
    .io_w_data_0(Mem1D_15_io_w_data_0),
    .io_w_en_0(Mem1D_15_io_w_en_0),
    .io_output(Mem1D_15_io_output)
  );
  StickySelects StickySelects ( // @[MemPrimitives.scala 121:29:@8491.4]
    .clock(StickySelects_clock),
    .reset(StickySelects_reset),
    .io_ins_0(StickySelects_io_ins_0),
    .io_ins_1(StickySelects_io_ins_1),
    .io_ins_2(StickySelects_io_ins_2),
    .io_outs_0(StickySelects_io_outs_0),
    .io_outs_1(StickySelects_io_outs_1),
    .io_outs_2(StickySelects_io_outs_2)
  );
  StickySelects StickySelects_1 ( // @[MemPrimitives.scala 121:29:@8523.4]
    .clock(StickySelects_1_clock),
    .reset(StickySelects_1_reset),
    .io_ins_0(StickySelects_1_io_ins_0),
    .io_ins_1(StickySelects_1_io_ins_1),
    .io_ins_2(StickySelects_1_io_ins_2),
    .io_outs_0(StickySelects_1_io_outs_0),
    .io_outs_1(StickySelects_1_io_outs_1),
    .io_outs_2(StickySelects_1_io_outs_2)
  );
  StickySelects_2 StickySelects_2 ( // @[MemPrimitives.scala 121:29:@8564.4]
    .clock(StickySelects_2_clock),
    .reset(StickySelects_2_reset),
    .io_ins_0(StickySelects_2_io_ins_0),
    .io_ins_1(StickySelects_2_io_ins_1),
    .io_ins_2(StickySelects_2_io_ins_2),
    .io_ins_3(StickySelects_2_io_ins_3),
    .io_ins_4(StickySelects_2_io_ins_4),
    .io_ins_5(StickySelects_2_io_ins_5),
    .io_outs_0(StickySelects_2_io_outs_0),
    .io_outs_1(StickySelects_2_io_outs_1),
    .io_outs_2(StickySelects_2_io_outs_2),
    .io_outs_3(StickySelects_2_io_outs_3),
    .io_outs_4(StickySelects_2_io_outs_4),
    .io_outs_5(StickySelects_2_io_outs_5)
  );
  StickySelects_2 StickySelects_3 ( // @[MemPrimitives.scala 121:29:@8620.4]
    .clock(StickySelects_3_clock),
    .reset(StickySelects_3_reset),
    .io_ins_0(StickySelects_3_io_ins_0),
    .io_ins_1(StickySelects_3_io_ins_1),
    .io_ins_2(StickySelects_3_io_ins_2),
    .io_ins_3(StickySelects_3_io_ins_3),
    .io_ins_4(StickySelects_3_io_ins_4),
    .io_ins_5(StickySelects_3_io_ins_5),
    .io_outs_0(StickySelects_3_io_outs_0),
    .io_outs_1(StickySelects_3_io_outs_1),
    .io_outs_2(StickySelects_3_io_outs_2),
    .io_outs_3(StickySelects_3_io_outs_3),
    .io_outs_4(StickySelects_3_io_outs_4),
    .io_outs_5(StickySelects_3_io_outs_5)
  );
  StickySelects StickySelects_4 ( // @[MemPrimitives.scala 121:29:@8667.4]
    .clock(StickySelects_4_clock),
    .reset(StickySelects_4_reset),
    .io_ins_0(StickySelects_4_io_ins_0),
    .io_ins_1(StickySelects_4_io_ins_1),
    .io_ins_2(StickySelects_4_io_ins_2),
    .io_outs_0(StickySelects_4_io_outs_0),
    .io_outs_1(StickySelects_4_io_outs_1),
    .io_outs_2(StickySelects_4_io_outs_2)
  );
  StickySelects StickySelects_5 ( // @[MemPrimitives.scala 121:29:@8699.4]
    .clock(StickySelects_5_clock),
    .reset(StickySelects_5_reset),
    .io_ins_0(StickySelects_5_io_ins_0),
    .io_ins_1(StickySelects_5_io_ins_1),
    .io_ins_2(StickySelects_5_io_ins_2),
    .io_outs_0(StickySelects_5_io_outs_0),
    .io_outs_1(StickySelects_5_io_outs_1),
    .io_outs_2(StickySelects_5_io_outs_2)
  );
  StickySelects_2 StickySelects_6 ( // @[MemPrimitives.scala 121:29:@8740.4]
    .clock(StickySelects_6_clock),
    .reset(StickySelects_6_reset),
    .io_ins_0(StickySelects_6_io_ins_0),
    .io_ins_1(StickySelects_6_io_ins_1),
    .io_ins_2(StickySelects_6_io_ins_2),
    .io_ins_3(StickySelects_6_io_ins_3),
    .io_ins_4(StickySelects_6_io_ins_4),
    .io_ins_5(StickySelects_6_io_ins_5),
    .io_outs_0(StickySelects_6_io_outs_0),
    .io_outs_1(StickySelects_6_io_outs_1),
    .io_outs_2(StickySelects_6_io_outs_2),
    .io_outs_3(StickySelects_6_io_outs_3),
    .io_outs_4(StickySelects_6_io_outs_4),
    .io_outs_5(StickySelects_6_io_outs_5)
  );
  StickySelects_2 StickySelects_7 ( // @[MemPrimitives.scala 121:29:@8796.4]
    .clock(StickySelects_7_clock),
    .reset(StickySelects_7_reset),
    .io_ins_0(StickySelects_7_io_ins_0),
    .io_ins_1(StickySelects_7_io_ins_1),
    .io_ins_2(StickySelects_7_io_ins_2),
    .io_ins_3(StickySelects_7_io_ins_3),
    .io_ins_4(StickySelects_7_io_ins_4),
    .io_ins_5(StickySelects_7_io_ins_5),
    .io_outs_0(StickySelects_7_io_outs_0),
    .io_outs_1(StickySelects_7_io_outs_1),
    .io_outs_2(StickySelects_7_io_outs_2),
    .io_outs_3(StickySelects_7_io_outs_3),
    .io_outs_4(StickySelects_7_io_outs_4),
    .io_outs_5(StickySelects_7_io_outs_5)
  );
  StickySelects StickySelects_8 ( // @[MemPrimitives.scala 121:29:@8843.4]
    .clock(StickySelects_8_clock),
    .reset(StickySelects_8_reset),
    .io_ins_0(StickySelects_8_io_ins_0),
    .io_ins_1(StickySelects_8_io_ins_1),
    .io_ins_2(StickySelects_8_io_ins_2),
    .io_outs_0(StickySelects_8_io_outs_0),
    .io_outs_1(StickySelects_8_io_outs_1),
    .io_outs_2(StickySelects_8_io_outs_2)
  );
  StickySelects StickySelects_9 ( // @[MemPrimitives.scala 121:29:@8875.4]
    .clock(StickySelects_9_clock),
    .reset(StickySelects_9_reset),
    .io_ins_0(StickySelects_9_io_ins_0),
    .io_ins_1(StickySelects_9_io_ins_1),
    .io_ins_2(StickySelects_9_io_ins_2),
    .io_outs_0(StickySelects_9_io_outs_0),
    .io_outs_1(StickySelects_9_io_outs_1),
    .io_outs_2(StickySelects_9_io_outs_2)
  );
  StickySelects_2 StickySelects_10 ( // @[MemPrimitives.scala 121:29:@8916.4]
    .clock(StickySelects_10_clock),
    .reset(StickySelects_10_reset),
    .io_ins_0(StickySelects_10_io_ins_0),
    .io_ins_1(StickySelects_10_io_ins_1),
    .io_ins_2(StickySelects_10_io_ins_2),
    .io_ins_3(StickySelects_10_io_ins_3),
    .io_ins_4(StickySelects_10_io_ins_4),
    .io_ins_5(StickySelects_10_io_ins_5),
    .io_outs_0(StickySelects_10_io_outs_0),
    .io_outs_1(StickySelects_10_io_outs_1),
    .io_outs_2(StickySelects_10_io_outs_2),
    .io_outs_3(StickySelects_10_io_outs_3),
    .io_outs_4(StickySelects_10_io_outs_4),
    .io_outs_5(StickySelects_10_io_outs_5)
  );
  StickySelects_2 StickySelects_11 ( // @[MemPrimitives.scala 121:29:@8972.4]
    .clock(StickySelects_11_clock),
    .reset(StickySelects_11_reset),
    .io_ins_0(StickySelects_11_io_ins_0),
    .io_ins_1(StickySelects_11_io_ins_1),
    .io_ins_2(StickySelects_11_io_ins_2),
    .io_ins_3(StickySelects_11_io_ins_3),
    .io_ins_4(StickySelects_11_io_ins_4),
    .io_ins_5(StickySelects_11_io_ins_5),
    .io_outs_0(StickySelects_11_io_outs_0),
    .io_outs_1(StickySelects_11_io_outs_1),
    .io_outs_2(StickySelects_11_io_outs_2),
    .io_outs_3(StickySelects_11_io_outs_3),
    .io_outs_4(StickySelects_11_io_outs_4),
    .io_outs_5(StickySelects_11_io_outs_5)
  );
  StickySelects StickySelects_12 ( // @[MemPrimitives.scala 121:29:@9019.4]
    .clock(StickySelects_12_clock),
    .reset(StickySelects_12_reset),
    .io_ins_0(StickySelects_12_io_ins_0),
    .io_ins_1(StickySelects_12_io_ins_1),
    .io_ins_2(StickySelects_12_io_ins_2),
    .io_outs_0(StickySelects_12_io_outs_0),
    .io_outs_1(StickySelects_12_io_outs_1),
    .io_outs_2(StickySelects_12_io_outs_2)
  );
  StickySelects StickySelects_13 ( // @[MemPrimitives.scala 121:29:@9051.4]
    .clock(StickySelects_13_clock),
    .reset(StickySelects_13_reset),
    .io_ins_0(StickySelects_13_io_ins_0),
    .io_ins_1(StickySelects_13_io_ins_1),
    .io_ins_2(StickySelects_13_io_ins_2),
    .io_outs_0(StickySelects_13_io_outs_0),
    .io_outs_1(StickySelects_13_io_outs_1),
    .io_outs_2(StickySelects_13_io_outs_2)
  );
  StickySelects_2 StickySelects_14 ( // @[MemPrimitives.scala 121:29:@9092.4]
    .clock(StickySelects_14_clock),
    .reset(StickySelects_14_reset),
    .io_ins_0(StickySelects_14_io_ins_0),
    .io_ins_1(StickySelects_14_io_ins_1),
    .io_ins_2(StickySelects_14_io_ins_2),
    .io_ins_3(StickySelects_14_io_ins_3),
    .io_ins_4(StickySelects_14_io_ins_4),
    .io_ins_5(StickySelects_14_io_ins_5),
    .io_outs_0(StickySelects_14_io_outs_0),
    .io_outs_1(StickySelects_14_io_outs_1),
    .io_outs_2(StickySelects_14_io_outs_2),
    .io_outs_3(StickySelects_14_io_outs_3),
    .io_outs_4(StickySelects_14_io_outs_4),
    .io_outs_5(StickySelects_14_io_outs_5)
  );
  StickySelects_2 StickySelects_15 ( // @[MemPrimitives.scala 121:29:@9148.4]
    .clock(StickySelects_15_clock),
    .reset(StickySelects_15_reset),
    .io_ins_0(StickySelects_15_io_ins_0),
    .io_ins_1(StickySelects_15_io_ins_1),
    .io_ins_2(StickySelects_15_io_ins_2),
    .io_ins_3(StickySelects_15_io_ins_3),
    .io_ins_4(StickySelects_15_io_ins_4),
    .io_ins_5(StickySelects_15_io_ins_5),
    .io_outs_0(StickySelects_15_io_outs_0),
    .io_outs_1(StickySelects_15_io_outs_1),
    .io_outs_2(StickySelects_15_io_outs_2),
    .io_outs_3(StickySelects_15_io_outs_3),
    .io_outs_4(StickySelects_15_io_outs_4),
    .io_outs_5(StickySelects_15_io_outs_5)
  );
  RetimeWrapper_52 RetimeWrapper ( // @[package.scala 93:22:@9199.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_1 ( // @[package.scala 93:22:@9207.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_2 ( // @[package.scala 93:22:@9215.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_3 ( // @[package.scala 93:22:@9223.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_4 ( // @[package.scala 93:22:@9247.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_5 ( // @[package.scala 93:22:@9255.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_6 ( // @[package.scala 93:22:@9263.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_7 ( // @[package.scala 93:22:@9271.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_8 ( // @[package.scala 93:22:@9295.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_9 ( // @[package.scala 93:22:@9303.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_10 ( // @[package.scala 93:22:@9311.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_11 ( // @[package.scala 93:22:@9319.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_12 ( // @[package.scala 93:22:@9343.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_13 ( // @[package.scala 93:22:@9351.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_14 ( // @[package.scala 93:22:@9359.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_15 ( // @[package.scala 93:22:@9367.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_16 ( // @[package.scala 93:22:@9391.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_17 ( // @[package.scala 93:22:@9399.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_18 ( // @[package.scala 93:22:@9407.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_19 ( // @[package.scala 93:22:@9415.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_20 ( // @[package.scala 93:22:@9439.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_21 ( // @[package.scala 93:22:@9447.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_22 ( // @[package.scala 93:22:@9455.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_23 ( // @[package.scala 93:22:@9463.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_24 ( // @[package.scala 93:22:@9487.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_25 ( // @[package.scala 93:22:@9495.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_26 ( // @[package.scala 93:22:@9503.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_27 ( // @[package.scala 93:22:@9511.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_28 ( // @[package.scala 93:22:@9535.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_29 ( // @[package.scala 93:22:@9543.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_30 ( // @[package.scala 93:22:@9551.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_31 ( // @[package.scala 93:22:@9559.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_32 ( // @[package.scala 93:22:@9583.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_33 ( // @[package.scala 93:22:@9591.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_34 ( // @[package.scala 93:22:@9599.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_35 ( // @[package.scala 93:22:@9607.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_36 ( // @[package.scala 93:22:@9631.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_37 ( // @[package.scala 93:22:@9639.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_38 ( // @[package.scala 93:22:@9647.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_39 ( // @[package.scala 93:22:@9655.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_40 ( // @[package.scala 93:22:@9679.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_41 ( // @[package.scala 93:22:@9687.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_42 ( // @[package.scala 93:22:@9695.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_43 ( // @[package.scala 93:22:@9703.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_44 ( // @[package.scala 93:22:@9727.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_45 ( // @[package.scala 93:22:@9735.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_46 ( // @[package.scala 93:22:@9743.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_47 ( // @[package.scala 93:22:@9751.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_48 ( // @[package.scala 93:22:@9775.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_49 ( // @[package.scala 93:22:@9783.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_50 ( // @[package.scala 93:22:@9791.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_51 ( // @[package.scala 93:22:@9799.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_52 ( // @[package.scala 93:22:@9823.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_53 ( // @[package.scala 93:22:@9831.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_54 ( // @[package.scala 93:22:@9839.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_55 ( // @[package.scala 93:22:@9847.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_56 ( // @[package.scala 93:22:@9871.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_57 ( // @[package.scala 93:22:@9879.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_58 ( // @[package.scala 93:22:@9887.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_59 ( // @[package.scala 93:22:@9895.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_60 ( // @[package.scala 93:22:@9919.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_61 ( // @[package.scala 93:22:@9927.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_62 ( // @[package.scala 93:22:@9935.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_63 ( // @[package.scala 93:22:@9943.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_64 ( // @[package.scala 93:22:@9967.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_65 ( // @[package.scala 93:22:@9975.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_66 ( // @[package.scala 93:22:@9983.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_67 ( // @[package.scala 93:22:@9991.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_68 ( // @[package.scala 93:22:@10015.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_69 ( // @[package.scala 93:22:@10023.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_70 ( // @[package.scala 93:22:@10031.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_71 ( // @[package.scala 93:22:@10039.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  assign _T_700 = io_wPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@8306.4]
  assign _T_703 = io_wPort_0_en_0 & _T_700; // @[MemPrimitives.scala 83:102:@8308.4]
  assign _T_705 = {_T_703,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@8310.4]
  assign _T_710 = io_wPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@8317.4]
  assign _T_713 = io_wPort_1_en_0 & _T_710; // @[MemPrimitives.scala 83:102:@8319.4]
  assign _T_715 = {_T_713,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@8321.4]
  assign _T_720 = io_wPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@8328.4]
  assign _T_723 = io_wPort_2_en_0 & _T_720; // @[MemPrimitives.scala 83:102:@8330.4]
  assign _T_725 = {_T_723,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@8332.4]
  assign _T_730 = io_wPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@8339.4]
  assign _T_733 = io_wPort_3_en_0 & _T_730; // @[MemPrimitives.scala 83:102:@8341.4]
  assign _T_735 = {_T_733,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@8343.4]
  assign _T_740 = io_wPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@8350.4]
  assign _T_743 = io_wPort_0_en_0 & _T_740; // @[MemPrimitives.scala 83:102:@8352.4]
  assign _T_745 = {_T_743,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@8354.4]
  assign _T_750 = io_wPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@8361.4]
  assign _T_753 = io_wPort_1_en_0 & _T_750; // @[MemPrimitives.scala 83:102:@8363.4]
  assign _T_755 = {_T_753,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@8365.4]
  assign _T_760 = io_wPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@8372.4]
  assign _T_763 = io_wPort_2_en_0 & _T_760; // @[MemPrimitives.scala 83:102:@8374.4]
  assign _T_765 = {_T_763,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@8376.4]
  assign _T_770 = io_wPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@8383.4]
  assign _T_773 = io_wPort_3_en_0 & _T_770; // @[MemPrimitives.scala 83:102:@8385.4]
  assign _T_775 = {_T_773,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@8387.4]
  assign _T_780 = io_wPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@8394.4]
  assign _T_783 = io_wPort_0_en_0 & _T_780; // @[MemPrimitives.scala 83:102:@8396.4]
  assign _T_785 = {_T_783,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@8398.4]
  assign _T_790 = io_wPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@8405.4]
  assign _T_793 = io_wPort_1_en_0 & _T_790; // @[MemPrimitives.scala 83:102:@8407.4]
  assign _T_795 = {_T_793,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@8409.4]
  assign _T_800 = io_wPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@8416.4]
  assign _T_803 = io_wPort_2_en_0 & _T_800; // @[MemPrimitives.scala 83:102:@8418.4]
  assign _T_805 = {_T_803,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@8420.4]
  assign _T_810 = io_wPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@8427.4]
  assign _T_813 = io_wPort_3_en_0 & _T_810; // @[MemPrimitives.scala 83:102:@8429.4]
  assign _T_815 = {_T_813,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@8431.4]
  assign _T_820 = io_wPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@8438.4]
  assign _T_823 = io_wPort_0_en_0 & _T_820; // @[MemPrimitives.scala 83:102:@8440.4]
  assign _T_825 = {_T_823,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@8442.4]
  assign _T_830 = io_wPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@8449.4]
  assign _T_833 = io_wPort_1_en_0 & _T_830; // @[MemPrimitives.scala 83:102:@8451.4]
  assign _T_835 = {_T_833,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@8453.4]
  assign _T_840 = io_wPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@8460.4]
  assign _T_843 = io_wPort_2_en_0 & _T_840; // @[MemPrimitives.scala 83:102:@8462.4]
  assign _T_845 = {_T_843,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@8464.4]
  assign _T_850 = io_wPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@8471.4]
  assign _T_853 = io_wPort_3_en_0 & _T_850; // @[MemPrimitives.scala 83:102:@8473.4]
  assign _T_855 = {_T_853,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@8475.4]
  assign _T_860 = io_rPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@8482.4]
  assign _T_865 = io_rPort_11_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@8485.4]
  assign _T_870 = io_rPort_15_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@8488.4]
  assign _T_874 = StickySelects_io_outs_0; // @[MemPrimitives.scala 123:41:@8497.4]
  assign _T_875 = StickySelects_io_outs_1; // @[MemPrimitives.scala 123:41:@8498.4]
  assign _T_876 = StickySelects_io_outs_2; // @[MemPrimitives.scala 123:41:@8499.4]
  assign _T_878 = {_T_874,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@8501.4]
  assign _T_880 = {_T_875,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@8503.4]
  assign _T_882 = {_T_876,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@8505.4]
  assign _T_883 = _T_875 ? _T_880 : _T_882; // @[Mux.scala 31:69:@8506.4]
  assign _T_884 = _T_874 ? _T_878 : _T_883; // @[Mux.scala 31:69:@8507.4]
  assign _T_889 = io_rPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@8514.4]
  assign _T_894 = io_rPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@8517.4]
  assign _T_899 = io_rPort_14_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@8520.4]
  assign _T_903 = StickySelects_1_io_outs_0; // @[MemPrimitives.scala 123:41:@8529.4]
  assign _T_904 = StickySelects_1_io_outs_1; // @[MemPrimitives.scala 123:41:@8530.4]
  assign _T_905 = StickySelects_1_io_outs_2; // @[MemPrimitives.scala 123:41:@8531.4]
  assign _T_907 = {_T_903,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@8533.4]
  assign _T_909 = {_T_904,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@8535.4]
  assign _T_911 = {_T_905,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@8537.4]
  assign _T_912 = _T_904 ? _T_909 : _T_911; // @[Mux.scala 31:69:@8538.4]
  assign _T_913 = _T_903 ? _T_907 : _T_912; // @[Mux.scala 31:69:@8539.4]
  assign _T_918 = io_rPort_4_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@8546.4]
  assign _T_923 = io_rPort_5_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@8549.4]
  assign _T_928 = io_rPort_6_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@8552.4]
  assign _T_933 = io_rPort_8_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@8555.4]
  assign _T_938 = io_rPort_9_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@8558.4]
  assign _T_943 = io_rPort_17_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@8561.4]
  assign _T_947 = StickySelects_2_io_outs_0; // @[MemPrimitives.scala 123:41:@8573.4]
  assign _T_948 = StickySelects_2_io_outs_1; // @[MemPrimitives.scala 123:41:@8574.4]
  assign _T_949 = StickySelects_2_io_outs_2; // @[MemPrimitives.scala 123:41:@8575.4]
  assign _T_950 = StickySelects_2_io_outs_3; // @[MemPrimitives.scala 123:41:@8576.4]
  assign _T_951 = StickySelects_2_io_outs_4; // @[MemPrimitives.scala 123:41:@8577.4]
  assign _T_952 = StickySelects_2_io_outs_5; // @[MemPrimitives.scala 123:41:@8578.4]
  assign _T_954 = {_T_947,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@8580.4]
  assign _T_956 = {_T_948,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@8582.4]
  assign _T_958 = {_T_949,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@8584.4]
  assign _T_960 = {_T_950,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@8586.4]
  assign _T_962 = {_T_951,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@8588.4]
  assign _T_964 = {_T_952,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@8590.4]
  assign _T_965 = _T_951 ? _T_962 : _T_964; // @[Mux.scala 31:69:@8591.4]
  assign _T_966 = _T_950 ? _T_960 : _T_965; // @[Mux.scala 31:69:@8592.4]
  assign _T_967 = _T_949 ? _T_958 : _T_966; // @[Mux.scala 31:69:@8593.4]
  assign _T_968 = _T_948 ? _T_956 : _T_967; // @[Mux.scala 31:69:@8594.4]
  assign _T_969 = _T_947 ? _T_954 : _T_968; // @[Mux.scala 31:69:@8595.4]
  assign _T_974 = io_rPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@8602.4]
  assign _T_979 = io_rPort_7_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@8605.4]
  assign _T_984 = io_rPort_10_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@8608.4]
  assign _T_989 = io_rPort_12_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@8611.4]
  assign _T_994 = io_rPort_13_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@8614.4]
  assign _T_999 = io_rPort_16_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@8617.4]
  assign _T_1003 = StickySelects_3_io_outs_0; // @[MemPrimitives.scala 123:41:@8629.4]
  assign _T_1004 = StickySelects_3_io_outs_1; // @[MemPrimitives.scala 123:41:@8630.4]
  assign _T_1005 = StickySelects_3_io_outs_2; // @[MemPrimitives.scala 123:41:@8631.4]
  assign _T_1006 = StickySelects_3_io_outs_3; // @[MemPrimitives.scala 123:41:@8632.4]
  assign _T_1007 = StickySelects_3_io_outs_4; // @[MemPrimitives.scala 123:41:@8633.4]
  assign _T_1008 = StickySelects_3_io_outs_5; // @[MemPrimitives.scala 123:41:@8634.4]
  assign _T_1010 = {_T_1003,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@8636.4]
  assign _T_1012 = {_T_1004,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@8638.4]
  assign _T_1014 = {_T_1005,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@8640.4]
  assign _T_1016 = {_T_1006,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@8642.4]
  assign _T_1018 = {_T_1007,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@8644.4]
  assign _T_1020 = {_T_1008,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@8646.4]
  assign _T_1021 = _T_1007 ? _T_1018 : _T_1020; // @[Mux.scala 31:69:@8647.4]
  assign _T_1022 = _T_1006 ? _T_1016 : _T_1021; // @[Mux.scala 31:69:@8648.4]
  assign _T_1023 = _T_1005 ? _T_1014 : _T_1022; // @[Mux.scala 31:69:@8649.4]
  assign _T_1024 = _T_1004 ? _T_1012 : _T_1023; // @[Mux.scala 31:69:@8650.4]
  assign _T_1025 = _T_1003 ? _T_1010 : _T_1024; // @[Mux.scala 31:69:@8651.4]
  assign _T_1030 = io_rPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@8658.4]
  assign _T_1035 = io_rPort_11_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@8661.4]
  assign _T_1040 = io_rPort_15_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@8664.4]
  assign _T_1044 = StickySelects_4_io_outs_0; // @[MemPrimitives.scala 123:41:@8673.4]
  assign _T_1045 = StickySelects_4_io_outs_1; // @[MemPrimitives.scala 123:41:@8674.4]
  assign _T_1046 = StickySelects_4_io_outs_2; // @[MemPrimitives.scala 123:41:@8675.4]
  assign _T_1048 = {_T_1044,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@8677.4]
  assign _T_1050 = {_T_1045,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@8679.4]
  assign _T_1052 = {_T_1046,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@8681.4]
  assign _T_1053 = _T_1045 ? _T_1050 : _T_1052; // @[Mux.scala 31:69:@8682.4]
  assign _T_1054 = _T_1044 ? _T_1048 : _T_1053; // @[Mux.scala 31:69:@8683.4]
  assign _T_1059 = io_rPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@8690.4]
  assign _T_1064 = io_rPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@8693.4]
  assign _T_1069 = io_rPort_14_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@8696.4]
  assign _T_1073 = StickySelects_5_io_outs_0; // @[MemPrimitives.scala 123:41:@8705.4]
  assign _T_1074 = StickySelects_5_io_outs_1; // @[MemPrimitives.scala 123:41:@8706.4]
  assign _T_1075 = StickySelects_5_io_outs_2; // @[MemPrimitives.scala 123:41:@8707.4]
  assign _T_1077 = {_T_1073,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@8709.4]
  assign _T_1079 = {_T_1074,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@8711.4]
  assign _T_1081 = {_T_1075,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@8713.4]
  assign _T_1082 = _T_1074 ? _T_1079 : _T_1081; // @[Mux.scala 31:69:@8714.4]
  assign _T_1083 = _T_1073 ? _T_1077 : _T_1082; // @[Mux.scala 31:69:@8715.4]
  assign _T_1088 = io_rPort_4_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@8722.4]
  assign _T_1093 = io_rPort_5_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@8725.4]
  assign _T_1098 = io_rPort_6_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@8728.4]
  assign _T_1103 = io_rPort_8_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@8731.4]
  assign _T_1108 = io_rPort_9_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@8734.4]
  assign _T_1113 = io_rPort_17_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@8737.4]
  assign _T_1117 = StickySelects_6_io_outs_0; // @[MemPrimitives.scala 123:41:@8749.4]
  assign _T_1118 = StickySelects_6_io_outs_1; // @[MemPrimitives.scala 123:41:@8750.4]
  assign _T_1119 = StickySelects_6_io_outs_2; // @[MemPrimitives.scala 123:41:@8751.4]
  assign _T_1120 = StickySelects_6_io_outs_3; // @[MemPrimitives.scala 123:41:@8752.4]
  assign _T_1121 = StickySelects_6_io_outs_4; // @[MemPrimitives.scala 123:41:@8753.4]
  assign _T_1122 = StickySelects_6_io_outs_5; // @[MemPrimitives.scala 123:41:@8754.4]
  assign _T_1124 = {_T_1117,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@8756.4]
  assign _T_1126 = {_T_1118,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@8758.4]
  assign _T_1128 = {_T_1119,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@8760.4]
  assign _T_1130 = {_T_1120,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@8762.4]
  assign _T_1132 = {_T_1121,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@8764.4]
  assign _T_1134 = {_T_1122,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@8766.4]
  assign _T_1135 = _T_1121 ? _T_1132 : _T_1134; // @[Mux.scala 31:69:@8767.4]
  assign _T_1136 = _T_1120 ? _T_1130 : _T_1135; // @[Mux.scala 31:69:@8768.4]
  assign _T_1137 = _T_1119 ? _T_1128 : _T_1136; // @[Mux.scala 31:69:@8769.4]
  assign _T_1138 = _T_1118 ? _T_1126 : _T_1137; // @[Mux.scala 31:69:@8770.4]
  assign _T_1139 = _T_1117 ? _T_1124 : _T_1138; // @[Mux.scala 31:69:@8771.4]
  assign _T_1144 = io_rPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@8778.4]
  assign _T_1149 = io_rPort_7_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@8781.4]
  assign _T_1154 = io_rPort_10_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@8784.4]
  assign _T_1159 = io_rPort_12_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@8787.4]
  assign _T_1164 = io_rPort_13_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@8790.4]
  assign _T_1169 = io_rPort_16_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@8793.4]
  assign _T_1173 = StickySelects_7_io_outs_0; // @[MemPrimitives.scala 123:41:@8805.4]
  assign _T_1174 = StickySelects_7_io_outs_1; // @[MemPrimitives.scala 123:41:@8806.4]
  assign _T_1175 = StickySelects_7_io_outs_2; // @[MemPrimitives.scala 123:41:@8807.4]
  assign _T_1176 = StickySelects_7_io_outs_3; // @[MemPrimitives.scala 123:41:@8808.4]
  assign _T_1177 = StickySelects_7_io_outs_4; // @[MemPrimitives.scala 123:41:@8809.4]
  assign _T_1178 = StickySelects_7_io_outs_5; // @[MemPrimitives.scala 123:41:@8810.4]
  assign _T_1180 = {_T_1173,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@8812.4]
  assign _T_1182 = {_T_1174,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@8814.4]
  assign _T_1184 = {_T_1175,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@8816.4]
  assign _T_1186 = {_T_1176,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@8818.4]
  assign _T_1188 = {_T_1177,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@8820.4]
  assign _T_1190 = {_T_1178,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@8822.4]
  assign _T_1191 = _T_1177 ? _T_1188 : _T_1190; // @[Mux.scala 31:69:@8823.4]
  assign _T_1192 = _T_1176 ? _T_1186 : _T_1191; // @[Mux.scala 31:69:@8824.4]
  assign _T_1193 = _T_1175 ? _T_1184 : _T_1192; // @[Mux.scala 31:69:@8825.4]
  assign _T_1194 = _T_1174 ? _T_1182 : _T_1193; // @[Mux.scala 31:69:@8826.4]
  assign _T_1195 = _T_1173 ? _T_1180 : _T_1194; // @[Mux.scala 31:69:@8827.4]
  assign _T_1200 = io_rPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@8834.4]
  assign _T_1205 = io_rPort_11_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@8837.4]
  assign _T_1210 = io_rPort_15_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@8840.4]
  assign _T_1214 = StickySelects_8_io_outs_0; // @[MemPrimitives.scala 123:41:@8849.4]
  assign _T_1215 = StickySelects_8_io_outs_1; // @[MemPrimitives.scala 123:41:@8850.4]
  assign _T_1216 = StickySelects_8_io_outs_2; // @[MemPrimitives.scala 123:41:@8851.4]
  assign _T_1218 = {_T_1214,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@8853.4]
  assign _T_1220 = {_T_1215,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@8855.4]
  assign _T_1222 = {_T_1216,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@8857.4]
  assign _T_1223 = _T_1215 ? _T_1220 : _T_1222; // @[Mux.scala 31:69:@8858.4]
  assign _T_1224 = _T_1214 ? _T_1218 : _T_1223; // @[Mux.scala 31:69:@8859.4]
  assign _T_1229 = io_rPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@8866.4]
  assign _T_1234 = io_rPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@8869.4]
  assign _T_1239 = io_rPort_14_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@8872.4]
  assign _T_1243 = StickySelects_9_io_outs_0; // @[MemPrimitives.scala 123:41:@8881.4]
  assign _T_1244 = StickySelects_9_io_outs_1; // @[MemPrimitives.scala 123:41:@8882.4]
  assign _T_1245 = StickySelects_9_io_outs_2; // @[MemPrimitives.scala 123:41:@8883.4]
  assign _T_1247 = {_T_1243,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@8885.4]
  assign _T_1249 = {_T_1244,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@8887.4]
  assign _T_1251 = {_T_1245,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@8889.4]
  assign _T_1252 = _T_1244 ? _T_1249 : _T_1251; // @[Mux.scala 31:69:@8890.4]
  assign _T_1253 = _T_1243 ? _T_1247 : _T_1252; // @[Mux.scala 31:69:@8891.4]
  assign _T_1258 = io_rPort_4_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@8898.4]
  assign _T_1263 = io_rPort_5_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@8901.4]
  assign _T_1268 = io_rPort_6_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@8904.4]
  assign _T_1273 = io_rPort_8_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@8907.4]
  assign _T_1278 = io_rPort_9_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@8910.4]
  assign _T_1283 = io_rPort_17_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@8913.4]
  assign _T_1287 = StickySelects_10_io_outs_0; // @[MemPrimitives.scala 123:41:@8925.4]
  assign _T_1288 = StickySelects_10_io_outs_1; // @[MemPrimitives.scala 123:41:@8926.4]
  assign _T_1289 = StickySelects_10_io_outs_2; // @[MemPrimitives.scala 123:41:@8927.4]
  assign _T_1290 = StickySelects_10_io_outs_3; // @[MemPrimitives.scala 123:41:@8928.4]
  assign _T_1291 = StickySelects_10_io_outs_4; // @[MemPrimitives.scala 123:41:@8929.4]
  assign _T_1292 = StickySelects_10_io_outs_5; // @[MemPrimitives.scala 123:41:@8930.4]
  assign _T_1294 = {_T_1287,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@8932.4]
  assign _T_1296 = {_T_1288,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@8934.4]
  assign _T_1298 = {_T_1289,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@8936.4]
  assign _T_1300 = {_T_1290,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@8938.4]
  assign _T_1302 = {_T_1291,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@8940.4]
  assign _T_1304 = {_T_1292,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@8942.4]
  assign _T_1305 = _T_1291 ? _T_1302 : _T_1304; // @[Mux.scala 31:69:@8943.4]
  assign _T_1306 = _T_1290 ? _T_1300 : _T_1305; // @[Mux.scala 31:69:@8944.4]
  assign _T_1307 = _T_1289 ? _T_1298 : _T_1306; // @[Mux.scala 31:69:@8945.4]
  assign _T_1308 = _T_1288 ? _T_1296 : _T_1307; // @[Mux.scala 31:69:@8946.4]
  assign _T_1309 = _T_1287 ? _T_1294 : _T_1308; // @[Mux.scala 31:69:@8947.4]
  assign _T_1314 = io_rPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@8954.4]
  assign _T_1319 = io_rPort_7_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@8957.4]
  assign _T_1324 = io_rPort_10_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@8960.4]
  assign _T_1329 = io_rPort_12_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@8963.4]
  assign _T_1334 = io_rPort_13_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@8966.4]
  assign _T_1339 = io_rPort_16_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@8969.4]
  assign _T_1343 = StickySelects_11_io_outs_0; // @[MemPrimitives.scala 123:41:@8981.4]
  assign _T_1344 = StickySelects_11_io_outs_1; // @[MemPrimitives.scala 123:41:@8982.4]
  assign _T_1345 = StickySelects_11_io_outs_2; // @[MemPrimitives.scala 123:41:@8983.4]
  assign _T_1346 = StickySelects_11_io_outs_3; // @[MemPrimitives.scala 123:41:@8984.4]
  assign _T_1347 = StickySelects_11_io_outs_4; // @[MemPrimitives.scala 123:41:@8985.4]
  assign _T_1348 = StickySelects_11_io_outs_5; // @[MemPrimitives.scala 123:41:@8986.4]
  assign _T_1350 = {_T_1343,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@8988.4]
  assign _T_1352 = {_T_1344,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@8990.4]
  assign _T_1354 = {_T_1345,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@8992.4]
  assign _T_1356 = {_T_1346,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@8994.4]
  assign _T_1358 = {_T_1347,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@8996.4]
  assign _T_1360 = {_T_1348,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@8998.4]
  assign _T_1361 = _T_1347 ? _T_1358 : _T_1360; // @[Mux.scala 31:69:@8999.4]
  assign _T_1362 = _T_1346 ? _T_1356 : _T_1361; // @[Mux.scala 31:69:@9000.4]
  assign _T_1363 = _T_1345 ? _T_1354 : _T_1362; // @[Mux.scala 31:69:@9001.4]
  assign _T_1364 = _T_1344 ? _T_1352 : _T_1363; // @[Mux.scala 31:69:@9002.4]
  assign _T_1365 = _T_1343 ? _T_1350 : _T_1364; // @[Mux.scala 31:69:@9003.4]
  assign _T_1370 = io_rPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@9010.4]
  assign _T_1375 = io_rPort_11_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@9013.4]
  assign _T_1380 = io_rPort_15_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@9016.4]
  assign _T_1384 = StickySelects_12_io_outs_0; // @[MemPrimitives.scala 123:41:@9025.4]
  assign _T_1385 = StickySelects_12_io_outs_1; // @[MemPrimitives.scala 123:41:@9026.4]
  assign _T_1386 = StickySelects_12_io_outs_2; // @[MemPrimitives.scala 123:41:@9027.4]
  assign _T_1388 = {_T_1384,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@9029.4]
  assign _T_1390 = {_T_1385,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@9031.4]
  assign _T_1392 = {_T_1386,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@9033.4]
  assign _T_1393 = _T_1385 ? _T_1390 : _T_1392; // @[Mux.scala 31:69:@9034.4]
  assign _T_1394 = _T_1384 ? _T_1388 : _T_1393; // @[Mux.scala 31:69:@9035.4]
  assign _T_1399 = io_rPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@9042.4]
  assign _T_1404 = io_rPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@9045.4]
  assign _T_1409 = io_rPort_14_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@9048.4]
  assign _T_1413 = StickySelects_13_io_outs_0; // @[MemPrimitives.scala 123:41:@9057.4]
  assign _T_1414 = StickySelects_13_io_outs_1; // @[MemPrimitives.scala 123:41:@9058.4]
  assign _T_1415 = StickySelects_13_io_outs_2; // @[MemPrimitives.scala 123:41:@9059.4]
  assign _T_1417 = {_T_1413,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@9061.4]
  assign _T_1419 = {_T_1414,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@9063.4]
  assign _T_1421 = {_T_1415,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@9065.4]
  assign _T_1422 = _T_1414 ? _T_1419 : _T_1421; // @[Mux.scala 31:69:@9066.4]
  assign _T_1423 = _T_1413 ? _T_1417 : _T_1422; // @[Mux.scala 31:69:@9067.4]
  assign _T_1428 = io_rPort_4_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@9074.4]
  assign _T_1433 = io_rPort_5_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@9077.4]
  assign _T_1438 = io_rPort_6_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@9080.4]
  assign _T_1443 = io_rPort_8_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@9083.4]
  assign _T_1448 = io_rPort_9_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@9086.4]
  assign _T_1453 = io_rPort_17_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@9089.4]
  assign _T_1457 = StickySelects_14_io_outs_0; // @[MemPrimitives.scala 123:41:@9101.4]
  assign _T_1458 = StickySelects_14_io_outs_1; // @[MemPrimitives.scala 123:41:@9102.4]
  assign _T_1459 = StickySelects_14_io_outs_2; // @[MemPrimitives.scala 123:41:@9103.4]
  assign _T_1460 = StickySelects_14_io_outs_3; // @[MemPrimitives.scala 123:41:@9104.4]
  assign _T_1461 = StickySelects_14_io_outs_4; // @[MemPrimitives.scala 123:41:@9105.4]
  assign _T_1462 = StickySelects_14_io_outs_5; // @[MemPrimitives.scala 123:41:@9106.4]
  assign _T_1464 = {_T_1457,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@9108.4]
  assign _T_1466 = {_T_1458,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@9110.4]
  assign _T_1468 = {_T_1459,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@9112.4]
  assign _T_1470 = {_T_1460,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@9114.4]
  assign _T_1472 = {_T_1461,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@9116.4]
  assign _T_1474 = {_T_1462,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@9118.4]
  assign _T_1475 = _T_1461 ? _T_1472 : _T_1474; // @[Mux.scala 31:69:@9119.4]
  assign _T_1476 = _T_1460 ? _T_1470 : _T_1475; // @[Mux.scala 31:69:@9120.4]
  assign _T_1477 = _T_1459 ? _T_1468 : _T_1476; // @[Mux.scala 31:69:@9121.4]
  assign _T_1478 = _T_1458 ? _T_1466 : _T_1477; // @[Mux.scala 31:69:@9122.4]
  assign _T_1479 = _T_1457 ? _T_1464 : _T_1478; // @[Mux.scala 31:69:@9123.4]
  assign _T_1484 = io_rPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@9130.4]
  assign _T_1489 = io_rPort_7_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@9133.4]
  assign _T_1494 = io_rPort_10_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@9136.4]
  assign _T_1499 = io_rPort_12_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@9139.4]
  assign _T_1504 = io_rPort_13_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@9142.4]
  assign _T_1509 = io_rPort_16_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@9145.4]
  assign _T_1513 = StickySelects_15_io_outs_0; // @[MemPrimitives.scala 123:41:@9157.4]
  assign _T_1514 = StickySelects_15_io_outs_1; // @[MemPrimitives.scala 123:41:@9158.4]
  assign _T_1515 = StickySelects_15_io_outs_2; // @[MemPrimitives.scala 123:41:@9159.4]
  assign _T_1516 = StickySelects_15_io_outs_3; // @[MemPrimitives.scala 123:41:@9160.4]
  assign _T_1517 = StickySelects_15_io_outs_4; // @[MemPrimitives.scala 123:41:@9161.4]
  assign _T_1518 = StickySelects_15_io_outs_5; // @[MemPrimitives.scala 123:41:@9162.4]
  assign _T_1520 = {_T_1513,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@9164.4]
  assign _T_1522 = {_T_1514,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@9166.4]
  assign _T_1524 = {_T_1515,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@9168.4]
  assign _T_1526 = {_T_1516,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@9170.4]
  assign _T_1528 = {_T_1517,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@9172.4]
  assign _T_1530 = {_T_1518,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@9174.4]
  assign _T_1531 = _T_1517 ? _T_1528 : _T_1530; // @[Mux.scala 31:69:@9175.4]
  assign _T_1532 = _T_1516 ? _T_1526 : _T_1531; // @[Mux.scala 31:69:@9176.4]
  assign _T_1533 = _T_1515 ? _T_1524 : _T_1532; // @[Mux.scala 31:69:@9177.4]
  assign _T_1534 = _T_1514 ? _T_1522 : _T_1533; // @[Mux.scala 31:69:@9178.4]
  assign _T_1535 = _T_1513 ? _T_1520 : _T_1534; // @[Mux.scala 31:69:@9179.4]
  assign _T_1567 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@9220.4 package.scala 96:25:@9221.4]
  assign _T_1571 = _T_1567 ? Mem1D_8_io_output : Mem1D_12_io_output; // @[Mux.scala 31:69:@9230.4]
  assign _T_1564 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@9212.4 package.scala 96:25:@9213.4]
  assign _T_1572 = _T_1564 ? Mem1D_4_io_output : _T_1571; // @[Mux.scala 31:69:@9231.4]
  assign _T_1561 = RetimeWrapper_io_out; // @[package.scala 96:25:@9204.4 package.scala 96:25:@9205.4]
  assign _T_1602 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@9268.4 package.scala 96:25:@9269.4]
  assign _T_1606 = _T_1602 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@9278.4]
  assign _T_1599 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@9260.4 package.scala 96:25:@9261.4]
  assign _T_1607 = _T_1599 ? Mem1D_7_io_output : _T_1606; // @[Mux.scala 31:69:@9279.4]
  assign _T_1596 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@9252.4 package.scala 96:25:@9253.4]
  assign _T_1637 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@9316.4 package.scala 96:25:@9317.4]
  assign _T_1641 = _T_1637 ? Mem1D_9_io_output : Mem1D_13_io_output; // @[Mux.scala 31:69:@9326.4]
  assign _T_1634 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@9308.4 package.scala 96:25:@9309.4]
  assign _T_1642 = _T_1634 ? Mem1D_5_io_output : _T_1641; // @[Mux.scala 31:69:@9327.4]
  assign _T_1631 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@9300.4 package.scala 96:25:@9301.4]
  assign _T_1672 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@9364.4 package.scala 96:25:@9365.4]
  assign _T_1676 = _T_1672 ? Mem1D_9_io_output : Mem1D_13_io_output; // @[Mux.scala 31:69:@9374.4]
  assign _T_1669 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@9356.4 package.scala 96:25:@9357.4]
  assign _T_1677 = _T_1669 ? Mem1D_5_io_output : _T_1676; // @[Mux.scala 31:69:@9375.4]
  assign _T_1666 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@9348.4 package.scala 96:25:@9349.4]
  assign _T_1707 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@9412.4 package.scala 96:25:@9413.4]
  assign _T_1711 = _T_1707 ? Mem1D_10_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@9422.4]
  assign _T_1704 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@9404.4 package.scala 96:25:@9405.4]
  assign _T_1712 = _T_1704 ? Mem1D_6_io_output : _T_1711; // @[Mux.scala 31:69:@9423.4]
  assign _T_1701 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@9396.4 package.scala 96:25:@9397.4]
  assign _T_1742 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@9460.4 package.scala 96:25:@9461.4]
  assign _T_1746 = _T_1742 ? Mem1D_10_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@9470.4]
  assign _T_1739 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@9452.4 package.scala 96:25:@9453.4]
  assign _T_1747 = _T_1739 ? Mem1D_6_io_output : _T_1746; // @[Mux.scala 31:69:@9471.4]
  assign _T_1736 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@9444.4 package.scala 96:25:@9445.4]
  assign _T_1777 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@9508.4 package.scala 96:25:@9509.4]
  assign _T_1781 = _T_1777 ? Mem1D_10_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@9518.4]
  assign _T_1774 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@9500.4 package.scala 96:25:@9501.4]
  assign _T_1782 = _T_1774 ? Mem1D_6_io_output : _T_1781; // @[Mux.scala 31:69:@9519.4]
  assign _T_1771 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@9492.4 package.scala 96:25:@9493.4]
  assign _T_1812 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@9556.4 package.scala 96:25:@9557.4]
  assign _T_1816 = _T_1812 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@9566.4]
  assign _T_1809 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@9548.4 package.scala 96:25:@9549.4]
  assign _T_1817 = _T_1809 ? Mem1D_7_io_output : _T_1816; // @[Mux.scala 31:69:@9567.4]
  assign _T_1806 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@9540.4 package.scala 96:25:@9541.4]
  assign _T_1847 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@9604.4 package.scala 96:25:@9605.4]
  assign _T_1851 = _T_1847 ? Mem1D_10_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@9614.4]
  assign _T_1844 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@9596.4 package.scala 96:25:@9597.4]
  assign _T_1852 = _T_1844 ? Mem1D_6_io_output : _T_1851; // @[Mux.scala 31:69:@9615.4]
  assign _T_1841 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@9588.4 package.scala 96:25:@9589.4]
  assign _T_1882 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@9652.4 package.scala 96:25:@9653.4]
  assign _T_1886 = _T_1882 ? Mem1D_10_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@9662.4]
  assign _T_1879 = RetimeWrapper_37_io_out; // @[package.scala 96:25:@9644.4 package.scala 96:25:@9645.4]
  assign _T_1887 = _T_1879 ? Mem1D_6_io_output : _T_1886; // @[Mux.scala 31:69:@9663.4]
  assign _T_1876 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@9636.4 package.scala 96:25:@9637.4]
  assign _T_1917 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@9700.4 package.scala 96:25:@9701.4]
  assign _T_1921 = _T_1917 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@9710.4]
  assign _T_1914 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@9692.4 package.scala 96:25:@9693.4]
  assign _T_1922 = _T_1914 ? Mem1D_7_io_output : _T_1921; // @[Mux.scala 31:69:@9711.4]
  assign _T_1911 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@9684.4 package.scala 96:25:@9685.4]
  assign _T_1952 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@9748.4 package.scala 96:25:@9749.4]
  assign _T_1956 = _T_1952 ? Mem1D_8_io_output : Mem1D_12_io_output; // @[Mux.scala 31:69:@9758.4]
  assign _T_1949 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@9740.4 package.scala 96:25:@9741.4]
  assign _T_1957 = _T_1949 ? Mem1D_4_io_output : _T_1956; // @[Mux.scala 31:69:@9759.4]
  assign _T_1946 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@9732.4 package.scala 96:25:@9733.4]
  assign _T_1987 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@9796.4 package.scala 96:25:@9797.4]
  assign _T_1991 = _T_1987 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@9806.4]
  assign _T_1984 = RetimeWrapper_49_io_out; // @[package.scala 96:25:@9788.4 package.scala 96:25:@9789.4]
  assign _T_1992 = _T_1984 ? Mem1D_7_io_output : _T_1991; // @[Mux.scala 31:69:@9807.4]
  assign _T_1981 = RetimeWrapper_48_io_out; // @[package.scala 96:25:@9780.4 package.scala 96:25:@9781.4]
  assign _T_2022 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@9844.4 package.scala 96:25:@9845.4]
  assign _T_2026 = _T_2022 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@9854.4]
  assign _T_2019 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@9836.4 package.scala 96:25:@9837.4]
  assign _T_2027 = _T_2019 ? Mem1D_7_io_output : _T_2026; // @[Mux.scala 31:69:@9855.4]
  assign _T_2016 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@9828.4 package.scala 96:25:@9829.4]
  assign _T_2057 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@9892.4 package.scala 96:25:@9893.4]
  assign _T_2061 = _T_2057 ? Mem1D_9_io_output : Mem1D_13_io_output; // @[Mux.scala 31:69:@9902.4]
  assign _T_2054 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@9884.4 package.scala 96:25:@9885.4]
  assign _T_2062 = _T_2054 ? Mem1D_5_io_output : _T_2061; // @[Mux.scala 31:69:@9903.4]
  assign _T_2051 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@9876.4 package.scala 96:25:@9877.4]
  assign _T_2092 = RetimeWrapper_62_io_out; // @[package.scala 96:25:@9940.4 package.scala 96:25:@9941.4]
  assign _T_2096 = _T_2092 ? Mem1D_8_io_output : Mem1D_12_io_output; // @[Mux.scala 31:69:@9950.4]
  assign _T_2089 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@9932.4 package.scala 96:25:@9933.4]
  assign _T_2097 = _T_2089 ? Mem1D_4_io_output : _T_2096; // @[Mux.scala 31:69:@9951.4]
  assign _T_2086 = RetimeWrapper_60_io_out; // @[package.scala 96:25:@9924.4 package.scala 96:25:@9925.4]
  assign _T_2127 = RetimeWrapper_66_io_out; // @[package.scala 96:25:@9988.4 package.scala 96:25:@9989.4]
  assign _T_2131 = _T_2127 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@9998.4]
  assign _T_2124 = RetimeWrapper_65_io_out; // @[package.scala 96:25:@9980.4 package.scala 96:25:@9981.4]
  assign _T_2132 = _T_2124 ? Mem1D_7_io_output : _T_2131; // @[Mux.scala 31:69:@9999.4]
  assign _T_2121 = RetimeWrapper_64_io_out; // @[package.scala 96:25:@9972.4 package.scala 96:25:@9973.4]
  assign _T_2162 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@10036.4 package.scala 96:25:@10037.4]
  assign _T_2166 = _T_2162 ? Mem1D_10_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@10046.4]
  assign _T_2159 = RetimeWrapper_69_io_out; // @[package.scala 96:25:@10028.4 package.scala 96:25:@10029.4]
  assign _T_2167 = _T_2159 ? Mem1D_6_io_output : _T_2166; // @[Mux.scala 31:69:@10047.4]
  assign _T_2156 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@10020.4 package.scala 96:25:@10021.4]
  assign io_rPort_17_output_0 = _T_2156 ? Mem1D_2_io_output : _T_2167; // @[MemPrimitives.scala 148:13:@10049.4]
  assign io_rPort_16_output_0 = _T_2121 ? Mem1D_3_io_output : _T_2132; // @[MemPrimitives.scala 148:13:@10001.4]
  assign io_rPort_15_output_0 = _T_2086 ? Mem1D_io_output : _T_2097; // @[MemPrimitives.scala 148:13:@9953.4]
  assign io_rPort_14_output_0 = _T_2051 ? Mem1D_1_io_output : _T_2062; // @[MemPrimitives.scala 148:13:@9905.4]
  assign io_rPort_13_output_0 = _T_2016 ? Mem1D_3_io_output : _T_2027; // @[MemPrimitives.scala 148:13:@9857.4]
  assign io_rPort_12_output_0 = _T_1981 ? Mem1D_3_io_output : _T_1992; // @[MemPrimitives.scala 148:13:@9809.4]
  assign io_rPort_11_output_0 = _T_1946 ? Mem1D_io_output : _T_1957; // @[MemPrimitives.scala 148:13:@9761.4]
  assign io_rPort_10_output_0 = _T_1911 ? Mem1D_3_io_output : _T_1922; // @[MemPrimitives.scala 148:13:@9713.4]
  assign io_rPort_9_output_0 = _T_1876 ? Mem1D_2_io_output : _T_1887; // @[MemPrimitives.scala 148:13:@9665.4]
  assign io_rPort_8_output_0 = _T_1841 ? Mem1D_2_io_output : _T_1852; // @[MemPrimitives.scala 148:13:@9617.4]
  assign io_rPort_7_output_0 = _T_1806 ? Mem1D_3_io_output : _T_1817; // @[MemPrimitives.scala 148:13:@9569.4]
  assign io_rPort_6_output_0 = _T_1771 ? Mem1D_2_io_output : _T_1782; // @[MemPrimitives.scala 148:13:@9521.4]
  assign io_rPort_5_output_0 = _T_1736 ? Mem1D_2_io_output : _T_1747; // @[MemPrimitives.scala 148:13:@9473.4]
  assign io_rPort_4_output_0 = _T_1701 ? Mem1D_2_io_output : _T_1712; // @[MemPrimitives.scala 148:13:@9425.4]
  assign io_rPort_3_output_0 = _T_1666 ? Mem1D_1_io_output : _T_1677; // @[MemPrimitives.scala 148:13:@9377.4]
  assign io_rPort_2_output_0 = _T_1631 ? Mem1D_1_io_output : _T_1642; // @[MemPrimitives.scala 148:13:@9329.4]
  assign io_rPort_1_output_0 = _T_1596 ? Mem1D_3_io_output : _T_1607; // @[MemPrimitives.scala 148:13:@9281.4]
  assign io_rPort_0_output_0 = _T_1561 ? Mem1D_io_output : _T_1572; // @[MemPrimitives.scala 148:13:@9233.4]
  assign Mem1D_clock = clock; // @[:@8051.4]
  assign Mem1D_reset = reset; // @[:@8052.4]
  assign Mem1D_io_r_ofs_0 = _T_884[0]; // @[MemPrimitives.scala 127:28:@8511.4]
  assign Mem1D_io_r_backpressure = _T_884[1]; // @[MemPrimitives.scala 128:32:@8512.4]
  assign Mem1D_io_w_ofs_0 = _T_705[0]; // @[MemPrimitives.scala 94:28:@8314.4]
  assign Mem1D_io_w_data_0 = _T_705[8:1]; // @[MemPrimitives.scala 95:29:@8315.4]
  assign Mem1D_io_w_en_0 = _T_705[9]; // @[MemPrimitives.scala 96:27:@8316.4]
  assign Mem1D_1_clock = clock; // @[:@8067.4]
  assign Mem1D_1_reset = reset; // @[:@8068.4]
  assign Mem1D_1_io_r_ofs_0 = _T_913[0]; // @[MemPrimitives.scala 127:28:@8543.4]
  assign Mem1D_1_io_r_backpressure = _T_913[1]; // @[MemPrimitives.scala 128:32:@8544.4]
  assign Mem1D_1_io_w_ofs_0 = _T_715[0]; // @[MemPrimitives.scala 94:28:@8325.4]
  assign Mem1D_1_io_w_data_0 = _T_715[8:1]; // @[MemPrimitives.scala 95:29:@8326.4]
  assign Mem1D_1_io_w_en_0 = _T_715[9]; // @[MemPrimitives.scala 96:27:@8327.4]
  assign Mem1D_2_clock = clock; // @[:@8083.4]
  assign Mem1D_2_reset = reset; // @[:@8084.4]
  assign Mem1D_2_io_r_ofs_0 = _T_969[0]; // @[MemPrimitives.scala 127:28:@8599.4]
  assign Mem1D_2_io_r_backpressure = _T_969[1]; // @[MemPrimitives.scala 128:32:@8600.4]
  assign Mem1D_2_io_w_ofs_0 = _T_725[0]; // @[MemPrimitives.scala 94:28:@8336.4]
  assign Mem1D_2_io_w_data_0 = _T_725[8:1]; // @[MemPrimitives.scala 95:29:@8337.4]
  assign Mem1D_2_io_w_en_0 = _T_725[9]; // @[MemPrimitives.scala 96:27:@8338.4]
  assign Mem1D_3_clock = clock; // @[:@8099.4]
  assign Mem1D_3_reset = reset; // @[:@8100.4]
  assign Mem1D_3_io_r_ofs_0 = _T_1025[0]; // @[MemPrimitives.scala 127:28:@8655.4]
  assign Mem1D_3_io_r_backpressure = _T_1025[1]; // @[MemPrimitives.scala 128:32:@8656.4]
  assign Mem1D_3_io_w_ofs_0 = _T_735[0]; // @[MemPrimitives.scala 94:28:@8347.4]
  assign Mem1D_3_io_w_data_0 = _T_735[8:1]; // @[MemPrimitives.scala 95:29:@8348.4]
  assign Mem1D_3_io_w_en_0 = _T_735[9]; // @[MemPrimitives.scala 96:27:@8349.4]
  assign Mem1D_4_clock = clock; // @[:@8115.4]
  assign Mem1D_4_reset = reset; // @[:@8116.4]
  assign Mem1D_4_io_r_ofs_0 = _T_1054[0]; // @[MemPrimitives.scala 127:28:@8687.4]
  assign Mem1D_4_io_r_backpressure = _T_1054[1]; // @[MemPrimitives.scala 128:32:@8688.4]
  assign Mem1D_4_io_w_ofs_0 = _T_745[0]; // @[MemPrimitives.scala 94:28:@8358.4]
  assign Mem1D_4_io_w_data_0 = _T_745[8:1]; // @[MemPrimitives.scala 95:29:@8359.4]
  assign Mem1D_4_io_w_en_0 = _T_745[9]; // @[MemPrimitives.scala 96:27:@8360.4]
  assign Mem1D_5_clock = clock; // @[:@8131.4]
  assign Mem1D_5_reset = reset; // @[:@8132.4]
  assign Mem1D_5_io_r_ofs_0 = _T_1083[0]; // @[MemPrimitives.scala 127:28:@8719.4]
  assign Mem1D_5_io_r_backpressure = _T_1083[1]; // @[MemPrimitives.scala 128:32:@8720.4]
  assign Mem1D_5_io_w_ofs_0 = _T_755[0]; // @[MemPrimitives.scala 94:28:@8369.4]
  assign Mem1D_5_io_w_data_0 = _T_755[8:1]; // @[MemPrimitives.scala 95:29:@8370.4]
  assign Mem1D_5_io_w_en_0 = _T_755[9]; // @[MemPrimitives.scala 96:27:@8371.4]
  assign Mem1D_6_clock = clock; // @[:@8147.4]
  assign Mem1D_6_reset = reset; // @[:@8148.4]
  assign Mem1D_6_io_r_ofs_0 = _T_1139[0]; // @[MemPrimitives.scala 127:28:@8775.4]
  assign Mem1D_6_io_r_backpressure = _T_1139[1]; // @[MemPrimitives.scala 128:32:@8776.4]
  assign Mem1D_6_io_w_ofs_0 = _T_765[0]; // @[MemPrimitives.scala 94:28:@8380.4]
  assign Mem1D_6_io_w_data_0 = _T_765[8:1]; // @[MemPrimitives.scala 95:29:@8381.4]
  assign Mem1D_6_io_w_en_0 = _T_765[9]; // @[MemPrimitives.scala 96:27:@8382.4]
  assign Mem1D_7_clock = clock; // @[:@8163.4]
  assign Mem1D_7_reset = reset; // @[:@8164.4]
  assign Mem1D_7_io_r_ofs_0 = _T_1195[0]; // @[MemPrimitives.scala 127:28:@8831.4]
  assign Mem1D_7_io_r_backpressure = _T_1195[1]; // @[MemPrimitives.scala 128:32:@8832.4]
  assign Mem1D_7_io_w_ofs_0 = _T_775[0]; // @[MemPrimitives.scala 94:28:@8391.4]
  assign Mem1D_7_io_w_data_0 = _T_775[8:1]; // @[MemPrimitives.scala 95:29:@8392.4]
  assign Mem1D_7_io_w_en_0 = _T_775[9]; // @[MemPrimitives.scala 96:27:@8393.4]
  assign Mem1D_8_clock = clock; // @[:@8179.4]
  assign Mem1D_8_reset = reset; // @[:@8180.4]
  assign Mem1D_8_io_r_ofs_0 = _T_1224[0]; // @[MemPrimitives.scala 127:28:@8863.4]
  assign Mem1D_8_io_r_backpressure = _T_1224[1]; // @[MemPrimitives.scala 128:32:@8864.4]
  assign Mem1D_8_io_w_ofs_0 = _T_785[0]; // @[MemPrimitives.scala 94:28:@8402.4]
  assign Mem1D_8_io_w_data_0 = _T_785[8:1]; // @[MemPrimitives.scala 95:29:@8403.4]
  assign Mem1D_8_io_w_en_0 = _T_785[9]; // @[MemPrimitives.scala 96:27:@8404.4]
  assign Mem1D_9_clock = clock; // @[:@8195.4]
  assign Mem1D_9_reset = reset; // @[:@8196.4]
  assign Mem1D_9_io_r_ofs_0 = _T_1253[0]; // @[MemPrimitives.scala 127:28:@8895.4]
  assign Mem1D_9_io_r_backpressure = _T_1253[1]; // @[MemPrimitives.scala 128:32:@8896.4]
  assign Mem1D_9_io_w_ofs_0 = _T_795[0]; // @[MemPrimitives.scala 94:28:@8413.4]
  assign Mem1D_9_io_w_data_0 = _T_795[8:1]; // @[MemPrimitives.scala 95:29:@8414.4]
  assign Mem1D_9_io_w_en_0 = _T_795[9]; // @[MemPrimitives.scala 96:27:@8415.4]
  assign Mem1D_10_clock = clock; // @[:@8211.4]
  assign Mem1D_10_reset = reset; // @[:@8212.4]
  assign Mem1D_10_io_r_ofs_0 = _T_1309[0]; // @[MemPrimitives.scala 127:28:@8951.4]
  assign Mem1D_10_io_r_backpressure = _T_1309[1]; // @[MemPrimitives.scala 128:32:@8952.4]
  assign Mem1D_10_io_w_ofs_0 = _T_805[0]; // @[MemPrimitives.scala 94:28:@8424.4]
  assign Mem1D_10_io_w_data_0 = _T_805[8:1]; // @[MemPrimitives.scala 95:29:@8425.4]
  assign Mem1D_10_io_w_en_0 = _T_805[9]; // @[MemPrimitives.scala 96:27:@8426.4]
  assign Mem1D_11_clock = clock; // @[:@8227.4]
  assign Mem1D_11_reset = reset; // @[:@8228.4]
  assign Mem1D_11_io_r_ofs_0 = _T_1365[0]; // @[MemPrimitives.scala 127:28:@9007.4]
  assign Mem1D_11_io_r_backpressure = _T_1365[1]; // @[MemPrimitives.scala 128:32:@9008.4]
  assign Mem1D_11_io_w_ofs_0 = _T_815[0]; // @[MemPrimitives.scala 94:28:@8435.4]
  assign Mem1D_11_io_w_data_0 = _T_815[8:1]; // @[MemPrimitives.scala 95:29:@8436.4]
  assign Mem1D_11_io_w_en_0 = _T_815[9]; // @[MemPrimitives.scala 96:27:@8437.4]
  assign Mem1D_12_clock = clock; // @[:@8243.4]
  assign Mem1D_12_reset = reset; // @[:@8244.4]
  assign Mem1D_12_io_r_ofs_0 = _T_1394[0]; // @[MemPrimitives.scala 127:28:@9039.4]
  assign Mem1D_12_io_r_backpressure = _T_1394[1]; // @[MemPrimitives.scala 128:32:@9040.4]
  assign Mem1D_12_io_w_ofs_0 = _T_825[0]; // @[MemPrimitives.scala 94:28:@8446.4]
  assign Mem1D_12_io_w_data_0 = _T_825[8:1]; // @[MemPrimitives.scala 95:29:@8447.4]
  assign Mem1D_12_io_w_en_0 = _T_825[9]; // @[MemPrimitives.scala 96:27:@8448.4]
  assign Mem1D_13_clock = clock; // @[:@8259.4]
  assign Mem1D_13_reset = reset; // @[:@8260.4]
  assign Mem1D_13_io_r_ofs_0 = _T_1423[0]; // @[MemPrimitives.scala 127:28:@9071.4]
  assign Mem1D_13_io_r_backpressure = _T_1423[1]; // @[MemPrimitives.scala 128:32:@9072.4]
  assign Mem1D_13_io_w_ofs_0 = _T_835[0]; // @[MemPrimitives.scala 94:28:@8457.4]
  assign Mem1D_13_io_w_data_0 = _T_835[8:1]; // @[MemPrimitives.scala 95:29:@8458.4]
  assign Mem1D_13_io_w_en_0 = _T_835[9]; // @[MemPrimitives.scala 96:27:@8459.4]
  assign Mem1D_14_clock = clock; // @[:@8275.4]
  assign Mem1D_14_reset = reset; // @[:@8276.4]
  assign Mem1D_14_io_r_ofs_0 = _T_1479[0]; // @[MemPrimitives.scala 127:28:@9127.4]
  assign Mem1D_14_io_r_backpressure = _T_1479[1]; // @[MemPrimitives.scala 128:32:@9128.4]
  assign Mem1D_14_io_w_ofs_0 = _T_845[0]; // @[MemPrimitives.scala 94:28:@8468.4]
  assign Mem1D_14_io_w_data_0 = _T_845[8:1]; // @[MemPrimitives.scala 95:29:@8469.4]
  assign Mem1D_14_io_w_en_0 = _T_845[9]; // @[MemPrimitives.scala 96:27:@8470.4]
  assign Mem1D_15_clock = clock; // @[:@8291.4]
  assign Mem1D_15_reset = reset; // @[:@8292.4]
  assign Mem1D_15_io_r_ofs_0 = _T_1535[0]; // @[MemPrimitives.scala 127:28:@9183.4]
  assign Mem1D_15_io_r_backpressure = _T_1535[1]; // @[MemPrimitives.scala 128:32:@9184.4]
  assign Mem1D_15_io_w_ofs_0 = _T_855[0]; // @[MemPrimitives.scala 94:28:@8479.4]
  assign Mem1D_15_io_w_data_0 = _T_855[8:1]; // @[MemPrimitives.scala 95:29:@8480.4]
  assign Mem1D_15_io_w_en_0 = _T_855[9]; // @[MemPrimitives.scala 96:27:@8481.4]
  assign StickySelects_clock = clock; // @[:@8492.4]
  assign StickySelects_reset = reset; // @[:@8493.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0 & _T_860; // @[MemPrimitives.scala 122:60:@8494.4]
  assign StickySelects_io_ins_1 = io_rPort_11_en_0 & _T_865; // @[MemPrimitives.scala 122:60:@8495.4]
  assign StickySelects_io_ins_2 = io_rPort_15_en_0 & _T_870; // @[MemPrimitives.scala 122:60:@8496.4]
  assign StickySelects_1_clock = clock; // @[:@8524.4]
  assign StickySelects_1_reset = reset; // @[:@8525.4]
  assign StickySelects_1_io_ins_0 = io_rPort_2_en_0 & _T_889; // @[MemPrimitives.scala 122:60:@8526.4]
  assign StickySelects_1_io_ins_1 = io_rPort_3_en_0 & _T_894; // @[MemPrimitives.scala 122:60:@8527.4]
  assign StickySelects_1_io_ins_2 = io_rPort_14_en_0 & _T_899; // @[MemPrimitives.scala 122:60:@8528.4]
  assign StickySelects_2_clock = clock; // @[:@8565.4]
  assign StickySelects_2_reset = reset; // @[:@8566.4]
  assign StickySelects_2_io_ins_0 = io_rPort_4_en_0 & _T_918; // @[MemPrimitives.scala 122:60:@8567.4]
  assign StickySelects_2_io_ins_1 = io_rPort_5_en_0 & _T_923; // @[MemPrimitives.scala 122:60:@8568.4]
  assign StickySelects_2_io_ins_2 = io_rPort_6_en_0 & _T_928; // @[MemPrimitives.scala 122:60:@8569.4]
  assign StickySelects_2_io_ins_3 = io_rPort_8_en_0 & _T_933; // @[MemPrimitives.scala 122:60:@8570.4]
  assign StickySelects_2_io_ins_4 = io_rPort_9_en_0 & _T_938; // @[MemPrimitives.scala 122:60:@8571.4]
  assign StickySelects_2_io_ins_5 = io_rPort_17_en_0 & _T_943; // @[MemPrimitives.scala 122:60:@8572.4]
  assign StickySelects_3_clock = clock; // @[:@8621.4]
  assign StickySelects_3_reset = reset; // @[:@8622.4]
  assign StickySelects_3_io_ins_0 = io_rPort_1_en_0 & _T_974; // @[MemPrimitives.scala 122:60:@8623.4]
  assign StickySelects_3_io_ins_1 = io_rPort_7_en_0 & _T_979; // @[MemPrimitives.scala 122:60:@8624.4]
  assign StickySelects_3_io_ins_2 = io_rPort_10_en_0 & _T_984; // @[MemPrimitives.scala 122:60:@8625.4]
  assign StickySelects_3_io_ins_3 = io_rPort_12_en_0 & _T_989; // @[MemPrimitives.scala 122:60:@8626.4]
  assign StickySelects_3_io_ins_4 = io_rPort_13_en_0 & _T_994; // @[MemPrimitives.scala 122:60:@8627.4]
  assign StickySelects_3_io_ins_5 = io_rPort_16_en_0 & _T_999; // @[MemPrimitives.scala 122:60:@8628.4]
  assign StickySelects_4_clock = clock; // @[:@8668.4]
  assign StickySelects_4_reset = reset; // @[:@8669.4]
  assign StickySelects_4_io_ins_0 = io_rPort_0_en_0 & _T_1030; // @[MemPrimitives.scala 122:60:@8670.4]
  assign StickySelects_4_io_ins_1 = io_rPort_11_en_0 & _T_1035; // @[MemPrimitives.scala 122:60:@8671.4]
  assign StickySelects_4_io_ins_2 = io_rPort_15_en_0 & _T_1040; // @[MemPrimitives.scala 122:60:@8672.4]
  assign StickySelects_5_clock = clock; // @[:@8700.4]
  assign StickySelects_5_reset = reset; // @[:@8701.4]
  assign StickySelects_5_io_ins_0 = io_rPort_2_en_0 & _T_1059; // @[MemPrimitives.scala 122:60:@8702.4]
  assign StickySelects_5_io_ins_1 = io_rPort_3_en_0 & _T_1064; // @[MemPrimitives.scala 122:60:@8703.4]
  assign StickySelects_5_io_ins_2 = io_rPort_14_en_0 & _T_1069; // @[MemPrimitives.scala 122:60:@8704.4]
  assign StickySelects_6_clock = clock; // @[:@8741.4]
  assign StickySelects_6_reset = reset; // @[:@8742.4]
  assign StickySelects_6_io_ins_0 = io_rPort_4_en_0 & _T_1088; // @[MemPrimitives.scala 122:60:@8743.4]
  assign StickySelects_6_io_ins_1 = io_rPort_5_en_0 & _T_1093; // @[MemPrimitives.scala 122:60:@8744.4]
  assign StickySelects_6_io_ins_2 = io_rPort_6_en_0 & _T_1098; // @[MemPrimitives.scala 122:60:@8745.4]
  assign StickySelects_6_io_ins_3 = io_rPort_8_en_0 & _T_1103; // @[MemPrimitives.scala 122:60:@8746.4]
  assign StickySelects_6_io_ins_4 = io_rPort_9_en_0 & _T_1108; // @[MemPrimitives.scala 122:60:@8747.4]
  assign StickySelects_6_io_ins_5 = io_rPort_17_en_0 & _T_1113; // @[MemPrimitives.scala 122:60:@8748.4]
  assign StickySelects_7_clock = clock; // @[:@8797.4]
  assign StickySelects_7_reset = reset; // @[:@8798.4]
  assign StickySelects_7_io_ins_0 = io_rPort_1_en_0 & _T_1144; // @[MemPrimitives.scala 122:60:@8799.4]
  assign StickySelects_7_io_ins_1 = io_rPort_7_en_0 & _T_1149; // @[MemPrimitives.scala 122:60:@8800.4]
  assign StickySelects_7_io_ins_2 = io_rPort_10_en_0 & _T_1154; // @[MemPrimitives.scala 122:60:@8801.4]
  assign StickySelects_7_io_ins_3 = io_rPort_12_en_0 & _T_1159; // @[MemPrimitives.scala 122:60:@8802.4]
  assign StickySelects_7_io_ins_4 = io_rPort_13_en_0 & _T_1164; // @[MemPrimitives.scala 122:60:@8803.4]
  assign StickySelects_7_io_ins_5 = io_rPort_16_en_0 & _T_1169; // @[MemPrimitives.scala 122:60:@8804.4]
  assign StickySelects_8_clock = clock; // @[:@8844.4]
  assign StickySelects_8_reset = reset; // @[:@8845.4]
  assign StickySelects_8_io_ins_0 = io_rPort_0_en_0 & _T_1200; // @[MemPrimitives.scala 122:60:@8846.4]
  assign StickySelects_8_io_ins_1 = io_rPort_11_en_0 & _T_1205; // @[MemPrimitives.scala 122:60:@8847.4]
  assign StickySelects_8_io_ins_2 = io_rPort_15_en_0 & _T_1210; // @[MemPrimitives.scala 122:60:@8848.4]
  assign StickySelects_9_clock = clock; // @[:@8876.4]
  assign StickySelects_9_reset = reset; // @[:@8877.4]
  assign StickySelects_9_io_ins_0 = io_rPort_2_en_0 & _T_1229; // @[MemPrimitives.scala 122:60:@8878.4]
  assign StickySelects_9_io_ins_1 = io_rPort_3_en_0 & _T_1234; // @[MemPrimitives.scala 122:60:@8879.4]
  assign StickySelects_9_io_ins_2 = io_rPort_14_en_0 & _T_1239; // @[MemPrimitives.scala 122:60:@8880.4]
  assign StickySelects_10_clock = clock; // @[:@8917.4]
  assign StickySelects_10_reset = reset; // @[:@8918.4]
  assign StickySelects_10_io_ins_0 = io_rPort_4_en_0 & _T_1258; // @[MemPrimitives.scala 122:60:@8919.4]
  assign StickySelects_10_io_ins_1 = io_rPort_5_en_0 & _T_1263; // @[MemPrimitives.scala 122:60:@8920.4]
  assign StickySelects_10_io_ins_2 = io_rPort_6_en_0 & _T_1268; // @[MemPrimitives.scala 122:60:@8921.4]
  assign StickySelects_10_io_ins_3 = io_rPort_8_en_0 & _T_1273; // @[MemPrimitives.scala 122:60:@8922.4]
  assign StickySelects_10_io_ins_4 = io_rPort_9_en_0 & _T_1278; // @[MemPrimitives.scala 122:60:@8923.4]
  assign StickySelects_10_io_ins_5 = io_rPort_17_en_0 & _T_1283; // @[MemPrimitives.scala 122:60:@8924.4]
  assign StickySelects_11_clock = clock; // @[:@8973.4]
  assign StickySelects_11_reset = reset; // @[:@8974.4]
  assign StickySelects_11_io_ins_0 = io_rPort_1_en_0 & _T_1314; // @[MemPrimitives.scala 122:60:@8975.4]
  assign StickySelects_11_io_ins_1 = io_rPort_7_en_0 & _T_1319; // @[MemPrimitives.scala 122:60:@8976.4]
  assign StickySelects_11_io_ins_2 = io_rPort_10_en_0 & _T_1324; // @[MemPrimitives.scala 122:60:@8977.4]
  assign StickySelects_11_io_ins_3 = io_rPort_12_en_0 & _T_1329; // @[MemPrimitives.scala 122:60:@8978.4]
  assign StickySelects_11_io_ins_4 = io_rPort_13_en_0 & _T_1334; // @[MemPrimitives.scala 122:60:@8979.4]
  assign StickySelects_11_io_ins_5 = io_rPort_16_en_0 & _T_1339; // @[MemPrimitives.scala 122:60:@8980.4]
  assign StickySelects_12_clock = clock; // @[:@9020.4]
  assign StickySelects_12_reset = reset; // @[:@9021.4]
  assign StickySelects_12_io_ins_0 = io_rPort_0_en_0 & _T_1370; // @[MemPrimitives.scala 122:60:@9022.4]
  assign StickySelects_12_io_ins_1 = io_rPort_11_en_0 & _T_1375; // @[MemPrimitives.scala 122:60:@9023.4]
  assign StickySelects_12_io_ins_2 = io_rPort_15_en_0 & _T_1380; // @[MemPrimitives.scala 122:60:@9024.4]
  assign StickySelects_13_clock = clock; // @[:@9052.4]
  assign StickySelects_13_reset = reset; // @[:@9053.4]
  assign StickySelects_13_io_ins_0 = io_rPort_2_en_0 & _T_1399; // @[MemPrimitives.scala 122:60:@9054.4]
  assign StickySelects_13_io_ins_1 = io_rPort_3_en_0 & _T_1404; // @[MemPrimitives.scala 122:60:@9055.4]
  assign StickySelects_13_io_ins_2 = io_rPort_14_en_0 & _T_1409; // @[MemPrimitives.scala 122:60:@9056.4]
  assign StickySelects_14_clock = clock; // @[:@9093.4]
  assign StickySelects_14_reset = reset; // @[:@9094.4]
  assign StickySelects_14_io_ins_0 = io_rPort_4_en_0 & _T_1428; // @[MemPrimitives.scala 122:60:@9095.4]
  assign StickySelects_14_io_ins_1 = io_rPort_5_en_0 & _T_1433; // @[MemPrimitives.scala 122:60:@9096.4]
  assign StickySelects_14_io_ins_2 = io_rPort_6_en_0 & _T_1438; // @[MemPrimitives.scala 122:60:@9097.4]
  assign StickySelects_14_io_ins_3 = io_rPort_8_en_0 & _T_1443; // @[MemPrimitives.scala 122:60:@9098.4]
  assign StickySelects_14_io_ins_4 = io_rPort_9_en_0 & _T_1448; // @[MemPrimitives.scala 122:60:@9099.4]
  assign StickySelects_14_io_ins_5 = io_rPort_17_en_0 & _T_1453; // @[MemPrimitives.scala 122:60:@9100.4]
  assign StickySelects_15_clock = clock; // @[:@9149.4]
  assign StickySelects_15_reset = reset; // @[:@9150.4]
  assign StickySelects_15_io_ins_0 = io_rPort_1_en_0 & _T_1484; // @[MemPrimitives.scala 122:60:@9151.4]
  assign StickySelects_15_io_ins_1 = io_rPort_7_en_0 & _T_1489; // @[MemPrimitives.scala 122:60:@9152.4]
  assign StickySelects_15_io_ins_2 = io_rPort_10_en_0 & _T_1494; // @[MemPrimitives.scala 122:60:@9153.4]
  assign StickySelects_15_io_ins_3 = io_rPort_12_en_0 & _T_1499; // @[MemPrimitives.scala 122:60:@9154.4]
  assign StickySelects_15_io_ins_4 = io_rPort_13_en_0 & _T_1504; // @[MemPrimitives.scala 122:60:@9155.4]
  assign StickySelects_15_io_ins_5 = io_rPort_16_en_0 & _T_1509; // @[MemPrimitives.scala 122:60:@9156.4]
  assign RetimeWrapper_clock = clock; // @[:@9200.4]
  assign RetimeWrapper_reset = reset; // @[:@9201.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@9203.4]
  assign RetimeWrapper_io_in = _T_860 & io_rPort_0_en_0; // @[package.scala 94:16:@9202.4]
  assign RetimeWrapper_1_clock = clock; // @[:@9208.4]
  assign RetimeWrapper_1_reset = reset; // @[:@9209.4]
  assign RetimeWrapper_1_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@9211.4]
  assign RetimeWrapper_1_io_in = _T_1030 & io_rPort_0_en_0; // @[package.scala 94:16:@9210.4]
  assign RetimeWrapper_2_clock = clock; // @[:@9216.4]
  assign RetimeWrapper_2_reset = reset; // @[:@9217.4]
  assign RetimeWrapper_2_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@9219.4]
  assign RetimeWrapper_2_io_in = _T_1200 & io_rPort_0_en_0; // @[package.scala 94:16:@9218.4]
  assign RetimeWrapper_3_clock = clock; // @[:@9224.4]
  assign RetimeWrapper_3_reset = reset; // @[:@9225.4]
  assign RetimeWrapper_3_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@9227.4]
  assign RetimeWrapper_3_io_in = _T_1370 & io_rPort_0_en_0; // @[package.scala 94:16:@9226.4]
  assign RetimeWrapper_4_clock = clock; // @[:@9248.4]
  assign RetimeWrapper_4_reset = reset; // @[:@9249.4]
  assign RetimeWrapper_4_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@9251.4]
  assign RetimeWrapper_4_io_in = _T_974 & io_rPort_1_en_0; // @[package.scala 94:16:@9250.4]
  assign RetimeWrapper_5_clock = clock; // @[:@9256.4]
  assign RetimeWrapper_5_reset = reset; // @[:@9257.4]
  assign RetimeWrapper_5_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@9259.4]
  assign RetimeWrapper_5_io_in = _T_1144 & io_rPort_1_en_0; // @[package.scala 94:16:@9258.4]
  assign RetimeWrapper_6_clock = clock; // @[:@9264.4]
  assign RetimeWrapper_6_reset = reset; // @[:@9265.4]
  assign RetimeWrapper_6_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@9267.4]
  assign RetimeWrapper_6_io_in = _T_1314 & io_rPort_1_en_0; // @[package.scala 94:16:@9266.4]
  assign RetimeWrapper_7_clock = clock; // @[:@9272.4]
  assign RetimeWrapper_7_reset = reset; // @[:@9273.4]
  assign RetimeWrapper_7_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@9275.4]
  assign RetimeWrapper_7_io_in = _T_1484 & io_rPort_1_en_0; // @[package.scala 94:16:@9274.4]
  assign RetimeWrapper_8_clock = clock; // @[:@9296.4]
  assign RetimeWrapper_8_reset = reset; // @[:@9297.4]
  assign RetimeWrapper_8_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@9299.4]
  assign RetimeWrapper_8_io_in = _T_889 & io_rPort_2_en_0; // @[package.scala 94:16:@9298.4]
  assign RetimeWrapper_9_clock = clock; // @[:@9304.4]
  assign RetimeWrapper_9_reset = reset; // @[:@9305.4]
  assign RetimeWrapper_9_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@9307.4]
  assign RetimeWrapper_9_io_in = _T_1059 & io_rPort_2_en_0; // @[package.scala 94:16:@9306.4]
  assign RetimeWrapper_10_clock = clock; // @[:@9312.4]
  assign RetimeWrapper_10_reset = reset; // @[:@9313.4]
  assign RetimeWrapper_10_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@9315.4]
  assign RetimeWrapper_10_io_in = _T_1229 & io_rPort_2_en_0; // @[package.scala 94:16:@9314.4]
  assign RetimeWrapper_11_clock = clock; // @[:@9320.4]
  assign RetimeWrapper_11_reset = reset; // @[:@9321.4]
  assign RetimeWrapper_11_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@9323.4]
  assign RetimeWrapper_11_io_in = _T_1399 & io_rPort_2_en_0; // @[package.scala 94:16:@9322.4]
  assign RetimeWrapper_12_clock = clock; // @[:@9344.4]
  assign RetimeWrapper_12_reset = reset; // @[:@9345.4]
  assign RetimeWrapper_12_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@9347.4]
  assign RetimeWrapper_12_io_in = _T_894 & io_rPort_3_en_0; // @[package.scala 94:16:@9346.4]
  assign RetimeWrapper_13_clock = clock; // @[:@9352.4]
  assign RetimeWrapper_13_reset = reset; // @[:@9353.4]
  assign RetimeWrapper_13_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@9355.4]
  assign RetimeWrapper_13_io_in = _T_1064 & io_rPort_3_en_0; // @[package.scala 94:16:@9354.4]
  assign RetimeWrapper_14_clock = clock; // @[:@9360.4]
  assign RetimeWrapper_14_reset = reset; // @[:@9361.4]
  assign RetimeWrapper_14_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@9363.4]
  assign RetimeWrapper_14_io_in = _T_1234 & io_rPort_3_en_0; // @[package.scala 94:16:@9362.4]
  assign RetimeWrapper_15_clock = clock; // @[:@9368.4]
  assign RetimeWrapper_15_reset = reset; // @[:@9369.4]
  assign RetimeWrapper_15_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@9371.4]
  assign RetimeWrapper_15_io_in = _T_1404 & io_rPort_3_en_0; // @[package.scala 94:16:@9370.4]
  assign RetimeWrapper_16_clock = clock; // @[:@9392.4]
  assign RetimeWrapper_16_reset = reset; // @[:@9393.4]
  assign RetimeWrapper_16_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@9395.4]
  assign RetimeWrapper_16_io_in = _T_918 & io_rPort_4_en_0; // @[package.scala 94:16:@9394.4]
  assign RetimeWrapper_17_clock = clock; // @[:@9400.4]
  assign RetimeWrapper_17_reset = reset; // @[:@9401.4]
  assign RetimeWrapper_17_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@9403.4]
  assign RetimeWrapper_17_io_in = _T_1088 & io_rPort_4_en_0; // @[package.scala 94:16:@9402.4]
  assign RetimeWrapper_18_clock = clock; // @[:@9408.4]
  assign RetimeWrapper_18_reset = reset; // @[:@9409.4]
  assign RetimeWrapper_18_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@9411.4]
  assign RetimeWrapper_18_io_in = _T_1258 & io_rPort_4_en_0; // @[package.scala 94:16:@9410.4]
  assign RetimeWrapper_19_clock = clock; // @[:@9416.4]
  assign RetimeWrapper_19_reset = reset; // @[:@9417.4]
  assign RetimeWrapper_19_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@9419.4]
  assign RetimeWrapper_19_io_in = _T_1428 & io_rPort_4_en_0; // @[package.scala 94:16:@9418.4]
  assign RetimeWrapper_20_clock = clock; // @[:@9440.4]
  assign RetimeWrapper_20_reset = reset; // @[:@9441.4]
  assign RetimeWrapper_20_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@9443.4]
  assign RetimeWrapper_20_io_in = _T_923 & io_rPort_5_en_0; // @[package.scala 94:16:@9442.4]
  assign RetimeWrapper_21_clock = clock; // @[:@9448.4]
  assign RetimeWrapper_21_reset = reset; // @[:@9449.4]
  assign RetimeWrapper_21_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@9451.4]
  assign RetimeWrapper_21_io_in = _T_1093 & io_rPort_5_en_0; // @[package.scala 94:16:@9450.4]
  assign RetimeWrapper_22_clock = clock; // @[:@9456.4]
  assign RetimeWrapper_22_reset = reset; // @[:@9457.4]
  assign RetimeWrapper_22_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@9459.4]
  assign RetimeWrapper_22_io_in = _T_1263 & io_rPort_5_en_0; // @[package.scala 94:16:@9458.4]
  assign RetimeWrapper_23_clock = clock; // @[:@9464.4]
  assign RetimeWrapper_23_reset = reset; // @[:@9465.4]
  assign RetimeWrapper_23_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@9467.4]
  assign RetimeWrapper_23_io_in = _T_1433 & io_rPort_5_en_0; // @[package.scala 94:16:@9466.4]
  assign RetimeWrapper_24_clock = clock; // @[:@9488.4]
  assign RetimeWrapper_24_reset = reset; // @[:@9489.4]
  assign RetimeWrapper_24_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@9491.4]
  assign RetimeWrapper_24_io_in = _T_928 & io_rPort_6_en_0; // @[package.scala 94:16:@9490.4]
  assign RetimeWrapper_25_clock = clock; // @[:@9496.4]
  assign RetimeWrapper_25_reset = reset; // @[:@9497.4]
  assign RetimeWrapper_25_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@9499.4]
  assign RetimeWrapper_25_io_in = _T_1098 & io_rPort_6_en_0; // @[package.scala 94:16:@9498.4]
  assign RetimeWrapper_26_clock = clock; // @[:@9504.4]
  assign RetimeWrapper_26_reset = reset; // @[:@9505.4]
  assign RetimeWrapper_26_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@9507.4]
  assign RetimeWrapper_26_io_in = _T_1268 & io_rPort_6_en_0; // @[package.scala 94:16:@9506.4]
  assign RetimeWrapper_27_clock = clock; // @[:@9512.4]
  assign RetimeWrapper_27_reset = reset; // @[:@9513.4]
  assign RetimeWrapper_27_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@9515.4]
  assign RetimeWrapper_27_io_in = _T_1438 & io_rPort_6_en_0; // @[package.scala 94:16:@9514.4]
  assign RetimeWrapper_28_clock = clock; // @[:@9536.4]
  assign RetimeWrapper_28_reset = reset; // @[:@9537.4]
  assign RetimeWrapper_28_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@9539.4]
  assign RetimeWrapper_28_io_in = _T_979 & io_rPort_7_en_0; // @[package.scala 94:16:@9538.4]
  assign RetimeWrapper_29_clock = clock; // @[:@9544.4]
  assign RetimeWrapper_29_reset = reset; // @[:@9545.4]
  assign RetimeWrapper_29_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@9547.4]
  assign RetimeWrapper_29_io_in = _T_1149 & io_rPort_7_en_0; // @[package.scala 94:16:@9546.4]
  assign RetimeWrapper_30_clock = clock; // @[:@9552.4]
  assign RetimeWrapper_30_reset = reset; // @[:@9553.4]
  assign RetimeWrapper_30_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@9555.4]
  assign RetimeWrapper_30_io_in = _T_1319 & io_rPort_7_en_0; // @[package.scala 94:16:@9554.4]
  assign RetimeWrapper_31_clock = clock; // @[:@9560.4]
  assign RetimeWrapper_31_reset = reset; // @[:@9561.4]
  assign RetimeWrapper_31_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@9563.4]
  assign RetimeWrapper_31_io_in = _T_1489 & io_rPort_7_en_0; // @[package.scala 94:16:@9562.4]
  assign RetimeWrapper_32_clock = clock; // @[:@9584.4]
  assign RetimeWrapper_32_reset = reset; // @[:@9585.4]
  assign RetimeWrapper_32_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@9587.4]
  assign RetimeWrapper_32_io_in = _T_933 & io_rPort_8_en_0; // @[package.scala 94:16:@9586.4]
  assign RetimeWrapper_33_clock = clock; // @[:@9592.4]
  assign RetimeWrapper_33_reset = reset; // @[:@9593.4]
  assign RetimeWrapper_33_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@9595.4]
  assign RetimeWrapper_33_io_in = _T_1103 & io_rPort_8_en_0; // @[package.scala 94:16:@9594.4]
  assign RetimeWrapper_34_clock = clock; // @[:@9600.4]
  assign RetimeWrapper_34_reset = reset; // @[:@9601.4]
  assign RetimeWrapper_34_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@9603.4]
  assign RetimeWrapper_34_io_in = _T_1273 & io_rPort_8_en_0; // @[package.scala 94:16:@9602.4]
  assign RetimeWrapper_35_clock = clock; // @[:@9608.4]
  assign RetimeWrapper_35_reset = reset; // @[:@9609.4]
  assign RetimeWrapper_35_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@9611.4]
  assign RetimeWrapper_35_io_in = _T_1443 & io_rPort_8_en_0; // @[package.scala 94:16:@9610.4]
  assign RetimeWrapper_36_clock = clock; // @[:@9632.4]
  assign RetimeWrapper_36_reset = reset; // @[:@9633.4]
  assign RetimeWrapper_36_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@9635.4]
  assign RetimeWrapper_36_io_in = _T_938 & io_rPort_9_en_0; // @[package.scala 94:16:@9634.4]
  assign RetimeWrapper_37_clock = clock; // @[:@9640.4]
  assign RetimeWrapper_37_reset = reset; // @[:@9641.4]
  assign RetimeWrapper_37_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@9643.4]
  assign RetimeWrapper_37_io_in = _T_1108 & io_rPort_9_en_0; // @[package.scala 94:16:@9642.4]
  assign RetimeWrapper_38_clock = clock; // @[:@9648.4]
  assign RetimeWrapper_38_reset = reset; // @[:@9649.4]
  assign RetimeWrapper_38_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@9651.4]
  assign RetimeWrapper_38_io_in = _T_1278 & io_rPort_9_en_0; // @[package.scala 94:16:@9650.4]
  assign RetimeWrapper_39_clock = clock; // @[:@9656.4]
  assign RetimeWrapper_39_reset = reset; // @[:@9657.4]
  assign RetimeWrapper_39_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@9659.4]
  assign RetimeWrapper_39_io_in = _T_1448 & io_rPort_9_en_0; // @[package.scala 94:16:@9658.4]
  assign RetimeWrapper_40_clock = clock; // @[:@9680.4]
  assign RetimeWrapper_40_reset = reset; // @[:@9681.4]
  assign RetimeWrapper_40_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@9683.4]
  assign RetimeWrapper_40_io_in = _T_984 & io_rPort_10_en_0; // @[package.scala 94:16:@9682.4]
  assign RetimeWrapper_41_clock = clock; // @[:@9688.4]
  assign RetimeWrapper_41_reset = reset; // @[:@9689.4]
  assign RetimeWrapper_41_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@9691.4]
  assign RetimeWrapper_41_io_in = _T_1154 & io_rPort_10_en_0; // @[package.scala 94:16:@9690.4]
  assign RetimeWrapper_42_clock = clock; // @[:@9696.4]
  assign RetimeWrapper_42_reset = reset; // @[:@9697.4]
  assign RetimeWrapper_42_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@9699.4]
  assign RetimeWrapper_42_io_in = _T_1324 & io_rPort_10_en_0; // @[package.scala 94:16:@9698.4]
  assign RetimeWrapper_43_clock = clock; // @[:@9704.4]
  assign RetimeWrapper_43_reset = reset; // @[:@9705.4]
  assign RetimeWrapper_43_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@9707.4]
  assign RetimeWrapper_43_io_in = _T_1494 & io_rPort_10_en_0; // @[package.scala 94:16:@9706.4]
  assign RetimeWrapper_44_clock = clock; // @[:@9728.4]
  assign RetimeWrapper_44_reset = reset; // @[:@9729.4]
  assign RetimeWrapper_44_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@9731.4]
  assign RetimeWrapper_44_io_in = _T_865 & io_rPort_11_en_0; // @[package.scala 94:16:@9730.4]
  assign RetimeWrapper_45_clock = clock; // @[:@9736.4]
  assign RetimeWrapper_45_reset = reset; // @[:@9737.4]
  assign RetimeWrapper_45_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@9739.4]
  assign RetimeWrapper_45_io_in = _T_1035 & io_rPort_11_en_0; // @[package.scala 94:16:@9738.4]
  assign RetimeWrapper_46_clock = clock; // @[:@9744.4]
  assign RetimeWrapper_46_reset = reset; // @[:@9745.4]
  assign RetimeWrapper_46_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@9747.4]
  assign RetimeWrapper_46_io_in = _T_1205 & io_rPort_11_en_0; // @[package.scala 94:16:@9746.4]
  assign RetimeWrapper_47_clock = clock; // @[:@9752.4]
  assign RetimeWrapper_47_reset = reset; // @[:@9753.4]
  assign RetimeWrapper_47_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@9755.4]
  assign RetimeWrapper_47_io_in = _T_1375 & io_rPort_11_en_0; // @[package.scala 94:16:@9754.4]
  assign RetimeWrapper_48_clock = clock; // @[:@9776.4]
  assign RetimeWrapper_48_reset = reset; // @[:@9777.4]
  assign RetimeWrapper_48_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@9779.4]
  assign RetimeWrapper_48_io_in = _T_989 & io_rPort_12_en_0; // @[package.scala 94:16:@9778.4]
  assign RetimeWrapper_49_clock = clock; // @[:@9784.4]
  assign RetimeWrapper_49_reset = reset; // @[:@9785.4]
  assign RetimeWrapper_49_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@9787.4]
  assign RetimeWrapper_49_io_in = _T_1159 & io_rPort_12_en_0; // @[package.scala 94:16:@9786.4]
  assign RetimeWrapper_50_clock = clock; // @[:@9792.4]
  assign RetimeWrapper_50_reset = reset; // @[:@9793.4]
  assign RetimeWrapper_50_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@9795.4]
  assign RetimeWrapper_50_io_in = _T_1329 & io_rPort_12_en_0; // @[package.scala 94:16:@9794.4]
  assign RetimeWrapper_51_clock = clock; // @[:@9800.4]
  assign RetimeWrapper_51_reset = reset; // @[:@9801.4]
  assign RetimeWrapper_51_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@9803.4]
  assign RetimeWrapper_51_io_in = _T_1499 & io_rPort_12_en_0; // @[package.scala 94:16:@9802.4]
  assign RetimeWrapper_52_clock = clock; // @[:@9824.4]
  assign RetimeWrapper_52_reset = reset; // @[:@9825.4]
  assign RetimeWrapper_52_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@9827.4]
  assign RetimeWrapper_52_io_in = _T_994 & io_rPort_13_en_0; // @[package.scala 94:16:@9826.4]
  assign RetimeWrapper_53_clock = clock; // @[:@9832.4]
  assign RetimeWrapper_53_reset = reset; // @[:@9833.4]
  assign RetimeWrapper_53_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@9835.4]
  assign RetimeWrapper_53_io_in = _T_1164 & io_rPort_13_en_0; // @[package.scala 94:16:@9834.4]
  assign RetimeWrapper_54_clock = clock; // @[:@9840.4]
  assign RetimeWrapper_54_reset = reset; // @[:@9841.4]
  assign RetimeWrapper_54_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@9843.4]
  assign RetimeWrapper_54_io_in = _T_1334 & io_rPort_13_en_0; // @[package.scala 94:16:@9842.4]
  assign RetimeWrapper_55_clock = clock; // @[:@9848.4]
  assign RetimeWrapper_55_reset = reset; // @[:@9849.4]
  assign RetimeWrapper_55_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@9851.4]
  assign RetimeWrapper_55_io_in = _T_1504 & io_rPort_13_en_0; // @[package.scala 94:16:@9850.4]
  assign RetimeWrapper_56_clock = clock; // @[:@9872.4]
  assign RetimeWrapper_56_reset = reset; // @[:@9873.4]
  assign RetimeWrapper_56_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@9875.4]
  assign RetimeWrapper_56_io_in = _T_899 & io_rPort_14_en_0; // @[package.scala 94:16:@9874.4]
  assign RetimeWrapper_57_clock = clock; // @[:@9880.4]
  assign RetimeWrapper_57_reset = reset; // @[:@9881.4]
  assign RetimeWrapper_57_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@9883.4]
  assign RetimeWrapper_57_io_in = _T_1069 & io_rPort_14_en_0; // @[package.scala 94:16:@9882.4]
  assign RetimeWrapper_58_clock = clock; // @[:@9888.4]
  assign RetimeWrapper_58_reset = reset; // @[:@9889.4]
  assign RetimeWrapper_58_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@9891.4]
  assign RetimeWrapper_58_io_in = _T_1239 & io_rPort_14_en_0; // @[package.scala 94:16:@9890.4]
  assign RetimeWrapper_59_clock = clock; // @[:@9896.4]
  assign RetimeWrapper_59_reset = reset; // @[:@9897.4]
  assign RetimeWrapper_59_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@9899.4]
  assign RetimeWrapper_59_io_in = _T_1409 & io_rPort_14_en_0; // @[package.scala 94:16:@9898.4]
  assign RetimeWrapper_60_clock = clock; // @[:@9920.4]
  assign RetimeWrapper_60_reset = reset; // @[:@9921.4]
  assign RetimeWrapper_60_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@9923.4]
  assign RetimeWrapper_60_io_in = _T_870 & io_rPort_15_en_0; // @[package.scala 94:16:@9922.4]
  assign RetimeWrapper_61_clock = clock; // @[:@9928.4]
  assign RetimeWrapper_61_reset = reset; // @[:@9929.4]
  assign RetimeWrapper_61_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@9931.4]
  assign RetimeWrapper_61_io_in = _T_1040 & io_rPort_15_en_0; // @[package.scala 94:16:@9930.4]
  assign RetimeWrapper_62_clock = clock; // @[:@9936.4]
  assign RetimeWrapper_62_reset = reset; // @[:@9937.4]
  assign RetimeWrapper_62_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@9939.4]
  assign RetimeWrapper_62_io_in = _T_1210 & io_rPort_15_en_0; // @[package.scala 94:16:@9938.4]
  assign RetimeWrapper_63_clock = clock; // @[:@9944.4]
  assign RetimeWrapper_63_reset = reset; // @[:@9945.4]
  assign RetimeWrapper_63_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@9947.4]
  assign RetimeWrapper_63_io_in = _T_1380 & io_rPort_15_en_0; // @[package.scala 94:16:@9946.4]
  assign RetimeWrapper_64_clock = clock; // @[:@9968.4]
  assign RetimeWrapper_64_reset = reset; // @[:@9969.4]
  assign RetimeWrapper_64_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@9971.4]
  assign RetimeWrapper_64_io_in = _T_999 & io_rPort_16_en_0; // @[package.scala 94:16:@9970.4]
  assign RetimeWrapper_65_clock = clock; // @[:@9976.4]
  assign RetimeWrapper_65_reset = reset; // @[:@9977.4]
  assign RetimeWrapper_65_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@9979.4]
  assign RetimeWrapper_65_io_in = _T_1169 & io_rPort_16_en_0; // @[package.scala 94:16:@9978.4]
  assign RetimeWrapper_66_clock = clock; // @[:@9984.4]
  assign RetimeWrapper_66_reset = reset; // @[:@9985.4]
  assign RetimeWrapper_66_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@9987.4]
  assign RetimeWrapper_66_io_in = _T_1339 & io_rPort_16_en_0; // @[package.scala 94:16:@9986.4]
  assign RetimeWrapper_67_clock = clock; // @[:@9992.4]
  assign RetimeWrapper_67_reset = reset; // @[:@9993.4]
  assign RetimeWrapper_67_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@9995.4]
  assign RetimeWrapper_67_io_in = _T_1509 & io_rPort_16_en_0; // @[package.scala 94:16:@9994.4]
  assign RetimeWrapper_68_clock = clock; // @[:@10016.4]
  assign RetimeWrapper_68_reset = reset; // @[:@10017.4]
  assign RetimeWrapper_68_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@10019.4]
  assign RetimeWrapper_68_io_in = _T_943 & io_rPort_17_en_0; // @[package.scala 94:16:@10018.4]
  assign RetimeWrapper_69_clock = clock; // @[:@10024.4]
  assign RetimeWrapper_69_reset = reset; // @[:@10025.4]
  assign RetimeWrapper_69_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@10027.4]
  assign RetimeWrapper_69_io_in = _T_1113 & io_rPort_17_en_0; // @[package.scala 94:16:@10026.4]
  assign RetimeWrapper_70_clock = clock; // @[:@10032.4]
  assign RetimeWrapper_70_reset = reset; // @[:@10033.4]
  assign RetimeWrapper_70_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@10035.4]
  assign RetimeWrapper_70_io_in = _T_1283 & io_rPort_17_en_0; // @[package.scala 94:16:@10034.4]
  assign RetimeWrapper_71_clock = clock; // @[:@10040.4]
  assign RetimeWrapper_71_reset = reset; // @[:@10041.4]
  assign RetimeWrapper_71_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@10043.4]
  assign RetimeWrapper_71_io_in = _T_1453 & io_rPort_17_en_0; // @[package.scala 94:16:@10042.4]
endmodule
module RetimeWrapper_124( // @[:@10063.2]
  input         clock, // @[:@10064.4]
  input         reset, // @[:@10065.4]
  input         io_flow, // @[:@10066.4]
  input  [31:0] io_in, // @[:@10066.4]
  output [31:0] io_out // @[:@10066.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@10068.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@10068.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@10068.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@10068.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@10068.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@10068.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@10068.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@10081.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@10080.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@10079.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@10078.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@10077.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@10075.4]
endmodule
module SimBlackBoxesfix2fixBox_2( // @[:@10083.2]
  input  [31:0] io_a, // @[:@10086.4]
  output [32:0] io_b // @[:@10086.4]
);
  wire  _T_20; // @[implicits.scala 69:16:@10093.4]
  assign _T_20 = io_a[31]; // @[implicits.scala 69:16:@10093.4]
  assign io_b = {_T_20,io_a}; // @[SimBlackBoxes.scala 99:40:@10098.4]
endmodule
module __2( // @[:@10100.2]
  input  [31:0] io_b, // @[:@10103.4]
  output [32:0] io_result // @[:@10103.4]
);
  wire [31:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@10108.4]
  wire [32:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@10108.4]
  SimBlackBoxesfix2fixBox_2 SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@10108.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@10121.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@10116.4]
endmodule
module fix2fixBox( // @[:@10195.2]
  input         clock, // @[:@10196.4]
  input         reset, // @[:@10197.4]
  input  [32:0] io_a, // @[:@10198.4]
  input         io_flow, // @[:@10198.4]
  output [31:0] io_b // @[:@10198.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@10208.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@10208.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@10208.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@10208.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@10208.4]
  RetimeWrapper_124 RetimeWrapper ( // @[package.scala 93:22:@10208.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@10215.4]
  assign RetimeWrapper_clock = clock; // @[:@10209.4]
  assign RetimeWrapper_reset = reset; // @[:@10210.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@10212.4]
  assign RetimeWrapper_io_in = io_a[31:0]; // @[package.scala 94:16:@10211.4]
endmodule
module x343_sum( // @[:@10217.2]
  input         clock, // @[:@10218.4]
  input         reset, // @[:@10219.4]
  input  [31:0] io_a, // @[:@10220.4]
  input  [31:0] io_b, // @[:@10220.4]
  input         io_flow, // @[:@10220.4]
  output [31:0] io_result // @[:@10220.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@10228.4]
  wire [32:0] __io_result; // @[Math.scala 709:24:@10228.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@10235.4]
  wire [32:0] __1_io_result; // @[Math.scala 709:24:@10235.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@10253.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@10253.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@10253.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@10253.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@10253.4]
  wire [32:0] a_upcast_number; // @[Math.scala 712:22:@10233.4 Math.scala 713:14:@10234.4]
  wire [32:0] b_upcast_number; // @[Math.scala 712:22:@10240.4 Math.scala 713:14:@10241.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@10242.4]
  __2 _ ( // @[Math.scala 709:24:@10228.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 709:24:@10235.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox fix2fixBox ( // @[Math.scala 141:30:@10253.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@10233.4 Math.scala 713:14:@10234.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@10240.4 Math.scala 713:14:@10241.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@10242.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@10261.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@10231.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@10238.4]
  assign fix2fixBox_clock = clock; // @[:@10254.4]
  assign fix2fixBox_reset = reset; // @[:@10255.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@10256.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@10259.4]
endmodule
module RetimeWrapper_126( // @[:@10275.2]
  input         clock, // @[:@10276.4]
  input         reset, // @[:@10277.4]
  input         io_flow, // @[:@10278.4]
  input  [31:0] io_in, // @[:@10278.4]
  output [31:0] io_out // @[:@10278.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@10280.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@10280.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@10280.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@10280.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@10280.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@10280.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(4)) sr ( // @[RetimeShiftRegister.scala 15:20:@10280.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@10293.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@10292.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@10291.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@10290.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@10289.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@10287.4]
endmodule
module RetimeWrapper_127( // @[:@10307.2]
  input   clock, // @[:@10308.4]
  input   reset, // @[:@10309.4]
  input   io_flow, // @[:@10310.4]
  input   io_in, // @[:@10310.4]
  output  io_out // @[:@10310.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@10312.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@10312.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@10312.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@10312.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@10312.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@10312.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(4)) sr ( // @[RetimeShiftRegister.scala 15:20:@10312.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@10325.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@10324.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@10323.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@10322.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@10321.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@10319.4]
endmodule
module RetimeWrapper_128( // @[:@10339.2]
  input         clock, // @[:@10340.4]
  input         reset, // @[:@10341.4]
  input         io_flow, // @[:@10342.4]
  input  [31:0] io_in, // @[:@10342.4]
  output [31:0] io_out // @[:@10342.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@10344.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@10344.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@10344.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@10344.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@10344.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@10344.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@10344.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@10357.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@10356.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@10355.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@10354.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@10353.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@10351.4]
endmodule
module RetimeWrapper_130( // @[:@10403.2]
  input        clock, // @[:@10404.4]
  input        reset, // @[:@10405.4]
  input        io_flow, // @[:@10406.4]
  input  [7:0] io_in, // @[:@10406.4]
  output [7:0] io_out // @[:@10406.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@10408.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@10408.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@10408.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@10408.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@10408.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@10408.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@10408.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@10421.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@10420.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@10419.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@10418.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@10417.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@10415.4]
endmodule
module RetimeWrapper_135( // @[:@10859.2]
  input         clock, // @[:@10860.4]
  input         reset, // @[:@10861.4]
  input         io_flow, // @[:@10862.4]
  input  [31:0] io_in, // @[:@10862.4]
  output [31:0] io_out // @[:@10862.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@10864.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@10864.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@10864.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@10864.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@10864.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@10864.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@10864.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@10877.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@10876.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@10875.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@10874.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@10873.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@10871.4]
endmodule
module RetimeWrapper_148( // @[:@11867.2]
  input         clock, // @[:@11868.4]
  input         reset, // @[:@11869.4]
  input         io_flow, // @[:@11870.4]
  input  [31:0] io_in, // @[:@11870.4]
  output [31:0] io_out // @[:@11870.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@11872.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@11872.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@11872.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@11872.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@11872.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@11872.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(6)) sr ( // @[RetimeShiftRegister.scala 15:20:@11872.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@11885.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@11884.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@11883.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@11882.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@11881.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@11879.4]
endmodule
module RetimeWrapper_155( // @[:@12239.2]
  input   clock, // @[:@12240.4]
  input   reset, // @[:@12241.4]
  input   io_flow, // @[:@12242.4]
  input   io_in, // @[:@12242.4]
  output  io_out // @[:@12242.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@12244.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@12244.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@12244.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@12244.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@12244.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@12244.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(8)) sr ( // @[RetimeShiftRegister.scala 15:20:@12244.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@12257.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@12256.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@12255.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@12254.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@12253.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@12251.4]
endmodule
module x438_rdrow( // @[:@14293.2]
  input         clock, // @[:@14294.4]
  input         reset, // @[:@14295.4]
  input  [31:0] io_a, // @[:@14296.4]
  input  [31:0] io_b, // @[:@14296.4]
  input         io_flow, // @[:@14296.4]
  output [31:0] io_result // @[:@14296.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@14304.4]
  wire [32:0] __io_result; // @[Math.scala 709:24:@14304.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@14311.4]
  wire [32:0] __1_io_result; // @[Math.scala 709:24:@14311.4]
  wire  fix2fixBox_clock; // @[Math.scala 182:30:@14330.4]
  wire  fix2fixBox_reset; // @[Math.scala 182:30:@14330.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 182:30:@14330.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 182:30:@14330.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 182:30:@14330.4]
  wire [32:0] a_upcast_number; // @[Math.scala 712:22:@14309.4 Math.scala 713:14:@14310.4]
  wire [32:0] b_upcast_number; // @[Math.scala 712:22:@14316.4 Math.scala 713:14:@14317.4]
  wire [33:0] _T_21; // @[Math.scala 177:37:@14318.4]
  wire [33:0] _T_22; // @[Math.scala 177:37:@14319.4]
  __2 _ ( // @[Math.scala 709:24:@14304.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 709:24:@14311.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox fix2fixBox ( // @[Math.scala 182:30:@14330.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@14309.4 Math.scala 713:14:@14310.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@14316.4 Math.scala 713:14:@14317.4]
  assign _T_21 = a_upcast_number - b_upcast_number; // @[Math.scala 177:37:@14318.4]
  assign _T_22 = $unsigned(_T_21); // @[Math.scala 177:37:@14319.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 188:17:@14338.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@14307.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@14314.4]
  assign fix2fixBox_clock = clock; // @[:@14331.4]
  assign fix2fixBox_reset = reset; // @[:@14332.4]
  assign fix2fixBox_io_a = _T_22[32:0]; // @[Math.scala 183:23:@14333.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 186:26:@14336.4]
endmodule
module RetimeWrapper_195( // @[:@15148.2]
  input         clock, // @[:@15149.4]
  input         reset, // @[:@15150.4]
  input         io_flow, // @[:@15151.4]
  input  [31:0] io_in, // @[:@15151.4]
  output [31:0] io_out // @[:@15151.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@15153.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@15153.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@15153.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@15153.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@15153.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@15153.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(7)) sr ( // @[RetimeShiftRegister.scala 15:20:@15153.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@15166.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@15165.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@15164.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@15163.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@15162.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@15160.4]
endmodule
module SimBlackBoxesfix2fixBox_60( // @[:@17577.2]
  input  [7:0] io_a, // @[:@17580.4]
  output [8:0] io_b // @[:@17580.4]
);
  assign io_b = {1'h0,io_a}; // @[SimBlackBoxes.scala 99:40:@17591.4]
endmodule
module __60( // @[:@17593.2]
  input  [7:0] io_b, // @[:@17596.4]
  output [8:0] io_result // @[:@17596.4]
);
  wire [7:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@17601.4]
  wire [8:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@17601.4]
  SimBlackBoxesfix2fixBox_60 SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@17601.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@17614.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@17609.4]
endmodule
module fix2fixBox_29( // @[:@17687.2]
  input        clock, // @[:@17688.4]
  input        reset, // @[:@17689.4]
  input  [8:0] io_a, // @[:@17690.4]
  input        io_flow, // @[:@17690.4]
  output [7:0] io_b // @[:@17690.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@17700.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@17700.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@17700.4]
  wire [7:0] RetimeWrapper_io_in; // @[package.scala 93:22:@17700.4]
  wire [7:0] RetimeWrapper_io_out; // @[package.scala 93:22:@17700.4]
  RetimeWrapper_21 RetimeWrapper ( // @[package.scala 93:22:@17700.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@17707.4]
  assign RetimeWrapper_clock = clock; // @[:@17701.4]
  assign RetimeWrapper_reset = reset; // @[:@17702.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@17704.4]
  assign RetimeWrapper_io_in = io_a[7:0]; // @[package.scala 94:16:@17703.4]
endmodule
module x539_x11( // @[:@17709.2]
  input        clock, // @[:@17710.4]
  input        reset, // @[:@17711.4]
  input  [7:0] io_a, // @[:@17712.4]
  input  [7:0] io_b, // @[:@17712.4]
  input        io_flow, // @[:@17712.4]
  output [7:0] io_result // @[:@17712.4]
);
  wire [7:0] __io_b; // @[Math.scala 709:24:@17720.4]
  wire [8:0] __io_result; // @[Math.scala 709:24:@17720.4]
  wire [7:0] __1_io_b; // @[Math.scala 709:24:@17727.4]
  wire [8:0] __1_io_result; // @[Math.scala 709:24:@17727.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@17737.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@17737.4]
  wire [8:0] fix2fixBox_io_a; // @[Math.scala 141:30:@17737.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@17737.4]
  wire [7:0] fix2fixBox_io_b; // @[Math.scala 141:30:@17737.4]
  wire [8:0] a_upcast_number; // @[Math.scala 712:22:@17725.4 Math.scala 713:14:@17726.4]
  wire [8:0] b_upcast_number; // @[Math.scala 712:22:@17732.4 Math.scala 713:14:@17733.4]
  wire [9:0] _T_21; // @[Math.scala 136:37:@17734.4]
  __60 _ ( // @[Math.scala 709:24:@17720.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __60 __1 ( // @[Math.scala 709:24:@17727.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_29 fix2fixBox ( // @[Math.scala 141:30:@17737.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@17725.4 Math.scala 713:14:@17726.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@17732.4 Math.scala 713:14:@17733.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@17734.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@17745.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@17723.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@17730.4]
  assign fix2fixBox_clock = clock; // @[:@17738.4]
  assign fix2fixBox_reset = reset; // @[:@17739.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@17740.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@17743.4]
endmodule
module fix2fixBox_33( // @[:@18335.2]
  input  [8:0] io_a, // @[:@18338.4]
  output [7:0] io_b // @[:@18338.4]
);
  assign io_b = io_a[7:0]; // @[Converter.scala 95:38:@18348.4]
endmodule
module x543_x11( // @[:@18350.2]
  input  [7:0] io_a, // @[:@18353.4]
  input  [7:0] io_b, // @[:@18353.4]
  output [7:0] io_result // @[:@18353.4]
);
  wire [7:0] __io_b; // @[Math.scala 709:24:@18361.4]
  wire [8:0] __io_result; // @[Math.scala 709:24:@18361.4]
  wire [7:0] __1_io_b; // @[Math.scala 709:24:@18368.4]
  wire [8:0] __1_io_result; // @[Math.scala 709:24:@18368.4]
  wire [8:0] fix2fixBox_io_a; // @[Math.scala 141:30:@18378.4]
  wire [7:0] fix2fixBox_io_b; // @[Math.scala 141:30:@18378.4]
  wire [8:0] a_upcast_number; // @[Math.scala 712:22:@18366.4 Math.scala 713:14:@18367.4]
  wire [8:0] b_upcast_number; // @[Math.scala 712:22:@18373.4 Math.scala 713:14:@18374.4]
  wire [9:0] _T_21; // @[Math.scala 136:37:@18375.4]
  __60 _ ( // @[Math.scala 709:24:@18361.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __60 __1 ( // @[Math.scala 709:24:@18368.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_33 fix2fixBox ( // @[Math.scala 141:30:@18378.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@18366.4 Math.scala 713:14:@18367.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@18373.4 Math.scala 713:14:@18374.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@18375.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@18386.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@18364.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@18371.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@18381.4]
endmodule
module x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1( // @[:@22777.2]
  input          clock, // @[:@22778.4]
  input          reset, // @[:@22779.4]
  output         io_in_x316_TREADY, // @[:@22780.4]
  input  [255:0] io_in_x316_TDATA, // @[:@22780.4]
  input  [7:0]   io_in_x316_TID, // @[:@22780.4]
  input  [7:0]   io_in_x316_TDEST, // @[:@22780.4]
  output         io_in_x317_TVALID, // @[:@22780.4]
  input          io_in_x317_TREADY, // @[:@22780.4]
  output [255:0] io_in_x317_TDATA, // @[:@22780.4]
  input          io_sigsIn_backpressure, // @[:@22780.4]
  input          io_sigsIn_datapathEn, // @[:@22780.4]
  input          io_sigsIn_break, // @[:@22780.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_1, // @[:@22780.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_0, // @[:@22780.4]
  input          io_sigsIn_cchainOutputs_0_oobs_0, // @[:@22780.4]
  input          io_sigsIn_cchainOutputs_0_oobs_1, // @[:@22780.4]
  input          io_rr // @[:@22780.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@22794.4]
  wire [31:0] __io_result; // @[Math.scala 709:24:@22794.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@22806.4]
  wire [31:0] __1_io_result; // @[Math.scala 709:24:@22806.4]
  wire  x329_lb_0_clock; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_reset; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [2:0] x329_lb_0_io_rPort_17_banks_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_17_ofs_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_17_en_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_17_backpressure; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [7:0] x329_lb_0_io_rPort_17_output_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [2:0] x329_lb_0_io_rPort_16_banks_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_16_ofs_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_16_en_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_16_backpressure; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [7:0] x329_lb_0_io_rPort_16_output_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [2:0] x329_lb_0_io_rPort_15_banks_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_15_ofs_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_15_en_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_15_backpressure; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [7:0] x329_lb_0_io_rPort_15_output_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [2:0] x329_lb_0_io_rPort_14_banks_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_14_ofs_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_14_en_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_14_backpressure; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [7:0] x329_lb_0_io_rPort_14_output_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [2:0] x329_lb_0_io_rPort_13_banks_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_13_ofs_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_13_en_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_13_backpressure; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [7:0] x329_lb_0_io_rPort_13_output_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [2:0] x329_lb_0_io_rPort_12_banks_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_12_ofs_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_12_en_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_12_backpressure; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [7:0] x329_lb_0_io_rPort_12_output_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [2:0] x329_lb_0_io_rPort_11_banks_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_11_ofs_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_11_en_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_11_backpressure; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [7:0] x329_lb_0_io_rPort_11_output_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [2:0] x329_lb_0_io_rPort_10_banks_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_10_ofs_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_10_en_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_10_backpressure; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [7:0] x329_lb_0_io_rPort_10_output_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [2:0] x329_lb_0_io_rPort_9_banks_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_9_ofs_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_9_en_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_9_backpressure; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [7:0] x329_lb_0_io_rPort_9_output_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [2:0] x329_lb_0_io_rPort_8_banks_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_8_ofs_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_8_en_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_8_backpressure; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [7:0] x329_lb_0_io_rPort_8_output_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [2:0] x329_lb_0_io_rPort_7_banks_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_7_ofs_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_7_en_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_7_backpressure; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [7:0] x329_lb_0_io_rPort_7_output_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [2:0] x329_lb_0_io_rPort_6_banks_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_6_ofs_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_6_en_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_6_backpressure; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [7:0] x329_lb_0_io_rPort_6_output_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [2:0] x329_lb_0_io_rPort_5_banks_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_5_ofs_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_5_en_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_5_backpressure; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [7:0] x329_lb_0_io_rPort_5_output_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [2:0] x329_lb_0_io_rPort_4_banks_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_4_ofs_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_4_en_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_4_backpressure; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [7:0] x329_lb_0_io_rPort_4_output_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [2:0] x329_lb_0_io_rPort_3_banks_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_3_ofs_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_3_en_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_3_backpressure; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [7:0] x329_lb_0_io_rPort_3_output_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [2:0] x329_lb_0_io_rPort_2_banks_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_2_ofs_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_2_en_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_2_backpressure; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [7:0] x329_lb_0_io_rPort_2_output_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [2:0] x329_lb_0_io_rPort_1_banks_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_1_ofs_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_1_en_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_1_backpressure; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [7:0] x329_lb_0_io_rPort_1_output_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [2:0] x329_lb_0_io_rPort_0_banks_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_0_ofs_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_0_en_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_rPort_0_backpressure; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [7:0] x329_lb_0_io_rPort_0_output_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [2:0] x329_lb_0_io_wPort_3_banks_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_wPort_3_ofs_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [7:0] x329_lb_0_io_wPort_3_data_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_wPort_3_en_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [2:0] x329_lb_0_io_wPort_2_banks_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_wPort_2_ofs_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [7:0] x329_lb_0_io_wPort_2_data_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_wPort_2_en_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [2:0] x329_lb_0_io_wPort_1_banks_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_wPort_1_ofs_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [7:0] x329_lb_0_io_wPort_1_data_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_wPort_1_en_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [2:0] x329_lb_0_io_wPort_0_banks_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_wPort_0_ofs_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire [7:0] x329_lb_0_io_wPort_0_data_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  x329_lb_0_io_wPort_0_en_0; // @[m_x329_lb_0.scala 47:17:@22816.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@22974.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@22974.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@22974.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@22974.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@22974.4]
  wire  x343_sum_1_clock; // @[Math.scala 150:24:@23074.4]
  wire  x343_sum_1_reset; // @[Math.scala 150:24:@23074.4]
  wire [31:0] x343_sum_1_io_a; // @[Math.scala 150:24:@23074.4]
  wire [31:0] x343_sum_1_io_b; // @[Math.scala 150:24:@23074.4]
  wire  x343_sum_1_io_flow; // @[Math.scala 150:24:@23074.4]
  wire [31:0] x343_sum_1_io_result; // @[Math.scala 150:24:@23074.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@23084.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@23084.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@23084.4]
  wire [31:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@23084.4]
  wire [31:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@23084.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@23093.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@23093.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@23093.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@23093.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@23093.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@23102.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@23102.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@23102.4]
  wire [31:0] RetimeWrapper_3_io_in; // @[package.scala 93:22:@23102.4]
  wire [31:0] RetimeWrapper_3_io_out; // @[package.scala 93:22:@23102.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@23111.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@23111.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@23111.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@23111.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@23111.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@23120.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@23120.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@23120.4]
  wire [7:0] RetimeWrapper_5_io_in; // @[package.scala 93:22:@23120.4]
  wire [7:0] RetimeWrapper_5_io_out; // @[package.scala 93:22:@23120.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@23133.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@23133.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@23133.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@23133.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@23133.4]
  wire  x349_rdcol_1_clock; // @[Math.scala 150:24:@23156.4]
  wire  x349_rdcol_1_reset; // @[Math.scala 150:24:@23156.4]
  wire [31:0] x349_rdcol_1_io_a; // @[Math.scala 150:24:@23156.4]
  wire [31:0] x349_rdcol_1_io_b; // @[Math.scala 150:24:@23156.4]
  wire  x349_rdcol_1_io_flow; // @[Math.scala 150:24:@23156.4]
  wire [31:0] x349_rdcol_1_io_result; // @[Math.scala 150:24:@23156.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@23177.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@23177.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@23177.4]
  wire [31:0] RetimeWrapper_7_io_in; // @[package.scala 93:22:@23177.4]
  wire [31:0] RetimeWrapper_7_io_out; // @[package.scala 93:22:@23177.4]
  wire  x353_sum_1_clock; // @[Math.scala 150:24:@23186.4]
  wire  x353_sum_1_reset; // @[Math.scala 150:24:@23186.4]
  wire [31:0] x353_sum_1_io_a; // @[Math.scala 150:24:@23186.4]
  wire [31:0] x353_sum_1_io_b; // @[Math.scala 150:24:@23186.4]
  wire  x353_sum_1_io_flow; // @[Math.scala 150:24:@23186.4]
  wire [31:0] x353_sum_1_io_result; // @[Math.scala 150:24:@23186.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@23196.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@23196.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@23196.4]
  wire [31:0] RetimeWrapper_8_io_in; // @[package.scala 93:22:@23196.4]
  wire [31:0] RetimeWrapper_8_io_out; // @[package.scala 93:22:@23196.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@23205.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@23205.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@23205.4]
  wire [7:0] RetimeWrapper_9_io_in; // @[package.scala 93:22:@23205.4]
  wire [7:0] RetimeWrapper_9_io_out; // @[package.scala 93:22:@23205.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@23218.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@23218.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@23218.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@23218.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@23218.4]
  wire  x358_rdcol_1_clock; // @[Math.scala 150:24:@23241.4]
  wire  x358_rdcol_1_reset; // @[Math.scala 150:24:@23241.4]
  wire [31:0] x358_rdcol_1_io_a; // @[Math.scala 150:24:@23241.4]
  wire [31:0] x358_rdcol_1_io_b; // @[Math.scala 150:24:@23241.4]
  wire  x358_rdcol_1_io_flow; // @[Math.scala 150:24:@23241.4]
  wire [31:0] x358_rdcol_1_io_result; // @[Math.scala 150:24:@23241.4]
  wire  x362_sum_1_clock; // @[Math.scala 150:24:@23262.4]
  wire  x362_sum_1_reset; // @[Math.scala 150:24:@23262.4]
  wire [31:0] x362_sum_1_io_a; // @[Math.scala 150:24:@23262.4]
  wire [31:0] x362_sum_1_io_b; // @[Math.scala 150:24:@23262.4]
  wire  x362_sum_1_io_flow; // @[Math.scala 150:24:@23262.4]
  wire [31:0] x362_sum_1_io_result; // @[Math.scala 150:24:@23262.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@23272.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@23272.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@23272.4]
  wire [31:0] RetimeWrapper_11_io_in; // @[package.scala 93:22:@23272.4]
  wire [31:0] RetimeWrapper_11_io_out; // @[package.scala 93:22:@23272.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@23281.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@23281.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@23281.4]
  wire [7:0] RetimeWrapper_12_io_in; // @[package.scala 93:22:@23281.4]
  wire [7:0] RetimeWrapper_12_io_out; // @[package.scala 93:22:@23281.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@23294.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@23294.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@23294.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@23294.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@23294.4]
  wire  x367_rdcol_1_clock; // @[Math.scala 150:24:@23317.4]
  wire  x367_rdcol_1_reset; // @[Math.scala 150:24:@23317.4]
  wire [31:0] x367_rdcol_1_io_a; // @[Math.scala 150:24:@23317.4]
  wire [31:0] x367_rdcol_1_io_b; // @[Math.scala 150:24:@23317.4]
  wire  x367_rdcol_1_io_flow; // @[Math.scala 150:24:@23317.4]
  wire [31:0] x367_rdcol_1_io_result; // @[Math.scala 150:24:@23317.4]
  wire  x371_sum_1_clock; // @[Math.scala 150:24:@23338.4]
  wire  x371_sum_1_reset; // @[Math.scala 150:24:@23338.4]
  wire [31:0] x371_sum_1_io_a; // @[Math.scala 150:24:@23338.4]
  wire [31:0] x371_sum_1_io_b; // @[Math.scala 150:24:@23338.4]
  wire  x371_sum_1_io_flow; // @[Math.scala 150:24:@23338.4]
  wire [31:0] x371_sum_1_io_result; // @[Math.scala 150:24:@23338.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@23348.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@23348.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@23348.4]
  wire [31:0] RetimeWrapper_14_io_in; // @[package.scala 93:22:@23348.4]
  wire [31:0] RetimeWrapper_14_io_out; // @[package.scala 93:22:@23348.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@23357.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@23357.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@23357.4]
  wire [7:0] RetimeWrapper_15_io_in; // @[package.scala 93:22:@23357.4]
  wire [7:0] RetimeWrapper_15_io_out; // @[package.scala 93:22:@23357.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@23370.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@23370.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@23370.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@23370.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@23370.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@23391.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@23391.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@23391.4]
  wire [31:0] RetimeWrapper_17_io_in; // @[package.scala 93:22:@23391.4]
  wire [31:0] RetimeWrapper_17_io_out; // @[package.scala 93:22:@23391.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@23418.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@23418.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@23418.4]
  wire [31:0] RetimeWrapper_18_io_in; // @[package.scala 93:22:@23418.4]
  wire [31:0] RetimeWrapper_18_io_out; // @[package.scala 93:22:@23418.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@23434.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@23434.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@23434.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@23434.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@23434.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@23471.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@23471.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@23471.4]
  wire [31:0] RetimeWrapper_20_io_in; // @[package.scala 93:22:@23471.4]
  wire [31:0] RetimeWrapper_20_io_out; // @[package.scala 93:22:@23471.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@23480.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@23480.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@23480.4]
  wire [31:0] RetimeWrapper_21_io_in; // @[package.scala 93:22:@23480.4]
  wire [31:0] RetimeWrapper_21_io_out; // @[package.scala 93:22:@23480.4]
  wire  x384_sum_1_clock; // @[Math.scala 150:24:@23489.4]
  wire  x384_sum_1_reset; // @[Math.scala 150:24:@23489.4]
  wire [31:0] x384_sum_1_io_a; // @[Math.scala 150:24:@23489.4]
  wire [31:0] x384_sum_1_io_b; // @[Math.scala 150:24:@23489.4]
  wire  x384_sum_1_io_flow; // @[Math.scala 150:24:@23489.4]
  wire [31:0] x384_sum_1_io_result; // @[Math.scala 150:24:@23489.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@23499.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@23499.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@23499.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@23499.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@23499.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@23508.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@23508.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@23508.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@23508.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@23508.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@23517.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@23517.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@23517.4]
  wire [31:0] RetimeWrapper_24_io_in; // @[package.scala 93:22:@23517.4]
  wire [31:0] RetimeWrapper_24_io_out; // @[package.scala 93:22:@23517.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@23526.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@23526.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@23526.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@23526.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@23526.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@23540.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@23540.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@23540.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@23540.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@23540.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@23561.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@23561.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@23561.4]
  wire [31:0] RetimeWrapper_27_io_in; // @[package.scala 93:22:@23561.4]
  wire [31:0] RetimeWrapper_27_io_out; // @[package.scala 93:22:@23561.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@23583.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@23583.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@23583.4]
  wire [31:0] RetimeWrapper_28_io_in; // @[package.scala 93:22:@23583.4]
  wire [31:0] RetimeWrapper_28_io_out; // @[package.scala 93:22:@23583.4]
  wire  x393_sum_1_clock; // @[Math.scala 150:24:@23592.4]
  wire  x393_sum_1_reset; // @[Math.scala 150:24:@23592.4]
  wire [31:0] x393_sum_1_io_a; // @[Math.scala 150:24:@23592.4]
  wire [31:0] x393_sum_1_io_b; // @[Math.scala 150:24:@23592.4]
  wire  x393_sum_1_io_flow; // @[Math.scala 150:24:@23592.4]
  wire [31:0] x393_sum_1_io_result; // @[Math.scala 150:24:@23592.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@23602.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@23602.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@23602.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@23602.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@23602.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@23616.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@23616.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@23616.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@23616.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@23616.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@23637.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@23637.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@23637.4]
  wire [31:0] RetimeWrapper_31_io_in; // @[package.scala 93:22:@23637.4]
  wire [31:0] RetimeWrapper_31_io_out; // @[package.scala 93:22:@23637.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@23659.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@23659.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@23659.4]
  wire [31:0] RetimeWrapper_32_io_in; // @[package.scala 93:22:@23659.4]
  wire [31:0] RetimeWrapper_32_io_out; // @[package.scala 93:22:@23659.4]
  wire  x401_sum_1_clock; // @[Math.scala 150:24:@23668.4]
  wire  x401_sum_1_reset; // @[Math.scala 150:24:@23668.4]
  wire [31:0] x401_sum_1_io_a; // @[Math.scala 150:24:@23668.4]
  wire [31:0] x401_sum_1_io_b; // @[Math.scala 150:24:@23668.4]
  wire  x401_sum_1_io_flow; // @[Math.scala 150:24:@23668.4]
  wire [31:0] x401_sum_1_io_result; // @[Math.scala 150:24:@23668.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@23678.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@23678.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@23678.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@23678.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@23678.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@23692.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@23692.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@23692.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@23692.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@23692.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@23713.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@23713.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@23713.4]
  wire [31:0] RetimeWrapper_35_io_in; // @[package.scala 93:22:@23713.4]
  wire [31:0] RetimeWrapper_35_io_out; // @[package.scala 93:22:@23713.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@23735.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@23735.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@23735.4]
  wire [31:0] RetimeWrapper_36_io_in; // @[package.scala 93:22:@23735.4]
  wire [31:0] RetimeWrapper_36_io_out; // @[package.scala 93:22:@23735.4]
  wire  x409_sum_1_clock; // @[Math.scala 150:24:@23744.4]
  wire  x409_sum_1_reset; // @[Math.scala 150:24:@23744.4]
  wire [31:0] x409_sum_1_io_a; // @[Math.scala 150:24:@23744.4]
  wire [31:0] x409_sum_1_io_b; // @[Math.scala 150:24:@23744.4]
  wire  x409_sum_1_io_flow; // @[Math.scala 150:24:@23744.4]
  wire [31:0] x409_sum_1_io_result; // @[Math.scala 150:24:@23744.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@23754.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@23754.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@23754.4]
  wire  RetimeWrapper_37_io_in; // @[package.scala 93:22:@23754.4]
  wire  RetimeWrapper_37_io_out; // @[package.scala 93:22:@23754.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@23763.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@23763.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@23763.4]
  wire [31:0] RetimeWrapper_38_io_in; // @[package.scala 93:22:@23763.4]
  wire [31:0] RetimeWrapper_38_io_out; // @[package.scala 93:22:@23763.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@23777.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@23777.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@23777.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@23777.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@23777.4]
  wire  x414_rdcol_1_clock; // @[Math.scala 150:24:@23800.4]
  wire  x414_rdcol_1_reset; // @[Math.scala 150:24:@23800.4]
  wire [31:0] x414_rdcol_1_io_a; // @[Math.scala 150:24:@23800.4]
  wire [31:0] x414_rdcol_1_io_b; // @[Math.scala 150:24:@23800.4]
  wire  x414_rdcol_1_io_flow; // @[Math.scala 150:24:@23800.4]
  wire [31:0] x414_rdcol_1_io_result; // @[Math.scala 150:24:@23800.4]
  wire  x420_sum_1_clock; // @[Math.scala 150:24:@23832.4]
  wire  x420_sum_1_reset; // @[Math.scala 150:24:@23832.4]
  wire [31:0] x420_sum_1_io_a; // @[Math.scala 150:24:@23832.4]
  wire [31:0] x420_sum_1_io_b; // @[Math.scala 150:24:@23832.4]
  wire  x420_sum_1_io_flow; // @[Math.scala 150:24:@23832.4]
  wire [31:0] x420_sum_1_io_result; // @[Math.scala 150:24:@23832.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@23842.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@23842.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@23842.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@23842.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@23842.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@23856.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@23856.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@23856.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@23856.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@23856.4]
  wire  x426_rdcol_1_clock; // @[Math.scala 150:24:@23881.4]
  wire  x426_rdcol_1_reset; // @[Math.scala 150:24:@23881.4]
  wire [31:0] x426_rdcol_1_io_a; // @[Math.scala 150:24:@23881.4]
  wire [31:0] x426_rdcol_1_io_b; // @[Math.scala 150:24:@23881.4]
  wire  x426_rdcol_1_io_flow; // @[Math.scala 150:24:@23881.4]
  wire [31:0] x426_rdcol_1_io_result; // @[Math.scala 150:24:@23881.4]
  wire  x432_sum_1_clock; // @[Math.scala 150:24:@23913.4]
  wire  x432_sum_1_reset; // @[Math.scala 150:24:@23913.4]
  wire [31:0] x432_sum_1_io_a; // @[Math.scala 150:24:@23913.4]
  wire [31:0] x432_sum_1_io_b; // @[Math.scala 150:24:@23913.4]
  wire  x432_sum_1_io_flow; // @[Math.scala 150:24:@23913.4]
  wire [31:0] x432_sum_1_io_result; // @[Math.scala 150:24:@23913.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@23923.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@23923.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@23923.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@23923.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@23923.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@23937.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@23937.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@23937.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@23937.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@23937.4]
  wire  x438_rdrow_1_clock; // @[Math.scala 191:24:@23960.4]
  wire  x438_rdrow_1_reset; // @[Math.scala 191:24:@23960.4]
  wire [31:0] x438_rdrow_1_io_a; // @[Math.scala 191:24:@23960.4]
  wire [31:0] x438_rdrow_1_io_b; // @[Math.scala 191:24:@23960.4]
  wire  x438_rdrow_1_io_flow; // @[Math.scala 191:24:@23960.4]
  wire [31:0] x438_rdrow_1_io_result; // @[Math.scala 191:24:@23960.4]
  wire  x445_sum_1_clock; // @[Math.scala 150:24:@24014.4]
  wire  x445_sum_1_reset; // @[Math.scala 150:24:@24014.4]
  wire [31:0] x445_sum_1_io_a; // @[Math.scala 150:24:@24014.4]
  wire [31:0] x445_sum_1_io_b; // @[Math.scala 150:24:@24014.4]
  wire  x445_sum_1_io_flow; // @[Math.scala 150:24:@24014.4]
  wire [31:0] x445_sum_1_io_result; // @[Math.scala 150:24:@24014.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@24024.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@24024.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@24024.4]
  wire [31:0] RetimeWrapper_44_io_in; // @[package.scala 93:22:@24024.4]
  wire [31:0] RetimeWrapper_44_io_out; // @[package.scala 93:22:@24024.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@24033.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@24033.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@24033.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@24033.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@24033.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@24047.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@24047.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@24047.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@24047.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@24047.4]
  wire  x453_sum_1_clock; // @[Math.scala 150:24:@24074.4]
  wire  x453_sum_1_reset; // @[Math.scala 150:24:@24074.4]
  wire [31:0] x453_sum_1_io_a; // @[Math.scala 150:24:@24074.4]
  wire [31:0] x453_sum_1_io_b; // @[Math.scala 150:24:@24074.4]
  wire  x453_sum_1_io_flow; // @[Math.scala 150:24:@24074.4]
  wire [31:0] x453_sum_1_io_result; // @[Math.scala 150:24:@24074.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@24084.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@24084.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@24084.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@24084.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@24084.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@24098.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@24098.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@24098.4]
  wire  RetimeWrapper_48_io_in; // @[package.scala 93:22:@24098.4]
  wire  RetimeWrapper_48_io_out; // @[package.scala 93:22:@24098.4]
  wire  x460_sum_1_clock; // @[Math.scala 150:24:@24125.4]
  wire  x460_sum_1_reset; // @[Math.scala 150:24:@24125.4]
  wire [31:0] x460_sum_1_io_a; // @[Math.scala 150:24:@24125.4]
  wire [31:0] x460_sum_1_io_b; // @[Math.scala 150:24:@24125.4]
  wire  x460_sum_1_io_flow; // @[Math.scala 150:24:@24125.4]
  wire [31:0] x460_sum_1_io_result; // @[Math.scala 150:24:@24125.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@24135.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@24135.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@24135.4]
  wire  RetimeWrapper_49_io_in; // @[package.scala 93:22:@24135.4]
  wire  RetimeWrapper_49_io_out; // @[package.scala 93:22:@24135.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@24149.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@24149.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@24149.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@24149.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@24149.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@24170.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@24170.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@24170.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@24170.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@24170.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@24185.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@24185.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@24185.4]
  wire [31:0] RetimeWrapper_52_io_in; // @[package.scala 93:22:@24185.4]
  wire [31:0] RetimeWrapper_52_io_out; // @[package.scala 93:22:@24185.4]
  wire  x467_sum_1_clock; // @[Math.scala 150:24:@24194.4]
  wire  x467_sum_1_reset; // @[Math.scala 150:24:@24194.4]
  wire [31:0] x467_sum_1_io_a; // @[Math.scala 150:24:@24194.4]
  wire [31:0] x467_sum_1_io_b; // @[Math.scala 150:24:@24194.4]
  wire  x467_sum_1_io_flow; // @[Math.scala 150:24:@24194.4]
  wire [31:0] x467_sum_1_io_result; // @[Math.scala 150:24:@24194.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@24204.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@24204.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@24204.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@24204.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@24204.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@24218.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@24218.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@24218.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@24218.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@24218.4]
  wire  x474_sum_1_clock; // @[Math.scala 150:24:@24245.4]
  wire  x474_sum_1_reset; // @[Math.scala 150:24:@24245.4]
  wire [31:0] x474_sum_1_io_a; // @[Math.scala 150:24:@24245.4]
  wire [31:0] x474_sum_1_io_b; // @[Math.scala 150:24:@24245.4]
  wire  x474_sum_1_io_flow; // @[Math.scala 150:24:@24245.4]
  wire [31:0] x474_sum_1_io_result; // @[Math.scala 150:24:@24245.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@24255.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@24255.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@24255.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@24255.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@24255.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@24269.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@24269.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@24269.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@24269.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@24269.4]
  wire  x481_sum_1_clock; // @[Math.scala 150:24:@24298.4]
  wire  x481_sum_1_reset; // @[Math.scala 150:24:@24298.4]
  wire [31:0] x481_sum_1_io_a; // @[Math.scala 150:24:@24298.4]
  wire [31:0] x481_sum_1_io_b; // @[Math.scala 150:24:@24298.4]
  wire  x481_sum_1_io_flow; // @[Math.scala 150:24:@24298.4]
  wire [31:0] x481_sum_1_io_result; // @[Math.scala 150:24:@24298.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@24308.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@24308.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@24308.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@24308.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@24308.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@24322.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@24322.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@24322.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@24322.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@24322.4]
  wire  x486_rdrow_1_clock; // @[Math.scala 191:24:@24345.4]
  wire  x486_rdrow_1_reset; // @[Math.scala 191:24:@24345.4]
  wire [31:0] x486_rdrow_1_io_a; // @[Math.scala 191:24:@24345.4]
  wire [31:0] x486_rdrow_1_io_b; // @[Math.scala 191:24:@24345.4]
  wire  x486_rdrow_1_io_flow; // @[Math.scala 191:24:@24345.4]
  wire [31:0] x486_rdrow_1_io_result; // @[Math.scala 191:24:@24345.4]
  wire  x493_sum_1_clock; // @[Math.scala 150:24:@24399.4]
  wire  x493_sum_1_reset; // @[Math.scala 150:24:@24399.4]
  wire [31:0] x493_sum_1_io_a; // @[Math.scala 150:24:@24399.4]
  wire [31:0] x493_sum_1_io_b; // @[Math.scala 150:24:@24399.4]
  wire  x493_sum_1_io_flow; // @[Math.scala 150:24:@24399.4]
  wire [31:0] x493_sum_1_io_result; // @[Math.scala 150:24:@24399.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@24409.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@24409.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@24409.4]
  wire [31:0] RetimeWrapper_59_io_in; // @[package.scala 93:22:@24409.4]
  wire [31:0] RetimeWrapper_59_io_out; // @[package.scala 93:22:@24409.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@24418.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@24418.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@24418.4]
  wire  RetimeWrapper_60_io_in; // @[package.scala 93:22:@24418.4]
  wire  RetimeWrapper_60_io_out; // @[package.scala 93:22:@24418.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@24432.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@24432.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@24432.4]
  wire  RetimeWrapper_61_io_in; // @[package.scala 93:22:@24432.4]
  wire  RetimeWrapper_61_io_out; // @[package.scala 93:22:@24432.4]
  wire  x501_sum_1_clock; // @[Math.scala 150:24:@24459.4]
  wire  x501_sum_1_reset; // @[Math.scala 150:24:@24459.4]
  wire [31:0] x501_sum_1_io_a; // @[Math.scala 150:24:@24459.4]
  wire [31:0] x501_sum_1_io_b; // @[Math.scala 150:24:@24459.4]
  wire  x501_sum_1_io_flow; // @[Math.scala 150:24:@24459.4]
  wire [31:0] x501_sum_1_io_result; // @[Math.scala 150:24:@24459.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@24469.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@24469.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@24469.4]
  wire  RetimeWrapper_62_io_in; // @[package.scala 93:22:@24469.4]
  wire  RetimeWrapper_62_io_out; // @[package.scala 93:22:@24469.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@24483.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@24483.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@24483.4]
  wire  RetimeWrapper_63_io_in; // @[package.scala 93:22:@24483.4]
  wire  RetimeWrapper_63_io_out; // @[package.scala 93:22:@24483.4]
  wire  x508_sum_1_clock; // @[Math.scala 150:24:@24510.4]
  wire  x508_sum_1_reset; // @[Math.scala 150:24:@24510.4]
  wire [31:0] x508_sum_1_io_a; // @[Math.scala 150:24:@24510.4]
  wire [31:0] x508_sum_1_io_b; // @[Math.scala 150:24:@24510.4]
  wire  x508_sum_1_io_flow; // @[Math.scala 150:24:@24510.4]
  wire [31:0] x508_sum_1_io_result; // @[Math.scala 150:24:@24510.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@24520.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@24520.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@24520.4]
  wire  RetimeWrapper_64_io_in; // @[package.scala 93:22:@24520.4]
  wire  RetimeWrapper_64_io_out; // @[package.scala 93:22:@24520.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@24534.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@24534.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@24534.4]
  wire  RetimeWrapper_65_io_in; // @[package.scala 93:22:@24534.4]
  wire  RetimeWrapper_65_io_out; // @[package.scala 93:22:@24534.4]
  wire  x515_sum_1_clock; // @[Math.scala 150:24:@24561.4]
  wire  x515_sum_1_reset; // @[Math.scala 150:24:@24561.4]
  wire [31:0] x515_sum_1_io_a; // @[Math.scala 150:24:@24561.4]
  wire [31:0] x515_sum_1_io_b; // @[Math.scala 150:24:@24561.4]
  wire  x515_sum_1_io_flow; // @[Math.scala 150:24:@24561.4]
  wire [31:0] x515_sum_1_io_result; // @[Math.scala 150:24:@24561.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@24571.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@24571.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@24571.4]
  wire  RetimeWrapper_66_io_in; // @[package.scala 93:22:@24571.4]
  wire  RetimeWrapper_66_io_out; // @[package.scala 93:22:@24571.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@24585.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@24585.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@24585.4]
  wire  RetimeWrapper_67_io_in; // @[package.scala 93:22:@24585.4]
  wire  RetimeWrapper_67_io_out; // @[package.scala 93:22:@24585.4]
  wire  x522_sum_1_clock; // @[Math.scala 150:24:@24612.4]
  wire  x522_sum_1_reset; // @[Math.scala 150:24:@24612.4]
  wire [31:0] x522_sum_1_io_a; // @[Math.scala 150:24:@24612.4]
  wire [31:0] x522_sum_1_io_b; // @[Math.scala 150:24:@24612.4]
  wire  x522_sum_1_io_flow; // @[Math.scala 150:24:@24612.4]
  wire [31:0] x522_sum_1_io_result; // @[Math.scala 150:24:@24612.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@24622.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@24622.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@24622.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@24622.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@24622.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@24636.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@24636.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@24636.4]
  wire  RetimeWrapper_69_io_in; // @[package.scala 93:22:@24636.4]
  wire  RetimeWrapper_69_io_out; // @[package.scala 93:22:@24636.4]
  wire  x529_sum_1_clock; // @[Math.scala 150:24:@24663.4]
  wire  x529_sum_1_reset; // @[Math.scala 150:24:@24663.4]
  wire [31:0] x529_sum_1_io_a; // @[Math.scala 150:24:@24663.4]
  wire [31:0] x529_sum_1_io_b; // @[Math.scala 150:24:@24663.4]
  wire  x529_sum_1_io_flow; // @[Math.scala 150:24:@24663.4]
  wire [31:0] x529_sum_1_io_result; // @[Math.scala 150:24:@24663.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@24673.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@24673.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@24673.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@24673.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@24673.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@24687.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@24687.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@24687.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@24687.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@24687.4]
  wire  x539_x11_1_clock; // @[Math.scala 150:24:@24735.4]
  wire  x539_x11_1_reset; // @[Math.scala 150:24:@24735.4]
  wire [7:0] x539_x11_1_io_a; // @[Math.scala 150:24:@24735.4]
  wire [7:0] x539_x11_1_io_b; // @[Math.scala 150:24:@24735.4]
  wire  x539_x11_1_io_flow; // @[Math.scala 150:24:@24735.4]
  wire [7:0] x539_x11_1_io_result; // @[Math.scala 150:24:@24735.4]
  wire  x540_x12_1_clock; // @[Math.scala 150:24:@24745.4]
  wire  x540_x12_1_reset; // @[Math.scala 150:24:@24745.4]
  wire [7:0] x540_x12_1_io_a; // @[Math.scala 150:24:@24745.4]
  wire [7:0] x540_x12_1_io_b; // @[Math.scala 150:24:@24745.4]
  wire  x540_x12_1_io_flow; // @[Math.scala 150:24:@24745.4]
  wire [7:0] x540_x12_1_io_result; // @[Math.scala 150:24:@24745.4]
  wire  x541_x11_1_clock; // @[Math.scala 150:24:@24755.4]
  wire  x541_x11_1_reset; // @[Math.scala 150:24:@24755.4]
  wire [7:0] x541_x11_1_io_a; // @[Math.scala 150:24:@24755.4]
  wire [7:0] x541_x11_1_io_b; // @[Math.scala 150:24:@24755.4]
  wire  x541_x11_1_io_flow; // @[Math.scala 150:24:@24755.4]
  wire [7:0] x541_x11_1_io_result; // @[Math.scala 150:24:@24755.4]
  wire  x542_x12_1_clock; // @[Math.scala 150:24:@24765.4]
  wire  x542_x12_1_reset; // @[Math.scala 150:24:@24765.4]
  wire [7:0] x542_x12_1_io_a; // @[Math.scala 150:24:@24765.4]
  wire [7:0] x542_x12_1_io_b; // @[Math.scala 150:24:@24765.4]
  wire  x542_x12_1_io_flow; // @[Math.scala 150:24:@24765.4]
  wire [7:0] x542_x12_1_io_result; // @[Math.scala 150:24:@24765.4]
  wire [7:0] x543_x11_1_io_a; // @[Math.scala 150:24:@24775.4]
  wire [7:0] x543_x11_1_io_b; // @[Math.scala 150:24:@24775.4]
  wire [7:0] x543_x11_1_io_result; // @[Math.scala 150:24:@24775.4]
  wire [7:0] x544_x12_1_io_a; // @[Math.scala 150:24:@24785.4]
  wire [7:0] x544_x12_1_io_b; // @[Math.scala 150:24:@24785.4]
  wire [7:0] x544_x12_1_io_result; // @[Math.scala 150:24:@24785.4]
  wire [7:0] x545_x11_1_io_a; // @[Math.scala 150:24:@24795.4]
  wire [7:0] x545_x11_1_io_b; // @[Math.scala 150:24:@24795.4]
  wire [7:0] x545_x11_1_io_result; // @[Math.scala 150:24:@24795.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@24805.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@24805.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@24805.4]
  wire [7:0] RetimeWrapper_72_io_in; // @[package.scala 93:22:@24805.4]
  wire [7:0] RetimeWrapper_72_io_out; // @[package.scala 93:22:@24805.4]
  wire [7:0] x546_sum_1_io_a; // @[Math.scala 150:24:@24814.4]
  wire [7:0] x546_sum_1_io_b; // @[Math.scala 150:24:@24814.4]
  wire [7:0] x546_sum_1_io_result; // @[Math.scala 150:24:@24814.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@24828.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@24828.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@24828.4]
  wire [7:0] RetimeWrapper_73_io_in; // @[package.scala 93:22:@24828.4]
  wire [7:0] RetimeWrapper_73_io_out; // @[package.scala 93:22:@24828.4]
  wire  x553_x11_1_clock; // @[Math.scala 150:24:@24863.4]
  wire  x553_x11_1_reset; // @[Math.scala 150:24:@24863.4]
  wire [7:0] x553_x11_1_io_a; // @[Math.scala 150:24:@24863.4]
  wire [7:0] x553_x11_1_io_b; // @[Math.scala 150:24:@24863.4]
  wire  x553_x11_1_io_flow; // @[Math.scala 150:24:@24863.4]
  wire [7:0] x553_x11_1_io_result; // @[Math.scala 150:24:@24863.4]
  wire  x554_x12_1_clock; // @[Math.scala 150:24:@24873.4]
  wire  x554_x12_1_reset; // @[Math.scala 150:24:@24873.4]
  wire [7:0] x554_x12_1_io_a; // @[Math.scala 150:24:@24873.4]
  wire [7:0] x554_x12_1_io_b; // @[Math.scala 150:24:@24873.4]
  wire  x554_x12_1_io_flow; // @[Math.scala 150:24:@24873.4]
  wire [7:0] x554_x12_1_io_result; // @[Math.scala 150:24:@24873.4]
  wire  x555_x11_1_clock; // @[Math.scala 150:24:@24883.4]
  wire  x555_x11_1_reset; // @[Math.scala 150:24:@24883.4]
  wire [7:0] x555_x11_1_io_a; // @[Math.scala 150:24:@24883.4]
  wire [7:0] x555_x11_1_io_b; // @[Math.scala 150:24:@24883.4]
  wire  x555_x11_1_io_flow; // @[Math.scala 150:24:@24883.4]
  wire [7:0] x555_x11_1_io_result; // @[Math.scala 150:24:@24883.4]
  wire  x556_x12_1_clock; // @[Math.scala 150:24:@24893.4]
  wire  x556_x12_1_reset; // @[Math.scala 150:24:@24893.4]
  wire [7:0] x556_x12_1_io_a; // @[Math.scala 150:24:@24893.4]
  wire [7:0] x556_x12_1_io_b; // @[Math.scala 150:24:@24893.4]
  wire  x556_x12_1_io_flow; // @[Math.scala 150:24:@24893.4]
  wire [7:0] x556_x12_1_io_result; // @[Math.scala 150:24:@24893.4]
  wire [7:0] x557_x11_1_io_a; // @[Math.scala 150:24:@24903.4]
  wire [7:0] x557_x11_1_io_b; // @[Math.scala 150:24:@24903.4]
  wire [7:0] x557_x11_1_io_result; // @[Math.scala 150:24:@24903.4]
  wire [7:0] x558_x12_1_io_a; // @[Math.scala 150:24:@24913.4]
  wire [7:0] x558_x12_1_io_b; // @[Math.scala 150:24:@24913.4]
  wire [7:0] x558_x12_1_io_result; // @[Math.scala 150:24:@24913.4]
  wire [7:0] x559_x11_1_io_a; // @[Math.scala 150:24:@24923.4]
  wire [7:0] x559_x11_1_io_b; // @[Math.scala 150:24:@24923.4]
  wire [7:0] x559_x11_1_io_result; // @[Math.scala 150:24:@24923.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@24933.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@24933.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@24933.4]
  wire [7:0] RetimeWrapper_74_io_in; // @[package.scala 93:22:@24933.4]
  wire [7:0] RetimeWrapper_74_io_out; // @[package.scala 93:22:@24933.4]
  wire [7:0] x560_sum_1_io_a; // @[Math.scala 150:24:@24942.4]
  wire [7:0] x560_sum_1_io_b; // @[Math.scala 150:24:@24942.4]
  wire [7:0] x560_sum_1_io_result; // @[Math.scala 150:24:@24942.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@24956.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@24956.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@24956.4]
  wire [7:0] RetimeWrapper_75_io_in; // @[package.scala 93:22:@24956.4]
  wire [7:0] RetimeWrapper_75_io_out; // @[package.scala 93:22:@24956.4]
  wire  x566_x11_1_clock; // @[Math.scala 150:24:@24986.4]
  wire  x566_x11_1_reset; // @[Math.scala 150:24:@24986.4]
  wire [7:0] x566_x11_1_io_a; // @[Math.scala 150:24:@24986.4]
  wire [7:0] x566_x11_1_io_b; // @[Math.scala 150:24:@24986.4]
  wire  x566_x11_1_io_flow; // @[Math.scala 150:24:@24986.4]
  wire [7:0] x566_x11_1_io_result; // @[Math.scala 150:24:@24986.4]
  wire  x567_x12_1_clock; // @[Math.scala 150:24:@24996.4]
  wire  x567_x12_1_reset; // @[Math.scala 150:24:@24996.4]
  wire [7:0] x567_x12_1_io_a; // @[Math.scala 150:24:@24996.4]
  wire [7:0] x567_x12_1_io_b; // @[Math.scala 150:24:@24996.4]
  wire  x567_x12_1_io_flow; // @[Math.scala 150:24:@24996.4]
  wire [7:0] x567_x12_1_io_result; // @[Math.scala 150:24:@24996.4]
  wire  x568_x11_1_clock; // @[Math.scala 150:24:@25006.4]
  wire  x568_x11_1_reset; // @[Math.scala 150:24:@25006.4]
  wire [7:0] x568_x11_1_io_a; // @[Math.scala 150:24:@25006.4]
  wire [7:0] x568_x11_1_io_b; // @[Math.scala 150:24:@25006.4]
  wire  x568_x11_1_io_flow; // @[Math.scala 150:24:@25006.4]
  wire [7:0] x568_x11_1_io_result; // @[Math.scala 150:24:@25006.4]
  wire  x569_x12_1_clock; // @[Math.scala 150:24:@25016.4]
  wire  x569_x12_1_reset; // @[Math.scala 150:24:@25016.4]
  wire [7:0] x569_x12_1_io_a; // @[Math.scala 150:24:@25016.4]
  wire [7:0] x569_x12_1_io_b; // @[Math.scala 150:24:@25016.4]
  wire  x569_x12_1_io_flow; // @[Math.scala 150:24:@25016.4]
  wire [7:0] x569_x12_1_io_result; // @[Math.scala 150:24:@25016.4]
  wire [7:0] x570_x11_1_io_a; // @[Math.scala 150:24:@25026.4]
  wire [7:0] x570_x11_1_io_b; // @[Math.scala 150:24:@25026.4]
  wire [7:0] x570_x11_1_io_result; // @[Math.scala 150:24:@25026.4]
  wire [7:0] x571_x12_1_io_a; // @[Math.scala 150:24:@25036.4]
  wire [7:0] x571_x12_1_io_b; // @[Math.scala 150:24:@25036.4]
  wire [7:0] x571_x12_1_io_result; // @[Math.scala 150:24:@25036.4]
  wire [7:0] x572_x11_1_io_a; // @[Math.scala 150:24:@25046.4]
  wire [7:0] x572_x11_1_io_b; // @[Math.scala 150:24:@25046.4]
  wire [7:0] x572_x11_1_io_result; // @[Math.scala 150:24:@25046.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@25056.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@25056.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@25056.4]
  wire [7:0] RetimeWrapper_76_io_in; // @[package.scala 93:22:@25056.4]
  wire [7:0] RetimeWrapper_76_io_out; // @[package.scala 93:22:@25056.4]
  wire [7:0] x573_sum_1_io_a; // @[Math.scala 150:24:@25065.4]
  wire [7:0] x573_sum_1_io_b; // @[Math.scala 150:24:@25065.4]
  wire [7:0] x573_sum_1_io_result; // @[Math.scala 150:24:@25065.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@25079.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@25079.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@25079.4]
  wire [7:0] RetimeWrapper_77_io_in; // @[package.scala 93:22:@25079.4]
  wire [7:0] RetimeWrapper_77_io_out; // @[package.scala 93:22:@25079.4]
  wire  x579_x11_1_clock; // @[Math.scala 150:24:@25109.4]
  wire  x579_x11_1_reset; // @[Math.scala 150:24:@25109.4]
  wire [7:0] x579_x11_1_io_a; // @[Math.scala 150:24:@25109.4]
  wire [7:0] x579_x11_1_io_b; // @[Math.scala 150:24:@25109.4]
  wire  x579_x11_1_io_flow; // @[Math.scala 150:24:@25109.4]
  wire [7:0] x579_x11_1_io_result; // @[Math.scala 150:24:@25109.4]
  wire  x580_x12_1_clock; // @[Math.scala 150:24:@25119.4]
  wire  x580_x12_1_reset; // @[Math.scala 150:24:@25119.4]
  wire [7:0] x580_x12_1_io_a; // @[Math.scala 150:24:@25119.4]
  wire [7:0] x580_x12_1_io_b; // @[Math.scala 150:24:@25119.4]
  wire  x580_x12_1_io_flow; // @[Math.scala 150:24:@25119.4]
  wire [7:0] x580_x12_1_io_result; // @[Math.scala 150:24:@25119.4]
  wire  x581_x11_1_clock; // @[Math.scala 150:24:@25131.4]
  wire  x581_x11_1_reset; // @[Math.scala 150:24:@25131.4]
  wire [7:0] x581_x11_1_io_a; // @[Math.scala 150:24:@25131.4]
  wire [7:0] x581_x11_1_io_b; // @[Math.scala 150:24:@25131.4]
  wire  x581_x11_1_io_flow; // @[Math.scala 150:24:@25131.4]
  wire [7:0] x581_x11_1_io_result; // @[Math.scala 150:24:@25131.4]
  wire  x582_x12_1_clock; // @[Math.scala 150:24:@25141.4]
  wire  x582_x12_1_reset; // @[Math.scala 150:24:@25141.4]
  wire [7:0] x582_x12_1_io_a; // @[Math.scala 150:24:@25141.4]
  wire [7:0] x582_x12_1_io_b; // @[Math.scala 150:24:@25141.4]
  wire  x582_x12_1_io_flow; // @[Math.scala 150:24:@25141.4]
  wire [7:0] x582_x12_1_io_result; // @[Math.scala 150:24:@25141.4]
  wire [7:0] x583_x11_1_io_a; // @[Math.scala 150:24:@25151.4]
  wire [7:0] x583_x11_1_io_b; // @[Math.scala 150:24:@25151.4]
  wire [7:0] x583_x11_1_io_result; // @[Math.scala 150:24:@25151.4]
  wire [7:0] x584_x12_1_io_a; // @[Math.scala 150:24:@25161.4]
  wire [7:0] x584_x12_1_io_b; // @[Math.scala 150:24:@25161.4]
  wire [7:0] x584_x12_1_io_result; // @[Math.scala 150:24:@25161.4]
  wire [7:0] x585_x11_1_io_a; // @[Math.scala 150:24:@25171.4]
  wire [7:0] x585_x11_1_io_b; // @[Math.scala 150:24:@25171.4]
  wire [7:0] x585_x11_1_io_result; // @[Math.scala 150:24:@25171.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@25181.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@25181.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@25181.4]
  wire [7:0] RetimeWrapper_78_io_in; // @[package.scala 93:22:@25181.4]
  wire [7:0] RetimeWrapper_78_io_out; // @[package.scala 93:22:@25181.4]
  wire [7:0] x586_sum_1_io_a; // @[Math.scala 150:24:@25190.4]
  wire [7:0] x586_sum_1_io_b; // @[Math.scala 150:24:@25190.4]
  wire [7:0] x586_sum_1_io_result; // @[Math.scala 150:24:@25190.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@25204.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@25204.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@25204.4]
  wire [7:0] RetimeWrapper_79_io_in; // @[package.scala 93:22:@25204.4]
  wire [7:0] RetimeWrapper_79_io_out; // @[package.scala 93:22:@25204.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@25224.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@25224.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@25224.4]
  wire [31:0] RetimeWrapper_80_io_in; // @[package.scala 93:22:@25224.4]
  wire [31:0] RetimeWrapper_80_io_out; // @[package.scala 93:22:@25224.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@25233.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@25233.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@25233.4]
  wire  RetimeWrapper_81_io_in; // @[package.scala 93:22:@25233.4]
  wire  RetimeWrapper_81_io_out; // @[package.scala 93:22:@25233.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@25242.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@25242.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@25242.4]
  wire  RetimeWrapper_82_io_in; // @[package.scala 93:22:@25242.4]
  wire  RetimeWrapper_82_io_out; // @[package.scala 93:22:@25242.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@25251.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@25251.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@25251.4]
  wire  RetimeWrapper_83_io_in; // @[package.scala 93:22:@25251.4]
  wire  RetimeWrapper_83_io_out; // @[package.scala 93:22:@25251.4]
  wire  b327; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 62:18:@22814.4]
  wire  b328; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 63:18:@22815.4]
  wire  _T_206; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 68:30:@22962.4]
  wire  _T_207; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 68:37:@22963.4]
  wire  _T_211; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 70:76:@22968.4]
  wire  _T_212; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 70:62:@22969.4]
  wire  _T_214; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 70:101:@22970.4]
  wire [31:0] x667_x330_D1_0_number; // @[package.scala 96:25:@22979.4 package.scala 96:25:@22980.4]
  wire [31:0] b325_number; // @[Math.scala 712:22:@22799.4 Math.scala 713:14:@22800.4]
  wire [31:0] _T_246; // @[Math.scala 499:52:@22999.4]
  wire  x334; // @[Math.scala 499:44:@23007.4]
  wire  x335; // @[Math.scala 499:44:@23014.4]
  wire  x336; // @[Math.scala 499:44:@23021.4]
  wire [31:0] _T_293; // @[Mux.scala 19:72:@23033.4]
  wire [31:0] _T_295; // @[Mux.scala 19:72:@23034.4]
  wire [31:0] _T_297; // @[Mux.scala 19:72:@23035.4]
  wire [31:0] _T_299; // @[Mux.scala 19:72:@23037.4]
  wire [31:0] x337_number; // @[Mux.scala 19:72:@23038.4]
  wire [31:0] _T_311; // @[Math.scala 406:49:@23048.4]
  wire [31:0] _T_313; // @[Math.scala 406:56:@23050.4]
  wire [31:0] _T_314; // @[Math.scala 406:56:@23051.4]
  wire  _T_319; // @[FixedPoint.scala 50:25:@23057.4]
  wire [1:0] _T_323; // @[Bitwise.scala 72:12:@23059.4]
  wire [29:0] _T_324; // @[FixedPoint.scala 18:52:@23060.4]
  wire [31:0] b326_number; // @[Math.scala 712:22:@22811.4 Math.scala 713:14:@22812.4]
  wire  _T_329; // @[FixedPoint.scala 50:25:@23066.4]
  wire [1:0] _T_333; // @[Bitwise.scala 72:12:@23068.4]
  wire [29:0] _T_334; // @[FixedPoint.scala 18:52:@23069.4]
  wire  _T_359; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 113:101:@23130.4]
  wire  _T_363; // @[package.scala 96:25:@23138.4 package.scala 96:25:@23139.4]
  wire  _T_365; // @[implicits.scala 55:10:@23140.4]
  wire  _T_366; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 113:118:@23141.4]
  wire  _T_368; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 113:205:@23143.4]
  wire  _T_369; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 113:224:@23144.4]
  wire  x671_b327_D4; // @[package.scala 96:25:@23116.4 package.scala 96:25:@23117.4]
  wire  _T_370; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 113:250:@23145.4]
  wire  x669_b328_D4; // @[package.scala 96:25:@23098.4 package.scala 96:25:@23099.4]
  wire [31:0] x349_rdcol_number; // @[Math.scala 154:22:@23162.4 Math.scala 155:14:@23163.4]
  wire  _T_383; // @[FixedPoint.scala 50:25:@23169.4]
  wire [1:0] _T_387; // @[Bitwise.scala 72:12:@23171.4]
  wire [29:0] _T_388; // @[FixedPoint.scala 18:52:@23172.4]
  wire  _T_411; // @[package.scala 96:25:@23223.4 package.scala 96:25:@23224.4]
  wire  _T_413; // @[implicits.scala 55:10:@23225.4]
  wire  _T_414; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 132:118:@23226.4]
  wire  _T_416; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 132:205:@23228.4]
  wire  _T_417; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 132:224:@23229.4]
  wire  _T_418; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 132:250:@23230.4]
  wire [31:0] x358_rdcol_number; // @[Math.scala 154:22:@23247.4 Math.scala 155:14:@23248.4]
  wire  _T_431; // @[FixedPoint.scala 50:25:@23254.4]
  wire [1:0] _T_435; // @[Bitwise.scala 72:12:@23256.4]
  wire [29:0] _T_436; // @[FixedPoint.scala 18:52:@23257.4]
  wire  _T_456; // @[package.scala 96:25:@23299.4 package.scala 96:25:@23300.4]
  wire  _T_458; // @[implicits.scala 55:10:@23301.4]
  wire  _T_459; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 149:118:@23302.4]
  wire  _T_461; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 149:205:@23304.4]
  wire  _T_462; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 149:224:@23305.4]
  wire  _T_463; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 149:250:@23306.4]
  wire [31:0] x367_rdcol_number; // @[Math.scala 154:22:@23323.4 Math.scala 155:14:@23324.4]
  wire  _T_476; // @[FixedPoint.scala 50:25:@23330.4]
  wire [1:0] _T_480; // @[Bitwise.scala 72:12:@23332.4]
  wire [29:0] _T_481; // @[FixedPoint.scala 18:52:@23333.4]
  wire  _T_501; // @[package.scala 96:25:@23375.4 package.scala 96:25:@23376.4]
  wire  _T_503; // @[implicits.scala 55:10:@23377.4]
  wire  _T_504; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 166:118:@23378.4]
  wire  _T_506; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 166:205:@23380.4]
  wire  _T_507; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 166:224:@23381.4]
  wire  _T_508; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 166:250:@23382.4]
  wire [31:0] x680_b325_D6_number; // @[package.scala 96:25:@23396.4 package.scala 96:25:@23397.4]
  wire [31:0] _T_520; // @[Math.scala 406:49:@23403.4]
  wire [31:0] _T_522; // @[Math.scala 406:56:@23405.4]
  wire [31:0] _T_523; // @[Math.scala 406:56:@23406.4]
  wire [31:0] x661_number; // @[implicits.scala 133:21:@23407.4]
  wire  x378; // @[Math.scala 465:44:@23415.4]
  wire [31:0] x681_x367_rdcol_D6_number; // @[package.scala 96:25:@23423.4 package.scala 96:25:@23424.4]
  wire [31:0] _T_541; // @[Math.scala 465:37:@23429.4]
  wire  x379; // @[Math.scala 465:44:@23431.4]
  wire  x682_x378_D1; // @[package.scala 96:25:@23439.4 package.scala 96:25:@23440.4]
  wire  x380; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 187:24:@23443.4]
  wire [31:0] _T_560; // @[Math.scala 406:49:@23454.4]
  wire [31:0] _T_562; // @[Math.scala 406:56:@23456.4]
  wire [31:0] _T_563; // @[Math.scala 406:56:@23457.4]
  wire  _T_568; // @[FixedPoint.scala 50:25:@23463.4]
  wire [1:0] _T_572; // @[Bitwise.scala 72:12:@23465.4]
  wire [29:0] _T_573; // @[FixedPoint.scala 18:52:@23466.4]
  wire  _T_611; // @[package.scala 96:25:@23545.4 package.scala 96:25:@23546.4]
  wire  _T_613; // @[implicits.scala 55:10:@23547.4]
  wire  _T_614; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 214:194:@23548.4]
  wire  x685_x381_D1; // @[package.scala 96:25:@23504.4 package.scala 96:25:@23505.4]
  wire  _T_615; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 214:281:@23549.4]
  wire  x688_b327_D8; // @[package.scala 96:25:@23531.4 package.scala 96:25:@23532.4]
  wire  _T_616; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 214:289:@23550.4]
  wire  x686_b328_D8; // @[package.scala 96:25:@23513.4 package.scala 96:25:@23514.4]
  wire [31:0] x689_x358_rdcol_D6_number; // @[package.scala 96:25:@23566.4 package.scala 96:25:@23567.4]
  wire [31:0] _T_627; // @[Math.scala 465:37:@23572.4]
  wire  x390; // @[Math.scala 465:44:@23574.4]
  wire  x391; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 222:24:@23577.4]
  wire  _T_658; // @[package.scala 96:25:@23621.4 package.scala 96:25:@23622.4]
  wire  _T_660; // @[implicits.scala 55:10:@23623.4]
  wire  _T_661; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 235:194:@23624.4]
  wire  x691_x392_D1; // @[package.scala 96:25:@23607.4 package.scala 96:25:@23608.4]
  wire  _T_662; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 235:281:@23625.4]
  wire  _T_663; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 235:289:@23626.4]
  wire [31:0] x692_x349_rdcol_D6_number; // @[package.scala 96:25:@23642.4 package.scala 96:25:@23643.4]
  wire [31:0] _T_674; // @[Math.scala 465:37:@23648.4]
  wire  x398; // @[Math.scala 465:44:@23650.4]
  wire  x399; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 243:24:@23653.4]
  wire  _T_705; // @[package.scala 96:25:@23697.4 package.scala 96:25:@23698.4]
  wire  _T_707; // @[implicits.scala 55:10:@23699.4]
  wire  _T_708; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 256:194:@23700.4]
  wire  x694_x400_D1; // @[package.scala 96:25:@23683.4 package.scala 96:25:@23684.4]
  wire  _T_709; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 256:281:@23701.4]
  wire  _T_710; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 256:289:@23702.4]
  wire [31:0] x695_b326_D6_number; // @[package.scala 96:25:@23718.4 package.scala 96:25:@23719.4]
  wire [31:0] _T_721; // @[Math.scala 465:37:@23724.4]
  wire  x406; // @[Math.scala 465:44:@23726.4]
  wire  x407; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 264:59:@23729.4]
  wire  _T_755; // @[package.scala 96:25:@23782.4 package.scala 96:25:@23783.4]
  wire  _T_757; // @[implicits.scala 55:10:@23784.4]
  wire  _T_758; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 279:194:@23785.4]
  wire  x697_x408_D2; // @[package.scala 96:25:@23759.4 package.scala 96:25:@23760.4]
  wire  _T_759; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 279:281:@23786.4]
  wire  _T_760; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 279:289:@23787.4]
  wire [31:0] x414_rdcol_number; // @[Math.scala 154:22:@23806.4 Math.scala 155:14:@23807.4]
  wire [31:0] _T_775; // @[Math.scala 465:37:@23812.4]
  wire  x415; // @[Math.scala 465:44:@23814.4]
  wire  x416; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 287:24:@23817.4]
  wire  _T_785; // @[FixedPoint.scala 50:25:@23824.4]
  wire [1:0] _T_789; // @[Bitwise.scala 72:12:@23826.4]
  wire [29:0] _T_790; // @[FixedPoint.scala 18:52:@23827.4]
  wire  _T_813; // @[package.scala 96:25:@23861.4 package.scala 96:25:@23862.4]
  wire  _T_815; // @[implicits.scala 55:10:@23863.4]
  wire  _T_816; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 306:194:@23864.4]
  wire  x699_x417_D1; // @[package.scala 96:25:@23847.4 package.scala 96:25:@23848.4]
  wire  _T_817; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 306:281:@23865.4]
  wire  _T_818; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 306:324:@23866.4]
  wire [31:0] x426_rdcol_number; // @[Math.scala 154:22:@23887.4 Math.scala 155:14:@23888.4]
  wire [31:0] _T_835; // @[Math.scala 465:37:@23893.4]
  wire  x427; // @[Math.scala 465:44:@23895.4]
  wire  x428; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 316:59:@23898.4]
  wire  _T_845; // @[FixedPoint.scala 50:25:@23905.4]
  wire [1:0] _T_849; // @[Bitwise.scala 72:12:@23907.4]
  wire [29:0] _T_850; // @[FixedPoint.scala 18:52:@23908.4]
  wire  _T_873; // @[package.scala 96:25:@23942.4 package.scala 96:25:@23943.4]
  wire  _T_875; // @[implicits.scala 55:10:@23944.4]
  wire  _T_876; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 329:194:@23945.4]
  wire  x700_x429_D1; // @[package.scala 96:25:@23928.4 package.scala 96:25:@23929.4]
  wire  _T_877; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 329:281:@23946.4]
  wire  _T_878; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 329:289:@23947.4]
  wire [31:0] x438_rdrow_number; // @[Math.scala 195:22:@23966.4 Math.scala 196:14:@23967.4]
  wire [31:0] _T_895; // @[Math.scala 406:49:@23973.4]
  wire [31:0] _T_897; // @[Math.scala 406:56:@23975.4]
  wire [31:0] _T_898; // @[Math.scala 406:56:@23976.4]
  wire [31:0] x663_number; // @[implicits.scala 133:21:@23977.4]
  wire  x440; // @[Math.scala 465:44:@23985.4]
  wire  x441; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 339:24:@23988.4]
  wire [31:0] _T_919; // @[Math.scala 406:49:@23997.4]
  wire [31:0] _T_921; // @[Math.scala 406:56:@23999.4]
  wire [31:0] _T_922; // @[Math.scala 406:56:@24000.4]
  wire  _T_927; // @[FixedPoint.scala 50:25:@24006.4]
  wire [1:0] _T_931; // @[Bitwise.scala 72:12:@24008.4]
  wire [29:0] _T_932; // @[FixedPoint.scala 18:52:@24009.4]
  wire  _T_958; // @[package.scala 96:25:@24052.4 package.scala 96:25:@24053.4]
  wire  _T_960; // @[implicits.scala 55:10:@24054.4]
  wire  _T_961; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 356:194:@24055.4]
  wire  x702_x442_D1; // @[package.scala 96:25:@24038.4 package.scala 96:25:@24039.4]
  wire  _T_962; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 356:281:@24056.4]
  wire  _T_963; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 356:289:@24057.4]
  wire  x451; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 360:24:@24068.4]
  wire  _T_991; // @[package.scala 96:25:@24103.4 package.scala 96:25:@24104.4]
  wire  _T_993; // @[implicits.scala 55:10:@24105.4]
  wire  _T_994; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 371:194:@24106.4]
  wire  x703_x452_D1; // @[package.scala 96:25:@24089.4 package.scala 96:25:@24090.4]
  wire  _T_995; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 371:281:@24107.4]
  wire  _T_996; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 371:289:@24108.4]
  wire  x458; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 375:24:@24119.4]
  wire  _T_1024; // @[package.scala 96:25:@24154.4 package.scala 96:25:@24155.4]
  wire  _T_1026; // @[implicits.scala 55:10:@24156.4]
  wire  _T_1027; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 386:194:@24157.4]
  wire  x704_x459_D1; // @[package.scala 96:25:@24140.4 package.scala 96:25:@24141.4]
  wire  _T_1028; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 386:281:@24158.4]
  wire  _T_1029; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 386:289:@24159.4]
  wire  x705_x406_D1; // @[package.scala 96:25:@24175.4 package.scala 96:25:@24176.4]
  wire  x465; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 392:24:@24179.4]
  wire  _T_1063; // @[package.scala 96:25:@24223.4 package.scala 96:25:@24224.4]
  wire  _T_1065; // @[implicits.scala 55:10:@24225.4]
  wire  _T_1066; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 405:194:@24226.4]
  wire  x707_x466_D1; // @[package.scala 96:25:@24209.4 package.scala 96:25:@24210.4]
  wire  _T_1067; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 405:281:@24227.4]
  wire  _T_1068; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 405:289:@24228.4]
  wire  x472; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 409:24:@24239.4]
  wire  _T_1096; // @[package.scala 96:25:@24274.4 package.scala 96:25:@24275.4]
  wire  _T_1098; // @[implicits.scala 55:10:@24276.4]
  wire  _T_1099; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 420:194:@24277.4]
  wire  x708_x473_D1; // @[package.scala 96:25:@24260.4 package.scala 96:25:@24261.4]
  wire  _T_1100; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 420:281:@24278.4]
  wire  _T_1101; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 420:289:@24279.4]
  wire  x479; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 430:59:@24290.4]
  wire  _T_1131; // @[package.scala 96:25:@24327.4 package.scala 96:25:@24328.4]
  wire  _T_1133; // @[implicits.scala 55:10:@24329.4]
  wire  _T_1134; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 443:194:@24330.4]
  wire  x709_x480_D1; // @[package.scala 96:25:@24313.4 package.scala 96:25:@24314.4]
  wire  _T_1135; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 443:281:@24331.4]
  wire  _T_1136; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 443:289:@24332.4]
  wire [31:0] x486_rdrow_number; // @[Math.scala 195:22:@24351.4 Math.scala 196:14:@24352.4]
  wire [31:0] _T_1153; // @[Math.scala 406:49:@24358.4]
  wire [31:0] _T_1155; // @[Math.scala 406:56:@24360.4]
  wire [31:0] _T_1156; // @[Math.scala 406:56:@24361.4]
  wire [31:0] x665_number; // @[implicits.scala 133:21:@24362.4]
  wire  x488; // @[Math.scala 465:44:@24370.4]
  wire  x489; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 453:24:@24373.4]
  wire [31:0] _T_1177; // @[Math.scala 406:49:@24382.4]
  wire [31:0] _T_1179; // @[Math.scala 406:56:@24384.4]
  wire [31:0] _T_1180; // @[Math.scala 406:56:@24385.4]
  wire  _T_1185; // @[FixedPoint.scala 50:25:@24391.4]
  wire [1:0] _T_1189; // @[Bitwise.scala 72:12:@24393.4]
  wire [29:0] _T_1190; // @[FixedPoint.scala 18:52:@24394.4]
  wire  _T_1216; // @[package.scala 96:25:@24437.4 package.scala 96:25:@24438.4]
  wire  _T_1218; // @[implicits.scala 55:10:@24439.4]
  wire  _T_1219; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 470:194:@24440.4]
  wire  x711_x490_D1; // @[package.scala 96:25:@24423.4 package.scala 96:25:@24424.4]
  wire  _T_1220; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 470:281:@24441.4]
  wire  _T_1221; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 470:289:@24442.4]
  wire  x499; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 474:24:@24453.4]
  wire  _T_1249; // @[package.scala 96:25:@24488.4 package.scala 96:25:@24489.4]
  wire  _T_1251; // @[implicits.scala 55:10:@24490.4]
  wire  _T_1252; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 485:194:@24491.4]
  wire  x712_x500_D1; // @[package.scala 96:25:@24474.4 package.scala 96:25:@24475.4]
  wire  _T_1253; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 485:281:@24492.4]
  wire  _T_1254; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 485:289:@24493.4]
  wire  x506; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 489:24:@24504.4]
  wire  _T_1282; // @[package.scala 96:25:@24539.4 package.scala 96:25:@24540.4]
  wire  _T_1284; // @[implicits.scala 55:10:@24541.4]
  wire  _T_1285; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 500:194:@24542.4]
  wire  x713_x507_D1; // @[package.scala 96:25:@24525.4 package.scala 96:25:@24526.4]
  wire  _T_1286; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 500:281:@24543.4]
  wire  _T_1287; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 500:289:@24544.4]
  wire  x513; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 504:24:@24555.4]
  wire  _T_1315; // @[package.scala 96:25:@24590.4 package.scala 96:25:@24591.4]
  wire  _T_1317; // @[implicits.scala 55:10:@24592.4]
  wire  _T_1318; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 515:194:@24593.4]
  wire  x714_x514_D1; // @[package.scala 96:25:@24576.4 package.scala 96:25:@24577.4]
  wire  _T_1319; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 515:281:@24594.4]
  wire  _T_1320; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 515:289:@24595.4]
  wire  x520; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 519:24:@24606.4]
  wire  _T_1348; // @[package.scala 96:25:@24641.4 package.scala 96:25:@24642.4]
  wire  _T_1350; // @[implicits.scala 55:10:@24643.4]
  wire  _T_1351; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 530:194:@24644.4]
  wire  x715_x521_D1; // @[package.scala 96:25:@24627.4 package.scala 96:25:@24628.4]
  wire  _T_1352; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 530:281:@24645.4]
  wire  _T_1353; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 530:289:@24646.4]
  wire  x527; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 534:24:@24657.4]
  wire  _T_1381; // @[package.scala 96:25:@24692.4 package.scala 96:25:@24693.4]
  wire  _T_1383; // @[implicits.scala 55:10:@24694.4]
  wire  _T_1384; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 545:194:@24695.4]
  wire  x716_x528_D1; // @[package.scala 96:25:@24678.4 package.scala 96:25:@24679.4]
  wire  _T_1385; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 545:281:@24696.4]
  wire  _T_1386; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 545:289:@24697.4]
  wire [7:0] x396_rd_0_number; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 231:29:@23610.4 sm_x592_inr_Foreach_SAMPLER_BOX.scala 235:336:@23633.4]
  wire [8:0] _GEN_0; // @[Math.scala 450:32:@24709.4]
  wire [8:0] _T_1392; // @[Math.scala 450:32:@24709.4]
  wire [7:0] x449_rd_0_number; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 352:29:@24041.4 sm_x592_inr_Foreach_SAMPLER_BOX.scala 356:406:@24064.4]
  wire [8:0] _GEN_1; // @[Math.scala 450:32:@24716.4]
  wire [8:0] _T_1398; // @[Math.scala 450:32:@24716.4]
  wire [7:0] x456_rd_0_number; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 367:29:@24092.4 sm_x592_inr_Foreach_SAMPLER_BOX.scala 371:406:@24115.4]
  wire [9:0] _GEN_2; // @[Math.scala 450:32:@24721.4]
  wire [9:0] _T_1402; // @[Math.scala 450:32:@24721.4]
  wire [7:0] x463_rd_0_number; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 382:29:@24143.4 sm_x592_inr_Foreach_SAMPLER_BOX.scala 386:406:@24166.4]
  wire [8:0] _GEN_3; // @[Math.scala 450:32:@24726.4]
  wire [8:0] _T_1406; // @[Math.scala 450:32:@24726.4]
  wire [7:0] x504_rd_0_number; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 481:29:@24477.4 sm_x592_inr_Foreach_SAMPLER_BOX.scala 485:406:@24500.4]
  wire [8:0] _GEN_4; // @[Math.scala 450:32:@24731.4]
  wire [8:0] _T_1410; // @[Math.scala 450:32:@24731.4]
  wire [7:0] x546_sum_number; // @[Math.scala 154:22:@24820.4 Math.scala 155:14:@24821.4]
  wire [3:0] _T_1446; // @[FixedPoint.scala 18:52:@24826.4]
  wire [7:0] x404_rd_0_number; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 252:29:@23686.4 sm_x592_inr_Foreach_SAMPLER_BOX.scala 256:336:@23709.4]
  wire [8:0] _GEN_5; // @[Math.scala 450:32:@24839.4]
  wire [8:0] _T_1453; // @[Math.scala 450:32:@24839.4]
  wire [8:0] _GEN_6; // @[Math.scala 450:32:@24844.4]
  wire [8:0] _T_1457; // @[Math.scala 450:32:@24844.4]
  wire [9:0] _GEN_7; // @[Math.scala 450:32:@24849.4]
  wire [9:0] _T_1461; // @[Math.scala 450:32:@24849.4]
  wire [7:0] x470_rd_0_number; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 401:29:@24212.4 sm_x592_inr_Foreach_SAMPLER_BOX.scala 405:406:@24235.4]
  wire [8:0] _GEN_8; // @[Math.scala 450:32:@24854.4]
  wire [8:0] _T_1465; // @[Math.scala 450:32:@24854.4]
  wire [7:0] x511_rd_0_number; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 496:29:@24528.4 sm_x592_inr_Foreach_SAMPLER_BOX.scala 500:406:@24551.4]
  wire [8:0] _GEN_9; // @[Math.scala 450:32:@24859.4]
  wire [8:0] _T_1469; // @[Math.scala 450:32:@24859.4]
  wire [7:0] x560_sum_number; // @[Math.scala 154:22:@24948.4 Math.scala 155:14:@24949.4]
  wire [3:0] _T_1505; // @[FixedPoint.scala 18:52:@24954.4]
  wire [7:0] x412_rd_0_number; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 275:29:@23771.4 sm_x592_inr_Foreach_SAMPLER_BOX.scala 279:336:@23794.4]
  wire [8:0] _GEN_10; // @[Math.scala 450:32:@24967.4]
  wire [8:0] _T_1512; // @[Math.scala 450:32:@24967.4]
  wire [9:0] _GEN_11; // @[Math.scala 450:32:@24972.4]
  wire [9:0] _T_1516; // @[Math.scala 450:32:@24972.4]
  wire [7:0] x477_rd_0_number; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 416:29:@24263.4 sm_x592_inr_Foreach_SAMPLER_BOX.scala 420:406:@24286.4]
  wire [8:0] _GEN_12; // @[Math.scala 450:32:@24977.4]
  wire [8:0] _T_1520; // @[Math.scala 450:32:@24977.4]
  wire [7:0] x518_rd_0_number; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 511:29:@24579.4 sm_x592_inr_Foreach_SAMPLER_BOX.scala 515:406:@24602.4]
  wire [8:0] _GEN_13; // @[Math.scala 450:32:@24982.4]
  wire [8:0] _T_1524; // @[Math.scala 450:32:@24982.4]
  wire [7:0] x573_sum_number; // @[Math.scala 154:22:@25071.4 Math.scala 155:14:@25072.4]
  wire [3:0] _T_1560; // @[FixedPoint.scala 18:52:@25077.4]
  wire [7:0] x424_rd_0_number; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 302:29:@23850.4 sm_x592_inr_Foreach_SAMPLER_BOX.scala 306:441:@23873.4]
  wire [8:0] _GEN_14; // @[Math.scala 450:32:@25090.4]
  wire [8:0] _T_1567; // @[Math.scala 450:32:@25090.4]
  wire [9:0] _GEN_15; // @[Math.scala 450:32:@25095.4]
  wire [9:0] _T_1571; // @[Math.scala 450:32:@25095.4]
  wire [7:0] x484_rd_0_number; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 439:29:@24316.4 sm_x592_inr_Foreach_SAMPLER_BOX.scala 443:406:@24339.4]
  wire [8:0] _GEN_16; // @[Math.scala 450:32:@25100.4]
  wire [8:0] _T_1575; // @[Math.scala 450:32:@25100.4]
  wire [7:0] x525_rd_0_number; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 526:29:@24630.4 sm_x592_inr_Foreach_SAMPLER_BOX.scala 530:406:@24653.4]
  wire [8:0] _GEN_17; // @[Math.scala 450:32:@25105.4]
  wire [8:0] _T_1579; // @[Math.scala 450:32:@25105.4]
  wire [7:0] x586_sum_number; // @[Math.scala 154:22:@25196.4 Math.scala 155:14:@25197.4]
  wire [3:0] _T_1617; // @[FixedPoint.scala 18:52:@25202.4]
  wire [7:0] x574_number; // @[package.scala 96:25:@25084.4 package.scala 96:25:@25085.4]
  wire [7:0] x587_number; // @[package.scala 96:25:@25209.4 package.scala 96:25:@25210.4]
  wire [15:0] _T_1632; // @[Cat.scala 30:58:@25219.4]
  wire [7:0] x547_number; // @[package.scala 96:25:@24833.4 package.scala 96:25:@24834.4]
  wire [7:0] x561_number; // @[package.scala 96:25:@24961.4 package.scala 96:25:@24962.4]
  wire [15:0] _T_1633; // @[Cat.scala 30:58:@25220.4]
  wire  _T_1646; // @[package.scala 96:25:@25256.4 package.scala 96:25:@25257.4]
  wire  _T_1648; // @[implicits.scala 55:10:@25258.4]
  wire  x721_b327_D15; // @[package.scala 96:25:@25238.4 package.scala 96:25:@25239.4]
  wire  _T_1649; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 689:116:@25259.4]
  wire  x722_b328_D15; // @[package.scala 96:25:@25247.4 package.scala 96:25:@25248.4]
  wire  _T_1650; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 689:122:@25260.4]
  wire [31:0] x668_x660_D4_number; // @[package.scala 96:25:@23089.4 package.scala 96:25:@23090.4]
  wire [31:0] x670_x343_sum_D3_number; // @[package.scala 96:25:@23107.4 package.scala 96:25:@23108.4]
  wire [31:0] x674_x353_sum_D2_number; // @[package.scala 96:25:@23201.4 package.scala 96:25:@23202.4]
  wire [31:0] x676_x362_sum_D2_number; // @[package.scala 96:25:@23277.4 package.scala 96:25:@23278.4]
  wire [31:0] x678_x371_sum_D2_number; // @[package.scala 96:25:@23353.4 package.scala 96:25:@23354.4]
  wire [31:0] x384_sum_number; // @[Math.scala 154:22:@23495.4 Math.scala 155:14:@23496.4]
  wire [31:0] x687_x662_D2_number; // @[package.scala 96:25:@23522.4 package.scala 96:25:@23523.4]
  wire [31:0] x393_sum_number; // @[Math.scala 154:22:@23598.4 Math.scala 155:14:@23599.4]
  wire [31:0] x401_sum_number; // @[Math.scala 154:22:@23674.4 Math.scala 155:14:@23675.4]
  wire [31:0] x698_x409_sum_D1_number; // @[package.scala 96:25:@23768.4 package.scala 96:25:@23769.4]
  wire [31:0] x420_sum_number; // @[Math.scala 154:22:@23838.4 Math.scala 155:14:@23839.4]
  wire [31:0] x432_sum_number; // @[Math.scala 154:22:@23919.4 Math.scala 155:14:@23920.4]
  wire [31:0] x445_sum_number; // @[Math.scala 154:22:@24020.4 Math.scala 155:14:@24021.4]
  wire [31:0] x701_x664_D1_number; // @[package.scala 96:25:@24029.4 package.scala 96:25:@24030.4]
  wire [31:0] x453_sum_number; // @[Math.scala 154:22:@24080.4 Math.scala 155:14:@24081.4]
  wire [31:0] x460_sum_number; // @[Math.scala 154:22:@24131.4 Math.scala 155:14:@24132.4]
  wire [31:0] x467_sum_number; // @[Math.scala 154:22:@24200.4 Math.scala 155:14:@24201.4]
  wire [31:0] x474_sum_number; // @[Math.scala 154:22:@24251.4 Math.scala 155:14:@24252.4]
  wire [31:0] x481_sum_number; // @[Math.scala 154:22:@24304.4 Math.scala 155:14:@24305.4]
  wire [31:0] x493_sum_number; // @[Math.scala 154:22:@24405.4 Math.scala 155:14:@24406.4]
  wire [31:0] x710_x666_D1_number; // @[package.scala 96:25:@24414.4 package.scala 96:25:@24415.4]
  wire [31:0] x501_sum_number; // @[Math.scala 154:22:@24465.4 Math.scala 155:14:@24466.4]
  wire [31:0] x508_sum_number; // @[Math.scala 154:22:@24516.4 Math.scala 155:14:@24517.4]
  wire [31:0] x515_sum_number; // @[Math.scala 154:22:@24567.4 Math.scala 155:14:@24568.4]
  wire [31:0] x522_sum_number; // @[Math.scala 154:22:@24618.4 Math.scala 155:14:@24619.4]
  wire [31:0] x529_sum_number; // @[Math.scala 154:22:@24669.4 Math.scala 155:14:@24670.4]
  _ _ ( // @[Math.scala 709:24:@22794.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 709:24:@22806.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  x329_lb_0 x329_lb_0 ( // @[m_x329_lb_0.scala 47:17:@22816.4]
    .clock(x329_lb_0_clock),
    .reset(x329_lb_0_reset),
    .io_rPort_17_banks_0(x329_lb_0_io_rPort_17_banks_0),
    .io_rPort_17_ofs_0(x329_lb_0_io_rPort_17_ofs_0),
    .io_rPort_17_en_0(x329_lb_0_io_rPort_17_en_0),
    .io_rPort_17_backpressure(x329_lb_0_io_rPort_17_backpressure),
    .io_rPort_17_output_0(x329_lb_0_io_rPort_17_output_0),
    .io_rPort_16_banks_0(x329_lb_0_io_rPort_16_banks_0),
    .io_rPort_16_ofs_0(x329_lb_0_io_rPort_16_ofs_0),
    .io_rPort_16_en_0(x329_lb_0_io_rPort_16_en_0),
    .io_rPort_16_backpressure(x329_lb_0_io_rPort_16_backpressure),
    .io_rPort_16_output_0(x329_lb_0_io_rPort_16_output_0),
    .io_rPort_15_banks_0(x329_lb_0_io_rPort_15_banks_0),
    .io_rPort_15_ofs_0(x329_lb_0_io_rPort_15_ofs_0),
    .io_rPort_15_en_0(x329_lb_0_io_rPort_15_en_0),
    .io_rPort_15_backpressure(x329_lb_0_io_rPort_15_backpressure),
    .io_rPort_15_output_0(x329_lb_0_io_rPort_15_output_0),
    .io_rPort_14_banks_0(x329_lb_0_io_rPort_14_banks_0),
    .io_rPort_14_ofs_0(x329_lb_0_io_rPort_14_ofs_0),
    .io_rPort_14_en_0(x329_lb_0_io_rPort_14_en_0),
    .io_rPort_14_backpressure(x329_lb_0_io_rPort_14_backpressure),
    .io_rPort_14_output_0(x329_lb_0_io_rPort_14_output_0),
    .io_rPort_13_banks_0(x329_lb_0_io_rPort_13_banks_0),
    .io_rPort_13_ofs_0(x329_lb_0_io_rPort_13_ofs_0),
    .io_rPort_13_en_0(x329_lb_0_io_rPort_13_en_0),
    .io_rPort_13_backpressure(x329_lb_0_io_rPort_13_backpressure),
    .io_rPort_13_output_0(x329_lb_0_io_rPort_13_output_0),
    .io_rPort_12_banks_0(x329_lb_0_io_rPort_12_banks_0),
    .io_rPort_12_ofs_0(x329_lb_0_io_rPort_12_ofs_0),
    .io_rPort_12_en_0(x329_lb_0_io_rPort_12_en_0),
    .io_rPort_12_backpressure(x329_lb_0_io_rPort_12_backpressure),
    .io_rPort_12_output_0(x329_lb_0_io_rPort_12_output_0),
    .io_rPort_11_banks_0(x329_lb_0_io_rPort_11_banks_0),
    .io_rPort_11_ofs_0(x329_lb_0_io_rPort_11_ofs_0),
    .io_rPort_11_en_0(x329_lb_0_io_rPort_11_en_0),
    .io_rPort_11_backpressure(x329_lb_0_io_rPort_11_backpressure),
    .io_rPort_11_output_0(x329_lb_0_io_rPort_11_output_0),
    .io_rPort_10_banks_0(x329_lb_0_io_rPort_10_banks_0),
    .io_rPort_10_ofs_0(x329_lb_0_io_rPort_10_ofs_0),
    .io_rPort_10_en_0(x329_lb_0_io_rPort_10_en_0),
    .io_rPort_10_backpressure(x329_lb_0_io_rPort_10_backpressure),
    .io_rPort_10_output_0(x329_lb_0_io_rPort_10_output_0),
    .io_rPort_9_banks_0(x329_lb_0_io_rPort_9_banks_0),
    .io_rPort_9_ofs_0(x329_lb_0_io_rPort_9_ofs_0),
    .io_rPort_9_en_0(x329_lb_0_io_rPort_9_en_0),
    .io_rPort_9_backpressure(x329_lb_0_io_rPort_9_backpressure),
    .io_rPort_9_output_0(x329_lb_0_io_rPort_9_output_0),
    .io_rPort_8_banks_0(x329_lb_0_io_rPort_8_banks_0),
    .io_rPort_8_ofs_0(x329_lb_0_io_rPort_8_ofs_0),
    .io_rPort_8_en_0(x329_lb_0_io_rPort_8_en_0),
    .io_rPort_8_backpressure(x329_lb_0_io_rPort_8_backpressure),
    .io_rPort_8_output_0(x329_lb_0_io_rPort_8_output_0),
    .io_rPort_7_banks_0(x329_lb_0_io_rPort_7_banks_0),
    .io_rPort_7_ofs_0(x329_lb_0_io_rPort_7_ofs_0),
    .io_rPort_7_en_0(x329_lb_0_io_rPort_7_en_0),
    .io_rPort_7_backpressure(x329_lb_0_io_rPort_7_backpressure),
    .io_rPort_7_output_0(x329_lb_0_io_rPort_7_output_0),
    .io_rPort_6_banks_0(x329_lb_0_io_rPort_6_banks_0),
    .io_rPort_6_ofs_0(x329_lb_0_io_rPort_6_ofs_0),
    .io_rPort_6_en_0(x329_lb_0_io_rPort_6_en_0),
    .io_rPort_6_backpressure(x329_lb_0_io_rPort_6_backpressure),
    .io_rPort_6_output_0(x329_lb_0_io_rPort_6_output_0),
    .io_rPort_5_banks_0(x329_lb_0_io_rPort_5_banks_0),
    .io_rPort_5_ofs_0(x329_lb_0_io_rPort_5_ofs_0),
    .io_rPort_5_en_0(x329_lb_0_io_rPort_5_en_0),
    .io_rPort_5_backpressure(x329_lb_0_io_rPort_5_backpressure),
    .io_rPort_5_output_0(x329_lb_0_io_rPort_5_output_0),
    .io_rPort_4_banks_0(x329_lb_0_io_rPort_4_banks_0),
    .io_rPort_4_ofs_0(x329_lb_0_io_rPort_4_ofs_0),
    .io_rPort_4_en_0(x329_lb_0_io_rPort_4_en_0),
    .io_rPort_4_backpressure(x329_lb_0_io_rPort_4_backpressure),
    .io_rPort_4_output_0(x329_lb_0_io_rPort_4_output_0),
    .io_rPort_3_banks_0(x329_lb_0_io_rPort_3_banks_0),
    .io_rPort_3_ofs_0(x329_lb_0_io_rPort_3_ofs_0),
    .io_rPort_3_en_0(x329_lb_0_io_rPort_3_en_0),
    .io_rPort_3_backpressure(x329_lb_0_io_rPort_3_backpressure),
    .io_rPort_3_output_0(x329_lb_0_io_rPort_3_output_0),
    .io_rPort_2_banks_0(x329_lb_0_io_rPort_2_banks_0),
    .io_rPort_2_ofs_0(x329_lb_0_io_rPort_2_ofs_0),
    .io_rPort_2_en_0(x329_lb_0_io_rPort_2_en_0),
    .io_rPort_2_backpressure(x329_lb_0_io_rPort_2_backpressure),
    .io_rPort_2_output_0(x329_lb_0_io_rPort_2_output_0),
    .io_rPort_1_banks_0(x329_lb_0_io_rPort_1_banks_0),
    .io_rPort_1_ofs_0(x329_lb_0_io_rPort_1_ofs_0),
    .io_rPort_1_en_0(x329_lb_0_io_rPort_1_en_0),
    .io_rPort_1_backpressure(x329_lb_0_io_rPort_1_backpressure),
    .io_rPort_1_output_0(x329_lb_0_io_rPort_1_output_0),
    .io_rPort_0_banks_0(x329_lb_0_io_rPort_0_banks_0),
    .io_rPort_0_ofs_0(x329_lb_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x329_lb_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x329_lb_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x329_lb_0_io_rPort_0_output_0),
    .io_wPort_3_banks_0(x329_lb_0_io_wPort_3_banks_0),
    .io_wPort_3_ofs_0(x329_lb_0_io_wPort_3_ofs_0),
    .io_wPort_3_data_0(x329_lb_0_io_wPort_3_data_0),
    .io_wPort_3_en_0(x329_lb_0_io_wPort_3_en_0),
    .io_wPort_2_banks_0(x329_lb_0_io_wPort_2_banks_0),
    .io_wPort_2_ofs_0(x329_lb_0_io_wPort_2_ofs_0),
    .io_wPort_2_data_0(x329_lb_0_io_wPort_2_data_0),
    .io_wPort_2_en_0(x329_lb_0_io_wPort_2_en_0),
    .io_wPort_1_banks_0(x329_lb_0_io_wPort_1_banks_0),
    .io_wPort_1_ofs_0(x329_lb_0_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(x329_lb_0_io_wPort_1_data_0),
    .io_wPort_1_en_0(x329_lb_0_io_wPort_1_en_0),
    .io_wPort_0_banks_0(x329_lb_0_io_wPort_0_banks_0),
    .io_wPort_0_ofs_0(x329_lb_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x329_lb_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x329_lb_0_io_wPort_0_en_0)
  );
  RetimeWrapper_124 RetimeWrapper ( // @[package.scala 93:22:@22974.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x343_sum x343_sum_1 ( // @[Math.scala 150:24:@23074.4]
    .clock(x343_sum_1_clock),
    .reset(x343_sum_1_reset),
    .io_a(x343_sum_1_io_a),
    .io_b(x343_sum_1_io_b),
    .io_flow(x343_sum_1_io_flow),
    .io_result(x343_sum_1_io_result)
  );
  RetimeWrapper_126 RetimeWrapper_1 ( // @[package.scala 93:22:@23084.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_127 RetimeWrapper_2 ( // @[package.scala 93:22:@23093.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_128 RetimeWrapper_3 ( // @[package.scala 93:22:@23102.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_127 RetimeWrapper_4 ( // @[package.scala 93:22:@23111.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_130 RetimeWrapper_5 ( // @[package.scala 93:22:@23120.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_127 RetimeWrapper_6 ( // @[package.scala 93:22:@23133.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  x343_sum x349_rdcol_1 ( // @[Math.scala 150:24:@23156.4]
    .clock(x349_rdcol_1_clock),
    .reset(x349_rdcol_1_reset),
    .io_a(x349_rdcol_1_io_a),
    .io_b(x349_rdcol_1_io_b),
    .io_flow(x349_rdcol_1_io_flow),
    .io_result(x349_rdcol_1_io_result)
  );
  RetimeWrapper_124 RetimeWrapper_7 ( // @[package.scala 93:22:@23177.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  x343_sum x353_sum_1 ( // @[Math.scala 150:24:@23186.4]
    .clock(x353_sum_1_clock),
    .reset(x353_sum_1_reset),
    .io_a(x353_sum_1_io_a),
    .io_b(x353_sum_1_io_b),
    .io_flow(x353_sum_1_io_flow),
    .io_result(x353_sum_1_io_result)
  );
  RetimeWrapper_135 RetimeWrapper_8 ( // @[package.scala 93:22:@23196.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_130 RetimeWrapper_9 ( // @[package.scala 93:22:@23205.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_127 RetimeWrapper_10 ( // @[package.scala 93:22:@23218.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  x343_sum x358_rdcol_1 ( // @[Math.scala 150:24:@23241.4]
    .clock(x358_rdcol_1_clock),
    .reset(x358_rdcol_1_reset),
    .io_a(x358_rdcol_1_io_a),
    .io_b(x358_rdcol_1_io_b),
    .io_flow(x358_rdcol_1_io_flow),
    .io_result(x358_rdcol_1_io_result)
  );
  x343_sum x362_sum_1 ( // @[Math.scala 150:24:@23262.4]
    .clock(x362_sum_1_clock),
    .reset(x362_sum_1_reset),
    .io_a(x362_sum_1_io_a),
    .io_b(x362_sum_1_io_b),
    .io_flow(x362_sum_1_io_flow),
    .io_result(x362_sum_1_io_result)
  );
  RetimeWrapper_135 RetimeWrapper_11 ( // @[package.scala 93:22:@23272.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_130 RetimeWrapper_12 ( // @[package.scala 93:22:@23281.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_127 RetimeWrapper_13 ( // @[package.scala 93:22:@23294.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  x343_sum x367_rdcol_1 ( // @[Math.scala 150:24:@23317.4]
    .clock(x367_rdcol_1_clock),
    .reset(x367_rdcol_1_reset),
    .io_a(x367_rdcol_1_io_a),
    .io_b(x367_rdcol_1_io_b),
    .io_flow(x367_rdcol_1_io_flow),
    .io_result(x367_rdcol_1_io_result)
  );
  x343_sum x371_sum_1 ( // @[Math.scala 150:24:@23338.4]
    .clock(x371_sum_1_clock),
    .reset(x371_sum_1_reset),
    .io_a(x371_sum_1_io_a),
    .io_b(x371_sum_1_io_b),
    .io_flow(x371_sum_1_io_flow),
    .io_result(x371_sum_1_io_result)
  );
  RetimeWrapper_135 RetimeWrapper_14 ( // @[package.scala 93:22:@23348.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_130 RetimeWrapper_15 ( // @[package.scala 93:22:@23357.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_127 RetimeWrapper_16 ( // @[package.scala 93:22:@23370.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_148 RetimeWrapper_17 ( // @[package.scala 93:22:@23391.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_148 RetimeWrapper_18 ( // @[package.scala 93:22:@23418.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper RetimeWrapper_19 ( // @[package.scala 93:22:@23434.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_124 RetimeWrapper_20 ( // @[package.scala 93:22:@23471.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_148 RetimeWrapper_21 ( // @[package.scala 93:22:@23480.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  x343_sum x384_sum_1 ( // @[Math.scala 150:24:@23489.4]
    .clock(x384_sum_1_clock),
    .reset(x384_sum_1_reset),
    .io_a(x384_sum_1_io_a),
    .io_b(x384_sum_1_io_b),
    .io_flow(x384_sum_1_io_flow),
    .io_result(x384_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_22 ( // @[package.scala 93:22:@23499.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_155 RetimeWrapper_23 ( // @[package.scala 93:22:@23508.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_135 RetimeWrapper_24 ( // @[package.scala 93:22:@23517.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_155 RetimeWrapper_25 ( // @[package.scala 93:22:@23526.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_155 RetimeWrapper_26 ( // @[package.scala 93:22:@23540.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_148 RetimeWrapper_27 ( // @[package.scala 93:22:@23561.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_148 RetimeWrapper_28 ( // @[package.scala 93:22:@23583.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  x343_sum x393_sum_1 ( // @[Math.scala 150:24:@23592.4]
    .clock(x393_sum_1_clock),
    .reset(x393_sum_1_reset),
    .io_a(x393_sum_1_io_a),
    .io_b(x393_sum_1_io_b),
    .io_flow(x393_sum_1_io_flow),
    .io_result(x393_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_29 ( // @[package.scala 93:22:@23602.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_155 RetimeWrapper_30 ( // @[package.scala 93:22:@23616.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_148 RetimeWrapper_31 ( // @[package.scala 93:22:@23637.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_148 RetimeWrapper_32 ( // @[package.scala 93:22:@23659.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  x343_sum x401_sum_1 ( // @[Math.scala 150:24:@23668.4]
    .clock(x401_sum_1_clock),
    .reset(x401_sum_1_reset),
    .io_a(x401_sum_1_io_a),
    .io_b(x401_sum_1_io_b),
    .io_flow(x401_sum_1_io_flow),
    .io_result(x401_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_33 ( // @[package.scala 93:22:@23678.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_155 RetimeWrapper_34 ( // @[package.scala 93:22:@23692.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_148 RetimeWrapper_35 ( // @[package.scala 93:22:@23713.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_148 RetimeWrapper_36 ( // @[package.scala 93:22:@23735.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  x343_sum x409_sum_1 ( // @[Math.scala 150:24:@23744.4]
    .clock(x409_sum_1_clock),
    .reset(x409_sum_1_reset),
    .io_a(x409_sum_1_io_a),
    .io_b(x409_sum_1_io_b),
    .io_flow(x409_sum_1_io_flow),
    .io_result(x409_sum_1_io_result)
  );
  RetimeWrapper_52 RetimeWrapper_37 ( // @[package.scala 93:22:@23754.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_124 RetimeWrapper_38 ( // @[package.scala 93:22:@23763.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_155 RetimeWrapper_39 ( // @[package.scala 93:22:@23777.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  x343_sum x414_rdcol_1 ( // @[Math.scala 150:24:@23800.4]
    .clock(x414_rdcol_1_clock),
    .reset(x414_rdcol_1_reset),
    .io_a(x414_rdcol_1_io_a),
    .io_b(x414_rdcol_1_io_b),
    .io_flow(x414_rdcol_1_io_flow),
    .io_result(x414_rdcol_1_io_result)
  );
  x343_sum x420_sum_1 ( // @[Math.scala 150:24:@23832.4]
    .clock(x420_sum_1_clock),
    .reset(x420_sum_1_reset),
    .io_a(x420_sum_1_io_a),
    .io_b(x420_sum_1_io_b),
    .io_flow(x420_sum_1_io_flow),
    .io_result(x420_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_40 ( // @[package.scala 93:22:@23842.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper_155 RetimeWrapper_41 ( // @[package.scala 93:22:@23856.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  x343_sum x426_rdcol_1 ( // @[Math.scala 150:24:@23881.4]
    .clock(x426_rdcol_1_clock),
    .reset(x426_rdcol_1_reset),
    .io_a(x426_rdcol_1_io_a),
    .io_b(x426_rdcol_1_io_b),
    .io_flow(x426_rdcol_1_io_flow),
    .io_result(x426_rdcol_1_io_result)
  );
  x343_sum x432_sum_1 ( // @[Math.scala 150:24:@23913.4]
    .clock(x432_sum_1_clock),
    .reset(x432_sum_1_reset),
    .io_a(x432_sum_1_io_a),
    .io_b(x432_sum_1_io_b),
    .io_flow(x432_sum_1_io_flow),
    .io_result(x432_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_42 ( // @[package.scala 93:22:@23923.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_155 RetimeWrapper_43 ( // @[package.scala 93:22:@23937.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  x438_rdrow x438_rdrow_1 ( // @[Math.scala 191:24:@23960.4]
    .clock(x438_rdrow_1_clock),
    .reset(x438_rdrow_1_reset),
    .io_a(x438_rdrow_1_io_a),
    .io_b(x438_rdrow_1_io_b),
    .io_flow(x438_rdrow_1_io_flow),
    .io_result(x438_rdrow_1_io_result)
  );
  x343_sum x445_sum_1 ( // @[Math.scala 150:24:@24014.4]
    .clock(x445_sum_1_clock),
    .reset(x445_sum_1_reset),
    .io_a(x445_sum_1_io_a),
    .io_b(x445_sum_1_io_b),
    .io_flow(x445_sum_1_io_flow),
    .io_result(x445_sum_1_io_result)
  );
  RetimeWrapper_124 RetimeWrapper_44 ( // @[package.scala 93:22:@24024.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper RetimeWrapper_45 ( // @[package.scala 93:22:@24033.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_155 RetimeWrapper_46 ( // @[package.scala 93:22:@24047.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  x343_sum x453_sum_1 ( // @[Math.scala 150:24:@24074.4]
    .clock(x453_sum_1_clock),
    .reset(x453_sum_1_reset),
    .io_a(x453_sum_1_io_a),
    .io_b(x453_sum_1_io_b),
    .io_flow(x453_sum_1_io_flow),
    .io_result(x453_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_47 ( // @[package.scala 93:22:@24084.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_155 RetimeWrapper_48 ( // @[package.scala 93:22:@24098.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  x343_sum x460_sum_1 ( // @[Math.scala 150:24:@24125.4]
    .clock(x460_sum_1_clock),
    .reset(x460_sum_1_reset),
    .io_a(x460_sum_1_io_a),
    .io_b(x460_sum_1_io_b),
    .io_flow(x460_sum_1_io_flow),
    .io_result(x460_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_49 ( // @[package.scala 93:22:@24135.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_155 RetimeWrapper_50 ( // @[package.scala 93:22:@24149.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper RetimeWrapper_51 ( // @[package.scala 93:22:@24170.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_195 RetimeWrapper_52 ( // @[package.scala 93:22:@24185.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  x343_sum x467_sum_1 ( // @[Math.scala 150:24:@24194.4]
    .clock(x467_sum_1_clock),
    .reset(x467_sum_1_reset),
    .io_a(x467_sum_1_io_a),
    .io_b(x467_sum_1_io_b),
    .io_flow(x467_sum_1_io_flow),
    .io_result(x467_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_53 ( // @[package.scala 93:22:@24204.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper_155 RetimeWrapper_54 ( // @[package.scala 93:22:@24218.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  x343_sum x474_sum_1 ( // @[Math.scala 150:24:@24245.4]
    .clock(x474_sum_1_clock),
    .reset(x474_sum_1_reset),
    .io_a(x474_sum_1_io_a),
    .io_b(x474_sum_1_io_b),
    .io_flow(x474_sum_1_io_flow),
    .io_result(x474_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_55 ( // @[package.scala 93:22:@24255.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper_155 RetimeWrapper_56 ( // @[package.scala 93:22:@24269.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  x343_sum x481_sum_1 ( // @[Math.scala 150:24:@24298.4]
    .clock(x481_sum_1_clock),
    .reset(x481_sum_1_reset),
    .io_a(x481_sum_1_io_a),
    .io_b(x481_sum_1_io_b),
    .io_flow(x481_sum_1_io_flow),
    .io_result(x481_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_57 ( // @[package.scala 93:22:@24308.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper_155 RetimeWrapper_58 ( // @[package.scala 93:22:@24322.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  x438_rdrow x486_rdrow_1 ( // @[Math.scala 191:24:@24345.4]
    .clock(x486_rdrow_1_clock),
    .reset(x486_rdrow_1_reset),
    .io_a(x486_rdrow_1_io_a),
    .io_b(x486_rdrow_1_io_b),
    .io_flow(x486_rdrow_1_io_flow),
    .io_result(x486_rdrow_1_io_result)
  );
  x343_sum x493_sum_1 ( // @[Math.scala 150:24:@24399.4]
    .clock(x493_sum_1_clock),
    .reset(x493_sum_1_reset),
    .io_a(x493_sum_1_io_a),
    .io_b(x493_sum_1_io_b),
    .io_flow(x493_sum_1_io_flow),
    .io_result(x493_sum_1_io_result)
  );
  RetimeWrapper_124 RetimeWrapper_59 ( // @[package.scala 93:22:@24409.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper RetimeWrapper_60 ( // @[package.scala 93:22:@24418.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_155 RetimeWrapper_61 ( // @[package.scala 93:22:@24432.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  x343_sum x501_sum_1 ( // @[Math.scala 150:24:@24459.4]
    .clock(x501_sum_1_clock),
    .reset(x501_sum_1_reset),
    .io_a(x501_sum_1_io_a),
    .io_b(x501_sum_1_io_b),
    .io_flow(x501_sum_1_io_flow),
    .io_result(x501_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_62 ( // @[package.scala 93:22:@24469.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_155 RetimeWrapper_63 ( // @[package.scala 93:22:@24483.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  x343_sum x508_sum_1 ( // @[Math.scala 150:24:@24510.4]
    .clock(x508_sum_1_clock),
    .reset(x508_sum_1_reset),
    .io_a(x508_sum_1_io_a),
    .io_b(x508_sum_1_io_b),
    .io_flow(x508_sum_1_io_flow),
    .io_result(x508_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_64 ( // @[package.scala 93:22:@24520.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_155 RetimeWrapper_65 ( // @[package.scala 93:22:@24534.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  x343_sum x515_sum_1 ( // @[Math.scala 150:24:@24561.4]
    .clock(x515_sum_1_clock),
    .reset(x515_sum_1_reset),
    .io_a(x515_sum_1_io_a),
    .io_b(x515_sum_1_io_b),
    .io_flow(x515_sum_1_io_flow),
    .io_result(x515_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_66 ( // @[package.scala 93:22:@24571.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper_155 RetimeWrapper_67 ( // @[package.scala 93:22:@24585.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  x343_sum x522_sum_1 ( // @[Math.scala 150:24:@24612.4]
    .clock(x522_sum_1_clock),
    .reset(x522_sum_1_reset),
    .io_a(x522_sum_1_io_a),
    .io_b(x522_sum_1_io_b),
    .io_flow(x522_sum_1_io_flow),
    .io_result(x522_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_68 ( // @[package.scala 93:22:@24622.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_155 RetimeWrapper_69 ( // @[package.scala 93:22:@24636.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  x343_sum x529_sum_1 ( // @[Math.scala 150:24:@24663.4]
    .clock(x529_sum_1_clock),
    .reset(x529_sum_1_reset),
    .io_a(x529_sum_1_io_a),
    .io_b(x529_sum_1_io_b),
    .io_flow(x529_sum_1_io_flow),
    .io_result(x529_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_70 ( // @[package.scala 93:22:@24673.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_155 RetimeWrapper_71 ( // @[package.scala 93:22:@24687.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  x539_x11 x539_x11_1 ( // @[Math.scala 150:24:@24735.4]
    .clock(x539_x11_1_clock),
    .reset(x539_x11_1_reset),
    .io_a(x539_x11_1_io_a),
    .io_b(x539_x11_1_io_b),
    .io_flow(x539_x11_1_io_flow),
    .io_result(x539_x11_1_io_result)
  );
  x539_x11 x540_x12_1 ( // @[Math.scala 150:24:@24745.4]
    .clock(x540_x12_1_clock),
    .reset(x540_x12_1_reset),
    .io_a(x540_x12_1_io_a),
    .io_b(x540_x12_1_io_b),
    .io_flow(x540_x12_1_io_flow),
    .io_result(x540_x12_1_io_result)
  );
  x539_x11 x541_x11_1 ( // @[Math.scala 150:24:@24755.4]
    .clock(x541_x11_1_clock),
    .reset(x541_x11_1_reset),
    .io_a(x541_x11_1_io_a),
    .io_b(x541_x11_1_io_b),
    .io_flow(x541_x11_1_io_flow),
    .io_result(x541_x11_1_io_result)
  );
  x539_x11 x542_x12_1 ( // @[Math.scala 150:24:@24765.4]
    .clock(x542_x12_1_clock),
    .reset(x542_x12_1_reset),
    .io_a(x542_x12_1_io_a),
    .io_b(x542_x12_1_io_b),
    .io_flow(x542_x12_1_io_flow),
    .io_result(x542_x12_1_io_result)
  );
  x543_x11 x543_x11_1 ( // @[Math.scala 150:24:@24775.4]
    .io_a(x543_x11_1_io_a),
    .io_b(x543_x11_1_io_b),
    .io_result(x543_x11_1_io_result)
  );
  x543_x11 x544_x12_1 ( // @[Math.scala 150:24:@24785.4]
    .io_a(x544_x12_1_io_a),
    .io_b(x544_x12_1_io_b),
    .io_result(x544_x12_1_io_result)
  );
  x543_x11 x545_x11_1 ( // @[Math.scala 150:24:@24795.4]
    .io_a(x545_x11_1_io_a),
    .io_b(x545_x11_1_io_b),
    .io_result(x545_x11_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_72 ( // @[package.scala 93:22:@24805.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  x543_x11 x546_sum_1 ( // @[Math.scala 150:24:@24814.4]
    .io_a(x546_sum_1_io_a),
    .io_b(x546_sum_1_io_b),
    .io_result(x546_sum_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_73 ( // @[package.scala 93:22:@24828.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  x539_x11 x553_x11_1 ( // @[Math.scala 150:24:@24863.4]
    .clock(x553_x11_1_clock),
    .reset(x553_x11_1_reset),
    .io_a(x553_x11_1_io_a),
    .io_b(x553_x11_1_io_b),
    .io_flow(x553_x11_1_io_flow),
    .io_result(x553_x11_1_io_result)
  );
  x539_x11 x554_x12_1 ( // @[Math.scala 150:24:@24873.4]
    .clock(x554_x12_1_clock),
    .reset(x554_x12_1_reset),
    .io_a(x554_x12_1_io_a),
    .io_b(x554_x12_1_io_b),
    .io_flow(x554_x12_1_io_flow),
    .io_result(x554_x12_1_io_result)
  );
  x539_x11 x555_x11_1 ( // @[Math.scala 150:24:@24883.4]
    .clock(x555_x11_1_clock),
    .reset(x555_x11_1_reset),
    .io_a(x555_x11_1_io_a),
    .io_b(x555_x11_1_io_b),
    .io_flow(x555_x11_1_io_flow),
    .io_result(x555_x11_1_io_result)
  );
  x539_x11 x556_x12_1 ( // @[Math.scala 150:24:@24893.4]
    .clock(x556_x12_1_clock),
    .reset(x556_x12_1_reset),
    .io_a(x556_x12_1_io_a),
    .io_b(x556_x12_1_io_b),
    .io_flow(x556_x12_1_io_flow),
    .io_result(x556_x12_1_io_result)
  );
  x543_x11 x557_x11_1 ( // @[Math.scala 150:24:@24903.4]
    .io_a(x557_x11_1_io_a),
    .io_b(x557_x11_1_io_b),
    .io_result(x557_x11_1_io_result)
  );
  x543_x11 x558_x12_1 ( // @[Math.scala 150:24:@24913.4]
    .io_a(x558_x12_1_io_a),
    .io_b(x558_x12_1_io_b),
    .io_result(x558_x12_1_io_result)
  );
  x543_x11 x559_x11_1 ( // @[Math.scala 150:24:@24923.4]
    .io_a(x559_x11_1_io_a),
    .io_b(x559_x11_1_io_b),
    .io_result(x559_x11_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_74 ( // @[package.scala 93:22:@24933.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  x543_x11 x560_sum_1 ( // @[Math.scala 150:24:@24942.4]
    .io_a(x560_sum_1_io_a),
    .io_b(x560_sum_1_io_b),
    .io_result(x560_sum_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_75 ( // @[package.scala 93:22:@24956.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  x539_x11 x566_x11_1 ( // @[Math.scala 150:24:@24986.4]
    .clock(x566_x11_1_clock),
    .reset(x566_x11_1_reset),
    .io_a(x566_x11_1_io_a),
    .io_b(x566_x11_1_io_b),
    .io_flow(x566_x11_1_io_flow),
    .io_result(x566_x11_1_io_result)
  );
  x539_x11 x567_x12_1 ( // @[Math.scala 150:24:@24996.4]
    .clock(x567_x12_1_clock),
    .reset(x567_x12_1_reset),
    .io_a(x567_x12_1_io_a),
    .io_b(x567_x12_1_io_b),
    .io_flow(x567_x12_1_io_flow),
    .io_result(x567_x12_1_io_result)
  );
  x539_x11 x568_x11_1 ( // @[Math.scala 150:24:@25006.4]
    .clock(x568_x11_1_clock),
    .reset(x568_x11_1_reset),
    .io_a(x568_x11_1_io_a),
    .io_b(x568_x11_1_io_b),
    .io_flow(x568_x11_1_io_flow),
    .io_result(x568_x11_1_io_result)
  );
  x539_x11 x569_x12_1 ( // @[Math.scala 150:24:@25016.4]
    .clock(x569_x12_1_clock),
    .reset(x569_x12_1_reset),
    .io_a(x569_x12_1_io_a),
    .io_b(x569_x12_1_io_b),
    .io_flow(x569_x12_1_io_flow),
    .io_result(x569_x12_1_io_result)
  );
  x543_x11 x570_x11_1 ( // @[Math.scala 150:24:@25026.4]
    .io_a(x570_x11_1_io_a),
    .io_b(x570_x11_1_io_b),
    .io_result(x570_x11_1_io_result)
  );
  x543_x11 x571_x12_1 ( // @[Math.scala 150:24:@25036.4]
    .io_a(x571_x12_1_io_a),
    .io_b(x571_x12_1_io_b),
    .io_result(x571_x12_1_io_result)
  );
  x543_x11 x572_x11_1 ( // @[Math.scala 150:24:@25046.4]
    .io_a(x572_x11_1_io_a),
    .io_b(x572_x11_1_io_b),
    .io_result(x572_x11_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_76 ( // @[package.scala 93:22:@25056.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  x543_x11 x573_sum_1 ( // @[Math.scala 150:24:@25065.4]
    .io_a(x573_sum_1_io_a),
    .io_b(x573_sum_1_io_b),
    .io_result(x573_sum_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_77 ( // @[package.scala 93:22:@25079.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  x539_x11 x579_x11_1 ( // @[Math.scala 150:24:@25109.4]
    .clock(x579_x11_1_clock),
    .reset(x579_x11_1_reset),
    .io_a(x579_x11_1_io_a),
    .io_b(x579_x11_1_io_b),
    .io_flow(x579_x11_1_io_flow),
    .io_result(x579_x11_1_io_result)
  );
  x539_x11 x580_x12_1 ( // @[Math.scala 150:24:@25119.4]
    .clock(x580_x12_1_clock),
    .reset(x580_x12_1_reset),
    .io_a(x580_x12_1_io_a),
    .io_b(x580_x12_1_io_b),
    .io_flow(x580_x12_1_io_flow),
    .io_result(x580_x12_1_io_result)
  );
  x539_x11 x581_x11_1 ( // @[Math.scala 150:24:@25131.4]
    .clock(x581_x11_1_clock),
    .reset(x581_x11_1_reset),
    .io_a(x581_x11_1_io_a),
    .io_b(x581_x11_1_io_b),
    .io_flow(x581_x11_1_io_flow),
    .io_result(x581_x11_1_io_result)
  );
  x539_x11 x582_x12_1 ( // @[Math.scala 150:24:@25141.4]
    .clock(x582_x12_1_clock),
    .reset(x582_x12_1_reset),
    .io_a(x582_x12_1_io_a),
    .io_b(x582_x12_1_io_b),
    .io_flow(x582_x12_1_io_flow),
    .io_result(x582_x12_1_io_result)
  );
  x543_x11 x583_x11_1 ( // @[Math.scala 150:24:@25151.4]
    .io_a(x583_x11_1_io_a),
    .io_b(x583_x11_1_io_b),
    .io_result(x583_x11_1_io_result)
  );
  x543_x11 x584_x12_1 ( // @[Math.scala 150:24:@25161.4]
    .io_a(x584_x12_1_io_a),
    .io_b(x584_x12_1_io_b),
    .io_result(x584_x12_1_io_result)
  );
  x543_x11 x585_x11_1 ( // @[Math.scala 150:24:@25171.4]
    .io_a(x585_x11_1_io_a),
    .io_b(x585_x11_1_io_b),
    .io_result(x585_x11_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_78 ( // @[package.scala 93:22:@25181.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  x543_x11 x586_sum_1 ( // @[Math.scala 150:24:@25190.4]
    .io_a(x586_sum_1_io_a),
    .io_b(x586_sum_1_io_b),
    .io_result(x586_sum_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_79 ( // @[package.scala 93:22:@25204.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper_128 RetimeWrapper_80 ( // @[package.scala 93:22:@25224.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  RetimeWrapper_12 RetimeWrapper_81 ( // @[package.scala 93:22:@25233.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_12 RetimeWrapper_82 ( // @[package.scala 93:22:@25242.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  RetimeWrapper_12 RetimeWrapper_83 ( // @[package.scala 93:22:@25251.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  assign b327 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 62:18:@22814.4]
  assign b328 = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 63:18:@22815.4]
  assign _T_206 = b327 & b328; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 68:30:@22962.4]
  assign _T_207 = _T_206 & io_sigsIn_datapathEn; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 68:37:@22963.4]
  assign _T_211 = io_in_x316_TID == 8'h0; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 70:76:@22968.4]
  assign _T_212 = _T_207 & _T_211; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 70:62:@22969.4]
  assign _T_214 = io_in_x316_TDEST == 8'h0; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 70:101:@22970.4]
  assign x667_x330_D1_0_number = RetimeWrapper_io_out; // @[package.scala 96:25:@22979.4 package.scala 96:25:@22980.4]
  assign b325_number = __io_result; // @[Math.scala 712:22:@22799.4 Math.scala 713:14:@22800.4]
  assign _T_246 = $signed(b325_number); // @[Math.scala 499:52:@22999.4]
  assign x334 = $signed(32'sh1) == $signed(_T_246); // @[Math.scala 499:44:@23007.4]
  assign x335 = $signed(32'sh2) == $signed(_T_246); // @[Math.scala 499:44:@23014.4]
  assign x336 = $signed(32'sh3) == $signed(_T_246); // @[Math.scala 499:44:@23021.4]
  assign _T_293 = x334 ? 32'h1 : 32'h0; // @[Mux.scala 19:72:@23033.4]
  assign _T_295 = x335 ? 32'h2 : 32'h0; // @[Mux.scala 19:72:@23034.4]
  assign _T_297 = x336 ? 32'h3 : 32'h0; // @[Mux.scala 19:72:@23035.4]
  assign _T_299 = _T_293 | _T_295; // @[Mux.scala 19:72:@23037.4]
  assign x337_number = _T_299 | _T_297; // @[Mux.scala 19:72:@23038.4]
  assign _T_311 = $signed(x337_number); // @[Math.scala 406:49:@23048.4]
  assign _T_313 = $signed(_T_311) & $signed(32'sh3); // @[Math.scala 406:56:@23050.4]
  assign _T_314 = $signed(_T_313); // @[Math.scala 406:56:@23051.4]
  assign _T_319 = x337_number[31]; // @[FixedPoint.scala 50:25:@23057.4]
  assign _T_323 = _T_319 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@23059.4]
  assign _T_324 = x337_number[31:2]; // @[FixedPoint.scala 18:52:@23060.4]
  assign b326_number = __1_io_result; // @[Math.scala 712:22:@22811.4 Math.scala 713:14:@22812.4]
  assign _T_329 = b326_number[31]; // @[FixedPoint.scala 50:25:@23066.4]
  assign _T_333 = _T_329 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@23068.4]
  assign _T_334 = b326_number[31:2]; // @[FixedPoint.scala 18:52:@23069.4]
  assign _T_359 = ~ io_sigsIn_break; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 113:101:@23130.4]
  assign _T_363 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@23138.4 package.scala 96:25:@23139.4]
  assign _T_365 = io_rr ? _T_363 : 1'h0; // @[implicits.scala 55:10:@23140.4]
  assign _T_366 = _T_359 & _T_365; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 113:118:@23141.4]
  assign _T_368 = _T_366 & _T_359; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 113:205:@23143.4]
  assign _T_369 = _T_368 & io_sigsIn_backpressure; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 113:224:@23144.4]
  assign x671_b327_D4 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@23116.4 package.scala 96:25:@23117.4]
  assign _T_370 = _T_369 & x671_b327_D4; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 113:250:@23145.4]
  assign x669_b328_D4 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@23098.4 package.scala 96:25:@23099.4]
  assign x349_rdcol_number = x349_rdcol_1_io_result; // @[Math.scala 154:22:@23162.4 Math.scala 155:14:@23163.4]
  assign _T_383 = x349_rdcol_number[31]; // @[FixedPoint.scala 50:25:@23169.4]
  assign _T_387 = _T_383 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@23171.4]
  assign _T_388 = x349_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@23172.4]
  assign _T_411 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@23223.4 package.scala 96:25:@23224.4]
  assign _T_413 = io_rr ? _T_411 : 1'h0; // @[implicits.scala 55:10:@23225.4]
  assign _T_414 = _T_359 & _T_413; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 132:118:@23226.4]
  assign _T_416 = _T_414 & _T_359; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 132:205:@23228.4]
  assign _T_417 = _T_416 & io_sigsIn_backpressure; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 132:224:@23229.4]
  assign _T_418 = _T_417 & x671_b327_D4; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 132:250:@23230.4]
  assign x358_rdcol_number = x358_rdcol_1_io_result; // @[Math.scala 154:22:@23247.4 Math.scala 155:14:@23248.4]
  assign _T_431 = x358_rdcol_number[31]; // @[FixedPoint.scala 50:25:@23254.4]
  assign _T_435 = _T_431 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@23256.4]
  assign _T_436 = x358_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@23257.4]
  assign _T_456 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@23299.4 package.scala 96:25:@23300.4]
  assign _T_458 = io_rr ? _T_456 : 1'h0; // @[implicits.scala 55:10:@23301.4]
  assign _T_459 = _T_359 & _T_458; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 149:118:@23302.4]
  assign _T_461 = _T_459 & _T_359; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 149:205:@23304.4]
  assign _T_462 = _T_461 & io_sigsIn_backpressure; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 149:224:@23305.4]
  assign _T_463 = _T_462 & x671_b327_D4; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 149:250:@23306.4]
  assign x367_rdcol_number = x367_rdcol_1_io_result; // @[Math.scala 154:22:@23323.4 Math.scala 155:14:@23324.4]
  assign _T_476 = x367_rdcol_number[31]; // @[FixedPoint.scala 50:25:@23330.4]
  assign _T_480 = _T_476 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@23332.4]
  assign _T_481 = x367_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@23333.4]
  assign _T_501 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@23375.4 package.scala 96:25:@23376.4]
  assign _T_503 = io_rr ? _T_501 : 1'h0; // @[implicits.scala 55:10:@23377.4]
  assign _T_504 = _T_359 & _T_503; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 166:118:@23378.4]
  assign _T_506 = _T_504 & _T_359; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 166:205:@23380.4]
  assign _T_507 = _T_506 & io_sigsIn_backpressure; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 166:224:@23381.4]
  assign _T_508 = _T_507 & x671_b327_D4; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 166:250:@23382.4]
  assign x680_b325_D6_number = RetimeWrapper_17_io_out; // @[package.scala 96:25:@23396.4 package.scala 96:25:@23397.4]
  assign _T_520 = $signed(x680_b325_D6_number); // @[Math.scala 406:49:@23403.4]
  assign _T_522 = $signed(_T_520) & $signed(32'sh3); // @[Math.scala 406:56:@23405.4]
  assign _T_523 = $signed(_T_522); // @[Math.scala 406:56:@23406.4]
  assign x661_number = $unsigned(_T_523); // @[implicits.scala 133:21:@23407.4]
  assign x378 = $signed(_T_520) < $signed(32'sh0); // @[Math.scala 465:44:@23415.4]
  assign x681_x367_rdcol_D6_number = RetimeWrapper_18_io_out; // @[package.scala 96:25:@23423.4 package.scala 96:25:@23424.4]
  assign _T_541 = $signed(x681_x367_rdcol_D6_number); // @[Math.scala 465:37:@23429.4]
  assign x379 = $signed(_T_541) < $signed(32'sh0); // @[Math.scala 465:44:@23431.4]
  assign x682_x378_D1 = RetimeWrapper_19_io_out; // @[package.scala 96:25:@23439.4 package.scala 96:25:@23440.4]
  assign x380 = x682_x378_D1 | x379; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 187:24:@23443.4]
  assign _T_560 = $signed(x661_number); // @[Math.scala 406:49:@23454.4]
  assign _T_562 = $signed(_T_560) & $signed(32'sh3); // @[Math.scala 406:56:@23456.4]
  assign _T_563 = $signed(_T_562); // @[Math.scala 406:56:@23457.4]
  assign _T_568 = x661_number[31]; // @[FixedPoint.scala 50:25:@23463.4]
  assign _T_572 = _T_568 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@23465.4]
  assign _T_573 = x661_number[31:2]; // @[FixedPoint.scala 18:52:@23466.4]
  assign _T_611 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@23545.4 package.scala 96:25:@23546.4]
  assign _T_613 = io_rr ? _T_611 : 1'h0; // @[implicits.scala 55:10:@23547.4]
  assign _T_614 = _T_359 & _T_613; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 214:194:@23548.4]
  assign x685_x381_D1 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@23504.4 package.scala 96:25:@23505.4]
  assign _T_615 = _T_614 & x685_x381_D1; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 214:281:@23549.4]
  assign x688_b327_D8 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@23531.4 package.scala 96:25:@23532.4]
  assign _T_616 = _T_615 & x688_b327_D8; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 214:289:@23550.4]
  assign x686_b328_D8 = RetimeWrapper_23_io_out; // @[package.scala 96:25:@23513.4 package.scala 96:25:@23514.4]
  assign x689_x358_rdcol_D6_number = RetimeWrapper_27_io_out; // @[package.scala 96:25:@23566.4 package.scala 96:25:@23567.4]
  assign _T_627 = $signed(x689_x358_rdcol_D6_number); // @[Math.scala 465:37:@23572.4]
  assign x390 = $signed(_T_627) < $signed(32'sh0); // @[Math.scala 465:44:@23574.4]
  assign x391 = x682_x378_D1 | x390; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 222:24:@23577.4]
  assign _T_658 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@23621.4 package.scala 96:25:@23622.4]
  assign _T_660 = io_rr ? _T_658 : 1'h0; // @[implicits.scala 55:10:@23623.4]
  assign _T_661 = _T_359 & _T_660; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 235:194:@23624.4]
  assign x691_x392_D1 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@23607.4 package.scala 96:25:@23608.4]
  assign _T_662 = _T_661 & x691_x392_D1; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 235:281:@23625.4]
  assign _T_663 = _T_662 & x688_b327_D8; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 235:289:@23626.4]
  assign x692_x349_rdcol_D6_number = RetimeWrapper_31_io_out; // @[package.scala 96:25:@23642.4 package.scala 96:25:@23643.4]
  assign _T_674 = $signed(x692_x349_rdcol_D6_number); // @[Math.scala 465:37:@23648.4]
  assign x398 = $signed(_T_674) < $signed(32'sh0); // @[Math.scala 465:44:@23650.4]
  assign x399 = x682_x378_D1 | x398; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 243:24:@23653.4]
  assign _T_705 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@23697.4 package.scala 96:25:@23698.4]
  assign _T_707 = io_rr ? _T_705 : 1'h0; // @[implicits.scala 55:10:@23699.4]
  assign _T_708 = _T_359 & _T_707; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 256:194:@23700.4]
  assign x694_x400_D1 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@23683.4 package.scala 96:25:@23684.4]
  assign _T_709 = _T_708 & x694_x400_D1; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 256:281:@23701.4]
  assign _T_710 = _T_709 & x688_b327_D8; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 256:289:@23702.4]
  assign x695_b326_D6_number = RetimeWrapper_35_io_out; // @[package.scala 96:25:@23718.4 package.scala 96:25:@23719.4]
  assign _T_721 = $signed(x695_b326_D6_number); // @[Math.scala 465:37:@23724.4]
  assign x406 = $signed(_T_721) < $signed(32'sh0); // @[Math.scala 465:44:@23726.4]
  assign x407 = x378 | x406; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 264:59:@23729.4]
  assign _T_755 = RetimeWrapper_39_io_out; // @[package.scala 96:25:@23782.4 package.scala 96:25:@23783.4]
  assign _T_757 = io_rr ? _T_755 : 1'h0; // @[implicits.scala 55:10:@23784.4]
  assign _T_758 = _T_359 & _T_757; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 279:194:@23785.4]
  assign x697_x408_D2 = RetimeWrapper_37_io_out; // @[package.scala 96:25:@23759.4 package.scala 96:25:@23760.4]
  assign _T_759 = _T_758 & x697_x408_D2; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 279:281:@23786.4]
  assign _T_760 = _T_759 & x688_b327_D8; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 279:289:@23787.4]
  assign x414_rdcol_number = x414_rdcol_1_io_result; // @[Math.scala 154:22:@23806.4 Math.scala 155:14:@23807.4]
  assign _T_775 = $signed(x414_rdcol_number); // @[Math.scala 465:37:@23812.4]
  assign x415 = $signed(_T_775) < $signed(32'sh0); // @[Math.scala 465:44:@23814.4]
  assign x416 = x682_x378_D1 | x415; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 287:24:@23817.4]
  assign _T_785 = x414_rdcol_number[31]; // @[FixedPoint.scala 50:25:@23824.4]
  assign _T_789 = _T_785 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@23826.4]
  assign _T_790 = x414_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@23827.4]
  assign _T_813 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@23861.4 package.scala 96:25:@23862.4]
  assign _T_815 = io_rr ? _T_813 : 1'h0; // @[implicits.scala 55:10:@23863.4]
  assign _T_816 = _T_359 & _T_815; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 306:194:@23864.4]
  assign x699_x417_D1 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@23847.4 package.scala 96:25:@23848.4]
  assign _T_817 = _T_816 & x699_x417_D1; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 306:281:@23865.4]
  assign _T_818 = _T_817 & x688_b327_D8; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 306:324:@23866.4]
  assign x426_rdcol_number = x426_rdcol_1_io_result; // @[Math.scala 154:22:@23887.4 Math.scala 155:14:@23888.4]
  assign _T_835 = $signed(x426_rdcol_number); // @[Math.scala 465:37:@23893.4]
  assign x427 = $signed(_T_835) < $signed(32'sh0); // @[Math.scala 465:44:@23895.4]
  assign x428 = x682_x378_D1 | x427; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 316:59:@23898.4]
  assign _T_845 = x426_rdcol_number[31]; // @[FixedPoint.scala 50:25:@23905.4]
  assign _T_849 = _T_845 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@23907.4]
  assign _T_850 = x426_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@23908.4]
  assign _T_873 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@23942.4 package.scala 96:25:@23943.4]
  assign _T_875 = io_rr ? _T_873 : 1'h0; // @[implicits.scala 55:10:@23944.4]
  assign _T_876 = _T_359 & _T_875; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 329:194:@23945.4]
  assign x700_x429_D1 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@23928.4 package.scala 96:25:@23929.4]
  assign _T_877 = _T_876 & x700_x429_D1; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 329:281:@23946.4]
  assign _T_878 = _T_877 & x688_b327_D8; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 329:289:@23947.4]
  assign x438_rdrow_number = x438_rdrow_1_io_result; // @[Math.scala 195:22:@23966.4 Math.scala 196:14:@23967.4]
  assign _T_895 = $signed(x438_rdrow_number); // @[Math.scala 406:49:@23973.4]
  assign _T_897 = $signed(_T_895) & $signed(32'sh3); // @[Math.scala 406:56:@23975.4]
  assign _T_898 = $signed(_T_897); // @[Math.scala 406:56:@23976.4]
  assign x663_number = $unsigned(_T_898); // @[implicits.scala 133:21:@23977.4]
  assign x440 = $signed(_T_895) < $signed(32'sh0); // @[Math.scala 465:44:@23985.4]
  assign x441 = x440 | x379; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 339:24:@23988.4]
  assign _T_919 = $signed(x663_number); // @[Math.scala 406:49:@23997.4]
  assign _T_921 = $signed(_T_919) & $signed(32'sh3); // @[Math.scala 406:56:@23999.4]
  assign _T_922 = $signed(_T_921); // @[Math.scala 406:56:@24000.4]
  assign _T_927 = x663_number[31]; // @[FixedPoint.scala 50:25:@24006.4]
  assign _T_931 = _T_927 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@24008.4]
  assign _T_932 = x663_number[31:2]; // @[FixedPoint.scala 18:52:@24009.4]
  assign _T_958 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@24052.4 package.scala 96:25:@24053.4]
  assign _T_960 = io_rr ? _T_958 : 1'h0; // @[implicits.scala 55:10:@24054.4]
  assign _T_961 = _T_359 & _T_960; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 356:194:@24055.4]
  assign x702_x442_D1 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@24038.4 package.scala 96:25:@24039.4]
  assign _T_962 = _T_961 & x702_x442_D1; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 356:281:@24056.4]
  assign _T_963 = _T_962 & x688_b327_D8; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 356:289:@24057.4]
  assign x451 = x440 | x390; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 360:24:@24068.4]
  assign _T_991 = RetimeWrapper_48_io_out; // @[package.scala 96:25:@24103.4 package.scala 96:25:@24104.4]
  assign _T_993 = io_rr ? _T_991 : 1'h0; // @[implicits.scala 55:10:@24105.4]
  assign _T_994 = _T_359 & _T_993; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 371:194:@24106.4]
  assign x703_x452_D1 = RetimeWrapper_47_io_out; // @[package.scala 96:25:@24089.4 package.scala 96:25:@24090.4]
  assign _T_995 = _T_994 & x703_x452_D1; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 371:281:@24107.4]
  assign _T_996 = _T_995 & x688_b327_D8; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 371:289:@24108.4]
  assign x458 = x440 | x398; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 375:24:@24119.4]
  assign _T_1024 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@24154.4 package.scala 96:25:@24155.4]
  assign _T_1026 = io_rr ? _T_1024 : 1'h0; // @[implicits.scala 55:10:@24156.4]
  assign _T_1027 = _T_359 & _T_1026; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 386:194:@24157.4]
  assign x704_x459_D1 = RetimeWrapper_49_io_out; // @[package.scala 96:25:@24140.4 package.scala 96:25:@24141.4]
  assign _T_1028 = _T_1027 & x704_x459_D1; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 386:281:@24158.4]
  assign _T_1029 = _T_1028 & x688_b327_D8; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 386:289:@24159.4]
  assign x705_x406_D1 = RetimeWrapper_51_io_out; // @[package.scala 96:25:@24175.4 package.scala 96:25:@24176.4]
  assign x465 = x440 | x705_x406_D1; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 392:24:@24179.4]
  assign _T_1063 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@24223.4 package.scala 96:25:@24224.4]
  assign _T_1065 = io_rr ? _T_1063 : 1'h0; // @[implicits.scala 55:10:@24225.4]
  assign _T_1066 = _T_359 & _T_1065; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 405:194:@24226.4]
  assign x707_x466_D1 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@24209.4 package.scala 96:25:@24210.4]
  assign _T_1067 = _T_1066 & x707_x466_D1; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 405:281:@24227.4]
  assign _T_1068 = _T_1067 & x688_b327_D8; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 405:289:@24228.4]
  assign x472 = x440 | x415; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 409:24:@24239.4]
  assign _T_1096 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@24274.4 package.scala 96:25:@24275.4]
  assign _T_1098 = io_rr ? _T_1096 : 1'h0; // @[implicits.scala 55:10:@24276.4]
  assign _T_1099 = _T_359 & _T_1098; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 420:194:@24277.4]
  assign x708_x473_D1 = RetimeWrapper_55_io_out; // @[package.scala 96:25:@24260.4 package.scala 96:25:@24261.4]
  assign _T_1100 = _T_1099 & x708_x473_D1; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 420:281:@24278.4]
  assign _T_1101 = _T_1100 & x688_b327_D8; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 420:289:@24279.4]
  assign x479 = x440 | x427; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 430:59:@24290.4]
  assign _T_1131 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@24327.4 package.scala 96:25:@24328.4]
  assign _T_1133 = io_rr ? _T_1131 : 1'h0; // @[implicits.scala 55:10:@24329.4]
  assign _T_1134 = _T_359 & _T_1133; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 443:194:@24330.4]
  assign x709_x480_D1 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@24313.4 package.scala 96:25:@24314.4]
  assign _T_1135 = _T_1134 & x709_x480_D1; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 443:281:@24331.4]
  assign _T_1136 = _T_1135 & x688_b327_D8; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 443:289:@24332.4]
  assign x486_rdrow_number = x486_rdrow_1_io_result; // @[Math.scala 195:22:@24351.4 Math.scala 196:14:@24352.4]
  assign _T_1153 = $signed(x486_rdrow_number); // @[Math.scala 406:49:@24358.4]
  assign _T_1155 = $signed(_T_1153) & $signed(32'sh3); // @[Math.scala 406:56:@24360.4]
  assign _T_1156 = $signed(_T_1155); // @[Math.scala 406:56:@24361.4]
  assign x665_number = $unsigned(_T_1156); // @[implicits.scala 133:21:@24362.4]
  assign x488 = $signed(_T_1153) < $signed(32'sh0); // @[Math.scala 465:44:@24370.4]
  assign x489 = x488 | x379; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 453:24:@24373.4]
  assign _T_1177 = $signed(x665_number); // @[Math.scala 406:49:@24382.4]
  assign _T_1179 = $signed(_T_1177) & $signed(32'sh3); // @[Math.scala 406:56:@24384.4]
  assign _T_1180 = $signed(_T_1179); // @[Math.scala 406:56:@24385.4]
  assign _T_1185 = x665_number[31]; // @[FixedPoint.scala 50:25:@24391.4]
  assign _T_1189 = _T_1185 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@24393.4]
  assign _T_1190 = x665_number[31:2]; // @[FixedPoint.scala 18:52:@24394.4]
  assign _T_1216 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@24437.4 package.scala 96:25:@24438.4]
  assign _T_1218 = io_rr ? _T_1216 : 1'h0; // @[implicits.scala 55:10:@24439.4]
  assign _T_1219 = _T_359 & _T_1218; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 470:194:@24440.4]
  assign x711_x490_D1 = RetimeWrapper_60_io_out; // @[package.scala 96:25:@24423.4 package.scala 96:25:@24424.4]
  assign _T_1220 = _T_1219 & x711_x490_D1; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 470:281:@24441.4]
  assign _T_1221 = _T_1220 & x688_b327_D8; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 470:289:@24442.4]
  assign x499 = x488 | x390; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 474:24:@24453.4]
  assign _T_1249 = RetimeWrapper_63_io_out; // @[package.scala 96:25:@24488.4 package.scala 96:25:@24489.4]
  assign _T_1251 = io_rr ? _T_1249 : 1'h0; // @[implicits.scala 55:10:@24490.4]
  assign _T_1252 = _T_359 & _T_1251; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 485:194:@24491.4]
  assign x712_x500_D1 = RetimeWrapper_62_io_out; // @[package.scala 96:25:@24474.4 package.scala 96:25:@24475.4]
  assign _T_1253 = _T_1252 & x712_x500_D1; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 485:281:@24492.4]
  assign _T_1254 = _T_1253 & x688_b327_D8; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 485:289:@24493.4]
  assign x506 = x488 | x398; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 489:24:@24504.4]
  assign _T_1282 = RetimeWrapper_65_io_out; // @[package.scala 96:25:@24539.4 package.scala 96:25:@24540.4]
  assign _T_1284 = io_rr ? _T_1282 : 1'h0; // @[implicits.scala 55:10:@24541.4]
  assign _T_1285 = _T_359 & _T_1284; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 500:194:@24542.4]
  assign x713_x507_D1 = RetimeWrapper_64_io_out; // @[package.scala 96:25:@24525.4 package.scala 96:25:@24526.4]
  assign _T_1286 = _T_1285 & x713_x507_D1; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 500:281:@24543.4]
  assign _T_1287 = _T_1286 & x688_b327_D8; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 500:289:@24544.4]
  assign x513 = x488 | x705_x406_D1; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 504:24:@24555.4]
  assign _T_1315 = RetimeWrapper_67_io_out; // @[package.scala 96:25:@24590.4 package.scala 96:25:@24591.4]
  assign _T_1317 = io_rr ? _T_1315 : 1'h0; // @[implicits.scala 55:10:@24592.4]
  assign _T_1318 = _T_359 & _T_1317; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 515:194:@24593.4]
  assign x714_x514_D1 = RetimeWrapper_66_io_out; // @[package.scala 96:25:@24576.4 package.scala 96:25:@24577.4]
  assign _T_1319 = _T_1318 & x714_x514_D1; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 515:281:@24594.4]
  assign _T_1320 = _T_1319 & x688_b327_D8; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 515:289:@24595.4]
  assign x520 = x488 | x415; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 519:24:@24606.4]
  assign _T_1348 = RetimeWrapper_69_io_out; // @[package.scala 96:25:@24641.4 package.scala 96:25:@24642.4]
  assign _T_1350 = io_rr ? _T_1348 : 1'h0; // @[implicits.scala 55:10:@24643.4]
  assign _T_1351 = _T_359 & _T_1350; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 530:194:@24644.4]
  assign x715_x521_D1 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@24627.4 package.scala 96:25:@24628.4]
  assign _T_1352 = _T_1351 & x715_x521_D1; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 530:281:@24645.4]
  assign _T_1353 = _T_1352 & x688_b327_D8; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 530:289:@24646.4]
  assign x527 = x488 | x427; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 534:24:@24657.4]
  assign _T_1381 = RetimeWrapper_71_io_out; // @[package.scala 96:25:@24692.4 package.scala 96:25:@24693.4]
  assign _T_1383 = io_rr ? _T_1381 : 1'h0; // @[implicits.scala 55:10:@24694.4]
  assign _T_1384 = _T_359 & _T_1383; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 545:194:@24695.4]
  assign x716_x528_D1 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@24678.4 package.scala 96:25:@24679.4]
  assign _T_1385 = _T_1384 & x716_x528_D1; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 545:281:@24696.4]
  assign _T_1386 = _T_1385 & x688_b327_D8; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 545:289:@24697.4]
  assign x396_rd_0_number = x329_lb_0_io_rPort_6_output_0; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 231:29:@23610.4 sm_x592_inr_Foreach_SAMPLER_BOX.scala 235:336:@23633.4]
  assign _GEN_0 = {{1'd0}, x396_rd_0_number}; // @[Math.scala 450:32:@24709.4]
  assign _T_1392 = _GEN_0 << 1; // @[Math.scala 450:32:@24709.4]
  assign x449_rd_0_number = x329_lb_0_io_rPort_1_output_0; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 352:29:@24041.4 sm_x592_inr_Foreach_SAMPLER_BOX.scala 356:406:@24064.4]
  assign _GEN_1 = {{1'd0}, x449_rd_0_number}; // @[Math.scala 450:32:@24716.4]
  assign _T_1398 = _GEN_1 << 1; // @[Math.scala 450:32:@24716.4]
  assign x456_rd_0_number = x329_lb_0_io_rPort_9_output_0; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 367:29:@24092.4 sm_x592_inr_Foreach_SAMPLER_BOX.scala 371:406:@24115.4]
  assign _GEN_2 = {{2'd0}, x456_rd_0_number}; // @[Math.scala 450:32:@24721.4]
  assign _T_1402 = _GEN_2 << 2; // @[Math.scala 450:32:@24721.4]
  assign x463_rd_0_number = x329_lb_0_io_rPort_14_output_0; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 382:29:@24143.4 sm_x592_inr_Foreach_SAMPLER_BOX.scala 386:406:@24166.4]
  assign _GEN_3 = {{1'd0}, x463_rd_0_number}; // @[Math.scala 450:32:@24726.4]
  assign _T_1406 = _GEN_3 << 1; // @[Math.scala 450:32:@24726.4]
  assign x504_rd_0_number = x329_lb_0_io_rPort_5_output_0; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 481:29:@24477.4 sm_x592_inr_Foreach_SAMPLER_BOX.scala 485:406:@24500.4]
  assign _GEN_4 = {{1'd0}, x504_rd_0_number}; // @[Math.scala 450:32:@24731.4]
  assign _T_1410 = _GEN_4 << 1; // @[Math.scala 450:32:@24731.4]
  assign x546_sum_number = x546_sum_1_io_result; // @[Math.scala 154:22:@24820.4 Math.scala 155:14:@24821.4]
  assign _T_1446 = x546_sum_number[7:4]; // @[FixedPoint.scala 18:52:@24826.4]
  assign x404_rd_0_number = x329_lb_0_io_rPort_3_output_0; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 252:29:@23686.4 sm_x592_inr_Foreach_SAMPLER_BOX.scala 256:336:@23709.4]
  assign _GEN_5 = {{1'd0}, x404_rd_0_number}; // @[Math.scala 450:32:@24839.4]
  assign _T_1453 = _GEN_5 << 1; // @[Math.scala 450:32:@24839.4]
  assign _GEN_6 = {{1'd0}, x456_rd_0_number}; // @[Math.scala 450:32:@24844.4]
  assign _T_1457 = _GEN_6 << 1; // @[Math.scala 450:32:@24844.4]
  assign _GEN_7 = {{2'd0}, x463_rd_0_number}; // @[Math.scala 450:32:@24849.4]
  assign _T_1461 = _GEN_7 << 2; // @[Math.scala 450:32:@24849.4]
  assign x470_rd_0_number = x329_lb_0_io_rPort_15_output_0; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 401:29:@24212.4 sm_x592_inr_Foreach_SAMPLER_BOX.scala 405:406:@24235.4]
  assign _GEN_8 = {{1'd0}, x470_rd_0_number}; // @[Math.scala 450:32:@24854.4]
  assign _T_1465 = _GEN_8 << 1; // @[Math.scala 450:32:@24854.4]
  assign x511_rd_0_number = x329_lb_0_io_rPort_2_output_0; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 496:29:@24528.4 sm_x592_inr_Foreach_SAMPLER_BOX.scala 500:406:@24551.4]
  assign _GEN_9 = {{1'd0}, x511_rd_0_number}; // @[Math.scala 450:32:@24859.4]
  assign _T_1469 = _GEN_9 << 1; // @[Math.scala 450:32:@24859.4]
  assign x560_sum_number = x560_sum_1_io_result; // @[Math.scala 154:22:@24948.4 Math.scala 155:14:@24949.4]
  assign _T_1505 = x560_sum_number[7:4]; // @[FixedPoint.scala 18:52:@24954.4]
  assign x412_rd_0_number = x329_lb_0_io_rPort_11_output_0; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 275:29:@23771.4 sm_x592_inr_Foreach_SAMPLER_BOX.scala 279:336:@23794.4]
  assign _GEN_10 = {{1'd0}, x412_rd_0_number}; // @[Math.scala 450:32:@24967.4]
  assign _T_1512 = _GEN_10 << 1; // @[Math.scala 450:32:@24967.4]
  assign _GEN_11 = {{2'd0}, x470_rd_0_number}; // @[Math.scala 450:32:@24972.4]
  assign _T_1516 = _GEN_11 << 2; // @[Math.scala 450:32:@24972.4]
  assign x477_rd_0_number = x329_lb_0_io_rPort_12_output_0; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 416:29:@24263.4 sm_x592_inr_Foreach_SAMPLER_BOX.scala 420:406:@24286.4]
  assign _GEN_12 = {{1'd0}, x477_rd_0_number}; // @[Math.scala 450:32:@24977.4]
  assign _T_1520 = _GEN_12 << 1; // @[Math.scala 450:32:@24977.4]
  assign x518_rd_0_number = x329_lb_0_io_rPort_0_output_0; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 511:29:@24579.4 sm_x592_inr_Foreach_SAMPLER_BOX.scala 515:406:@24602.4]
  assign _GEN_13 = {{1'd0}, x518_rd_0_number}; // @[Math.scala 450:32:@24982.4]
  assign _T_1524 = _GEN_13 << 1; // @[Math.scala 450:32:@24982.4]
  assign x573_sum_number = x573_sum_1_io_result; // @[Math.scala 154:22:@25071.4 Math.scala 155:14:@25072.4]
  assign _T_1560 = x573_sum_number[7:4]; // @[FixedPoint.scala 18:52:@25077.4]
  assign x424_rd_0_number = x329_lb_0_io_rPort_7_output_0; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 302:29:@23850.4 sm_x592_inr_Foreach_SAMPLER_BOX.scala 306:441:@23873.4]
  assign _GEN_14 = {{1'd0}, x424_rd_0_number}; // @[Math.scala 450:32:@25090.4]
  assign _T_1567 = _GEN_14 << 1; // @[Math.scala 450:32:@25090.4]
  assign _GEN_15 = {{2'd0}, x477_rd_0_number}; // @[Math.scala 450:32:@25095.4]
  assign _T_1571 = _GEN_15 << 2; // @[Math.scala 450:32:@25095.4]
  assign x484_rd_0_number = x329_lb_0_io_rPort_8_output_0; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 439:29:@24316.4 sm_x592_inr_Foreach_SAMPLER_BOX.scala 443:406:@24339.4]
  assign _GEN_16 = {{1'd0}, x484_rd_0_number}; // @[Math.scala 450:32:@25100.4]
  assign _T_1575 = _GEN_16 << 1; // @[Math.scala 450:32:@25100.4]
  assign x525_rd_0_number = x329_lb_0_io_rPort_13_output_0; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 526:29:@24630.4 sm_x592_inr_Foreach_SAMPLER_BOX.scala 530:406:@24653.4]
  assign _GEN_17 = {{1'd0}, x525_rd_0_number}; // @[Math.scala 450:32:@25105.4]
  assign _T_1579 = _GEN_17 << 1; // @[Math.scala 450:32:@25105.4]
  assign x586_sum_number = x586_sum_1_io_result; // @[Math.scala 154:22:@25196.4 Math.scala 155:14:@25197.4]
  assign _T_1617 = x586_sum_number[7:4]; // @[FixedPoint.scala 18:52:@25202.4]
  assign x574_number = RetimeWrapper_77_io_out; // @[package.scala 96:25:@25084.4 package.scala 96:25:@25085.4]
  assign x587_number = RetimeWrapper_79_io_out; // @[package.scala 96:25:@25209.4 package.scala 96:25:@25210.4]
  assign _T_1632 = {x574_number,x587_number}; // @[Cat.scala 30:58:@25219.4]
  assign x547_number = RetimeWrapper_73_io_out; // @[package.scala 96:25:@24833.4 package.scala 96:25:@24834.4]
  assign x561_number = RetimeWrapper_75_io_out; // @[package.scala 96:25:@24961.4 package.scala 96:25:@24962.4]
  assign _T_1633 = {x547_number,x561_number}; // @[Cat.scala 30:58:@25220.4]
  assign _T_1646 = RetimeWrapper_83_io_out; // @[package.scala 96:25:@25256.4 package.scala 96:25:@25257.4]
  assign _T_1648 = io_rr ? _T_1646 : 1'h0; // @[implicits.scala 55:10:@25258.4]
  assign x721_b327_D15 = RetimeWrapper_81_io_out; // @[package.scala 96:25:@25238.4 package.scala 96:25:@25239.4]
  assign _T_1649 = _T_1648 & x721_b327_D15; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 689:116:@25259.4]
  assign x722_b328_D15 = RetimeWrapper_82_io_out; // @[package.scala 96:25:@25247.4 package.scala 96:25:@25248.4]
  assign _T_1650 = _T_1649 & x722_b328_D15; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 689:122:@25260.4]
  assign x668_x660_D4_number = RetimeWrapper_1_io_out; // @[package.scala 96:25:@23089.4 package.scala 96:25:@23090.4]
  assign x670_x343_sum_D3_number = RetimeWrapper_3_io_out; // @[package.scala 96:25:@23107.4 package.scala 96:25:@23108.4]
  assign x674_x353_sum_D2_number = RetimeWrapper_8_io_out; // @[package.scala 96:25:@23201.4 package.scala 96:25:@23202.4]
  assign x676_x362_sum_D2_number = RetimeWrapper_11_io_out; // @[package.scala 96:25:@23277.4 package.scala 96:25:@23278.4]
  assign x678_x371_sum_D2_number = RetimeWrapper_14_io_out; // @[package.scala 96:25:@23353.4 package.scala 96:25:@23354.4]
  assign x384_sum_number = x384_sum_1_io_result; // @[Math.scala 154:22:@23495.4 Math.scala 155:14:@23496.4]
  assign x687_x662_D2_number = RetimeWrapper_24_io_out; // @[package.scala 96:25:@23522.4 package.scala 96:25:@23523.4]
  assign x393_sum_number = x393_sum_1_io_result; // @[Math.scala 154:22:@23598.4 Math.scala 155:14:@23599.4]
  assign x401_sum_number = x401_sum_1_io_result; // @[Math.scala 154:22:@23674.4 Math.scala 155:14:@23675.4]
  assign x698_x409_sum_D1_number = RetimeWrapper_38_io_out; // @[package.scala 96:25:@23768.4 package.scala 96:25:@23769.4]
  assign x420_sum_number = x420_sum_1_io_result; // @[Math.scala 154:22:@23838.4 Math.scala 155:14:@23839.4]
  assign x432_sum_number = x432_sum_1_io_result; // @[Math.scala 154:22:@23919.4 Math.scala 155:14:@23920.4]
  assign x445_sum_number = x445_sum_1_io_result; // @[Math.scala 154:22:@24020.4 Math.scala 155:14:@24021.4]
  assign x701_x664_D1_number = RetimeWrapper_44_io_out; // @[package.scala 96:25:@24029.4 package.scala 96:25:@24030.4]
  assign x453_sum_number = x453_sum_1_io_result; // @[Math.scala 154:22:@24080.4 Math.scala 155:14:@24081.4]
  assign x460_sum_number = x460_sum_1_io_result; // @[Math.scala 154:22:@24131.4 Math.scala 155:14:@24132.4]
  assign x467_sum_number = x467_sum_1_io_result; // @[Math.scala 154:22:@24200.4 Math.scala 155:14:@24201.4]
  assign x474_sum_number = x474_sum_1_io_result; // @[Math.scala 154:22:@24251.4 Math.scala 155:14:@24252.4]
  assign x481_sum_number = x481_sum_1_io_result; // @[Math.scala 154:22:@24304.4 Math.scala 155:14:@24305.4]
  assign x493_sum_number = x493_sum_1_io_result; // @[Math.scala 154:22:@24405.4 Math.scala 155:14:@24406.4]
  assign x710_x666_D1_number = RetimeWrapper_59_io_out; // @[package.scala 96:25:@24414.4 package.scala 96:25:@24415.4]
  assign x501_sum_number = x501_sum_1_io_result; // @[Math.scala 154:22:@24465.4 Math.scala 155:14:@24466.4]
  assign x508_sum_number = x508_sum_1_io_result; // @[Math.scala 154:22:@24516.4 Math.scala 155:14:@24517.4]
  assign x515_sum_number = x515_sum_1_io_result; // @[Math.scala 154:22:@24567.4 Math.scala 155:14:@24568.4]
  assign x522_sum_number = x522_sum_1_io_result; // @[Math.scala 154:22:@24618.4 Math.scala 155:14:@24619.4]
  assign x529_sum_number = x529_sum_1_io_result; // @[Math.scala 154:22:@24669.4 Math.scala 155:14:@24670.4]
  assign io_in_x316_TREADY = _T_212 & _T_214; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 68:22:@22964.4 sm_x592_inr_Foreach_SAMPLER_BOX.scala 70:22:@22972.4]
  assign io_in_x317_TVALID = _T_1650 & io_sigsIn_backpressure; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 689:22:@25262.4]
  assign io_in_x317_TDATA = {{224'd0}, RetimeWrapper_80_io_out}; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 690:24:@25263.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 710:17:@22797.4]
  assign __1_io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_1); // @[Math.scala 710:17:@22809.4]
  assign x329_lb_0_clock = clock; // @[:@22817.4]
  assign x329_lb_0_reset = reset; // @[:@22818.4]
  assign x329_lb_0_io_rPort_17_banks_0 = x710_x666_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@24699.4]
  assign x329_lb_0_io_rPort_17_ofs_0 = x529_sum_number[0]; // @[MemInterfaceType.scala 107:54:@24701.4]
  assign x329_lb_0_io_rPort_17_en_0 = _T_1386 & x686_b328_D8; // @[MemInterfaceType.scala 110:79:@24703.4]
  assign x329_lb_0_io_rPort_17_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@24702.4]
  assign x329_lb_0_io_rPort_16_banks_0 = x710_x666_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@24444.4]
  assign x329_lb_0_io_rPort_16_ofs_0 = x493_sum_number[0]; // @[MemInterfaceType.scala 107:54:@24446.4]
  assign x329_lb_0_io_rPort_16_en_0 = _T_1221 & x686_b328_D8; // @[MemInterfaceType.scala 110:79:@24448.4]
  assign x329_lb_0_io_rPort_16_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@24447.4]
  assign x329_lb_0_io_rPort_15_banks_0 = x701_x664_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@24230.4]
  assign x329_lb_0_io_rPort_15_ofs_0 = x467_sum_number[0]; // @[MemInterfaceType.scala 107:54:@24232.4]
  assign x329_lb_0_io_rPort_15_en_0 = _T_1068 & x686_b328_D8; // @[MemInterfaceType.scala 110:79:@24234.4]
  assign x329_lb_0_io_rPort_15_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@24233.4]
  assign x329_lb_0_io_rPort_14_banks_0 = x701_x664_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@24161.4]
  assign x329_lb_0_io_rPort_14_ofs_0 = x460_sum_number[0]; // @[MemInterfaceType.scala 107:54:@24163.4]
  assign x329_lb_0_io_rPort_14_en_0 = _T_1029 & x686_b328_D8; // @[MemInterfaceType.scala 110:79:@24165.4]
  assign x329_lb_0_io_rPort_14_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@24164.4]
  assign x329_lb_0_io_rPort_13_banks_0 = x710_x666_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@24648.4]
  assign x329_lb_0_io_rPort_13_ofs_0 = x522_sum_number[0]; // @[MemInterfaceType.scala 107:54:@24650.4]
  assign x329_lb_0_io_rPort_13_en_0 = _T_1353 & x686_b328_D8; // @[MemInterfaceType.scala 110:79:@24652.4]
  assign x329_lb_0_io_rPort_13_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@24651.4]
  assign x329_lb_0_io_rPort_12_banks_0 = x701_x664_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@24281.4]
  assign x329_lb_0_io_rPort_12_ofs_0 = x474_sum_number[0]; // @[MemInterfaceType.scala 107:54:@24283.4]
  assign x329_lb_0_io_rPort_12_en_0 = _T_1101 & x686_b328_D8; // @[MemInterfaceType.scala 110:79:@24285.4]
  assign x329_lb_0_io_rPort_12_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@24284.4]
  assign x329_lb_0_io_rPort_11_banks_0 = x687_x662_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@23789.4]
  assign x329_lb_0_io_rPort_11_ofs_0 = x698_x409_sum_D1_number[0]; // @[MemInterfaceType.scala 107:54:@23791.4]
  assign x329_lb_0_io_rPort_11_en_0 = _T_760 & x686_b328_D8; // @[MemInterfaceType.scala 110:79:@23793.4]
  assign x329_lb_0_io_rPort_11_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@23792.4]
  assign x329_lb_0_io_rPort_10_banks_0 = x687_x662_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@23552.4]
  assign x329_lb_0_io_rPort_10_ofs_0 = x384_sum_number[0]; // @[MemInterfaceType.scala 107:54:@23554.4]
  assign x329_lb_0_io_rPort_10_en_0 = _T_616 & x686_b328_D8; // @[MemInterfaceType.scala 110:79:@23556.4]
  assign x329_lb_0_io_rPort_10_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@23555.4]
  assign x329_lb_0_io_rPort_9_banks_0 = x701_x664_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@24110.4]
  assign x329_lb_0_io_rPort_9_ofs_0 = x453_sum_number[0]; // @[MemInterfaceType.scala 107:54:@24112.4]
  assign x329_lb_0_io_rPort_9_en_0 = _T_996 & x686_b328_D8; // @[MemInterfaceType.scala 110:79:@24114.4]
  assign x329_lb_0_io_rPort_9_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@24113.4]
  assign x329_lb_0_io_rPort_8_banks_0 = x701_x664_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@24334.4]
  assign x329_lb_0_io_rPort_8_ofs_0 = x481_sum_number[0]; // @[MemInterfaceType.scala 107:54:@24336.4]
  assign x329_lb_0_io_rPort_8_en_0 = _T_1136 & x686_b328_D8; // @[MemInterfaceType.scala 110:79:@24338.4]
  assign x329_lb_0_io_rPort_8_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@24337.4]
  assign x329_lb_0_io_rPort_7_banks_0 = x687_x662_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@23868.4]
  assign x329_lb_0_io_rPort_7_ofs_0 = x420_sum_number[0]; // @[MemInterfaceType.scala 107:54:@23870.4]
  assign x329_lb_0_io_rPort_7_en_0 = _T_818 & x686_b328_D8; // @[MemInterfaceType.scala 110:79:@23872.4]
  assign x329_lb_0_io_rPort_7_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@23871.4]
  assign x329_lb_0_io_rPort_6_banks_0 = x687_x662_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@23628.4]
  assign x329_lb_0_io_rPort_6_ofs_0 = x393_sum_number[0]; // @[MemInterfaceType.scala 107:54:@23630.4]
  assign x329_lb_0_io_rPort_6_en_0 = _T_663 & x686_b328_D8; // @[MemInterfaceType.scala 110:79:@23632.4]
  assign x329_lb_0_io_rPort_6_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@23631.4]
  assign x329_lb_0_io_rPort_5_banks_0 = x710_x666_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@24495.4]
  assign x329_lb_0_io_rPort_5_ofs_0 = x501_sum_number[0]; // @[MemInterfaceType.scala 107:54:@24497.4]
  assign x329_lb_0_io_rPort_5_en_0 = _T_1254 & x686_b328_D8; // @[MemInterfaceType.scala 110:79:@24499.4]
  assign x329_lb_0_io_rPort_5_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@24498.4]
  assign x329_lb_0_io_rPort_4_banks_0 = x687_x662_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@23949.4]
  assign x329_lb_0_io_rPort_4_ofs_0 = x432_sum_number[0]; // @[MemInterfaceType.scala 107:54:@23951.4]
  assign x329_lb_0_io_rPort_4_en_0 = _T_878 & x686_b328_D8; // @[MemInterfaceType.scala 110:79:@23953.4]
  assign x329_lb_0_io_rPort_4_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@23952.4]
  assign x329_lb_0_io_rPort_3_banks_0 = x687_x662_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@23704.4]
  assign x329_lb_0_io_rPort_3_ofs_0 = x401_sum_number[0]; // @[MemInterfaceType.scala 107:54:@23706.4]
  assign x329_lb_0_io_rPort_3_en_0 = _T_710 & x686_b328_D8; // @[MemInterfaceType.scala 110:79:@23708.4]
  assign x329_lb_0_io_rPort_3_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@23707.4]
  assign x329_lb_0_io_rPort_2_banks_0 = x710_x666_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@24546.4]
  assign x329_lb_0_io_rPort_2_ofs_0 = x508_sum_number[0]; // @[MemInterfaceType.scala 107:54:@24548.4]
  assign x329_lb_0_io_rPort_2_en_0 = _T_1287 & x686_b328_D8; // @[MemInterfaceType.scala 110:79:@24550.4]
  assign x329_lb_0_io_rPort_2_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@24549.4]
  assign x329_lb_0_io_rPort_1_banks_0 = x701_x664_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@24059.4]
  assign x329_lb_0_io_rPort_1_ofs_0 = x445_sum_number[0]; // @[MemInterfaceType.scala 107:54:@24061.4]
  assign x329_lb_0_io_rPort_1_en_0 = _T_963 & x686_b328_D8; // @[MemInterfaceType.scala 110:79:@24063.4]
  assign x329_lb_0_io_rPort_1_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@24062.4]
  assign x329_lb_0_io_rPort_0_banks_0 = x710_x666_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@24597.4]
  assign x329_lb_0_io_rPort_0_ofs_0 = x515_sum_number[0]; // @[MemInterfaceType.scala 107:54:@24599.4]
  assign x329_lb_0_io_rPort_0_en_0 = _T_1320 & x686_b328_D8; // @[MemInterfaceType.scala 110:79:@24601.4]
  assign x329_lb_0_io_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@24600.4]
  assign x329_lb_0_io_wPort_3_banks_0 = x668_x660_D4_number[2:0]; // @[MemInterfaceType.scala 88:58:@23384.4]
  assign x329_lb_0_io_wPort_3_ofs_0 = x678_x371_sum_D2_number[0]; // @[MemInterfaceType.scala 89:54:@23386.4]
  assign x329_lb_0_io_wPort_3_data_0 = RetimeWrapper_15_io_out; // @[MemInterfaceType.scala 90:56:@23387.4]
  assign x329_lb_0_io_wPort_3_en_0 = _T_508 & x669_b328_D4; // @[MemInterfaceType.scala 93:57:@23389.4]
  assign x329_lb_0_io_wPort_2_banks_0 = x668_x660_D4_number[2:0]; // @[MemInterfaceType.scala 88:58:@23308.4]
  assign x329_lb_0_io_wPort_2_ofs_0 = x676_x362_sum_D2_number[0]; // @[MemInterfaceType.scala 89:54:@23310.4]
  assign x329_lb_0_io_wPort_2_data_0 = RetimeWrapper_12_io_out; // @[MemInterfaceType.scala 90:56:@23311.4]
  assign x329_lb_0_io_wPort_2_en_0 = _T_463 & x669_b328_D4; // @[MemInterfaceType.scala 93:57:@23313.4]
  assign x329_lb_0_io_wPort_1_banks_0 = x668_x660_D4_number[2:0]; // @[MemInterfaceType.scala 88:58:@23232.4]
  assign x329_lb_0_io_wPort_1_ofs_0 = x674_x353_sum_D2_number[0]; // @[MemInterfaceType.scala 89:54:@23234.4]
  assign x329_lb_0_io_wPort_1_data_0 = RetimeWrapper_9_io_out; // @[MemInterfaceType.scala 90:56:@23235.4]
  assign x329_lb_0_io_wPort_1_en_0 = _T_418 & x669_b328_D4; // @[MemInterfaceType.scala 93:57:@23237.4]
  assign x329_lb_0_io_wPort_0_banks_0 = x668_x660_D4_number[2:0]; // @[MemInterfaceType.scala 88:58:@23147.4]
  assign x329_lb_0_io_wPort_0_ofs_0 = x670_x343_sum_D3_number[0]; // @[MemInterfaceType.scala 89:54:@23149.4]
  assign x329_lb_0_io_wPort_0_data_0 = RetimeWrapper_5_io_out; // @[MemInterfaceType.scala 90:56:@23150.4]
  assign x329_lb_0_io_wPort_0_en_0 = _T_370 & x669_b328_D4; // @[MemInterfaceType.scala 93:57:@23152.4]
  assign RetimeWrapper_clock = clock; // @[:@22975.4]
  assign RetimeWrapper_reset = reset; // @[:@22976.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22978.4]
  assign RetimeWrapper_io_in = io_in_x316_TDATA[31:0]; // @[package.scala 94:16:@22977.4]
  assign x343_sum_1_clock = clock; // @[:@23075.4]
  assign x343_sum_1_reset = reset; // @[:@23076.4]
  assign x343_sum_1_io_a = {_T_323,_T_324}; // @[Math.scala 151:17:@23077.4]
  assign x343_sum_1_io_b = {_T_333,_T_334}; // @[Math.scala 152:17:@23078.4]
  assign x343_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@23079.4]
  assign RetimeWrapper_1_clock = clock; // @[:@23085.4]
  assign RetimeWrapper_1_reset = reset; // @[:@23086.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@23088.4]
  assign RetimeWrapper_1_io_in = $unsigned(_T_314); // @[package.scala 94:16:@23087.4]
  assign RetimeWrapper_2_clock = clock; // @[:@23094.4]
  assign RetimeWrapper_2_reset = reset; // @[:@23095.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@23097.4]
  assign RetimeWrapper_2_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@23096.4]
  assign RetimeWrapper_3_clock = clock; // @[:@23103.4]
  assign RetimeWrapper_3_reset = reset; // @[:@23104.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@23106.4]
  assign RetimeWrapper_3_io_in = x343_sum_1_io_result; // @[package.scala 94:16:@23105.4]
  assign RetimeWrapper_4_clock = clock; // @[:@23112.4]
  assign RetimeWrapper_4_reset = reset; // @[:@23113.4]
  assign RetimeWrapper_4_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@23115.4]
  assign RetimeWrapper_4_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@23114.4]
  assign RetimeWrapper_5_clock = clock; // @[:@23121.4]
  assign RetimeWrapper_5_reset = reset; // @[:@23122.4]
  assign RetimeWrapper_5_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@23124.4]
  assign RetimeWrapper_5_io_in = x667_x330_D1_0_number[7:0]; // @[package.scala 94:16:@23123.4]
  assign RetimeWrapper_6_clock = clock; // @[:@23134.4]
  assign RetimeWrapper_6_reset = reset; // @[:@23135.4]
  assign RetimeWrapper_6_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@23137.4]
  assign RetimeWrapper_6_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@23136.4]
  assign x349_rdcol_1_clock = clock; // @[:@23157.4]
  assign x349_rdcol_1_reset = reset; // @[:@23158.4]
  assign x349_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@23159.4]
  assign x349_rdcol_1_io_b = 32'h1; // @[Math.scala 152:17:@23160.4]
  assign x349_rdcol_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@23161.4]
  assign RetimeWrapper_7_clock = clock; // @[:@23178.4]
  assign RetimeWrapper_7_reset = reset; // @[:@23179.4]
  assign RetimeWrapper_7_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@23181.4]
  assign RetimeWrapper_7_io_in = {_T_323,_T_324}; // @[package.scala 94:16:@23180.4]
  assign x353_sum_1_clock = clock; // @[:@23187.4]
  assign x353_sum_1_reset = reset; // @[:@23188.4]
  assign x353_sum_1_io_a = RetimeWrapper_7_io_out; // @[Math.scala 151:17:@23189.4]
  assign x353_sum_1_io_b = {_T_387,_T_388}; // @[Math.scala 152:17:@23190.4]
  assign x353_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@23191.4]
  assign RetimeWrapper_8_clock = clock; // @[:@23197.4]
  assign RetimeWrapper_8_reset = reset; // @[:@23198.4]
  assign RetimeWrapper_8_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@23200.4]
  assign RetimeWrapper_8_io_in = x353_sum_1_io_result; // @[package.scala 94:16:@23199.4]
  assign RetimeWrapper_9_clock = clock; // @[:@23206.4]
  assign RetimeWrapper_9_reset = reset; // @[:@23207.4]
  assign RetimeWrapper_9_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@23209.4]
  assign RetimeWrapper_9_io_in = x667_x330_D1_0_number[15:8]; // @[package.scala 94:16:@23208.4]
  assign RetimeWrapper_10_clock = clock; // @[:@23219.4]
  assign RetimeWrapper_10_reset = reset; // @[:@23220.4]
  assign RetimeWrapper_10_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@23222.4]
  assign RetimeWrapper_10_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@23221.4]
  assign x358_rdcol_1_clock = clock; // @[:@23242.4]
  assign x358_rdcol_1_reset = reset; // @[:@23243.4]
  assign x358_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@23244.4]
  assign x358_rdcol_1_io_b = 32'h2; // @[Math.scala 152:17:@23245.4]
  assign x358_rdcol_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@23246.4]
  assign x362_sum_1_clock = clock; // @[:@23263.4]
  assign x362_sum_1_reset = reset; // @[:@23264.4]
  assign x362_sum_1_io_a = RetimeWrapper_7_io_out; // @[Math.scala 151:17:@23265.4]
  assign x362_sum_1_io_b = {_T_435,_T_436}; // @[Math.scala 152:17:@23266.4]
  assign x362_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@23267.4]
  assign RetimeWrapper_11_clock = clock; // @[:@23273.4]
  assign RetimeWrapper_11_reset = reset; // @[:@23274.4]
  assign RetimeWrapper_11_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@23276.4]
  assign RetimeWrapper_11_io_in = x362_sum_1_io_result; // @[package.scala 94:16:@23275.4]
  assign RetimeWrapper_12_clock = clock; // @[:@23282.4]
  assign RetimeWrapper_12_reset = reset; // @[:@23283.4]
  assign RetimeWrapper_12_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@23285.4]
  assign RetimeWrapper_12_io_in = x667_x330_D1_0_number[23:16]; // @[package.scala 94:16:@23284.4]
  assign RetimeWrapper_13_clock = clock; // @[:@23295.4]
  assign RetimeWrapper_13_reset = reset; // @[:@23296.4]
  assign RetimeWrapper_13_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@23298.4]
  assign RetimeWrapper_13_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@23297.4]
  assign x367_rdcol_1_clock = clock; // @[:@23318.4]
  assign x367_rdcol_1_reset = reset; // @[:@23319.4]
  assign x367_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@23320.4]
  assign x367_rdcol_1_io_b = 32'h3; // @[Math.scala 152:17:@23321.4]
  assign x367_rdcol_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@23322.4]
  assign x371_sum_1_clock = clock; // @[:@23339.4]
  assign x371_sum_1_reset = reset; // @[:@23340.4]
  assign x371_sum_1_io_a = RetimeWrapper_7_io_out; // @[Math.scala 151:17:@23341.4]
  assign x371_sum_1_io_b = {_T_480,_T_481}; // @[Math.scala 152:17:@23342.4]
  assign x371_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@23343.4]
  assign RetimeWrapper_14_clock = clock; // @[:@23349.4]
  assign RetimeWrapper_14_reset = reset; // @[:@23350.4]
  assign RetimeWrapper_14_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@23352.4]
  assign RetimeWrapper_14_io_in = x371_sum_1_io_result; // @[package.scala 94:16:@23351.4]
  assign RetimeWrapper_15_clock = clock; // @[:@23358.4]
  assign RetimeWrapper_15_reset = reset; // @[:@23359.4]
  assign RetimeWrapper_15_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@23361.4]
  assign RetimeWrapper_15_io_in = x667_x330_D1_0_number[31:24]; // @[package.scala 94:16:@23360.4]
  assign RetimeWrapper_16_clock = clock; // @[:@23371.4]
  assign RetimeWrapper_16_reset = reset; // @[:@23372.4]
  assign RetimeWrapper_16_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@23374.4]
  assign RetimeWrapper_16_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@23373.4]
  assign RetimeWrapper_17_clock = clock; // @[:@23392.4]
  assign RetimeWrapper_17_reset = reset; // @[:@23393.4]
  assign RetimeWrapper_17_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@23395.4]
  assign RetimeWrapper_17_io_in = __io_result; // @[package.scala 94:16:@23394.4]
  assign RetimeWrapper_18_clock = clock; // @[:@23419.4]
  assign RetimeWrapper_18_reset = reset; // @[:@23420.4]
  assign RetimeWrapper_18_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@23422.4]
  assign RetimeWrapper_18_io_in = x367_rdcol_1_io_result; // @[package.scala 94:16:@23421.4]
  assign RetimeWrapper_19_clock = clock; // @[:@23435.4]
  assign RetimeWrapper_19_reset = reset; // @[:@23436.4]
  assign RetimeWrapper_19_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@23438.4]
  assign RetimeWrapper_19_io_in = $signed(_T_520) < $signed(32'sh0); // @[package.scala 94:16:@23437.4]
  assign RetimeWrapper_20_clock = clock; // @[:@23472.4]
  assign RetimeWrapper_20_reset = reset; // @[:@23473.4]
  assign RetimeWrapper_20_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@23475.4]
  assign RetimeWrapper_20_io_in = {_T_572,_T_573}; // @[package.scala 94:16:@23474.4]
  assign RetimeWrapper_21_clock = clock; // @[:@23481.4]
  assign RetimeWrapper_21_reset = reset; // @[:@23482.4]
  assign RetimeWrapper_21_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@23484.4]
  assign RetimeWrapper_21_io_in = {_T_480,_T_481}; // @[package.scala 94:16:@23483.4]
  assign x384_sum_1_clock = clock; // @[:@23490.4]
  assign x384_sum_1_reset = reset; // @[:@23491.4]
  assign x384_sum_1_io_a = RetimeWrapper_20_io_out; // @[Math.scala 151:17:@23492.4]
  assign x384_sum_1_io_b = RetimeWrapper_21_io_out; // @[Math.scala 152:17:@23493.4]
  assign x384_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@23494.4]
  assign RetimeWrapper_22_clock = clock; // @[:@23500.4]
  assign RetimeWrapper_22_reset = reset; // @[:@23501.4]
  assign RetimeWrapper_22_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@23503.4]
  assign RetimeWrapper_22_io_in = ~ x380; // @[package.scala 94:16:@23502.4]
  assign RetimeWrapper_23_clock = clock; // @[:@23509.4]
  assign RetimeWrapper_23_reset = reset; // @[:@23510.4]
  assign RetimeWrapper_23_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@23512.4]
  assign RetimeWrapper_23_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@23511.4]
  assign RetimeWrapper_24_clock = clock; // @[:@23518.4]
  assign RetimeWrapper_24_reset = reset; // @[:@23519.4]
  assign RetimeWrapper_24_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@23521.4]
  assign RetimeWrapper_24_io_in = $unsigned(_T_563); // @[package.scala 94:16:@23520.4]
  assign RetimeWrapper_25_clock = clock; // @[:@23527.4]
  assign RetimeWrapper_25_reset = reset; // @[:@23528.4]
  assign RetimeWrapper_25_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@23530.4]
  assign RetimeWrapper_25_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@23529.4]
  assign RetimeWrapper_26_clock = clock; // @[:@23541.4]
  assign RetimeWrapper_26_reset = reset; // @[:@23542.4]
  assign RetimeWrapper_26_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@23544.4]
  assign RetimeWrapper_26_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@23543.4]
  assign RetimeWrapper_27_clock = clock; // @[:@23562.4]
  assign RetimeWrapper_27_reset = reset; // @[:@23563.4]
  assign RetimeWrapper_27_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@23565.4]
  assign RetimeWrapper_27_io_in = x358_rdcol_1_io_result; // @[package.scala 94:16:@23564.4]
  assign RetimeWrapper_28_clock = clock; // @[:@23584.4]
  assign RetimeWrapper_28_reset = reset; // @[:@23585.4]
  assign RetimeWrapper_28_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@23587.4]
  assign RetimeWrapper_28_io_in = {_T_435,_T_436}; // @[package.scala 94:16:@23586.4]
  assign x393_sum_1_clock = clock; // @[:@23593.4]
  assign x393_sum_1_reset = reset; // @[:@23594.4]
  assign x393_sum_1_io_a = RetimeWrapper_20_io_out; // @[Math.scala 151:17:@23595.4]
  assign x393_sum_1_io_b = RetimeWrapper_28_io_out; // @[Math.scala 152:17:@23596.4]
  assign x393_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@23597.4]
  assign RetimeWrapper_29_clock = clock; // @[:@23603.4]
  assign RetimeWrapper_29_reset = reset; // @[:@23604.4]
  assign RetimeWrapper_29_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@23606.4]
  assign RetimeWrapper_29_io_in = ~ x391; // @[package.scala 94:16:@23605.4]
  assign RetimeWrapper_30_clock = clock; // @[:@23617.4]
  assign RetimeWrapper_30_reset = reset; // @[:@23618.4]
  assign RetimeWrapper_30_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@23620.4]
  assign RetimeWrapper_30_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@23619.4]
  assign RetimeWrapper_31_clock = clock; // @[:@23638.4]
  assign RetimeWrapper_31_reset = reset; // @[:@23639.4]
  assign RetimeWrapper_31_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@23641.4]
  assign RetimeWrapper_31_io_in = x349_rdcol_1_io_result; // @[package.scala 94:16:@23640.4]
  assign RetimeWrapper_32_clock = clock; // @[:@23660.4]
  assign RetimeWrapper_32_reset = reset; // @[:@23661.4]
  assign RetimeWrapper_32_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@23663.4]
  assign RetimeWrapper_32_io_in = {_T_387,_T_388}; // @[package.scala 94:16:@23662.4]
  assign x401_sum_1_clock = clock; // @[:@23669.4]
  assign x401_sum_1_reset = reset; // @[:@23670.4]
  assign x401_sum_1_io_a = RetimeWrapper_20_io_out; // @[Math.scala 151:17:@23671.4]
  assign x401_sum_1_io_b = RetimeWrapper_32_io_out; // @[Math.scala 152:17:@23672.4]
  assign x401_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@23673.4]
  assign RetimeWrapper_33_clock = clock; // @[:@23679.4]
  assign RetimeWrapper_33_reset = reset; // @[:@23680.4]
  assign RetimeWrapper_33_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@23682.4]
  assign RetimeWrapper_33_io_in = ~ x399; // @[package.scala 94:16:@23681.4]
  assign RetimeWrapper_34_clock = clock; // @[:@23693.4]
  assign RetimeWrapper_34_reset = reset; // @[:@23694.4]
  assign RetimeWrapper_34_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@23696.4]
  assign RetimeWrapper_34_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@23695.4]
  assign RetimeWrapper_35_clock = clock; // @[:@23714.4]
  assign RetimeWrapper_35_reset = reset; // @[:@23715.4]
  assign RetimeWrapper_35_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@23717.4]
  assign RetimeWrapper_35_io_in = __1_io_result; // @[package.scala 94:16:@23716.4]
  assign RetimeWrapper_36_clock = clock; // @[:@23736.4]
  assign RetimeWrapper_36_reset = reset; // @[:@23737.4]
  assign RetimeWrapper_36_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@23739.4]
  assign RetimeWrapper_36_io_in = {_T_333,_T_334}; // @[package.scala 94:16:@23738.4]
  assign x409_sum_1_clock = clock; // @[:@23745.4]
  assign x409_sum_1_reset = reset; // @[:@23746.4]
  assign x409_sum_1_io_a = {_T_572,_T_573}; // @[Math.scala 151:17:@23747.4]
  assign x409_sum_1_io_b = RetimeWrapper_36_io_out; // @[Math.scala 152:17:@23748.4]
  assign x409_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@23749.4]
  assign RetimeWrapper_37_clock = clock; // @[:@23755.4]
  assign RetimeWrapper_37_reset = reset; // @[:@23756.4]
  assign RetimeWrapper_37_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@23758.4]
  assign RetimeWrapper_37_io_in = ~ x407; // @[package.scala 94:16:@23757.4]
  assign RetimeWrapper_38_clock = clock; // @[:@23764.4]
  assign RetimeWrapper_38_reset = reset; // @[:@23765.4]
  assign RetimeWrapper_38_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@23767.4]
  assign RetimeWrapper_38_io_in = x409_sum_1_io_result; // @[package.scala 94:16:@23766.4]
  assign RetimeWrapper_39_clock = clock; // @[:@23778.4]
  assign RetimeWrapper_39_reset = reset; // @[:@23779.4]
  assign RetimeWrapper_39_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@23781.4]
  assign RetimeWrapper_39_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@23780.4]
  assign x414_rdcol_1_clock = clock; // @[:@23801.4]
  assign x414_rdcol_1_reset = reset; // @[:@23802.4]
  assign x414_rdcol_1_io_a = RetimeWrapper_35_io_out; // @[Math.scala 151:17:@23803.4]
  assign x414_rdcol_1_io_b = 32'hffffffff; // @[Math.scala 152:17:@23804.4]
  assign x414_rdcol_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@23805.4]
  assign x420_sum_1_clock = clock; // @[:@23833.4]
  assign x420_sum_1_reset = reset; // @[:@23834.4]
  assign x420_sum_1_io_a = RetimeWrapper_20_io_out; // @[Math.scala 151:17:@23835.4]
  assign x420_sum_1_io_b = {_T_789,_T_790}; // @[Math.scala 152:17:@23836.4]
  assign x420_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@23837.4]
  assign RetimeWrapper_40_clock = clock; // @[:@23843.4]
  assign RetimeWrapper_40_reset = reset; // @[:@23844.4]
  assign RetimeWrapper_40_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@23846.4]
  assign RetimeWrapper_40_io_in = ~ x416; // @[package.scala 94:16:@23845.4]
  assign RetimeWrapper_41_clock = clock; // @[:@23857.4]
  assign RetimeWrapper_41_reset = reset; // @[:@23858.4]
  assign RetimeWrapper_41_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@23860.4]
  assign RetimeWrapper_41_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@23859.4]
  assign x426_rdcol_1_clock = clock; // @[:@23882.4]
  assign x426_rdcol_1_reset = reset; // @[:@23883.4]
  assign x426_rdcol_1_io_a = RetimeWrapper_35_io_out; // @[Math.scala 151:17:@23884.4]
  assign x426_rdcol_1_io_b = 32'hfffffffe; // @[Math.scala 152:17:@23885.4]
  assign x426_rdcol_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@23886.4]
  assign x432_sum_1_clock = clock; // @[:@23914.4]
  assign x432_sum_1_reset = reset; // @[:@23915.4]
  assign x432_sum_1_io_a = RetimeWrapper_20_io_out; // @[Math.scala 151:17:@23916.4]
  assign x432_sum_1_io_b = {_T_849,_T_850}; // @[Math.scala 152:17:@23917.4]
  assign x432_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@23918.4]
  assign RetimeWrapper_42_clock = clock; // @[:@23924.4]
  assign RetimeWrapper_42_reset = reset; // @[:@23925.4]
  assign RetimeWrapper_42_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@23927.4]
  assign RetimeWrapper_42_io_in = ~ x428; // @[package.scala 94:16:@23926.4]
  assign RetimeWrapper_43_clock = clock; // @[:@23938.4]
  assign RetimeWrapper_43_reset = reset; // @[:@23939.4]
  assign RetimeWrapper_43_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@23941.4]
  assign RetimeWrapper_43_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@23940.4]
  assign x438_rdrow_1_clock = clock; // @[:@23961.4]
  assign x438_rdrow_1_reset = reset; // @[:@23962.4]
  assign x438_rdrow_1_io_a = RetimeWrapper_17_io_out; // @[Math.scala 192:17:@23963.4]
  assign x438_rdrow_1_io_b = 32'h1; // @[Math.scala 193:17:@23964.4]
  assign x438_rdrow_1_io_flow = io_in_x317_TREADY; // @[Math.scala 194:20:@23965.4]
  assign x445_sum_1_clock = clock; // @[:@24015.4]
  assign x445_sum_1_reset = reset; // @[:@24016.4]
  assign x445_sum_1_io_a = {_T_931,_T_932}; // @[Math.scala 151:17:@24017.4]
  assign x445_sum_1_io_b = RetimeWrapper_21_io_out; // @[Math.scala 152:17:@24018.4]
  assign x445_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@24019.4]
  assign RetimeWrapper_44_clock = clock; // @[:@24025.4]
  assign RetimeWrapper_44_reset = reset; // @[:@24026.4]
  assign RetimeWrapper_44_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24028.4]
  assign RetimeWrapper_44_io_in = $unsigned(_T_922); // @[package.scala 94:16:@24027.4]
  assign RetimeWrapper_45_clock = clock; // @[:@24034.4]
  assign RetimeWrapper_45_reset = reset; // @[:@24035.4]
  assign RetimeWrapper_45_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24037.4]
  assign RetimeWrapper_45_io_in = ~ x441; // @[package.scala 94:16:@24036.4]
  assign RetimeWrapper_46_clock = clock; // @[:@24048.4]
  assign RetimeWrapper_46_reset = reset; // @[:@24049.4]
  assign RetimeWrapper_46_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24051.4]
  assign RetimeWrapper_46_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@24050.4]
  assign x453_sum_1_clock = clock; // @[:@24075.4]
  assign x453_sum_1_reset = reset; // @[:@24076.4]
  assign x453_sum_1_io_a = {_T_931,_T_932}; // @[Math.scala 151:17:@24077.4]
  assign x453_sum_1_io_b = RetimeWrapper_28_io_out; // @[Math.scala 152:17:@24078.4]
  assign x453_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@24079.4]
  assign RetimeWrapper_47_clock = clock; // @[:@24085.4]
  assign RetimeWrapper_47_reset = reset; // @[:@24086.4]
  assign RetimeWrapper_47_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24088.4]
  assign RetimeWrapper_47_io_in = ~ x451; // @[package.scala 94:16:@24087.4]
  assign RetimeWrapper_48_clock = clock; // @[:@24099.4]
  assign RetimeWrapper_48_reset = reset; // @[:@24100.4]
  assign RetimeWrapper_48_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24102.4]
  assign RetimeWrapper_48_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@24101.4]
  assign x460_sum_1_clock = clock; // @[:@24126.4]
  assign x460_sum_1_reset = reset; // @[:@24127.4]
  assign x460_sum_1_io_a = {_T_931,_T_932}; // @[Math.scala 151:17:@24128.4]
  assign x460_sum_1_io_b = RetimeWrapper_32_io_out; // @[Math.scala 152:17:@24129.4]
  assign x460_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@24130.4]
  assign RetimeWrapper_49_clock = clock; // @[:@24136.4]
  assign RetimeWrapper_49_reset = reset; // @[:@24137.4]
  assign RetimeWrapper_49_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24139.4]
  assign RetimeWrapper_49_io_in = ~ x458; // @[package.scala 94:16:@24138.4]
  assign RetimeWrapper_50_clock = clock; // @[:@24150.4]
  assign RetimeWrapper_50_reset = reset; // @[:@24151.4]
  assign RetimeWrapper_50_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24153.4]
  assign RetimeWrapper_50_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@24152.4]
  assign RetimeWrapper_51_clock = clock; // @[:@24171.4]
  assign RetimeWrapper_51_reset = reset; // @[:@24172.4]
  assign RetimeWrapper_51_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24174.4]
  assign RetimeWrapper_51_io_in = $signed(_T_721) < $signed(32'sh0); // @[package.scala 94:16:@24173.4]
  assign RetimeWrapper_52_clock = clock; // @[:@24186.4]
  assign RetimeWrapper_52_reset = reset; // @[:@24187.4]
  assign RetimeWrapper_52_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24189.4]
  assign RetimeWrapper_52_io_in = {_T_333,_T_334}; // @[package.scala 94:16:@24188.4]
  assign x467_sum_1_clock = clock; // @[:@24195.4]
  assign x467_sum_1_reset = reset; // @[:@24196.4]
  assign x467_sum_1_io_a = {_T_931,_T_932}; // @[Math.scala 151:17:@24197.4]
  assign x467_sum_1_io_b = RetimeWrapper_52_io_out; // @[Math.scala 152:17:@24198.4]
  assign x467_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@24199.4]
  assign RetimeWrapper_53_clock = clock; // @[:@24205.4]
  assign RetimeWrapper_53_reset = reset; // @[:@24206.4]
  assign RetimeWrapper_53_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24208.4]
  assign RetimeWrapper_53_io_in = ~ x465; // @[package.scala 94:16:@24207.4]
  assign RetimeWrapper_54_clock = clock; // @[:@24219.4]
  assign RetimeWrapper_54_reset = reset; // @[:@24220.4]
  assign RetimeWrapper_54_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24222.4]
  assign RetimeWrapper_54_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@24221.4]
  assign x474_sum_1_clock = clock; // @[:@24246.4]
  assign x474_sum_1_reset = reset; // @[:@24247.4]
  assign x474_sum_1_io_a = {_T_931,_T_932}; // @[Math.scala 151:17:@24248.4]
  assign x474_sum_1_io_b = {_T_789,_T_790}; // @[Math.scala 152:17:@24249.4]
  assign x474_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@24250.4]
  assign RetimeWrapper_55_clock = clock; // @[:@24256.4]
  assign RetimeWrapper_55_reset = reset; // @[:@24257.4]
  assign RetimeWrapper_55_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24259.4]
  assign RetimeWrapper_55_io_in = ~ x472; // @[package.scala 94:16:@24258.4]
  assign RetimeWrapper_56_clock = clock; // @[:@24270.4]
  assign RetimeWrapper_56_reset = reset; // @[:@24271.4]
  assign RetimeWrapper_56_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24273.4]
  assign RetimeWrapper_56_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@24272.4]
  assign x481_sum_1_clock = clock; // @[:@24299.4]
  assign x481_sum_1_reset = reset; // @[:@24300.4]
  assign x481_sum_1_io_a = {_T_931,_T_932}; // @[Math.scala 151:17:@24301.4]
  assign x481_sum_1_io_b = {_T_849,_T_850}; // @[Math.scala 152:17:@24302.4]
  assign x481_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@24303.4]
  assign RetimeWrapper_57_clock = clock; // @[:@24309.4]
  assign RetimeWrapper_57_reset = reset; // @[:@24310.4]
  assign RetimeWrapper_57_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24312.4]
  assign RetimeWrapper_57_io_in = ~ x479; // @[package.scala 94:16:@24311.4]
  assign RetimeWrapper_58_clock = clock; // @[:@24323.4]
  assign RetimeWrapper_58_reset = reset; // @[:@24324.4]
  assign RetimeWrapper_58_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24326.4]
  assign RetimeWrapper_58_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@24325.4]
  assign x486_rdrow_1_clock = clock; // @[:@24346.4]
  assign x486_rdrow_1_reset = reset; // @[:@24347.4]
  assign x486_rdrow_1_io_a = RetimeWrapper_17_io_out; // @[Math.scala 192:17:@24348.4]
  assign x486_rdrow_1_io_b = 32'h2; // @[Math.scala 193:17:@24349.4]
  assign x486_rdrow_1_io_flow = io_in_x317_TREADY; // @[Math.scala 194:20:@24350.4]
  assign x493_sum_1_clock = clock; // @[:@24400.4]
  assign x493_sum_1_reset = reset; // @[:@24401.4]
  assign x493_sum_1_io_a = {_T_1189,_T_1190}; // @[Math.scala 151:17:@24402.4]
  assign x493_sum_1_io_b = RetimeWrapper_21_io_out; // @[Math.scala 152:17:@24403.4]
  assign x493_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@24404.4]
  assign RetimeWrapper_59_clock = clock; // @[:@24410.4]
  assign RetimeWrapper_59_reset = reset; // @[:@24411.4]
  assign RetimeWrapper_59_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24413.4]
  assign RetimeWrapper_59_io_in = $unsigned(_T_1180); // @[package.scala 94:16:@24412.4]
  assign RetimeWrapper_60_clock = clock; // @[:@24419.4]
  assign RetimeWrapper_60_reset = reset; // @[:@24420.4]
  assign RetimeWrapper_60_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24422.4]
  assign RetimeWrapper_60_io_in = ~ x489; // @[package.scala 94:16:@24421.4]
  assign RetimeWrapper_61_clock = clock; // @[:@24433.4]
  assign RetimeWrapper_61_reset = reset; // @[:@24434.4]
  assign RetimeWrapper_61_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24436.4]
  assign RetimeWrapper_61_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@24435.4]
  assign x501_sum_1_clock = clock; // @[:@24460.4]
  assign x501_sum_1_reset = reset; // @[:@24461.4]
  assign x501_sum_1_io_a = {_T_1189,_T_1190}; // @[Math.scala 151:17:@24462.4]
  assign x501_sum_1_io_b = RetimeWrapper_28_io_out; // @[Math.scala 152:17:@24463.4]
  assign x501_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@24464.4]
  assign RetimeWrapper_62_clock = clock; // @[:@24470.4]
  assign RetimeWrapper_62_reset = reset; // @[:@24471.4]
  assign RetimeWrapper_62_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24473.4]
  assign RetimeWrapper_62_io_in = ~ x499; // @[package.scala 94:16:@24472.4]
  assign RetimeWrapper_63_clock = clock; // @[:@24484.4]
  assign RetimeWrapper_63_reset = reset; // @[:@24485.4]
  assign RetimeWrapper_63_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24487.4]
  assign RetimeWrapper_63_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@24486.4]
  assign x508_sum_1_clock = clock; // @[:@24511.4]
  assign x508_sum_1_reset = reset; // @[:@24512.4]
  assign x508_sum_1_io_a = {_T_1189,_T_1190}; // @[Math.scala 151:17:@24513.4]
  assign x508_sum_1_io_b = RetimeWrapper_32_io_out; // @[Math.scala 152:17:@24514.4]
  assign x508_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@24515.4]
  assign RetimeWrapper_64_clock = clock; // @[:@24521.4]
  assign RetimeWrapper_64_reset = reset; // @[:@24522.4]
  assign RetimeWrapper_64_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24524.4]
  assign RetimeWrapper_64_io_in = ~ x506; // @[package.scala 94:16:@24523.4]
  assign RetimeWrapper_65_clock = clock; // @[:@24535.4]
  assign RetimeWrapper_65_reset = reset; // @[:@24536.4]
  assign RetimeWrapper_65_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24538.4]
  assign RetimeWrapper_65_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@24537.4]
  assign x515_sum_1_clock = clock; // @[:@24562.4]
  assign x515_sum_1_reset = reset; // @[:@24563.4]
  assign x515_sum_1_io_a = {_T_1189,_T_1190}; // @[Math.scala 151:17:@24564.4]
  assign x515_sum_1_io_b = RetimeWrapper_52_io_out; // @[Math.scala 152:17:@24565.4]
  assign x515_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@24566.4]
  assign RetimeWrapper_66_clock = clock; // @[:@24572.4]
  assign RetimeWrapper_66_reset = reset; // @[:@24573.4]
  assign RetimeWrapper_66_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24575.4]
  assign RetimeWrapper_66_io_in = ~ x513; // @[package.scala 94:16:@24574.4]
  assign RetimeWrapper_67_clock = clock; // @[:@24586.4]
  assign RetimeWrapper_67_reset = reset; // @[:@24587.4]
  assign RetimeWrapper_67_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24589.4]
  assign RetimeWrapper_67_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@24588.4]
  assign x522_sum_1_clock = clock; // @[:@24613.4]
  assign x522_sum_1_reset = reset; // @[:@24614.4]
  assign x522_sum_1_io_a = {_T_1189,_T_1190}; // @[Math.scala 151:17:@24615.4]
  assign x522_sum_1_io_b = {_T_789,_T_790}; // @[Math.scala 152:17:@24616.4]
  assign x522_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@24617.4]
  assign RetimeWrapper_68_clock = clock; // @[:@24623.4]
  assign RetimeWrapper_68_reset = reset; // @[:@24624.4]
  assign RetimeWrapper_68_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24626.4]
  assign RetimeWrapper_68_io_in = ~ x520; // @[package.scala 94:16:@24625.4]
  assign RetimeWrapper_69_clock = clock; // @[:@24637.4]
  assign RetimeWrapper_69_reset = reset; // @[:@24638.4]
  assign RetimeWrapper_69_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24640.4]
  assign RetimeWrapper_69_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@24639.4]
  assign x529_sum_1_clock = clock; // @[:@24664.4]
  assign x529_sum_1_reset = reset; // @[:@24665.4]
  assign x529_sum_1_io_a = {_T_1189,_T_1190}; // @[Math.scala 151:17:@24666.4]
  assign x529_sum_1_io_b = {_T_849,_T_850}; // @[Math.scala 152:17:@24667.4]
  assign x529_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@24668.4]
  assign RetimeWrapper_70_clock = clock; // @[:@24674.4]
  assign RetimeWrapper_70_reset = reset; // @[:@24675.4]
  assign RetimeWrapper_70_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24677.4]
  assign RetimeWrapper_70_io_in = ~ x527; // @[package.scala 94:16:@24676.4]
  assign RetimeWrapper_71_clock = clock; // @[:@24688.4]
  assign RetimeWrapper_71_reset = reset; // @[:@24689.4]
  assign RetimeWrapper_71_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24691.4]
  assign RetimeWrapper_71_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@24690.4]
  assign x539_x11_1_clock = clock; // @[:@24736.4]
  assign x539_x11_1_reset = reset; // @[:@24737.4]
  assign x539_x11_1_io_a = x329_lb_0_io_rPort_10_output_0; // @[Math.scala 151:17:@24738.4]
  assign x539_x11_1_io_b = _T_1392[7:0]; // @[Math.scala 152:17:@24739.4]
  assign x539_x11_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@24740.4]
  assign x540_x12_1_clock = clock; // @[:@24746.4]
  assign x540_x12_1_reset = reset; // @[:@24747.4]
  assign x540_x12_1_io_a = x329_lb_0_io_rPort_3_output_0; // @[Math.scala 151:17:@24748.4]
  assign x540_x12_1_io_b = _T_1398[7:0]; // @[Math.scala 152:17:@24749.4]
  assign x540_x12_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@24750.4]
  assign x541_x11_1_clock = clock; // @[:@24756.4]
  assign x541_x11_1_reset = reset; // @[:@24757.4]
  assign x541_x11_1_io_a = _T_1402[7:0]; // @[Math.scala 151:17:@24758.4]
  assign x541_x11_1_io_b = _T_1406[7:0]; // @[Math.scala 152:17:@24759.4]
  assign x541_x11_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@24760.4]
  assign x542_x12_1_clock = clock; // @[:@24766.4]
  assign x542_x12_1_reset = reset; // @[:@24767.4]
  assign x542_x12_1_io_a = x329_lb_0_io_rPort_16_output_0; // @[Math.scala 151:17:@24768.4]
  assign x542_x12_1_io_b = _T_1410[7:0]; // @[Math.scala 152:17:@24769.4]
  assign x542_x12_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@24770.4]
  assign x543_x11_1_io_a = x539_x11_1_io_result; // @[Math.scala 151:17:@24778.4]
  assign x543_x11_1_io_b = x540_x12_1_io_result; // @[Math.scala 152:17:@24779.4]
  assign x544_x12_1_io_a = x541_x11_1_io_result; // @[Math.scala 151:17:@24788.4]
  assign x544_x12_1_io_b = x542_x12_1_io_result; // @[Math.scala 152:17:@24789.4]
  assign x545_x11_1_io_a = x543_x11_1_io_result; // @[Math.scala 151:17:@24798.4]
  assign x545_x11_1_io_b = x544_x12_1_io_result; // @[Math.scala 152:17:@24799.4]
  assign RetimeWrapper_72_clock = clock; // @[:@24806.4]
  assign RetimeWrapper_72_reset = reset; // @[:@24807.4]
  assign RetimeWrapper_72_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24809.4]
  assign RetimeWrapper_72_io_in = x329_lb_0_io_rPort_2_output_0; // @[package.scala 94:16:@24808.4]
  assign x546_sum_1_io_a = x545_x11_1_io_result; // @[Math.scala 151:17:@24817.4]
  assign x546_sum_1_io_b = RetimeWrapper_72_io_out; // @[Math.scala 152:17:@24818.4]
  assign RetimeWrapper_73_clock = clock; // @[:@24829.4]
  assign RetimeWrapper_73_reset = reset; // @[:@24830.4]
  assign RetimeWrapper_73_io_flow = io_in_x317_TREADY; // @[package.scala 95:18:@24832.4]
  assign RetimeWrapper_73_io_in = {4'h0,_T_1446}; // @[package.scala 94:16:@24831.4]
  assign x553_x11_1_clock = clock; // @[:@24864.4]
  assign x553_x11_1_reset = reset; // @[:@24865.4]
  assign x553_x11_1_io_a = x329_lb_0_io_rPort_6_output_0; // @[Math.scala 151:17:@24866.4]
  assign x553_x11_1_io_b = _T_1453[7:0]; // @[Math.scala 152:17:@24867.4]
  assign x553_x11_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@24868.4]
  assign x554_x12_1_clock = clock; // @[:@24874.4]
  assign x554_x12_1_reset = reset; // @[:@24875.4]
  assign x554_x12_1_io_a = x329_lb_0_io_rPort_11_output_0; // @[Math.scala 151:17:@24876.4]
  assign x554_x12_1_io_b = _T_1457[7:0]; // @[Math.scala 152:17:@24877.4]
  assign x554_x12_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@24878.4]
  assign x555_x11_1_clock = clock; // @[:@24884.4]
  assign x555_x11_1_reset = reset; // @[:@24885.4]
  assign x555_x11_1_io_a = _T_1461[7:0]; // @[Math.scala 151:17:@24886.4]
  assign x555_x11_1_io_b = _T_1465[7:0]; // @[Math.scala 152:17:@24887.4]
  assign x555_x11_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@24888.4]
  assign x556_x12_1_clock = clock; // @[:@24894.4]
  assign x556_x12_1_reset = reset; // @[:@24895.4]
  assign x556_x12_1_io_a = x329_lb_0_io_rPort_5_output_0; // @[Math.scala 151:17:@24896.4]
  assign x556_x12_1_io_b = _T_1469[7:0]; // @[Math.scala 152:17:@24897.4]
  assign x556_x12_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@24898.4]
  assign x557_x11_1_io_a = x553_x11_1_io_result; // @[Math.scala 151:17:@24906.4]
  assign x557_x11_1_io_b = x554_x12_1_io_result; // @[Math.scala 152:17:@24907.4]
  assign x558_x12_1_io_a = x555_x11_1_io_result; // @[Math.scala 151:17:@24916.4]
  assign x558_x12_1_io_b = x556_x12_1_io_result; // @[Math.scala 152:17:@24917.4]
  assign x559_x11_1_io_a = x557_x11_1_io_result; // @[Math.scala 151:17:@24926.4]
  assign x559_x11_1_io_b = x558_x12_1_io_result; // @[Math.scala 152:17:@24927.4]
  assign RetimeWrapper_74_clock = clock; // @[:@24934.4]
  assign RetimeWrapper_74_reset = reset; // @[:@24935.4]
  assign RetimeWrapper_74_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@24937.4]
  assign RetimeWrapper_74_io_in = x329_lb_0_io_rPort_0_output_0; // @[package.scala 94:16:@24936.4]
  assign x560_sum_1_io_a = x559_x11_1_io_result; // @[Math.scala 151:17:@24945.4]
  assign x560_sum_1_io_b = RetimeWrapper_74_io_out; // @[Math.scala 152:17:@24946.4]
  assign RetimeWrapper_75_clock = clock; // @[:@24957.4]
  assign RetimeWrapper_75_reset = reset; // @[:@24958.4]
  assign RetimeWrapper_75_io_flow = io_in_x317_TREADY; // @[package.scala 95:18:@24960.4]
  assign RetimeWrapper_75_io_in = {4'h0,_T_1505}; // @[package.scala 94:16:@24959.4]
  assign x566_x11_1_clock = clock; // @[:@24987.4]
  assign x566_x11_1_reset = reset; // @[:@24988.4]
  assign x566_x11_1_io_a = x329_lb_0_io_rPort_3_output_0; // @[Math.scala 151:17:@24989.4]
  assign x566_x11_1_io_b = _T_1512[7:0]; // @[Math.scala 152:17:@24990.4]
  assign x566_x11_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@24991.4]
  assign x567_x12_1_clock = clock; // @[:@24997.4]
  assign x567_x12_1_reset = reset; // @[:@24998.4]
  assign x567_x12_1_io_a = x329_lb_0_io_rPort_7_output_0; // @[Math.scala 151:17:@24999.4]
  assign x567_x12_1_io_b = _T_1406[7:0]; // @[Math.scala 152:17:@25000.4]
  assign x567_x12_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@25001.4]
  assign x568_x11_1_clock = clock; // @[:@25007.4]
  assign x568_x11_1_reset = reset; // @[:@25008.4]
  assign x568_x11_1_io_a = _T_1516[7:0]; // @[Math.scala 151:17:@25009.4]
  assign x568_x11_1_io_b = _T_1520[7:0]; // @[Math.scala 152:17:@25010.4]
  assign x568_x11_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@25011.4]
  assign x569_x12_1_clock = clock; // @[:@25017.4]
  assign x569_x12_1_reset = reset; // @[:@25018.4]
  assign x569_x12_1_io_a = x329_lb_0_io_rPort_2_output_0; // @[Math.scala 151:17:@25019.4]
  assign x569_x12_1_io_b = _T_1524[7:0]; // @[Math.scala 152:17:@25020.4]
  assign x569_x12_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@25021.4]
  assign x570_x11_1_io_a = x566_x11_1_io_result; // @[Math.scala 151:17:@25029.4]
  assign x570_x11_1_io_b = x567_x12_1_io_result; // @[Math.scala 152:17:@25030.4]
  assign x571_x12_1_io_a = x568_x11_1_io_result; // @[Math.scala 151:17:@25039.4]
  assign x571_x12_1_io_b = x569_x12_1_io_result; // @[Math.scala 152:17:@25040.4]
  assign x572_x11_1_io_a = x570_x11_1_io_result; // @[Math.scala 151:17:@25049.4]
  assign x572_x11_1_io_b = x571_x12_1_io_result; // @[Math.scala 152:17:@25050.4]
  assign RetimeWrapper_76_clock = clock; // @[:@25057.4]
  assign RetimeWrapper_76_reset = reset; // @[:@25058.4]
  assign RetimeWrapper_76_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25060.4]
  assign RetimeWrapper_76_io_in = x329_lb_0_io_rPort_13_output_0; // @[package.scala 94:16:@25059.4]
  assign x573_sum_1_io_a = x572_x11_1_io_result; // @[Math.scala 151:17:@25068.4]
  assign x573_sum_1_io_b = RetimeWrapper_76_io_out; // @[Math.scala 152:17:@25069.4]
  assign RetimeWrapper_77_clock = clock; // @[:@25080.4]
  assign RetimeWrapper_77_reset = reset; // @[:@25081.4]
  assign RetimeWrapper_77_io_flow = io_in_x317_TREADY; // @[package.scala 95:18:@25083.4]
  assign RetimeWrapper_77_io_in = {4'h0,_T_1560}; // @[package.scala 94:16:@25082.4]
  assign x579_x11_1_clock = clock; // @[:@25110.4]
  assign x579_x11_1_reset = reset; // @[:@25111.4]
  assign x579_x11_1_io_a = x329_lb_0_io_rPort_11_output_0; // @[Math.scala 151:17:@25112.4]
  assign x579_x11_1_io_b = _T_1567[7:0]; // @[Math.scala 152:17:@25113.4]
  assign x579_x11_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@25114.4]
  assign x580_x12_1_clock = clock; // @[:@25120.4]
  assign x580_x12_1_reset = reset; // @[:@25121.4]
  assign x580_x12_1_io_a = x329_lb_0_io_rPort_4_output_0; // @[Math.scala 151:17:@25122.4]
  assign x580_x12_1_io_b = _T_1465[7:0]; // @[Math.scala 152:17:@25123.4]
  assign x580_x12_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@25124.4]
  assign x581_x11_1_clock = clock; // @[:@25132.4]
  assign x581_x11_1_reset = reset; // @[:@25133.4]
  assign x581_x11_1_io_a = _T_1571[7:0]; // @[Math.scala 151:17:@25134.4]
  assign x581_x11_1_io_b = _T_1575[7:0]; // @[Math.scala 152:17:@25135.4]
  assign x581_x11_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@25136.4]
  assign x582_x12_1_clock = clock; // @[:@25142.4]
  assign x582_x12_1_reset = reset; // @[:@25143.4]
  assign x582_x12_1_io_a = x329_lb_0_io_rPort_0_output_0; // @[Math.scala 151:17:@25144.4]
  assign x582_x12_1_io_b = _T_1579[7:0]; // @[Math.scala 152:17:@25145.4]
  assign x582_x12_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@25146.4]
  assign x583_x11_1_io_a = x579_x11_1_io_result; // @[Math.scala 151:17:@25154.4]
  assign x583_x11_1_io_b = x580_x12_1_io_result; // @[Math.scala 152:17:@25155.4]
  assign x584_x12_1_io_a = x581_x11_1_io_result; // @[Math.scala 151:17:@25164.4]
  assign x584_x12_1_io_b = x582_x12_1_io_result; // @[Math.scala 152:17:@25165.4]
  assign x585_x11_1_io_a = x583_x11_1_io_result; // @[Math.scala 151:17:@25174.4]
  assign x585_x11_1_io_b = x584_x12_1_io_result; // @[Math.scala 152:17:@25175.4]
  assign RetimeWrapper_78_clock = clock; // @[:@25182.4]
  assign RetimeWrapper_78_reset = reset; // @[:@25183.4]
  assign RetimeWrapper_78_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25185.4]
  assign RetimeWrapper_78_io_in = x329_lb_0_io_rPort_17_output_0; // @[package.scala 94:16:@25184.4]
  assign x586_sum_1_io_a = x585_x11_1_io_result; // @[Math.scala 151:17:@25193.4]
  assign x586_sum_1_io_b = RetimeWrapper_78_io_out; // @[Math.scala 152:17:@25194.4]
  assign RetimeWrapper_79_clock = clock; // @[:@25205.4]
  assign RetimeWrapper_79_reset = reset; // @[:@25206.4]
  assign RetimeWrapper_79_io_flow = io_in_x317_TREADY; // @[package.scala 95:18:@25208.4]
  assign RetimeWrapper_79_io_in = {4'h0,_T_1617}; // @[package.scala 94:16:@25207.4]
  assign RetimeWrapper_80_clock = clock; // @[:@25225.4]
  assign RetimeWrapper_80_reset = reset; // @[:@25226.4]
  assign RetimeWrapper_80_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25228.4]
  assign RetimeWrapper_80_io_in = {_T_1633,_T_1632}; // @[package.scala 94:16:@25227.4]
  assign RetimeWrapper_81_clock = clock; // @[:@25234.4]
  assign RetimeWrapper_81_reset = reset; // @[:@25235.4]
  assign RetimeWrapper_81_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25237.4]
  assign RetimeWrapper_81_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@25236.4]
  assign RetimeWrapper_82_clock = clock; // @[:@25243.4]
  assign RetimeWrapper_82_reset = reset; // @[:@25244.4]
  assign RetimeWrapper_82_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25246.4]
  assign RetimeWrapper_82_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@25245.4]
  assign RetimeWrapper_83_clock = clock; // @[:@25252.4]
  assign RetimeWrapper_83_reset = reset; // @[:@25253.4]
  assign RetimeWrapper_83_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25255.4]
  assign RetimeWrapper_83_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@25254.4]
endmodule
module x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1( // @[:@25273.2]
  input          clock, // @[:@25274.4]
  input          reset, // @[:@25275.4]
  input          io_in_x316_TVALID, // @[:@25276.4]
  output         io_in_x316_TREADY, // @[:@25276.4]
  input  [255:0] io_in_x316_TDATA, // @[:@25276.4]
  input  [7:0]   io_in_x316_TID, // @[:@25276.4]
  input  [7:0]   io_in_x316_TDEST, // @[:@25276.4]
  output         io_in_x317_TVALID, // @[:@25276.4]
  input          io_in_x317_TREADY, // @[:@25276.4]
  output [255:0] io_in_x317_TDATA, // @[:@25276.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@25276.4]
  input          io_sigsIn_smChildAcks_0, // @[:@25276.4]
  output         io_sigsOut_smDoneIn_0, // @[:@25276.4]
  output         io_sigsOut_smCtrCopyDone_0, // @[:@25276.4]
  input          io_rr // @[:@25276.4]
);
  wire  x324_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@25286.4]
  wire  x324_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@25286.4]
  wire  x324_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@25286.4]
  wire  x324_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@25286.4]
  wire [31:0] x324_ctrchain_io_output_counts_1; // @[SpatialBlocks.scala 37:22:@25286.4]
  wire [31:0] x324_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@25286.4]
  wire  x324_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@25286.4]
  wire  x324_ctrchain_io_output_oobs_1; // @[SpatialBlocks.scala 37:22:@25286.4]
  wire  x324_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@25286.4]
  wire  x592_inr_Foreach_SAMPLER_BOX_sm_clock; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 32:18:@25345.4]
  wire  x592_inr_Foreach_SAMPLER_BOX_sm_reset; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 32:18:@25345.4]
  wire  x592_inr_Foreach_SAMPLER_BOX_sm_io_enable; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 32:18:@25345.4]
  wire  x592_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 32:18:@25345.4]
  wire  x592_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 32:18:@25345.4]
  wire  x592_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 32:18:@25345.4]
  wire  x592_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 32:18:@25345.4]
  wire  x592_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 32:18:@25345.4]
  wire  x592_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 32:18:@25345.4]
  wire  x592_inr_Foreach_SAMPLER_BOX_sm_io_parentAck; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 32:18:@25345.4]
  wire  x592_inr_Foreach_SAMPLER_BOX_sm_io_backpressure; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 32:18:@25345.4]
  wire  x592_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 32:18:@25345.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@25373.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@25373.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@25373.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@25373.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@25373.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@25415.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@25415.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@25415.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@25415.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@25415.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@25423.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@25423.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@25423.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@25423.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@25423.4]
  wire  x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_clock; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 702:24:@25455.4]
  wire  x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_reset; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 702:24:@25455.4]
  wire  x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x316_TREADY; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 702:24:@25455.4]
  wire [255:0] x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x316_TDATA; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 702:24:@25455.4]
  wire [7:0] x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x316_TID; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 702:24:@25455.4]
  wire [7:0] x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x316_TDEST; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 702:24:@25455.4]
  wire  x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x317_TVALID; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 702:24:@25455.4]
  wire  x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x317_TREADY; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 702:24:@25455.4]
  wire [255:0] x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x317_TDATA; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 702:24:@25455.4]
  wire  x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 702:24:@25455.4]
  wire  x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 702:24:@25455.4]
  wire  x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 702:24:@25455.4]
  wire [31:0] x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 702:24:@25455.4]
  wire [31:0] x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 702:24:@25455.4]
  wire  x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 702:24:@25455.4]
  wire  x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 702:24:@25455.4]
  wire  x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_rr; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 702:24:@25455.4]
  wire  _T_239; // @[package.scala 96:25:@25378.4 package.scala 96:25:@25379.4]
  wire  x592_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[sm_x593_outr_UnitPipe.scala 68:66:@25384.4]
  wire  _T_252; // @[package.scala 96:25:@25420.4 package.scala 96:25:@25421.4]
  wire  _T_258; // @[package.scala 96:25:@25428.4 package.scala 96:25:@25429.4]
  wire  _T_261; // @[SpatialBlocks.scala 110:93:@25431.4]
  wire  x592_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn; // @[SpatialBlocks.scala 110:90:@25432.4]
  wire  _T_263; // @[SpatialBlocks.scala 128:36:@25440.4]
  wire  _T_264; // @[SpatialBlocks.scala 128:78:@25441.4]
  wire  _T_269; // @[SpatialBlocks.scala 130:61:@25450.4]
  x324_ctrchain x324_ctrchain ( // @[SpatialBlocks.scala 37:22:@25286.4]
    .clock(x324_ctrchain_clock),
    .reset(x324_ctrchain_reset),
    .io_input_reset(x324_ctrchain_io_input_reset),
    .io_input_enable(x324_ctrchain_io_input_enable),
    .io_output_counts_1(x324_ctrchain_io_output_counts_1),
    .io_output_counts_0(x324_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x324_ctrchain_io_output_oobs_0),
    .io_output_oobs_1(x324_ctrchain_io_output_oobs_1),
    .io_output_done(x324_ctrchain_io_output_done)
  );
  x592_inr_Foreach_SAMPLER_BOX_sm x592_inr_Foreach_SAMPLER_BOX_sm ( // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 32:18:@25345.4]
    .clock(x592_inr_Foreach_SAMPLER_BOX_sm_clock),
    .reset(x592_inr_Foreach_SAMPLER_BOX_sm_reset),
    .io_enable(x592_inr_Foreach_SAMPLER_BOX_sm_io_enable),
    .io_done(x592_inr_Foreach_SAMPLER_BOX_sm_io_done),
    .io_doneLatch(x592_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch),
    .io_ctrDone(x592_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone),
    .io_datapathEn(x592_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn),
    .io_ctrInc(x592_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc),
    .io_ctrRst(x592_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst),
    .io_parentAck(x592_inr_Foreach_SAMPLER_BOX_sm_io_parentAck),
    .io_backpressure(x592_inr_Foreach_SAMPLER_BOX_sm_io_backpressure),
    .io_break(x592_inr_Foreach_SAMPLER_BOX_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@25373.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@25415.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@25423.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1 x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1 ( // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 702:24:@25455.4]
    .clock(x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_clock),
    .reset(x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_reset),
    .io_in_x316_TREADY(x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x316_TREADY),
    .io_in_x316_TDATA(x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x316_TDATA),
    .io_in_x316_TID(x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x316_TID),
    .io_in_x316_TDEST(x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x316_TDEST),
    .io_in_x317_TVALID(x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x317_TVALID),
    .io_in_x317_TREADY(x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x317_TREADY),
    .io_in_x317_TDATA(x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x317_TDATA),
    .io_sigsIn_backpressure(x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_1(x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsIn_cchainOutputs_0_oobs_1(x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1),
    .io_rr(x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_rr)
  );
  assign _T_239 = RetimeWrapper_io_out; // @[package.scala 96:25:@25378.4 package.scala 96:25:@25379.4]
  assign x592_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure = io_in_x316_TVALID | x592_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x593_outr_UnitPipe.scala 68:66:@25384.4]
  assign _T_252 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@25420.4 package.scala 96:25:@25421.4]
  assign _T_258 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@25428.4 package.scala 96:25:@25429.4]
  assign _T_261 = ~ _T_258; // @[SpatialBlocks.scala 110:93:@25431.4]
  assign x592_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn = _T_252 & _T_261; // @[SpatialBlocks.scala 110:90:@25432.4]
  assign _T_263 = x592_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[SpatialBlocks.scala 128:36:@25440.4]
  assign _T_264 = ~ x592_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[SpatialBlocks.scala 128:78:@25441.4]
  assign _T_269 = x592_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[SpatialBlocks.scala 130:61:@25450.4]
  assign io_in_x316_TREADY = x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x316_TREADY; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 48:23:@25512.4]
  assign io_in_x317_TVALID = x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x317_TVALID; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 49:23:@25522.4]
  assign io_in_x317_TDATA = x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x317_TDATA; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 49:23:@25520.4]
  assign io_sigsOut_smDoneIn_0 = x592_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[SpatialBlocks.scala 127:53:@25438.4]
  assign io_sigsOut_smCtrCopyDone_0 = x592_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[SpatialBlocks.scala 139:125:@25454.4]
  assign x324_ctrchain_clock = clock; // @[:@25287.4]
  assign x324_ctrchain_reset = reset; // @[:@25288.4]
  assign x324_ctrchain_io_input_reset = x592_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[SpatialBlocks.scala 130:103:@25453.4]
  assign x324_ctrchain_io_input_enable = _T_269 & x592_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 104:75:@25408.4 SpatialBlocks.scala 130:45:@25452.4]
  assign x592_inr_Foreach_SAMPLER_BOX_sm_clock = clock; // @[:@25346.4]
  assign x592_inr_Foreach_SAMPLER_BOX_sm_reset = reset; // @[:@25347.4]
  assign x592_inr_Foreach_SAMPLER_BOX_sm_io_enable = x592_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn & x592_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 112:18:@25435.4]
  assign x592_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone = io_rr ? _T_239 : 1'h0; // @[sm_x593_outr_UnitPipe.scala 66:50:@25381.4]
  assign x592_inr_Foreach_SAMPLER_BOX_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 114:21:@25437.4]
  assign x592_inr_Foreach_SAMPLER_BOX_sm_io_backpressure = io_in_x317_TREADY | x592_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[SpatialBlocks.scala 105:24:@25409.4]
  assign x592_inr_Foreach_SAMPLER_BOX_sm_io_break = 1'h0; // @[sm_x593_outr_UnitPipe.scala 70:48:@25387.4]
  assign RetimeWrapper_clock = clock; // @[:@25374.4]
  assign RetimeWrapper_reset = reset; // @[:@25375.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@25377.4]
  assign RetimeWrapper_io_in = x324_ctrchain_io_output_done; // @[package.scala 94:16:@25376.4]
  assign RetimeWrapper_1_clock = clock; // @[:@25416.4]
  assign RetimeWrapper_1_reset = reset; // @[:@25417.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@25419.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@25418.4]
  assign RetimeWrapper_2_clock = clock; // @[:@25424.4]
  assign RetimeWrapper_2_reset = reset; // @[:@25425.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@25427.4]
  assign RetimeWrapper_2_io_in = x592_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[package.scala 94:16:@25426.4]
  assign x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_clock = clock; // @[:@25456.4]
  assign x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_reset = reset; // @[:@25457.4]
  assign x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x316_TDATA = io_in_x316_TDATA; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 48:23:@25511.4]
  assign x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x316_TID = io_in_x316_TID; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 48:23:@25507.4]
  assign x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x316_TDEST = io_in_x316_TDEST; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 48:23:@25506.4]
  assign x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x317_TREADY = io_in_x317_TREADY; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 49:23:@25521.4]
  assign x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure = io_in_x317_TREADY | x592_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 706:22:@25539.4]
  assign x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn = _T_263 & _T_264; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 706:22:@25537.4]
  assign x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break = x592_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 706:22:@25535.4]
  assign x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1 = x324_ctrchain_io_output_counts_1; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 706:22:@25530.4]
  assign x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = x324_ctrchain_io_output_counts_0; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 706:22:@25529.4]
  assign x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x324_ctrchain_io_output_oobs_0; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 706:22:@25527.4]
  assign x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1 = x324_ctrchain_io_output_oobs_1; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 706:22:@25528.4]
  assign x592_inr_Foreach_SAMPLER_BOX_kernelx592_inr_Foreach_SAMPLER_BOX_concrete1_io_rr = io_rr; // @[sm_x592_inr_Foreach_SAMPLER_BOX.scala 705:18:@25523.4]
endmodule
module RootController_kernelRootController_concrete1( // @[:@25552.2]
  input          clock, // @[:@25553.4]
  input          reset, // @[:@25554.4]
  input          io_in_x316_TVALID, // @[:@25555.4]
  output         io_in_x316_TREADY, // @[:@25555.4]
  input  [255:0] io_in_x316_TDATA, // @[:@25555.4]
  input  [7:0]   io_in_x316_TID, // @[:@25555.4]
  input  [7:0]   io_in_x316_TDEST, // @[:@25555.4]
  output         io_in_x317_TVALID, // @[:@25555.4]
  input          io_in_x317_TREADY, // @[:@25555.4]
  output [255:0] io_in_x317_TDATA, // @[:@25555.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@25555.4]
  input          io_sigsIn_smChildAcks_0, // @[:@25555.4]
  output         io_sigsOut_smDoneIn_0, // @[:@25555.4]
  input          io_rr // @[:@25555.4]
);
  wire  x593_outr_UnitPipe_sm_clock; // @[sm_x593_outr_UnitPipe.scala 32:18:@25696.4]
  wire  x593_outr_UnitPipe_sm_reset; // @[sm_x593_outr_UnitPipe.scala 32:18:@25696.4]
  wire  x593_outr_UnitPipe_sm_io_enable; // @[sm_x593_outr_UnitPipe.scala 32:18:@25696.4]
  wire  x593_outr_UnitPipe_sm_io_done; // @[sm_x593_outr_UnitPipe.scala 32:18:@25696.4]
  wire  x593_outr_UnitPipe_sm_io_parentAck; // @[sm_x593_outr_UnitPipe.scala 32:18:@25696.4]
  wire  x593_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x593_outr_UnitPipe.scala 32:18:@25696.4]
  wire  x593_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x593_outr_UnitPipe.scala 32:18:@25696.4]
  wire  x593_outr_UnitPipe_sm_io_childAck_0; // @[sm_x593_outr_UnitPipe.scala 32:18:@25696.4]
  wire  x593_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x593_outr_UnitPipe.scala 32:18:@25696.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@25748.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@25748.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@25748.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@25748.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@25748.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@25756.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@25756.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@25756.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@25756.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@25756.4]
  wire  x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_clock; // @[sm_x593_outr_UnitPipe.scala 75:24:@25783.4]
  wire  x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_reset; // @[sm_x593_outr_UnitPipe.scala 75:24:@25783.4]
  wire  x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_io_in_x316_TVALID; // @[sm_x593_outr_UnitPipe.scala 75:24:@25783.4]
  wire  x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_io_in_x316_TREADY; // @[sm_x593_outr_UnitPipe.scala 75:24:@25783.4]
  wire [255:0] x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_io_in_x316_TDATA; // @[sm_x593_outr_UnitPipe.scala 75:24:@25783.4]
  wire [7:0] x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_io_in_x316_TID; // @[sm_x593_outr_UnitPipe.scala 75:24:@25783.4]
  wire [7:0] x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_io_in_x316_TDEST; // @[sm_x593_outr_UnitPipe.scala 75:24:@25783.4]
  wire  x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_io_in_x317_TVALID; // @[sm_x593_outr_UnitPipe.scala 75:24:@25783.4]
  wire  x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_io_in_x317_TREADY; // @[sm_x593_outr_UnitPipe.scala 75:24:@25783.4]
  wire [255:0] x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_io_in_x317_TDATA; // @[sm_x593_outr_UnitPipe.scala 75:24:@25783.4]
  wire  x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x593_outr_UnitPipe.scala 75:24:@25783.4]
  wire  x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x593_outr_UnitPipe.scala 75:24:@25783.4]
  wire  x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x593_outr_UnitPipe.scala 75:24:@25783.4]
  wire  x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x593_outr_UnitPipe.scala 75:24:@25783.4]
  wire  x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_io_rr; // @[sm_x593_outr_UnitPipe.scala 75:24:@25783.4]
  wire  _T_246; // @[package.scala 96:25:@25753.4 package.scala 96:25:@25754.4]
  wire  _T_252; // @[package.scala 96:25:@25761.4 package.scala 96:25:@25762.4]
  wire  _T_255; // @[SpatialBlocks.scala 110:93:@25764.4]
  x593_outr_UnitPipe_sm x593_outr_UnitPipe_sm ( // @[sm_x593_outr_UnitPipe.scala 32:18:@25696.4]
    .clock(x593_outr_UnitPipe_sm_clock),
    .reset(x593_outr_UnitPipe_sm_reset),
    .io_enable(x593_outr_UnitPipe_sm_io_enable),
    .io_done(x593_outr_UnitPipe_sm_io_done),
    .io_parentAck(x593_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x593_outr_UnitPipe_sm_io_doneIn_0),
    .io_enableOut_0(x593_outr_UnitPipe_sm_io_enableOut_0),
    .io_childAck_0(x593_outr_UnitPipe_sm_io_childAck_0),
    .io_ctrCopyDone_0(x593_outr_UnitPipe_sm_io_ctrCopyDone_0)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@25748.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@25756.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1 x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1 ( // @[sm_x593_outr_UnitPipe.scala 75:24:@25783.4]
    .clock(x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_clock),
    .reset(x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_reset),
    .io_in_x316_TVALID(x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_io_in_x316_TVALID),
    .io_in_x316_TREADY(x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_io_in_x316_TREADY),
    .io_in_x316_TDATA(x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_io_in_x316_TDATA),
    .io_in_x316_TID(x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_io_in_x316_TID),
    .io_in_x316_TDEST(x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_io_in_x316_TDEST),
    .io_in_x317_TVALID(x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_io_in_x317_TVALID),
    .io_in_x317_TREADY(x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_io_in_x317_TREADY),
    .io_in_x317_TDATA(x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_io_in_x317_TDATA),
    .io_sigsIn_smEnableOuts_0(x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smCtrCopyDone_0(x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_rr(x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_246 = RetimeWrapper_io_out; // @[package.scala 96:25:@25753.4 package.scala 96:25:@25754.4]
  assign _T_252 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@25761.4 package.scala 96:25:@25762.4]
  assign _T_255 = ~ _T_252; // @[SpatialBlocks.scala 110:93:@25764.4]
  assign io_in_x316_TREADY = x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_io_in_x316_TREADY; // @[sm_x593_outr_UnitPipe.scala 48:23:@25838.4]
  assign io_in_x317_TVALID = x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_io_in_x317_TVALID; // @[sm_x593_outr_UnitPipe.scala 49:23:@25848.4]
  assign io_in_x317_TDATA = x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_io_in_x317_TDATA; // @[sm_x593_outr_UnitPipe.scala 49:23:@25846.4]
  assign io_sigsOut_smDoneIn_0 = x593_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 127:53:@25771.4]
  assign x593_outr_UnitPipe_sm_clock = clock; // @[:@25697.4]
  assign x593_outr_UnitPipe_sm_reset = reset; // @[:@25698.4]
  assign x593_outr_UnitPipe_sm_io_enable = _T_246 & _T_255; // @[SpatialBlocks.scala 112:18:@25768.4]
  assign x593_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 114:21:@25770.4]
  assign x593_outr_UnitPipe_sm_io_doneIn_0 = x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 102:67:@25740.4]
  assign x593_outr_UnitPipe_sm_io_ctrCopyDone_0 = x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 132:80:@25782.4]
  assign RetimeWrapper_clock = clock; // @[:@25749.4]
  assign RetimeWrapper_reset = reset; // @[:@25750.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@25752.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@25751.4]
  assign RetimeWrapper_1_clock = clock; // @[:@25757.4]
  assign RetimeWrapper_1_reset = reset; // @[:@25758.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@25760.4]
  assign RetimeWrapper_1_io_in = x593_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@25759.4]
  assign x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_clock = clock; // @[:@25784.4]
  assign x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_reset = reset; // @[:@25785.4]
  assign x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_io_in_x316_TVALID = io_in_x316_TVALID; // @[sm_x593_outr_UnitPipe.scala 48:23:@25839.4]
  assign x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_io_in_x316_TDATA = io_in_x316_TDATA; // @[sm_x593_outr_UnitPipe.scala 48:23:@25837.4]
  assign x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_io_in_x316_TID = io_in_x316_TID; // @[sm_x593_outr_UnitPipe.scala 48:23:@25833.4]
  assign x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_io_in_x316_TDEST = io_in_x316_TDEST; // @[sm_x593_outr_UnitPipe.scala 48:23:@25832.4]
  assign x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_io_in_x317_TREADY = io_in_x317_TREADY; // @[sm_x593_outr_UnitPipe.scala 49:23:@25847.4]
  assign x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x593_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x593_outr_UnitPipe.scala 79:22:@25857.4]
  assign x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x593_outr_UnitPipe_sm_io_childAck_0; // @[sm_x593_outr_UnitPipe.scala 79:22:@25855.4]
  assign x593_outr_UnitPipe_kernelx593_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x593_outr_UnitPipe.scala 78:18:@25849.4]
endmodule
module AccelUnit( // @[:@25876.2]
  input          clock, // @[:@25877.4]
  input          reset, // @[:@25878.4]
  input          io_enable, // @[:@25879.4]
  output         io_done, // @[:@25879.4]
  input          io_reset, // @[:@25879.4]
  input          io_memStreams_loads_0_cmd_ready, // @[:@25879.4]
  output         io_memStreams_loads_0_cmd_valid, // @[:@25879.4]
  output [63:0]  io_memStreams_loads_0_cmd_bits_addr, // @[:@25879.4]
  output [31:0]  io_memStreams_loads_0_cmd_bits_size, // @[:@25879.4]
  output         io_memStreams_loads_0_data_ready, // @[:@25879.4]
  input          io_memStreams_loads_0_data_valid, // @[:@25879.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_0, // @[:@25879.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_1, // @[:@25879.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_2, // @[:@25879.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_3, // @[:@25879.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_4, // @[:@25879.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_5, // @[:@25879.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_6, // @[:@25879.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_7, // @[:@25879.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_8, // @[:@25879.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_9, // @[:@25879.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_10, // @[:@25879.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_11, // @[:@25879.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_12, // @[:@25879.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_13, // @[:@25879.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_14, // @[:@25879.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_15, // @[:@25879.4]
  input          io_memStreams_stores_0_cmd_ready, // @[:@25879.4]
  output         io_memStreams_stores_0_cmd_valid, // @[:@25879.4]
  output [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@25879.4]
  output [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@25879.4]
  input          io_memStreams_stores_0_data_ready, // @[:@25879.4]
  output         io_memStreams_stores_0_data_valid, // @[:@25879.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_0, // @[:@25879.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_1, // @[:@25879.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_2, // @[:@25879.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_3, // @[:@25879.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_4, // @[:@25879.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_5, // @[:@25879.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_6, // @[:@25879.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_7, // @[:@25879.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_8, // @[:@25879.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_9, // @[:@25879.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_10, // @[:@25879.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_11, // @[:@25879.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_12, // @[:@25879.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_13, // @[:@25879.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_14, // @[:@25879.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_15, // @[:@25879.4]
  output [15:0]  io_memStreams_stores_0_data_bits_wstrb, // @[:@25879.4]
  output         io_memStreams_stores_0_wresp_ready, // @[:@25879.4]
  input          io_memStreams_stores_0_wresp_valid, // @[:@25879.4]
  input          io_memStreams_stores_0_wresp_bits, // @[:@25879.4]
  input          io_memStreams_gathers_0_cmd_ready, // @[:@25879.4]
  output         io_memStreams_gathers_0_cmd_valid, // @[:@25879.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_0, // @[:@25879.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_1, // @[:@25879.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_2, // @[:@25879.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_3, // @[:@25879.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_4, // @[:@25879.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_5, // @[:@25879.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_6, // @[:@25879.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_7, // @[:@25879.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_8, // @[:@25879.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_9, // @[:@25879.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_10, // @[:@25879.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_11, // @[:@25879.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_12, // @[:@25879.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_13, // @[:@25879.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_14, // @[:@25879.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_15, // @[:@25879.4]
  output         io_memStreams_gathers_0_data_ready, // @[:@25879.4]
  input          io_memStreams_gathers_0_data_valid, // @[:@25879.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_0, // @[:@25879.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_1, // @[:@25879.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_2, // @[:@25879.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_3, // @[:@25879.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_4, // @[:@25879.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_5, // @[:@25879.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_6, // @[:@25879.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_7, // @[:@25879.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_8, // @[:@25879.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_9, // @[:@25879.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_10, // @[:@25879.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_11, // @[:@25879.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_12, // @[:@25879.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_13, // @[:@25879.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_14, // @[:@25879.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_15, // @[:@25879.4]
  input          io_memStreams_scatters_0_cmd_ready, // @[:@25879.4]
  output         io_memStreams_scatters_0_cmd_valid, // @[:@25879.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_0, // @[:@25879.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_1, // @[:@25879.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_2, // @[:@25879.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_3, // @[:@25879.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_4, // @[:@25879.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_5, // @[:@25879.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_6, // @[:@25879.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_7, // @[:@25879.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_8, // @[:@25879.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_9, // @[:@25879.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_10, // @[:@25879.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_11, // @[:@25879.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_12, // @[:@25879.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_13, // @[:@25879.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_14, // @[:@25879.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_15, // @[:@25879.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_0, // @[:@25879.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_1, // @[:@25879.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_2, // @[:@25879.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_3, // @[:@25879.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_4, // @[:@25879.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_5, // @[:@25879.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_6, // @[:@25879.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_7, // @[:@25879.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_8, // @[:@25879.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_9, // @[:@25879.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_10, // @[:@25879.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_11, // @[:@25879.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_12, // @[:@25879.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_13, // @[:@25879.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_14, // @[:@25879.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_15, // @[:@25879.4]
  output         io_memStreams_scatters_0_wresp_ready, // @[:@25879.4]
  input          io_memStreams_scatters_0_wresp_valid, // @[:@25879.4]
  input          io_memStreams_scatters_0_wresp_bits, // @[:@25879.4]
  input          io_axiStreamsIn_0_TVALID, // @[:@25879.4]
  output         io_axiStreamsIn_0_TREADY, // @[:@25879.4]
  input  [255:0] io_axiStreamsIn_0_TDATA, // @[:@25879.4]
  input  [31:0]  io_axiStreamsIn_0_TSTRB, // @[:@25879.4]
  input  [31:0]  io_axiStreamsIn_0_TKEEP, // @[:@25879.4]
  input          io_axiStreamsIn_0_TLAST, // @[:@25879.4]
  input  [7:0]   io_axiStreamsIn_0_TID, // @[:@25879.4]
  input  [7:0]   io_axiStreamsIn_0_TDEST, // @[:@25879.4]
  input  [31:0]  io_axiStreamsIn_0_TUSER, // @[:@25879.4]
  output         io_axiStreamsOut_0_TVALID, // @[:@25879.4]
  input          io_axiStreamsOut_0_TREADY, // @[:@25879.4]
  output [255:0] io_axiStreamsOut_0_TDATA, // @[:@25879.4]
  output [31:0]  io_axiStreamsOut_0_TSTRB, // @[:@25879.4]
  output [31:0]  io_axiStreamsOut_0_TKEEP, // @[:@25879.4]
  output         io_axiStreamsOut_0_TLAST, // @[:@25879.4]
  output [7:0]   io_axiStreamsOut_0_TID, // @[:@25879.4]
  output [7:0]   io_axiStreamsOut_0_TDEST, // @[:@25879.4]
  output [31:0]  io_axiStreamsOut_0_TUSER, // @[:@25879.4]
  output         io_heap_0_req_valid, // @[:@25879.4]
  output         io_heap_0_req_bits_allocDealloc, // @[:@25879.4]
  output [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@25879.4]
  input          io_heap_0_resp_valid, // @[:@25879.4]
  input          io_heap_0_resp_bits_allocDealloc, // @[:@25879.4]
  input  [63:0]  io_heap_0_resp_bits_sizeAddr, // @[:@25879.4]
  input  [63:0]  io_argIns_0, // @[:@25879.4]
  input  [63:0]  io_argIns_1, // @[:@25879.4]
  input          io_argOuts_0_port_ready, // @[:@25879.4]
  output         io_argOuts_0_port_valid, // @[:@25879.4]
  output [63:0]  io_argOuts_0_port_bits, // @[:@25879.4]
  input  [63:0]  io_argOuts_0_echo // @[:@25879.4]
);
  wire  SingleCounter_clock; // @[Main.scala 35:32:@26042.4]
  wire  SingleCounter_reset; // @[Main.scala 35:32:@26042.4]
  wire  SingleCounter_io_input_reset; // @[Main.scala 35:32:@26042.4]
  wire  SingleCounter_io_output_done; // @[Main.scala 35:32:@26042.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@26060.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@26060.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@26060.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@26060.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@26060.4]
  wire  SRFF_clock; // @[Main.scala 39:28:@26069.4]
  wire  SRFF_reset; // @[Main.scala 39:28:@26069.4]
  wire  SRFF_io_input_set; // @[Main.scala 39:28:@26069.4]
  wire  SRFF_io_input_reset; // @[Main.scala 39:28:@26069.4]
  wire  SRFF_io_input_asyn_reset; // @[Main.scala 39:28:@26069.4]
  wire  SRFF_io_output; // @[Main.scala 39:28:@26069.4]
  wire  RootController_sm_clock; // @[sm_RootController.scala 32:18:@26107.4]
  wire  RootController_sm_reset; // @[sm_RootController.scala 32:18:@26107.4]
  wire  RootController_sm_io_enable; // @[sm_RootController.scala 32:18:@26107.4]
  wire  RootController_sm_io_done; // @[sm_RootController.scala 32:18:@26107.4]
  wire  RootController_sm_io_rst; // @[sm_RootController.scala 32:18:@26107.4]
  wire  RootController_sm_io_ctrDone; // @[sm_RootController.scala 32:18:@26107.4]
  wire  RootController_sm_io_ctrInc; // @[sm_RootController.scala 32:18:@26107.4]
  wire  RootController_sm_io_doneIn_0; // @[sm_RootController.scala 32:18:@26107.4]
  wire  RootController_sm_io_enableOut_0; // @[sm_RootController.scala 32:18:@26107.4]
  wire  RootController_sm_io_childAck_0; // @[sm_RootController.scala 32:18:@26107.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@26139.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@26139.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@26139.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@26139.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@26139.4]
  wire  RootController_kernelRootController_concrete1_clock; // @[sm_RootController.scala 73:24:@26198.4]
  wire  RootController_kernelRootController_concrete1_reset; // @[sm_RootController.scala 73:24:@26198.4]
  wire  RootController_kernelRootController_concrete1_io_in_x316_TVALID; // @[sm_RootController.scala 73:24:@26198.4]
  wire  RootController_kernelRootController_concrete1_io_in_x316_TREADY; // @[sm_RootController.scala 73:24:@26198.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x316_TDATA; // @[sm_RootController.scala 73:24:@26198.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x316_TID; // @[sm_RootController.scala 73:24:@26198.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x316_TDEST; // @[sm_RootController.scala 73:24:@26198.4]
  wire  RootController_kernelRootController_concrete1_io_in_x317_TVALID; // @[sm_RootController.scala 73:24:@26198.4]
  wire  RootController_kernelRootController_concrete1_io_in_x317_TREADY; // @[sm_RootController.scala 73:24:@26198.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x317_TDATA; // @[sm_RootController.scala 73:24:@26198.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_RootController.scala 73:24:@26198.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0; // @[sm_RootController.scala 73:24:@26198.4]
  wire  RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[sm_RootController.scala 73:24:@26198.4]
  wire  RootController_kernelRootController_concrete1_io_rr; // @[sm_RootController.scala 73:24:@26198.4]
  wire  _T_599; // @[package.scala 96:25:@26065.4 package.scala 96:25:@26066.4]
  wire  _T_664; // @[Main.scala 41:50:@26135.4]
  wire  _T_665; // @[Main.scala 41:59:@26136.4]
  wire  _T_677; // @[package.scala 100:49:@26156.4]
  reg  _T_680; // @[package.scala 48:56:@26157.4]
  reg [31:0] _RAND_0;
  SingleCounter SingleCounter ( // @[Main.scala 35:32:@26042.4]
    .clock(SingleCounter_clock),
    .reset(SingleCounter_reset),
    .io_input_reset(SingleCounter_io_input_reset),
    .io_output_done(SingleCounter_io_output_done)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@26060.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  SRFF SRFF ( // @[Main.scala 39:28:@26069.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  RootController_sm RootController_sm ( // @[sm_RootController.scala 32:18:@26107.4]
    .clock(RootController_sm_clock),
    .reset(RootController_sm_reset),
    .io_enable(RootController_sm_io_enable),
    .io_done(RootController_sm_io_done),
    .io_rst(RootController_sm_io_rst),
    .io_ctrDone(RootController_sm_io_ctrDone),
    .io_ctrInc(RootController_sm_io_ctrInc),
    .io_doneIn_0(RootController_sm_io_doneIn_0),
    .io_enableOut_0(RootController_sm_io_enableOut_0),
    .io_childAck_0(RootController_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@26139.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RootController_kernelRootController_concrete1 RootController_kernelRootController_concrete1 ( // @[sm_RootController.scala 73:24:@26198.4]
    .clock(RootController_kernelRootController_concrete1_clock),
    .reset(RootController_kernelRootController_concrete1_reset),
    .io_in_x316_TVALID(RootController_kernelRootController_concrete1_io_in_x316_TVALID),
    .io_in_x316_TREADY(RootController_kernelRootController_concrete1_io_in_x316_TREADY),
    .io_in_x316_TDATA(RootController_kernelRootController_concrete1_io_in_x316_TDATA),
    .io_in_x316_TID(RootController_kernelRootController_concrete1_io_in_x316_TID),
    .io_in_x316_TDEST(RootController_kernelRootController_concrete1_io_in_x316_TDEST),
    .io_in_x317_TVALID(RootController_kernelRootController_concrete1_io_in_x317_TVALID),
    .io_in_x317_TREADY(RootController_kernelRootController_concrete1_io_in_x317_TREADY),
    .io_in_x317_TDATA(RootController_kernelRootController_concrete1_io_in_x317_TDATA),
    .io_sigsIn_smEnableOuts_0(RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(RootController_kernelRootController_concrete1_io_rr)
  );
  assign _T_599 = RetimeWrapper_io_out; // @[package.scala 96:25:@26065.4 package.scala 96:25:@26066.4]
  assign _T_664 = io_enable & _T_599; // @[Main.scala 41:50:@26135.4]
  assign _T_665 = ~ SRFF_io_output; // @[Main.scala 41:59:@26136.4]
  assign _T_677 = RootController_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@26156.4]
  assign io_done = SRFF_io_output; // @[Main.scala 48:23:@26155.4]
  assign io_memStreams_loads_0_cmd_valid = 1'h0;
  assign io_memStreams_loads_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_loads_0_cmd_bits_size = 32'h0;
  assign io_memStreams_loads_0_data_ready = 1'h0;
  assign io_memStreams_stores_0_cmd_valid = 1'h0;
  assign io_memStreams_stores_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_stores_0_cmd_bits_size = 32'h0;
  assign io_memStreams_stores_0_data_valid = 1'h0;
  assign io_memStreams_stores_0_data_bits_wdata_0 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_1 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_2 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_3 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_4 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_5 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_6 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_7 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_8 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_9 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_10 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_11 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_12 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_13 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_14 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_15 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wstrb = 16'h0;
  assign io_memStreams_stores_0_wresp_ready = 1'h0;
  assign io_memStreams_gathers_0_cmd_valid = 1'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_0 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_1 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_2 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_3 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_4 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_5 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_6 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_7 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_8 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_9 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_10 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_11 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_12 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_13 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_14 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_15 = 64'h0;
  assign io_memStreams_gathers_0_data_ready = 1'h0;
  assign io_memStreams_scatters_0_cmd_valid = 1'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_0 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_1 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_2 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_3 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_4 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_5 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_6 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_7 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_8 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_9 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_10 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_11 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_12 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_13 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_14 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_15 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_0 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_1 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_2 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_3 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_4 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_5 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_6 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_7 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_8 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_9 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_10 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_11 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_12 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_13 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_14 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_15 = 32'h0;
  assign io_memStreams_scatters_0_wresp_ready = 1'h0;
  assign io_axiStreamsIn_0_TREADY = RootController_kernelRootController_concrete1_io_in_x316_TREADY; // @[sm_RootController.scala 48:23:@26253.4]
  assign io_axiStreamsOut_0_TVALID = RootController_kernelRootController_concrete1_io_in_x317_TVALID; // @[sm_RootController.scala 49:23:@26263.4]
  assign io_axiStreamsOut_0_TDATA = RootController_kernelRootController_concrete1_io_in_x317_TDATA; // @[sm_RootController.scala 49:23:@26261.4]
  assign io_axiStreamsOut_0_TSTRB = 32'hffffffff; // @[sm_RootController.scala 49:23:@26260.4]
  assign io_axiStreamsOut_0_TKEEP = 32'hffffffff; // @[sm_RootController.scala 49:23:@26259.4]
  assign io_axiStreamsOut_0_TLAST = 1'h0; // @[sm_RootController.scala 49:23:@26258.4]
  assign io_axiStreamsOut_0_TID = 8'h0; // @[sm_RootController.scala 49:23:@26257.4]
  assign io_axiStreamsOut_0_TDEST = 8'h0; // @[sm_RootController.scala 49:23:@26256.4]
  assign io_axiStreamsOut_0_TUSER = 32'h4; // @[sm_RootController.scala 49:23:@26255.4]
  assign io_heap_0_req_valid = 1'h0;
  assign io_heap_0_req_bits_allocDealloc = 1'h0;
  assign io_heap_0_req_bits_sizeAddr = 64'h0;
  assign io_argOuts_0_port_valid = 1'h0;
  assign io_argOuts_0_port_bits = 64'h0;
  assign SingleCounter_clock = clock; // @[:@26043.4]
  assign SingleCounter_reset = reset; // @[:@26044.4]
  assign SingleCounter_io_input_reset = reset; // @[Main.scala 36:79:@26058.4]
  assign RetimeWrapper_clock = clock; // @[:@26061.4]
  assign RetimeWrapper_reset = reset; // @[:@26062.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@26064.4]
  assign RetimeWrapper_io_in = SingleCounter_io_output_done; // @[package.scala 94:16:@26063.4]
  assign SRFF_clock = clock; // @[:@26070.4]
  assign SRFF_reset = reset; // @[:@26071.4]
  assign SRFF_io_input_set = RootController_sm_io_done; // @[Main.scala 57:29:@26290.4]
  assign SRFF_io_input_reset = RetimeWrapper_1_io_out; // @[Main.scala 46:31:@26153.4]
  assign SRFF_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[Main.scala 47:36:@26154.4]
  assign RootController_sm_clock = clock; // @[:@26108.4]
  assign RootController_sm_reset = reset; // @[:@26109.4]
  assign RootController_sm_io_enable = _T_664 & _T_665; // @[Main.scala 45:33:@26152.4 SpatialBlocks.scala 112:18:@26186.4]
  assign RootController_sm_io_rst = RetimeWrapper_1_io_out; // @[SpatialBlocks.scala 106:15:@26180.4]
  assign RootController_sm_io_ctrDone = RootController_sm_io_ctrInc & _T_680; // @[Main.scala 49:34:@26160.4]
  assign RootController_sm_io_doneIn_0 = RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 102:67:@26177.4]
  assign RetimeWrapper_1_clock = clock; // @[:@26140.4]
  assign RetimeWrapper_1_reset = reset; // @[:@26141.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@26143.4]
  assign RetimeWrapper_1_io_in = reset | io_reset; // @[package.scala 94:16:@26142.4]
  assign RootController_kernelRootController_concrete1_clock = clock; // @[:@26199.4]
  assign RootController_kernelRootController_concrete1_reset = reset; // @[:@26200.4]
  assign RootController_kernelRootController_concrete1_io_in_x316_TVALID = io_axiStreamsIn_0_TVALID; // @[sm_RootController.scala 48:23:@26254.4]
  assign RootController_kernelRootController_concrete1_io_in_x316_TDATA = io_axiStreamsIn_0_TDATA; // @[sm_RootController.scala 48:23:@26252.4]
  assign RootController_kernelRootController_concrete1_io_in_x316_TID = io_axiStreamsIn_0_TID; // @[sm_RootController.scala 48:23:@26248.4]
  assign RootController_kernelRootController_concrete1_io_in_x316_TDEST = io_axiStreamsIn_0_TDEST; // @[sm_RootController.scala 48:23:@26247.4]
  assign RootController_kernelRootController_concrete1_io_in_x317_TREADY = io_axiStreamsOut_0_TREADY; // @[sm_RootController.scala 49:23:@26262.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0 = RootController_sm_io_enableOut_0; // @[sm_RootController.scala 77:22:@26272.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0 = RootController_sm_io_childAck_0; // @[sm_RootController.scala 77:22:@26270.4]
  assign RootController_kernelRootController_concrete1_io_rr = RetimeWrapper_io_out; // @[sm_RootController.scala 76:18:@26264.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_680 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_680 <= 1'h0;
    end else begin
      _T_680 <= _T_677;
    end
  end
endmodule
module SpatialIP( // @[:@26292.2]
  input         clock, // @[:@26293.4]
  input         reset, // @[:@26294.4]
  input  [31:0] io_raddr, // @[:@26295.4]
  input         io_wen, // @[:@26295.4]
  input  [31:0] io_waddr, // @[:@26295.4]
  input  [63:0] io_wdata, // @[:@26295.4]
  output [63:0] io_rdata // @[:@26295.4]
);
  wire  accel_clock; // @[Instantiator.scala 53:44:@26297.4]
  wire  accel_reset; // @[Instantiator.scala 53:44:@26297.4]
  wire  accel_io_enable; // @[Instantiator.scala 53:44:@26297.4]
  wire  accel_io_done; // @[Instantiator.scala 53:44:@26297.4]
  wire  accel_io_reset; // @[Instantiator.scala 53:44:@26297.4]
  wire  accel_io_memStreams_loads_0_cmd_ready; // @[Instantiator.scala 53:44:@26297.4]
  wire  accel_io_memStreams_loads_0_cmd_valid; // @[Instantiator.scala 53:44:@26297.4]
  wire [63:0] accel_io_memStreams_loads_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_loads_0_cmd_bits_size; // @[Instantiator.scala 53:44:@26297.4]
  wire  accel_io_memStreams_loads_0_data_ready; // @[Instantiator.scala 53:44:@26297.4]
  wire  accel_io_memStreams_loads_0_data_valid; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_0; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_1; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_2; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_3; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_4; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_5; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_6; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_7; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_8; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_9; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_10; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_11; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_12; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_13; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_14; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_15; // @[Instantiator.scala 53:44:@26297.4]
  wire  accel_io_memStreams_stores_0_cmd_ready; // @[Instantiator.scala 53:44:@26297.4]
  wire  accel_io_memStreams_stores_0_cmd_valid; // @[Instantiator.scala 53:44:@26297.4]
  wire [63:0] accel_io_memStreams_stores_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_stores_0_cmd_bits_size; // @[Instantiator.scala 53:44:@26297.4]
  wire  accel_io_memStreams_stores_0_data_ready; // @[Instantiator.scala 53:44:@26297.4]
  wire  accel_io_memStreams_stores_0_data_valid; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_1; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_2; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_3; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_4; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_5; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_6; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_7; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_8; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_9; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_10; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_11; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_12; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_13; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_14; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_15; // @[Instantiator.scala 53:44:@26297.4]
  wire [15:0] accel_io_memStreams_stores_0_data_bits_wstrb; // @[Instantiator.scala 53:44:@26297.4]
  wire  accel_io_memStreams_stores_0_wresp_ready; // @[Instantiator.scala 53:44:@26297.4]
  wire  accel_io_memStreams_stores_0_wresp_valid; // @[Instantiator.scala 53:44:@26297.4]
  wire  accel_io_memStreams_stores_0_wresp_bits; // @[Instantiator.scala 53:44:@26297.4]
  wire  accel_io_memStreams_gathers_0_cmd_ready; // @[Instantiator.scala 53:44:@26297.4]
  wire  accel_io_memStreams_gathers_0_cmd_valid; // @[Instantiator.scala 53:44:@26297.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_0; // @[Instantiator.scala 53:44:@26297.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_1; // @[Instantiator.scala 53:44:@26297.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_2; // @[Instantiator.scala 53:44:@26297.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_3; // @[Instantiator.scala 53:44:@26297.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_4; // @[Instantiator.scala 53:44:@26297.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_5; // @[Instantiator.scala 53:44:@26297.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_6; // @[Instantiator.scala 53:44:@26297.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_7; // @[Instantiator.scala 53:44:@26297.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_8; // @[Instantiator.scala 53:44:@26297.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_9; // @[Instantiator.scala 53:44:@26297.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_10; // @[Instantiator.scala 53:44:@26297.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_11; // @[Instantiator.scala 53:44:@26297.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_12; // @[Instantiator.scala 53:44:@26297.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_13; // @[Instantiator.scala 53:44:@26297.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_14; // @[Instantiator.scala 53:44:@26297.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_15; // @[Instantiator.scala 53:44:@26297.4]
  wire  accel_io_memStreams_gathers_0_data_ready; // @[Instantiator.scala 53:44:@26297.4]
  wire  accel_io_memStreams_gathers_0_data_valid; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_0; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_1; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_2; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_3; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_4; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_5; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_6; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_7; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_8; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_9; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_10; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_11; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_12; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_13; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_14; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_15; // @[Instantiator.scala 53:44:@26297.4]
  wire  accel_io_memStreams_scatters_0_cmd_ready; // @[Instantiator.scala 53:44:@26297.4]
  wire  accel_io_memStreams_scatters_0_cmd_valid; // @[Instantiator.scala 53:44:@26297.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0; // @[Instantiator.scala 53:44:@26297.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1; // @[Instantiator.scala 53:44:@26297.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2; // @[Instantiator.scala 53:44:@26297.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3; // @[Instantiator.scala 53:44:@26297.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4; // @[Instantiator.scala 53:44:@26297.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5; // @[Instantiator.scala 53:44:@26297.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6; // @[Instantiator.scala 53:44:@26297.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7; // @[Instantiator.scala 53:44:@26297.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8; // @[Instantiator.scala 53:44:@26297.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9; // @[Instantiator.scala 53:44:@26297.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10; // @[Instantiator.scala 53:44:@26297.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11; // @[Instantiator.scala 53:44:@26297.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12; // @[Instantiator.scala 53:44:@26297.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13; // @[Instantiator.scala 53:44:@26297.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14; // @[Instantiator.scala 53:44:@26297.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_0; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_1; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_2; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_3; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_4; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_5; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_6; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_7; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_8; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_9; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_10; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_11; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_12; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_13; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_14; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_15; // @[Instantiator.scala 53:44:@26297.4]
  wire  accel_io_memStreams_scatters_0_wresp_ready; // @[Instantiator.scala 53:44:@26297.4]
  wire  accel_io_memStreams_scatters_0_wresp_valid; // @[Instantiator.scala 53:44:@26297.4]
  wire  accel_io_memStreams_scatters_0_wresp_bits; // @[Instantiator.scala 53:44:@26297.4]
  wire  accel_io_axiStreamsIn_0_TVALID; // @[Instantiator.scala 53:44:@26297.4]
  wire  accel_io_axiStreamsIn_0_TREADY; // @[Instantiator.scala 53:44:@26297.4]
  wire [255:0] accel_io_axiStreamsIn_0_TDATA; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_axiStreamsIn_0_TSTRB; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_axiStreamsIn_0_TKEEP; // @[Instantiator.scala 53:44:@26297.4]
  wire  accel_io_axiStreamsIn_0_TLAST; // @[Instantiator.scala 53:44:@26297.4]
  wire [7:0] accel_io_axiStreamsIn_0_TID; // @[Instantiator.scala 53:44:@26297.4]
  wire [7:0] accel_io_axiStreamsIn_0_TDEST; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_axiStreamsIn_0_TUSER; // @[Instantiator.scala 53:44:@26297.4]
  wire  accel_io_axiStreamsOut_0_TVALID; // @[Instantiator.scala 53:44:@26297.4]
  wire  accel_io_axiStreamsOut_0_TREADY; // @[Instantiator.scala 53:44:@26297.4]
  wire [255:0] accel_io_axiStreamsOut_0_TDATA; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_axiStreamsOut_0_TSTRB; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_axiStreamsOut_0_TKEEP; // @[Instantiator.scala 53:44:@26297.4]
  wire  accel_io_axiStreamsOut_0_TLAST; // @[Instantiator.scala 53:44:@26297.4]
  wire [7:0] accel_io_axiStreamsOut_0_TID; // @[Instantiator.scala 53:44:@26297.4]
  wire [7:0] accel_io_axiStreamsOut_0_TDEST; // @[Instantiator.scala 53:44:@26297.4]
  wire [31:0] accel_io_axiStreamsOut_0_TUSER; // @[Instantiator.scala 53:44:@26297.4]
  wire  accel_io_heap_0_req_valid; // @[Instantiator.scala 53:44:@26297.4]
  wire  accel_io_heap_0_req_bits_allocDealloc; // @[Instantiator.scala 53:44:@26297.4]
  wire [63:0] accel_io_heap_0_req_bits_sizeAddr; // @[Instantiator.scala 53:44:@26297.4]
  wire  accel_io_heap_0_resp_valid; // @[Instantiator.scala 53:44:@26297.4]
  wire  accel_io_heap_0_resp_bits_allocDealloc; // @[Instantiator.scala 53:44:@26297.4]
  wire [63:0] accel_io_heap_0_resp_bits_sizeAddr; // @[Instantiator.scala 53:44:@26297.4]
  wire [63:0] accel_io_argIns_0; // @[Instantiator.scala 53:44:@26297.4]
  wire [63:0] accel_io_argIns_1; // @[Instantiator.scala 53:44:@26297.4]
  wire  accel_io_argOuts_0_port_ready; // @[Instantiator.scala 53:44:@26297.4]
  wire  accel_io_argOuts_0_port_valid; // @[Instantiator.scala 53:44:@26297.4]
  wire [63:0] accel_io_argOuts_0_port_bits; // @[Instantiator.scala 53:44:@26297.4]
  wire [63:0] accel_io_argOuts_0_echo; // @[Instantiator.scala 53:44:@26297.4]
  AccelUnit accel ( // @[Instantiator.scala 53:44:@26297.4]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_enable(accel_io_enable),
    .io_done(accel_io_done),
    .io_reset(accel_io_reset),
    .io_memStreams_loads_0_cmd_ready(accel_io_memStreams_loads_0_cmd_ready),
    .io_memStreams_loads_0_cmd_valid(accel_io_memStreams_loads_0_cmd_valid),
    .io_memStreams_loads_0_cmd_bits_addr(accel_io_memStreams_loads_0_cmd_bits_addr),
    .io_memStreams_loads_0_cmd_bits_size(accel_io_memStreams_loads_0_cmd_bits_size),
    .io_memStreams_loads_0_data_ready(accel_io_memStreams_loads_0_data_ready),
    .io_memStreams_loads_0_data_valid(accel_io_memStreams_loads_0_data_valid),
    .io_memStreams_loads_0_data_bits_rdata_0(accel_io_memStreams_loads_0_data_bits_rdata_0),
    .io_memStreams_loads_0_data_bits_rdata_1(accel_io_memStreams_loads_0_data_bits_rdata_1),
    .io_memStreams_loads_0_data_bits_rdata_2(accel_io_memStreams_loads_0_data_bits_rdata_2),
    .io_memStreams_loads_0_data_bits_rdata_3(accel_io_memStreams_loads_0_data_bits_rdata_3),
    .io_memStreams_loads_0_data_bits_rdata_4(accel_io_memStreams_loads_0_data_bits_rdata_4),
    .io_memStreams_loads_0_data_bits_rdata_5(accel_io_memStreams_loads_0_data_bits_rdata_5),
    .io_memStreams_loads_0_data_bits_rdata_6(accel_io_memStreams_loads_0_data_bits_rdata_6),
    .io_memStreams_loads_0_data_bits_rdata_7(accel_io_memStreams_loads_0_data_bits_rdata_7),
    .io_memStreams_loads_0_data_bits_rdata_8(accel_io_memStreams_loads_0_data_bits_rdata_8),
    .io_memStreams_loads_0_data_bits_rdata_9(accel_io_memStreams_loads_0_data_bits_rdata_9),
    .io_memStreams_loads_0_data_bits_rdata_10(accel_io_memStreams_loads_0_data_bits_rdata_10),
    .io_memStreams_loads_0_data_bits_rdata_11(accel_io_memStreams_loads_0_data_bits_rdata_11),
    .io_memStreams_loads_0_data_bits_rdata_12(accel_io_memStreams_loads_0_data_bits_rdata_12),
    .io_memStreams_loads_0_data_bits_rdata_13(accel_io_memStreams_loads_0_data_bits_rdata_13),
    .io_memStreams_loads_0_data_bits_rdata_14(accel_io_memStreams_loads_0_data_bits_rdata_14),
    .io_memStreams_loads_0_data_bits_rdata_15(accel_io_memStreams_loads_0_data_bits_rdata_15),
    .io_memStreams_stores_0_cmd_ready(accel_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(accel_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(accel_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(accel_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(accel_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(accel_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(accel_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wdata_1(accel_io_memStreams_stores_0_data_bits_wdata_1),
    .io_memStreams_stores_0_data_bits_wdata_2(accel_io_memStreams_stores_0_data_bits_wdata_2),
    .io_memStreams_stores_0_data_bits_wdata_3(accel_io_memStreams_stores_0_data_bits_wdata_3),
    .io_memStreams_stores_0_data_bits_wdata_4(accel_io_memStreams_stores_0_data_bits_wdata_4),
    .io_memStreams_stores_0_data_bits_wdata_5(accel_io_memStreams_stores_0_data_bits_wdata_5),
    .io_memStreams_stores_0_data_bits_wdata_6(accel_io_memStreams_stores_0_data_bits_wdata_6),
    .io_memStreams_stores_0_data_bits_wdata_7(accel_io_memStreams_stores_0_data_bits_wdata_7),
    .io_memStreams_stores_0_data_bits_wdata_8(accel_io_memStreams_stores_0_data_bits_wdata_8),
    .io_memStreams_stores_0_data_bits_wdata_9(accel_io_memStreams_stores_0_data_bits_wdata_9),
    .io_memStreams_stores_0_data_bits_wdata_10(accel_io_memStreams_stores_0_data_bits_wdata_10),
    .io_memStreams_stores_0_data_bits_wdata_11(accel_io_memStreams_stores_0_data_bits_wdata_11),
    .io_memStreams_stores_0_data_bits_wdata_12(accel_io_memStreams_stores_0_data_bits_wdata_12),
    .io_memStreams_stores_0_data_bits_wdata_13(accel_io_memStreams_stores_0_data_bits_wdata_13),
    .io_memStreams_stores_0_data_bits_wdata_14(accel_io_memStreams_stores_0_data_bits_wdata_14),
    .io_memStreams_stores_0_data_bits_wdata_15(accel_io_memStreams_stores_0_data_bits_wdata_15),
    .io_memStreams_stores_0_data_bits_wstrb(accel_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(accel_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(accel_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(accel_io_memStreams_stores_0_wresp_bits),
    .io_memStreams_gathers_0_cmd_ready(accel_io_memStreams_gathers_0_cmd_ready),
    .io_memStreams_gathers_0_cmd_valid(accel_io_memStreams_gathers_0_cmd_valid),
    .io_memStreams_gathers_0_cmd_bits_addr_0(accel_io_memStreams_gathers_0_cmd_bits_addr_0),
    .io_memStreams_gathers_0_cmd_bits_addr_1(accel_io_memStreams_gathers_0_cmd_bits_addr_1),
    .io_memStreams_gathers_0_cmd_bits_addr_2(accel_io_memStreams_gathers_0_cmd_bits_addr_2),
    .io_memStreams_gathers_0_cmd_bits_addr_3(accel_io_memStreams_gathers_0_cmd_bits_addr_3),
    .io_memStreams_gathers_0_cmd_bits_addr_4(accel_io_memStreams_gathers_0_cmd_bits_addr_4),
    .io_memStreams_gathers_0_cmd_bits_addr_5(accel_io_memStreams_gathers_0_cmd_bits_addr_5),
    .io_memStreams_gathers_0_cmd_bits_addr_6(accel_io_memStreams_gathers_0_cmd_bits_addr_6),
    .io_memStreams_gathers_0_cmd_bits_addr_7(accel_io_memStreams_gathers_0_cmd_bits_addr_7),
    .io_memStreams_gathers_0_cmd_bits_addr_8(accel_io_memStreams_gathers_0_cmd_bits_addr_8),
    .io_memStreams_gathers_0_cmd_bits_addr_9(accel_io_memStreams_gathers_0_cmd_bits_addr_9),
    .io_memStreams_gathers_0_cmd_bits_addr_10(accel_io_memStreams_gathers_0_cmd_bits_addr_10),
    .io_memStreams_gathers_0_cmd_bits_addr_11(accel_io_memStreams_gathers_0_cmd_bits_addr_11),
    .io_memStreams_gathers_0_cmd_bits_addr_12(accel_io_memStreams_gathers_0_cmd_bits_addr_12),
    .io_memStreams_gathers_0_cmd_bits_addr_13(accel_io_memStreams_gathers_0_cmd_bits_addr_13),
    .io_memStreams_gathers_0_cmd_bits_addr_14(accel_io_memStreams_gathers_0_cmd_bits_addr_14),
    .io_memStreams_gathers_0_cmd_bits_addr_15(accel_io_memStreams_gathers_0_cmd_bits_addr_15),
    .io_memStreams_gathers_0_data_ready(accel_io_memStreams_gathers_0_data_ready),
    .io_memStreams_gathers_0_data_valid(accel_io_memStreams_gathers_0_data_valid),
    .io_memStreams_gathers_0_data_bits_0(accel_io_memStreams_gathers_0_data_bits_0),
    .io_memStreams_gathers_0_data_bits_1(accel_io_memStreams_gathers_0_data_bits_1),
    .io_memStreams_gathers_0_data_bits_2(accel_io_memStreams_gathers_0_data_bits_2),
    .io_memStreams_gathers_0_data_bits_3(accel_io_memStreams_gathers_0_data_bits_3),
    .io_memStreams_gathers_0_data_bits_4(accel_io_memStreams_gathers_0_data_bits_4),
    .io_memStreams_gathers_0_data_bits_5(accel_io_memStreams_gathers_0_data_bits_5),
    .io_memStreams_gathers_0_data_bits_6(accel_io_memStreams_gathers_0_data_bits_6),
    .io_memStreams_gathers_0_data_bits_7(accel_io_memStreams_gathers_0_data_bits_7),
    .io_memStreams_gathers_0_data_bits_8(accel_io_memStreams_gathers_0_data_bits_8),
    .io_memStreams_gathers_0_data_bits_9(accel_io_memStreams_gathers_0_data_bits_9),
    .io_memStreams_gathers_0_data_bits_10(accel_io_memStreams_gathers_0_data_bits_10),
    .io_memStreams_gathers_0_data_bits_11(accel_io_memStreams_gathers_0_data_bits_11),
    .io_memStreams_gathers_0_data_bits_12(accel_io_memStreams_gathers_0_data_bits_12),
    .io_memStreams_gathers_0_data_bits_13(accel_io_memStreams_gathers_0_data_bits_13),
    .io_memStreams_gathers_0_data_bits_14(accel_io_memStreams_gathers_0_data_bits_14),
    .io_memStreams_gathers_0_data_bits_15(accel_io_memStreams_gathers_0_data_bits_15),
    .io_memStreams_scatters_0_cmd_ready(accel_io_memStreams_scatters_0_cmd_ready),
    .io_memStreams_scatters_0_cmd_valid(accel_io_memStreams_scatters_0_cmd_valid),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_0(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_1(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_2(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_3(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_4(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_5(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_6(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_7(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_8(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_9(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_10(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_11(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_12(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_13(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_14(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_15(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15),
    .io_memStreams_scatters_0_cmd_bits_wdata_0(accel_io_memStreams_scatters_0_cmd_bits_wdata_0),
    .io_memStreams_scatters_0_cmd_bits_wdata_1(accel_io_memStreams_scatters_0_cmd_bits_wdata_1),
    .io_memStreams_scatters_0_cmd_bits_wdata_2(accel_io_memStreams_scatters_0_cmd_bits_wdata_2),
    .io_memStreams_scatters_0_cmd_bits_wdata_3(accel_io_memStreams_scatters_0_cmd_bits_wdata_3),
    .io_memStreams_scatters_0_cmd_bits_wdata_4(accel_io_memStreams_scatters_0_cmd_bits_wdata_4),
    .io_memStreams_scatters_0_cmd_bits_wdata_5(accel_io_memStreams_scatters_0_cmd_bits_wdata_5),
    .io_memStreams_scatters_0_cmd_bits_wdata_6(accel_io_memStreams_scatters_0_cmd_bits_wdata_6),
    .io_memStreams_scatters_0_cmd_bits_wdata_7(accel_io_memStreams_scatters_0_cmd_bits_wdata_7),
    .io_memStreams_scatters_0_cmd_bits_wdata_8(accel_io_memStreams_scatters_0_cmd_bits_wdata_8),
    .io_memStreams_scatters_0_cmd_bits_wdata_9(accel_io_memStreams_scatters_0_cmd_bits_wdata_9),
    .io_memStreams_scatters_0_cmd_bits_wdata_10(accel_io_memStreams_scatters_0_cmd_bits_wdata_10),
    .io_memStreams_scatters_0_cmd_bits_wdata_11(accel_io_memStreams_scatters_0_cmd_bits_wdata_11),
    .io_memStreams_scatters_0_cmd_bits_wdata_12(accel_io_memStreams_scatters_0_cmd_bits_wdata_12),
    .io_memStreams_scatters_0_cmd_bits_wdata_13(accel_io_memStreams_scatters_0_cmd_bits_wdata_13),
    .io_memStreams_scatters_0_cmd_bits_wdata_14(accel_io_memStreams_scatters_0_cmd_bits_wdata_14),
    .io_memStreams_scatters_0_cmd_bits_wdata_15(accel_io_memStreams_scatters_0_cmd_bits_wdata_15),
    .io_memStreams_scatters_0_wresp_ready(accel_io_memStreams_scatters_0_wresp_ready),
    .io_memStreams_scatters_0_wresp_valid(accel_io_memStreams_scatters_0_wresp_valid),
    .io_memStreams_scatters_0_wresp_bits(accel_io_memStreams_scatters_0_wresp_bits),
    .io_axiStreamsIn_0_TVALID(accel_io_axiStreamsIn_0_TVALID),
    .io_axiStreamsIn_0_TREADY(accel_io_axiStreamsIn_0_TREADY),
    .io_axiStreamsIn_0_TDATA(accel_io_axiStreamsIn_0_TDATA),
    .io_axiStreamsIn_0_TSTRB(accel_io_axiStreamsIn_0_TSTRB),
    .io_axiStreamsIn_0_TKEEP(accel_io_axiStreamsIn_0_TKEEP),
    .io_axiStreamsIn_0_TLAST(accel_io_axiStreamsIn_0_TLAST),
    .io_axiStreamsIn_0_TID(accel_io_axiStreamsIn_0_TID),
    .io_axiStreamsIn_0_TDEST(accel_io_axiStreamsIn_0_TDEST),
    .io_axiStreamsIn_0_TUSER(accel_io_axiStreamsIn_0_TUSER),
    .io_axiStreamsOut_0_TVALID(accel_io_axiStreamsOut_0_TVALID),
    .io_axiStreamsOut_0_TREADY(accel_io_axiStreamsOut_0_TREADY),
    .io_axiStreamsOut_0_TDATA(accel_io_axiStreamsOut_0_TDATA),
    .io_axiStreamsOut_0_TSTRB(accel_io_axiStreamsOut_0_TSTRB),
    .io_axiStreamsOut_0_TKEEP(accel_io_axiStreamsOut_0_TKEEP),
    .io_axiStreamsOut_0_TLAST(accel_io_axiStreamsOut_0_TLAST),
    .io_axiStreamsOut_0_TID(accel_io_axiStreamsOut_0_TID),
    .io_axiStreamsOut_0_TDEST(accel_io_axiStreamsOut_0_TDEST),
    .io_axiStreamsOut_0_TUSER(accel_io_axiStreamsOut_0_TUSER),
    .io_heap_0_req_valid(accel_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(accel_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(accel_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(accel_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(accel_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(accel_io_heap_0_resp_bits_sizeAddr),
    .io_argIns_0(accel_io_argIns_0),
    .io_argIns_1(accel_io_argIns_1),
    .io_argOuts_0_port_ready(accel_io_argOuts_0_port_ready),
    .io_argOuts_0_port_valid(accel_io_argOuts_0_port_valid),
    .io_argOuts_0_port_bits(accel_io_argOuts_0_port_bits),
    .io_argOuts_0_echo(accel_io_argOuts_0_echo)
  );
  assign io_rdata = 64'h0;
  assign accel_clock = clock; // @[:@26298.4]
  assign accel_reset = reset; // @[:@26299.4]
  assign accel_io_enable = 1'h0;
  assign accel_io_reset = 1'h0;
  assign accel_io_memStreams_loads_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_loads_0_data_valid = 1'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_0 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_1 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_2 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_3 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_4 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_5 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_6 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_7 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_8 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_9 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_10 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_11 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_12 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_13 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_14 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_15 = 32'h0;
  assign accel_io_memStreams_stores_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_stores_0_data_ready = 1'h0;
  assign accel_io_memStreams_stores_0_wresp_valid = 1'h0;
  assign accel_io_memStreams_stores_0_wresp_bits = 1'h0;
  assign accel_io_memStreams_gathers_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_gathers_0_data_valid = 1'h0;
  assign accel_io_memStreams_gathers_0_data_bits_0 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_1 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_2 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_3 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_4 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_5 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_6 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_7 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_8 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_9 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_10 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_11 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_12 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_13 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_14 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_15 = 32'h0;
  assign accel_io_memStreams_scatters_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_scatters_0_wresp_valid = 1'h0;
  assign accel_io_memStreams_scatters_0_wresp_bits = 1'h0;
  assign accel_io_axiStreamsIn_0_TVALID = 1'h0;
  assign accel_io_axiStreamsIn_0_TDATA = 256'h0;
  assign accel_io_axiStreamsIn_0_TSTRB = 32'h0;
  assign accel_io_axiStreamsIn_0_TKEEP = 32'h0;
  assign accel_io_axiStreamsIn_0_TLAST = 1'h0;
  assign accel_io_axiStreamsIn_0_TID = 8'h0;
  assign accel_io_axiStreamsIn_0_TDEST = 8'h0;
  assign accel_io_axiStreamsIn_0_TUSER = 32'h0;
  assign accel_io_axiStreamsOut_0_TREADY = 1'h0;
  assign accel_io_heap_0_resp_valid = 1'h0;
  assign accel_io_heap_0_resp_bits_allocDealloc = 1'h0;
  assign accel_io_heap_0_resp_bits_sizeAddr = 64'h0;
  assign accel_io_argIns_0 = 64'h0;
  assign accel_io_argIns_1 = 64'h0;
  assign accel_io_argOuts_0_port_ready = 1'h0;
  assign accel_io_argOuts_0_echo = 64'h0;
endmodule
