// Latency = 4
module Top(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  input  [7:0] I_2,
  input  [7:0] I_3,
  input  [7:0] I_4,
  input  [7:0] I_5,
  input  [7:0] I_6,
  input  [7:0] I_7,
  output [7:0] O_0_0_0,
  output [7:0] O_1_0_0,
  output [7:0] O_2_0_0,
  output [7:0] O_3_0_0,
  output [7:0] O_4_0_0,
  output [7:0] O_5_0_0,
  output [7:0] O_6_0_0,
  output [7:0] O_7_0_0
);
  wire dontcare;
  wire [31:0] io_output_counts_1;
  wire [31:0] io_output_counts_0;

  x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1 sampler_box ( // @[m_x55_ctr_0.scala 26:17:@1721.4]
    .clock(CLKclock), // @[:@1296.4]
    .reset('b0), // @[:@1297.4]
    .io_in_x426_TREADY(dontcare), // @[:@1298.4]
    .io_in_x426_TDATA({I_0,I_1,I_2,I_3,I_4,I_5,I_6,I_7}), // @[:@1298.4]
    .io_in_x426_TID(8'h0),
    .io_in_x426_TDEST(8'h0),
    .io_in_x427_TVALID(valid_down), // @[:@1298.4]
    .io_in_x427_TDATA({O_0_0_0,O_1_0_0,O_2_0_0,O_3_0_0,O_4_0_0,O_5_0_0,O_6_0_0,O_7_0_0}), // @[:@1298.4]
    .io_in_x427_TREADY(1'b1), // @[:@1298.4]
    .io_sigsIn_datapathEn(valid_up), // @[:@1298.4]
    .io_sigsIn_backpressure(1'b1), // @[:@20563.4]
    .io_sigsIn_break(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_1(io_output_counts_1), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_0(io_output_counts_0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_0(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_1(1'b0), // @[:@20563.4]
    .io_rr('b1) // @[:@1298.4]
  );

  wire dontcare2;

  wire io_output_oobs_0;
  wire io_output_oobs_1;
  x434_ctrchain cchain ( // @[:@2879.2]
    .clock(clock), // @[:@2880.4]
    .reset(1'b0), // @[:@2881.4]
    .io_input_reset(1'b0), // @[:@2882.4]
    .io_input_enable(valid_up), // @[:@2882.4]
    .io_output_counts_1(io_output_counts_1), // @[:@2882.4]
    .io_output_counts_0(io_output_counts_0), // @[:@2882.4]
    .io_output_oobs_0(io_output_oobs_0), // @[:@2882.4]
    .io_output_oobs_1(io_output_oobs_1), // @[:@2882.4]
    .io_output_done(dontcare2) // @[:@2882.4]
  );

endmodule

module SRAMVerilogSim
#(
    parameter WORDS = 1024,
    parameter AWIDTH = 10,
    parameter DWIDTH = 32)
(
    input clk,
    input [AWIDTH-1:0] raddr,
    input [AWIDTH-1:0] waddr,
    input raddrEn,
    input waddrEn,
    input wen,
    input [DWIDTH-1:0] wdata,
    input backpressure,
    output reg [DWIDTH-1:0] rdata
);

    reg [DWIDTH-1:0] mem [0:WORDS-1];

    always @(posedge clk) begin
      if (wen) mem[waddr] <= wdata;
      if (backpressure) rdata <= mem[raddr];
    end

endmodule
module RetimeShiftRegister
#(
    parameter WIDTH = 1,
    parameter STAGES = 1)
(
    input clock,
    input reset,
    input flow,
    input [WIDTH-1:0] init,
    input [WIDTH-1:0] in,
    output reg [WIDTH-1:0] out
);
  integer i;
  reg [WIDTH-1:0] sr[STAGES:0]; // Create 'STAGES' number of register, each 'WIDTH' bits wide

   /* synopsys dc_tcl_script_begin
    set_ungroup [current_design] true
    set_flatten true -effort high -phase true -design [current_design]
    set_dont_retime [current_design] false
    set_optimize_registers true -design [current_design]
    */
  always @(posedge clock) begin
    if (reset) begin
      for(i=0; i<STAGES; i=i+1) begin
        sr[i] <= init;
      end
    end else begin
      if (flow) begin 
        sr[0] <= in;
        for(i=1; i<STAGES; i=i+1) begin
          sr[i] <= sr[i-1];
        end
      end
    end
  end

  always @(*) begin
    out = sr[STAGES-1];
  end
endmodule
module FF( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  output [31:0] io_rPort_0_output_0, // @[:@6.4]
  input  [31:0] io_wPort_0_data_0, // @[:@6.4]
  input         io_wPort_0_reset, // @[:@6.4]
  input         io_wPort_0_en_0 // @[:@6.4]
);
  reg [31:0] ff; // @[MemPrimitives.scala 173:19:@21.4]
  reg [31:0] _RAND_0;
  wire [31:0] _T_68; // @[MemPrimitives.scala 177:32:@23.4]
  wire [31:0] _T_69; // @[MemPrimitives.scala 177:12:@24.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 177:32:@23.4]
  assign _T_69 = io_wPort_0_reset ? 32'h0 : _T_68; // @[MemPrimitives.scala 177:12:@24.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 178:34:@26.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 32'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 32'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SRFF( // @[:@28.2]
  input   clock, // @[:@29.4]
  input   reset, // @[:@30.4]
  input   io_input_set, // @[:@31.4]
  input   io_input_reset, // @[:@31.4]
  input   io_input_asyn_reset, // @[:@31.4]
  output  io_output // @[:@31.4]
);
  reg  _T_15; // @[SRFF.scala 20:21:@33.4]
  reg [31:0] _RAND_0;
  wire  _T_19; // @[SRFF.scala 21:74:@34.4]
  wire  _T_20; // @[SRFF.scala 21:48:@35.4]
  wire  _T_21; // @[SRFF.scala 21:14:@36.4]
  assign _T_19 = io_input_reset ? 1'h0 : _T_15; // @[SRFF.scala 21:74:@34.4]
  assign _T_20 = io_input_set ? 1'h1 : _T_19; // @[SRFF.scala 21:48:@35.4]
  assign _T_21 = io_input_asyn_reset ? 1'h0 : _T_20; // @[SRFF.scala 21:14:@36.4]
  assign io_output = io_input_asyn_reset ? 1'h0 : _T_15; // @[SRFF.scala 22:15:@39.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_15 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_15 <= 1'h0;
    end else begin
      if (io_input_asyn_reset) begin
        _T_15 <= 1'h0;
      end else begin
        if (io_input_set) begin
          _T_15 <= 1'h1;
        end else begin
          if (io_input_reset) begin
            _T_15 <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module SingleCounter( // @[:@41.2]
  input   clock, // @[:@42.4]
  input   reset, // @[:@43.4]
  input   io_input_reset, // @[:@44.4]
  output  io_output_done // @[:@44.4]
);
  wire  bases_0_clock; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_reset; // @[Counter.scala 253:53:@57.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 253:53:@57.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 253:53:@57.4]
  wire  SRFF_clock; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_set; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_output; // @[Counter.scala 255:22:@73.4]
  wire [12:0] _T_48; // @[Counter.scala 279:52:@101.4]
  wire [13:0] _T_50; // @[Counter.scala 283:33:@102.4]
  wire [12:0] _T_51; // @[Counter.scala 283:33:@103.4]
  wire [12:0] _T_52; // @[Counter.scala 283:33:@104.4]
  wire  _T_57; // @[Counter.scala 285:18:@106.4]
  wire [12:0] _T_68; // @[Counter.scala 291:115:@114.4]
  wire [12:0] _T_71; // @[Counter.scala 291:152:@117.4]
  wire [12:0] _T_72; // @[Counter.scala 291:74:@118.4]
  FF bases_0 ( // @[Counter.scala 253:53:@57.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 255:22:@73.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 279:52:@101.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@102.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@103.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 283:33:@104.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh13); // @[Counter.scala 285:18:@106.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 291:115:@114.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 291:152:@117.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 291:74:@118.4]
  assign io_output_done = $signed(_T_52) >= $signed(32'sh13); // @[Counter.scala 325:20:@127.4]
  assign bases_0_clock = clock; // @[:@58.4]
  assign bases_0_reset = reset; // @[:@59.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 291:31:@120.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 273:27:@99.4]
  assign bases_0_io_wPort_0_en_0 = 1'h1; // @[Counter.scala 276:29:@100.4]
  assign SRFF_clock = clock; // @[:@74.4]
  assign SRFF_reset = reset; // @[:@75.4]
  assign SRFF_io_input_set = io_input_reset == 1'h0; // @[Counter.scala 256:23:@78.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 257:25:@80.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 258:30:@81.4]
endmodule
module RetimeWrapper( // @[:@144.2]
  input   clock, // @[:@145.4]
  input   reset, // @[:@146.4]
  input   io_flow, // @[:@147.4]
  input   io_in, // @[:@147.4]
  output  io_out // @[:@147.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@149.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@149.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@162.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@161.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@160.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@159.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@158.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@156.4]
endmodule
module RootController_sm( // @[:@312.2]
  input   clock, // @[:@313.4]
  input   reset, // @[:@314.4]
  input   io_enable, // @[:@315.4]
  output  io_done, // @[:@315.4]
  input   io_rst, // @[:@315.4]
  input   io_ctrDone, // @[:@315.4]
  output  io_ctrInc, // @[:@315.4]
  input   io_doneIn_0, // @[:@315.4]
  output  io_enableOut_0, // @[:@315.4]
  output  io_childAck_0 // @[:@315.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@318.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@321.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@338.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@433.4]
  wire  finished; // @[Controllers.scala 81:26:@324.4]
  wire  synchronize; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  wire  _T_122; // @[Controllers.scala 128:33:@371.4]
  wire  _T_124; // @[Controllers.scala 128:54:@372.4]
  wire  _T_125; // @[Controllers.scala 128:52:@373.4]
  wire  _T_126; // @[Controllers.scala 128:66:@374.4]
  wire  _T_128; // @[Controllers.scala 128:98:@376.4]
  wire  _T_129; // @[Controllers.scala 128:96:@377.4]
  wire  _T_131; // @[Controllers.scala 128:123:@378.4]
  wire  _T_133; // @[Controllers.scala 129:48:@381.4]
  wire  _T_138; // @[Controllers.scala 130:52:@386.4]
  wire  _T_139; // @[Controllers.scala 130:50:@387.4]
  wire  _T_147; // @[Controllers.scala 130:129:@393.4]
  wire  _T_150; // @[Controllers.scala 131:45:@396.4]
  wire  _T_154; // @[Controllers.scala 213:68:@402.4]
  wire  _T_156; // @[Controllers.scala 213:90:@404.4]
  wire  _T_158; // @[Controllers.scala 213:132:@406.4]
  wire  _T_159; // @[Controllers.scala 213:130:@407.4]
  wire  _T_160; // @[Controllers.scala 213:156:@408.4]
  reg  _T_166; // @[package.scala 48:56:@412.4]
  reg [31:0] _RAND_0;
  reg  _T_180; // @[package.scala 48:56:@430.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@318.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@321.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@338.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@357.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@416.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@433.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  assign finished = done_0_io_output | io_done; // @[Controllers.scala 81:26:@324.4]
  assign synchronize = RetimeWrapper_io_out; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  assign _T_122 = done_0_io_output == 1'h0; // @[Controllers.scala 128:33:@371.4]
  assign _T_124 = io_ctrDone == 1'h0; // @[Controllers.scala 128:54:@372.4]
  assign _T_125 = _T_122 & _T_124; // @[Controllers.scala 128:52:@373.4]
  assign _T_126 = _T_125 & io_enable; // @[Controllers.scala 128:66:@374.4]
  assign _T_128 = ~ iterDone_0_io_output; // @[Controllers.scala 128:98:@376.4]
  assign _T_129 = _T_126 & _T_128; // @[Controllers.scala 128:96:@377.4]
  assign _T_131 = io_doneIn_0 == 1'h0; // @[Controllers.scala 128:123:@378.4]
  assign _T_133 = io_doneIn_0 | io_rst; // @[Controllers.scala 129:48:@381.4]
  assign _T_138 = synchronize == 1'h0; // @[Controllers.scala 130:52:@386.4]
  assign _T_139 = io_doneIn_0 & _T_138; // @[Controllers.scala 130:50:@387.4]
  assign _T_147 = finished == 1'h0; // @[Controllers.scala 130:129:@393.4]
  assign _T_150 = io_rst == 1'h0; // @[Controllers.scala 131:45:@396.4]
  assign _T_154 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@402.4]
  assign _T_156 = _T_154 & _T_128; // @[Controllers.scala 213:90:@404.4]
  assign _T_158 = ~ done_0_io_output; // @[Controllers.scala 213:132:@406.4]
  assign _T_159 = _T_156 & _T_158; // @[Controllers.scala 213:130:@407.4]
  assign _T_160 = ~ io_ctrDone; // @[Controllers.scala 213:156:@408.4]
  assign io_done = RetimeWrapper_2_io_out; // @[Controllers.scala 245:13:@440.4]
  assign io_ctrInc = io_doneIn_0; // @[Controllers.scala 122:17:@356.4]
  assign io_enableOut_0 = _T_159 & _T_160; // @[Controllers.scala 213:55:@410.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@401.4]
  assign active_0_clock = clock; // @[:@319.4]
  assign active_0_reset = reset; // @[:@320.4]
  assign active_0_io_input_set = _T_129 & _T_131; // @[Controllers.scala 128:30:@380.4]
  assign active_0_io_input_reset = _T_133 | done_0_io_output; // @[Controllers.scala 129:32:@385.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@326.4]
  assign done_0_clock = clock; // @[:@322.4]
  assign done_0_reset = reset; // @[:@323.4]
  assign done_0_io_input_set = io_ctrDone & _T_150; // @[Controllers.scala 131:28:@399.4]
  assign done_0_io_input_reset = io_rst | done_0_io_output; // @[Controllers.scala 86:33:@336.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@327.4]
  assign iterDone_0_clock = clock; // @[:@339.4]
  assign iterDone_0_reset = reset; // @[:@340.4]
  assign iterDone_0_io_input_set = _T_139 & _T_147; // @[Controllers.scala 130:32:@395.4]
  assign iterDone_0_io_input_reset = synchronize | io_rst; // @[Controllers.scala 92:37:@350.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@341.4]
  assign RetimeWrapper_clock = clock; // @[:@358.4]
  assign RetimeWrapper_reset = reset; // @[:@359.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@361.4]
  assign RetimeWrapper_io_in = io_doneIn_0; // @[package.scala 94:16:@360.4]
  assign RetimeWrapper_1_clock = clock; // @[:@417.4]
  assign RetimeWrapper_1_reset = reset; // @[:@418.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@420.4]
  assign RetimeWrapper_1_io_in = done_0_io_output & _T_166; // @[package.scala 94:16:@419.4]
  assign RetimeWrapper_2_clock = clock; // @[:@434.4]
  assign RetimeWrapper_2_reset = reset; // @[:@435.4]
  assign RetimeWrapper_2_io_flow = io_enable; // @[package.scala 95:18:@437.4]
  assign RetimeWrapper_2_io_in = done_0_io_output & _T_180; // @[package.scala 94:16:@436.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_166 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_180 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_166 <= 1'h0;
    end else begin
      _T_166 <= _T_122;
    end
    if (reset) begin
      _T_180 <= 1'h0;
    end else begin
      _T_180 <= _T_122;
    end
  end
endmodule
module x825_outr_UnitPipe_sm( // @[:@2389.2]
  input   clock, // @[:@2390.4]
  input   reset, // @[:@2391.4]
  input   io_enable, // @[:@2392.4]
  output  io_done, // @[:@2392.4]
  input   io_parentAck, // @[:@2392.4]
  input   io_doneIn_0, // @[:@2392.4]
  output  io_enableOut_0, // @[:@2392.4]
  output  io_childAck_0, // @[:@2392.4]
  input   io_ctrCopyDone_0 // @[:@2392.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@2395.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@2395.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@2395.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@2395.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@2395.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@2395.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@2398.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@2398.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@2398.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@2398.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@2398.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@2398.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@2415.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@2415.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@2415.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@2415.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@2415.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@2415.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@2446.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@2446.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@2446.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@2446.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@2446.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@2460.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@2460.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@2460.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@2460.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@2460.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@2478.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@2478.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@2478.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@2478.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@2478.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@2515.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@2515.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@2515.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@2515.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@2515.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@2532.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@2532.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@2532.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@2532.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@2532.4]
  wire  _T_105; // @[Controllers.scala 165:35:@2430.4]
  wire  _T_107; // @[Controllers.scala 165:60:@2431.4]
  wire  _T_108; // @[Controllers.scala 165:58:@2432.4]
  wire  _T_110; // @[Controllers.scala 165:76:@2433.4]
  wire  _T_111; // @[Controllers.scala 165:74:@2434.4]
  wire  _T_115; // @[Controllers.scala 165:109:@2437.4]
  wire  _T_118; // @[Controllers.scala 165:141:@2439.4]
  wire  _T_126; // @[package.scala 96:25:@2451.4 package.scala 96:25:@2452.4]
  wire  _T_130; // @[Controllers.scala 167:54:@2454.4]
  wire  _T_131; // @[Controllers.scala 167:52:@2455.4]
  wire  _T_138; // @[package.scala 96:25:@2465.4 package.scala 96:25:@2466.4]
  wire  _T_156; // @[package.scala 96:25:@2483.4 package.scala 96:25:@2484.4]
  wire  _T_160; // @[Controllers.scala 169:67:@2486.4]
  wire  _T_161; // @[Controllers.scala 169:86:@2487.4]
  wire  _T_174; // @[Controllers.scala 213:68:@2501.4]
  wire  _T_176; // @[Controllers.scala 213:90:@2503.4]
  wire  _T_178; // @[Controllers.scala 213:132:@2505.4]
  reg  _T_186; // @[package.scala 48:56:@2511.4]
  reg [31:0] _RAND_0;
  wire  _T_187; // @[package.scala 100:41:@2513.4]
  reg  _T_200; // @[package.scala 48:56:@2529.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@2395.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@2398.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@2415.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@2446.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@2460.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@2478.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@2515.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@2532.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_105 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@2430.4]
  assign _T_107 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@2431.4]
  assign _T_108 = _T_105 & _T_107; // @[Controllers.scala 165:58:@2432.4]
  assign _T_110 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@2433.4]
  assign _T_111 = _T_108 & _T_110; // @[Controllers.scala 165:74:@2434.4]
  assign _T_115 = _T_111 & io_enable; // @[Controllers.scala 165:109:@2437.4]
  assign _T_118 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@2439.4]
  assign _T_126 = RetimeWrapper_io_out; // @[package.scala 96:25:@2451.4 package.scala 96:25:@2452.4]
  assign _T_130 = _T_126 == 1'h0; // @[Controllers.scala 167:54:@2454.4]
  assign _T_131 = io_doneIn_0 | _T_130; // @[Controllers.scala 167:52:@2455.4]
  assign _T_138 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@2465.4 package.scala 96:25:@2466.4]
  assign _T_156 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@2483.4 package.scala 96:25:@2484.4]
  assign _T_160 = _T_156 == 1'h0; // @[Controllers.scala 169:67:@2486.4]
  assign _T_161 = _T_160 & io_enable; // @[Controllers.scala 169:86:@2487.4]
  assign _T_174 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@2501.4]
  assign _T_176 = _T_174 & _T_105; // @[Controllers.scala 213:90:@2503.4]
  assign _T_178 = ~ done_0_io_output; // @[Controllers.scala 213:132:@2505.4]
  assign _T_187 = done_0_io_output & _T_186; // @[package.scala 100:41:@2513.4]
  assign io_done = RetimeWrapper_4_io_out; // @[Controllers.scala 245:13:@2539.4]
  assign io_enableOut_0 = _T_176 & _T_178; // @[Controllers.scala 213:55:@2509.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@2500.4]
  assign active_0_clock = clock; // @[:@2396.4]
  assign active_0_reset = reset; // @[:@2397.4]
  assign active_0_io_input_set = _T_115 & _T_118; // @[Controllers.scala 165:32:@2441.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@2445.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@2403.4]
  assign done_0_clock = clock; // @[:@2399.4]
  assign done_0_reset = reset; // @[:@2400.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_161; // @[Controllers.scala 169:30:@2491.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@2413.4 Controllers.scala 170:32:@2498.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@2404.4]
  assign iterDone_0_clock = clock; // @[:@2416.4]
  assign iterDone_0_reset = reset; // @[:@2417.4]
  assign iterDone_0_io_input_set = _T_131 & io_enable; // @[Controllers.scala 167:34:@2459.4]
  assign iterDone_0_io_input_reset = _T_138 | io_parentAck; // @[Controllers.scala 92:37:@2427.4 Controllers.scala 168:36:@2475.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@2418.4]
  assign RetimeWrapper_clock = clock; // @[:@2447.4]
  assign RetimeWrapper_reset = reset; // @[:@2448.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@2450.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@2449.4]
  assign RetimeWrapper_1_clock = clock; // @[:@2461.4]
  assign RetimeWrapper_1_reset = reset; // @[:@2462.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@2464.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@2463.4]
  assign RetimeWrapper_2_clock = clock; // @[:@2479.4]
  assign RetimeWrapper_2_reset = reset; // @[:@2480.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@2482.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@2481.4]
  assign RetimeWrapper_3_clock = clock; // @[:@2516.4]
  assign RetimeWrapper_3_reset = reset; // @[:@2517.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@2519.4]
  assign RetimeWrapper_3_io_in = _T_187 | io_parentAck; // @[package.scala 94:16:@2518.4]
  assign RetimeWrapper_4_clock = clock; // @[:@2533.4]
  assign RetimeWrapper_4_reset = reset; // @[:@2534.4]
  assign RetimeWrapper_4_io_flow = io_enable; // @[package.scala 95:18:@2536.4]
  assign RetimeWrapper_4_io_in = done_0_io_output & _T_200; // @[package.scala 94:16:@2535.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_186 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_200 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_186 <= 1'h0;
    end else begin
      _T_186 <= _T_110;
    end
    if (reset) begin
      _T_200 <= 1'h0;
    end else begin
      _T_200 <= _T_110;
    end
  end
endmodule
module SingleCounter_1( // @[:@2659.2]
  input         clock, // @[:@2660.4]
  input         reset, // @[:@2661.4]
  input         io_input_reset, // @[:@2662.4]
  input         io_input_enable, // @[:@2662.4]
  output [31:0] io_output_count_0, // @[:@2662.4]
  output        io_output_oobs_0, // @[:@2662.4]
  output        io_output_done, // @[:@2662.4]
  output        io_output_saturated // @[:@2662.4]
);
  wire  bases_0_clock; // @[Counter.scala 253:53:@2675.4]
  wire  bases_0_reset; // @[Counter.scala 253:53:@2675.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 253:53:@2675.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 253:53:@2675.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 253:53:@2675.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 253:53:@2675.4]
  wire  SRFF_clock; // @[Counter.scala 255:22:@2691.4]
  wire  SRFF_reset; // @[Counter.scala 255:22:@2691.4]
  wire  SRFF_io_input_set; // @[Counter.scala 255:22:@2691.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 255:22:@2691.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 255:22:@2691.4]
  wire  SRFF_io_output; // @[Counter.scala 255:22:@2691.4]
  wire  _T_36; // @[Counter.scala 256:45:@2694.4]
  wire [12:0] _T_48; // @[Counter.scala 279:52:@2719.4]
  wire [13:0] _T_50; // @[Counter.scala 283:33:@2720.4]
  wire [12:0] _T_51; // @[Counter.scala 283:33:@2721.4]
  wire [12:0] _T_52; // @[Counter.scala 283:33:@2722.4]
  wire  _T_57; // @[Counter.scala 285:18:@2724.4]
  wire [12:0] _T_68; // @[Counter.scala 291:115:@2732.4]
  wire [12:0] _T_71; // @[Counter.scala 291:152:@2735.4]
  wire [12:0] _T_72; // @[Counter.scala 291:74:@2736.4]
  wire  _T_75; // @[Counter.scala 314:102:@2740.4]
  wire  _T_77; // @[Counter.scala 314:130:@2741.4]
  FF bases_0 ( // @[Counter.scala 253:53:@2675.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 255:22:@2691.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 256:45:@2694.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 279:52:@2719.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh2); // @[Counter.scala 283:33:@2720.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh2); // @[Counter.scala 283:33:@2721.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 283:33:@2722.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh4); // @[Counter.scala 285:18:@2724.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 291:115:@2732.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 291:152:@2735.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 291:74:@2736.4]
  assign _T_75 = $signed(_T_48) < $signed(32'sh0); // @[Counter.scala 314:102:@2740.4]
  assign _T_77 = $signed(_T_48) >= $signed(32'sh4); // @[Counter.scala 314:130:@2741.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 296:28:@2739.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 314:60:@2743.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 325:20:@2745.4]
  assign io_output_saturated = $signed(_T_52) >= $signed(32'sh4); // @[Counter.scala 332:25:@2748.4]
  assign bases_0_clock = clock; // @[:@2676.4]
  assign bases_0_reset = reset; // @[:@2677.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 291:31:@2738.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 273:27:@2717.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 276:29:@2718.4]
  assign SRFF_clock = clock; // @[:@2692.4]
  assign SRFF_reset = reset; // @[:@2693.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 256:23:@2696.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 257:25:@2698.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 258:30:@2699.4]
endmodule
module SingleCounter_2( // @[:@2788.2]
  input         clock, // @[:@2789.4]
  input         reset, // @[:@2790.4]
  input         io_setup_saturate, // @[:@2791.4]
  input         io_input_reset, // @[:@2791.4]
  input         io_input_enable, // @[:@2791.4]
  output [31:0] io_output_count_0, // @[:@2791.4]
  output        io_output_oobs_0, // @[:@2791.4]
  output        io_output_done // @[:@2791.4]
);
  wire  bases_0_clock; // @[Counter.scala 253:53:@2804.4]
  wire  bases_0_reset; // @[Counter.scala 253:53:@2804.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 253:53:@2804.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 253:53:@2804.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 253:53:@2804.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 253:53:@2804.4]
  wire  SRFF_clock; // @[Counter.scala 255:22:@2820.4]
  wire  SRFF_reset; // @[Counter.scala 255:22:@2820.4]
  wire  SRFF_io_input_set; // @[Counter.scala 255:22:@2820.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 255:22:@2820.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 255:22:@2820.4]
  wire  SRFF_io_output; // @[Counter.scala 255:22:@2820.4]
  wire  _T_36; // @[Counter.scala 256:45:@2823.4]
  wire [12:0] _T_48; // @[Counter.scala 279:52:@2848.4]
  wire [13:0] _T_50; // @[Counter.scala 283:33:@2849.4]
  wire [12:0] _T_51; // @[Counter.scala 283:33:@2850.4]
  wire [12:0] _T_52; // @[Counter.scala 283:33:@2851.4]
  wire  _T_57; // @[Counter.scala 285:18:@2853.4]
  wire [12:0] _T_68; // @[Counter.scala 291:115:@2861.4]
  wire [12:0] _T_70; // @[Counter.scala 291:85:@2863.4]
  wire [12:0] _T_71; // @[Counter.scala 291:152:@2864.4]
  wire [12:0] _T_72; // @[Counter.scala 291:74:@2865.4]
  wire  _T_75; // @[Counter.scala 314:102:@2869.4]
  wire  _T_77; // @[Counter.scala 314:130:@2870.4]
  FF bases_0 ( // @[Counter.scala 253:53:@2804.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 255:22:@2820.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 256:45:@2823.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 279:52:@2848.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh4); // @[Counter.scala 283:33:@2849.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh4); // @[Counter.scala 283:33:@2850.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 283:33:@2851.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh4); // @[Counter.scala 285:18:@2853.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 291:115:@2861.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 32'h0; // @[Counter.scala 291:85:@2863.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 291:152:@2864.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 291:74:@2865.4]
  assign _T_75 = $signed(_T_48) < $signed(32'sh0); // @[Counter.scala 314:102:@2869.4]
  assign _T_77 = $signed(_T_48) >= $signed(32'sh4); // @[Counter.scala 314:130:@2870.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 296:28:@2868.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 314:60:@2872.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 325:20:@2874.4]
  assign bases_0_clock = clock; // @[:@2805.4]
  assign bases_0_reset = reset; // @[:@2806.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 291:31:@2867.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 273:27:@2846.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 276:29:@2847.4]
  assign SRFF_clock = clock; // @[:@2821.4]
  assign SRFF_reset = reset; // @[:@2822.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 256:23:@2825.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 257:25:@2827.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 258:30:@2828.4]
endmodule
module x434_ctrchain( // @[:@2879.2]
  input         clock, // @[:@2880.4]
  input         reset, // @[:@2881.4]
  input         io_input_reset, // @[:@2882.4]
  input         io_input_enable, // @[:@2882.4]
  output [31:0] io_output_counts_1, // @[:@2882.4]
  output [31:0] io_output_counts_0, // @[:@2882.4]
  output        io_output_oobs_0, // @[:@2882.4]
  output        io_output_oobs_1, // @[:@2882.4]
  output        io_output_done // @[:@2882.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_reset; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 505:46:@2884.4]
  wire [31:0] ctrs_0_io_output_count_0; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_io_output_saturated; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_1_clock; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_reset; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_io_setup_saturate; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_io_input_reset; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_io_input_enable; // @[Counter.scala 505:46:@2887.4]
  wire [31:0] ctrs_1_io_output_count_0; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_io_output_oobs_0; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_io_output_done; // @[Counter.scala 505:46:@2887.4]
  wire  isDone; // @[Counter.scala 533:51:@2904.4]
  reg  wasDone; // @[Counter.scala 534:24:@2905.4]
  reg [31:0] _RAND_0;
  wire  _T_64; // @[Counter.scala 538:69:@2913.4]
  wire  _T_66; // @[Counter.scala 538:80:@2914.4]
  reg  doneLatch; // @[Counter.scala 542:26:@2919.4]
  reg [31:0] _RAND_1;
  wire  _T_73; // @[Counter.scala 543:48:@2920.4]
  wire  _T_74; // @[Counter.scala 543:19:@2921.4]
  SingleCounter_1 ctrs_0 ( // @[Counter.scala 505:46:@2884.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done),
    .io_output_saturated(ctrs_0_io_output_saturated)
  );
  SingleCounter_2 ctrs_1 ( // @[Counter.scala 505:46:@2887.4]
    .clock(ctrs_1_clock),
    .reset(ctrs_1_reset),
    .io_setup_saturate(ctrs_1_io_setup_saturate),
    .io_input_reset(ctrs_1_io_input_reset),
    .io_input_enable(ctrs_1_io_input_enable),
    .io_output_count_0(ctrs_1_io_output_count_0),
    .io_output_oobs_0(ctrs_1_io_output_oobs_0),
    .io_output_done(ctrs_1_io_output_done)
  );
  assign isDone = ctrs_0_io_output_done & ctrs_1_io_output_done; // @[Counter.scala 533:51:@2904.4]
  assign _T_64 = io_input_enable & isDone; // @[Counter.scala 538:69:@2913.4]
  assign _T_66 = wasDone == 1'h0; // @[Counter.scala 538:80:@2914.4]
  assign _T_73 = isDone ? 1'h1 : doneLatch; // @[Counter.scala 543:48:@2920.4]
  assign _T_74 = io_input_reset ? 1'h0 : _T_73; // @[Counter.scala 543:19:@2921.4]
  assign io_output_counts_1 = ctrs_1_io_output_count_0; // @[Counter.scala 549:32:@2926.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 549:32:@2923.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 550:30:@2925.4]
  assign io_output_oobs_1 = ctrs_1_io_output_oobs_0 | doneLatch; // @[Counter.scala 550:30:@2928.4]
  assign io_output_done = _T_64 & _T_66; // @[Counter.scala 538:18:@2916.4]
  assign ctrs_0_clock = clock; // @[:@2885.4]
  assign ctrs_0_reset = reset; // @[:@2886.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 512:24:@2893.4]
  assign ctrs_0_io_input_enable = ctrs_1_io_output_done & io_input_enable; // @[Counter.scala 518:29:@2900.4]
  assign ctrs_1_clock = clock; // @[:@2888.4]
  assign ctrs_1_reset = reset; // @[:@2889.4]
  assign ctrs_1_io_setup_saturate = ctrs_0_io_output_saturated; // @[Counter.scala 524:31:@2903.4]
  assign ctrs_1_io_input_reset = io_input_reset; // @[Counter.scala 512:24:@2897.4]
  assign ctrs_1_io_input_enable = io_input_enable; // @[Counter.scala 516:33:@2898.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= isDone;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (isDone) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module RetimeWrapper_12( // @[:@2968.2]
  input   clock, // @[:@2969.4]
  input   reset, // @[:@2970.4]
  input   io_flow, // @[:@2971.4]
  input   io_in, // @[:@2971.4]
  output  io_out // @[:@2971.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(19)) sr ( // @[RetimeShiftRegister.scala 15:20:@2973.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@2986.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@2985.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@2984.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@2983.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@2982.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@2980.4]
endmodule
module RetimeWrapper_16( // @[:@3096.2]
  input   clock, // @[:@3097.4]
  input   reset, // @[:@3098.4]
  input   io_flow, // @[:@3099.4]
  input   io_in, // @[:@3099.4]
  output  io_out // @[:@3099.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(18)) sr ( // @[RetimeShiftRegister.scala 15:20:@3101.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3114.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3113.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3112.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3111.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3110.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3108.4]
endmodule
module x824_inr_Foreach_SAMPLER_BOX_sm( // @[:@3116.2]
  input   clock, // @[:@3117.4]
  input   reset, // @[:@3118.4]
  input   io_enable, // @[:@3119.4]
  output  io_done, // @[:@3119.4]
  output  io_doneLatch, // @[:@3119.4]
  input   io_ctrDone, // @[:@3119.4]
  output  io_datapathEn, // @[:@3119.4]
  output  io_ctrInc, // @[:@3119.4]
  output  io_ctrRst, // @[:@3119.4]
  input   io_parentAck, // @[:@3119.4]
  input   io_backpressure, // @[:@3119.4]
  input   io_break // @[:@3119.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@3121.4]
  wire  active_reset; // @[Controllers.scala 261:22:@3121.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@3121.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@3121.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@3121.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@3121.4]
  wire  done_clock; // @[Controllers.scala 262:20:@3124.4]
  wire  done_reset; // @[Controllers.scala 262:20:@3124.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@3124.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@3124.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@3124.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@3124.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3158.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3158.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3158.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@3158.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@3158.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@3180.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@3180.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@3180.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@3180.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@3180.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@3192.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@3192.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@3192.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@3192.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@3192.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@3200.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@3200.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@3200.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@3200.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@3200.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@3216.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@3216.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@3216.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@3216.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@3216.4]
  wire  _T_80; // @[Controllers.scala 264:48:@3129.4]
  wire  _T_81; // @[Controllers.scala 264:46:@3130.4]
  wire  _T_82; // @[Controllers.scala 264:62:@3131.4]
  wire  _T_83; // @[Controllers.scala 264:60:@3132.4]
  wire  _T_100; // @[package.scala 100:49:@3149.4]
  reg  _T_103; // @[package.scala 48:56:@3150.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@3163.4 package.scala 96:25:@3164.4]
  wire  _T_110; // @[package.scala 100:49:@3165.4]
  reg  _T_113; // @[package.scala 48:56:@3166.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@3168.4]
  wire  _T_118; // @[Controllers.scala 283:41:@3173.4]
  wire  _T_119; // @[Controllers.scala 283:59:@3174.4]
  wire  _T_121; // @[Controllers.scala 284:37:@3177.4]
  wire  _T_124; // @[package.scala 96:25:@3185.4 package.scala 96:25:@3186.4]
  wire  _T_126; // @[package.scala 100:49:@3187.4]
  reg  _T_129; // @[package.scala 48:56:@3188.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@3210.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@3212.4]
  reg  _T_153; // @[package.scala 48:56:@3213.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@3221.4 package.scala 96:25:@3222.4]
  wire  _T_158; // @[Controllers.scala 292:61:@3223.4]
  wire  _T_159; // @[Controllers.scala 292:24:@3224.4]
  SRFF active ( // @[Controllers.scala 261:22:@3121.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@3124.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_12 RetimeWrapper ( // @[package.scala 93:22:@3158.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_12 RetimeWrapper_1 ( // @[package.scala 93:22:@3180.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@3192.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@3200.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_16 RetimeWrapper_4 ( // @[package.scala 93:22:@3216.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@3129.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@3130.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@3131.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@3132.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@3149.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@3163.4 package.scala 96:25:@3164.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@3165.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@3168.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@3173.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@3174.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@3177.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@3185.4 package.scala 96:25:@3186.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@3187.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@3212.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@3221.4 package.scala 96:25:@3222.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@3223.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@3224.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@3191.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@3226.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@3176.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@3179.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@3171.4]
  assign active_clock = clock; // @[:@3122.4]
  assign active_reset = reset; // @[:@3123.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@3134.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@3138.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@3139.4]
  assign done_clock = clock; // @[:@3125.4]
  assign done_reset = reset; // @[:@3126.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@3154.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@3147.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@3148.4]
  assign RetimeWrapper_clock = clock; // @[:@3159.4]
  assign RetimeWrapper_reset = reset; // @[:@3160.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@3162.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@3161.4]
  assign RetimeWrapper_1_clock = clock; // @[:@3181.4]
  assign RetimeWrapper_1_reset = reset; // @[:@3182.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@3184.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@3183.4]
  assign RetimeWrapper_2_clock = clock; // @[:@3193.4]
  assign RetimeWrapper_2_reset = reset; // @[:@3194.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@3196.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@3195.4]
  assign RetimeWrapper_3_clock = clock; // @[:@3201.4]
  assign RetimeWrapper_3_reset = reset; // @[:@3202.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@3204.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@3203.4]
  assign RetimeWrapper_4_clock = clock; // @[:@3217.4]
  assign RetimeWrapper_4_reset = reset; // @[:@3218.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@3220.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@3219.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module SimBlackBoxesfix2fixBox( // @[:@3332.2]
  input  [31:0] io_a, // @[:@3335.4]
  output [31:0] io_b // @[:@3335.4]
);
  assign io_b = io_a; // @[SimBlackBoxes.scala 99:40:@3345.4]
endmodule
module _( // @[:@3347.2]
  input  [31:0] io_b, // @[:@3350.4]
  output [31:0] io_result // @[:@3350.4]
);
  wire [31:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@3355.4]
  wire [31:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@3355.4]
  SimBlackBoxesfix2fixBox SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@3355.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@3368.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@3363.4]
endmodule
module RetimeWrapper_21( // @[:@3452.2]
  input        clock, // @[:@3453.4]
  input        reset, // @[:@3454.4]
  input        io_flow, // @[:@3455.4]
  input  [7:0] io_in, // @[:@3455.4]
  output [7:0] io_out // @[:@3455.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@3457.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3470.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3469.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@3468.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3467.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3466.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3464.4]
endmodule
module Mem1D_4( // @[:@3472.2]
  input        clock, // @[:@3473.4]
  input        reset, // @[:@3474.4]
  input        io_r_ofs_0, // @[:@3475.4]
  input        io_r_backpressure, // @[:@3475.4]
  input        io_w_ofs_0, // @[:@3475.4]
  input  [7:0] io_w_data_0, // @[:@3475.4]
  input        io_w_en_0, // @[:@3475.4]
  output [7:0] io_output // @[:@3475.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3485.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3485.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3485.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@3485.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@3485.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@3494.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@3494.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@3494.4]
  wire [7:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@3494.4]
  wire [7:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@3494.4]
  reg [7:0] _T_127; // @[MemPrimitives.scala 560:26:@3479.4]
  reg [31:0] _RAND_0;
  wire  _T_130; // @[MemPrimitives.scala 561:61:@3481.4]
  wire  _T_131; // @[MemPrimitives.scala 561:44:@3482.4]
  wire [7:0] _T_132; // @[MemPrimitives.scala 561:19:@3483.4]
  wire  _T_135; // @[package.scala 96:25:@3490.4 package.scala 96:25:@3491.4]
  wire  _T_137; // @[Mux.scala 46:19:@3492.4]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@3485.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_1 ( // @[package.scala 93:22:@3494.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign _T_130 = io_w_ofs_0 == 1'h0; // @[MemPrimitives.scala 561:61:@3481.4]
  assign _T_131 = io_w_en_0 & _T_130; // @[MemPrimitives.scala 561:44:@3482.4]
  assign _T_132 = _T_131 ? io_w_data_0 : _T_127; // @[MemPrimitives.scala 561:19:@3483.4]
  assign _T_135 = RetimeWrapper_io_out; // @[package.scala 96:25:@3490.4 package.scala 96:25:@3491.4]
  assign _T_137 = 1'h0 == _T_135; // @[Mux.scala 46:19:@3492.4]
  assign io_output = RetimeWrapper_1_io_out; // @[MemPrimitives.scala 565:17:@3501.4]
  assign RetimeWrapper_clock = clock; // @[:@3486.4]
  assign RetimeWrapper_reset = reset; // @[:@3487.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@3489.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@3488.4]
  assign RetimeWrapper_1_clock = clock; // @[:@3495.4]
  assign RetimeWrapper_1_reset = reset; // @[:@3496.4]
  assign RetimeWrapper_1_io_flow = io_r_backpressure; // @[package.scala 95:18:@3498.4]
  assign RetimeWrapper_1_io_in = _T_137 ? _T_127 : 8'h0; // @[package.scala 94:16:@3497.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_127 = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_127 <= 8'h0;
    end else begin
      if (_T_131) begin
        _T_127 <= io_w_data_0;
      end
    end
  end
endmodule
module StickySelects( // @[:@4928.2]
  input   clock, // @[:@4929.4]
  input   reset, // @[:@4930.4]
  input   io_ins_0, // @[:@4931.4]
  input   io_ins_1, // @[:@4931.4]
  input   io_ins_2, // @[:@4931.4]
  input   io_ins_3, // @[:@4931.4]
  output  io_outs_0, // @[:@4931.4]
  output  io_outs_1, // @[:@4931.4]
  output  io_outs_2, // @[:@4931.4]
  output  io_outs_3 // @[:@4931.4]
);
  reg  _T_19; // @[StickySelects.scala 21:22:@4933.4]
  reg [31:0] _RAND_0;
  wire  _T_20; // @[StickySelects.scala 22:54:@4934.4]
  wire  _T_21; // @[StickySelects.scala 22:54:@4935.4]
  wire  _T_23; // @[StickySelects.scala 24:52:@4936.4]
  wire  _T_24; // @[StickySelects.scala 24:21:@4937.4]
  reg  _T_27; // @[StickySelects.scala 21:22:@4939.4]
  reg [31:0] _RAND_1;
  wire  _T_28; // @[StickySelects.scala 22:54:@4940.4]
  wire  _T_29; // @[StickySelects.scala 22:54:@4941.4]
  wire  _T_31; // @[StickySelects.scala 24:52:@4942.4]
  wire  _T_32; // @[StickySelects.scala 24:21:@4943.4]
  reg  _T_35; // @[StickySelects.scala 21:22:@4945.4]
  reg [31:0] _RAND_2;
  wire  _T_36; // @[StickySelects.scala 22:54:@4946.4]
  wire  _T_37; // @[StickySelects.scala 22:54:@4947.4]
  wire  _T_39; // @[StickySelects.scala 24:52:@4948.4]
  wire  _T_40; // @[StickySelects.scala 24:21:@4949.4]
  reg  _T_43; // @[StickySelects.scala 21:22:@4951.4]
  reg [31:0] _RAND_3;
  wire  _T_45; // @[StickySelects.scala 22:54:@4953.4]
  wire  _T_47; // @[StickySelects.scala 24:52:@4954.4]
  wire  _T_48; // @[StickySelects.scala 24:21:@4955.4]
  assign _T_20 = io_ins_1 | io_ins_2; // @[StickySelects.scala 22:54:@4934.4]
  assign _T_21 = _T_20 | io_ins_3; // @[StickySelects.scala 22:54:@4935.4]
  assign _T_23 = io_ins_0 | _T_19; // @[StickySelects.scala 24:52:@4936.4]
  assign _T_24 = _T_21 ? 1'h0 : _T_23; // @[StickySelects.scala 24:21:@4937.4]
  assign _T_28 = io_ins_0 | io_ins_2; // @[StickySelects.scala 22:54:@4940.4]
  assign _T_29 = _T_28 | io_ins_3; // @[StickySelects.scala 22:54:@4941.4]
  assign _T_31 = io_ins_1 | _T_27; // @[StickySelects.scala 24:52:@4942.4]
  assign _T_32 = _T_29 ? 1'h0 : _T_31; // @[StickySelects.scala 24:21:@4943.4]
  assign _T_36 = io_ins_0 | io_ins_1; // @[StickySelects.scala 22:54:@4946.4]
  assign _T_37 = _T_36 | io_ins_3; // @[StickySelects.scala 22:54:@4947.4]
  assign _T_39 = io_ins_2 | _T_35; // @[StickySelects.scala 24:52:@4948.4]
  assign _T_40 = _T_37 ? 1'h0 : _T_39; // @[StickySelects.scala 24:21:@4949.4]
  assign _T_45 = _T_36 | io_ins_2; // @[StickySelects.scala 22:54:@4953.4]
  assign _T_47 = io_ins_3 | _T_43; // @[StickySelects.scala 24:52:@4954.4]
  assign _T_48 = _T_45 ? 1'h0 : _T_47; // @[StickySelects.scala 24:21:@4955.4]
  assign io_outs_0 = _T_21 ? 1'h0 : _T_23; // @[StickySelects.scala 28:52:@4957.4]
  assign io_outs_1 = _T_29 ? 1'h0 : _T_31; // @[StickySelects.scala 28:52:@4958.4]
  assign io_outs_2 = _T_37 ? 1'h0 : _T_39; // @[StickySelects.scala 28:52:@4959.4]
  assign io_outs_3 = _T_45 ? 1'h0 : _T_47; // @[StickySelects.scala 28:52:@4960.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_27 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_35 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_43 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (_T_21) begin
        _T_19 <= 1'h0;
      end else begin
        _T_19 <= _T_23;
      end
    end
    if (reset) begin
      _T_27 <= 1'h0;
    end else begin
      if (_T_29) begin
        _T_27 <= 1'h0;
      end else begin
        _T_27 <= _T_31;
      end
    end
    if (reset) begin
      _T_35 <= 1'h0;
    end else begin
      if (_T_37) begin
        _T_35 <= 1'h0;
      end else begin
        _T_35 <= _T_39;
      end
    end
    if (reset) begin
      _T_43 <= 1'h0;
    end else begin
      if (_T_45) begin
        _T_43 <= 1'h0;
      end else begin
        _T_43 <= _T_47;
      end
    end
  end
endmodule
module StickySelects_2( // @[:@4996.2]
  input   clock, // @[:@4997.4]
  input   reset, // @[:@4998.4]
  input   io_ins_0, // @[:@4999.4]
  input   io_ins_1, // @[:@4999.4]
  input   io_ins_2, // @[:@4999.4]
  input   io_ins_3, // @[:@4999.4]
  input   io_ins_4, // @[:@4999.4]
  input   io_ins_5, // @[:@4999.4]
  input   io_ins_6, // @[:@4999.4]
  input   io_ins_7, // @[:@4999.4]
  output  io_outs_0, // @[:@4999.4]
  output  io_outs_1, // @[:@4999.4]
  output  io_outs_2, // @[:@4999.4]
  output  io_outs_3, // @[:@4999.4]
  output  io_outs_4, // @[:@4999.4]
  output  io_outs_5, // @[:@4999.4]
  output  io_outs_6, // @[:@4999.4]
  output  io_outs_7 // @[:@4999.4]
);
  reg  _T_19; // @[StickySelects.scala 21:22:@5001.4]
  reg [31:0] _RAND_0;
  wire  _T_20; // @[StickySelects.scala 22:54:@5002.4]
  wire  _T_21; // @[StickySelects.scala 22:54:@5003.4]
  wire  _T_22; // @[StickySelects.scala 22:54:@5004.4]
  wire  _T_23; // @[StickySelects.scala 22:54:@5005.4]
  wire  _T_24; // @[StickySelects.scala 22:54:@5006.4]
  wire  _T_25; // @[StickySelects.scala 22:54:@5007.4]
  wire  _T_27; // @[StickySelects.scala 24:52:@5008.4]
  wire  _T_28; // @[StickySelects.scala 24:21:@5009.4]
  reg  _T_31; // @[StickySelects.scala 21:22:@5011.4]
  reg [31:0] _RAND_1;
  wire  _T_32; // @[StickySelects.scala 22:54:@5012.4]
  wire  _T_33; // @[StickySelects.scala 22:54:@5013.4]
  wire  _T_34; // @[StickySelects.scala 22:54:@5014.4]
  wire  _T_35; // @[StickySelects.scala 22:54:@5015.4]
  wire  _T_36; // @[StickySelects.scala 22:54:@5016.4]
  wire  _T_37; // @[StickySelects.scala 22:54:@5017.4]
  wire  _T_39; // @[StickySelects.scala 24:52:@5018.4]
  wire  _T_40; // @[StickySelects.scala 24:21:@5019.4]
  reg  _T_43; // @[StickySelects.scala 21:22:@5021.4]
  reg [31:0] _RAND_2;
  wire  _T_44; // @[StickySelects.scala 22:54:@5022.4]
  wire  _T_45; // @[StickySelects.scala 22:54:@5023.4]
  wire  _T_46; // @[StickySelects.scala 22:54:@5024.4]
  wire  _T_47; // @[StickySelects.scala 22:54:@5025.4]
  wire  _T_48; // @[StickySelects.scala 22:54:@5026.4]
  wire  _T_49; // @[StickySelects.scala 22:54:@5027.4]
  wire  _T_51; // @[StickySelects.scala 24:52:@5028.4]
  wire  _T_52; // @[StickySelects.scala 24:21:@5029.4]
  reg  _T_55; // @[StickySelects.scala 21:22:@5031.4]
  reg [31:0] _RAND_3;
  wire  _T_57; // @[StickySelects.scala 22:54:@5033.4]
  wire  _T_58; // @[StickySelects.scala 22:54:@5034.4]
  wire  _T_59; // @[StickySelects.scala 22:54:@5035.4]
  wire  _T_60; // @[StickySelects.scala 22:54:@5036.4]
  wire  _T_61; // @[StickySelects.scala 22:54:@5037.4]
  wire  _T_63; // @[StickySelects.scala 24:52:@5038.4]
  wire  _T_64; // @[StickySelects.scala 24:21:@5039.4]
  reg  _T_67; // @[StickySelects.scala 21:22:@5041.4]
  reg [31:0] _RAND_4;
  wire  _T_70; // @[StickySelects.scala 22:54:@5044.4]
  wire  _T_71; // @[StickySelects.scala 22:54:@5045.4]
  wire  _T_72; // @[StickySelects.scala 22:54:@5046.4]
  wire  _T_73; // @[StickySelects.scala 22:54:@5047.4]
  wire  _T_75; // @[StickySelects.scala 24:52:@5048.4]
  wire  _T_76; // @[StickySelects.scala 24:21:@5049.4]
  reg  _T_79; // @[StickySelects.scala 21:22:@5051.4]
  reg [31:0] _RAND_5;
  wire  _T_83; // @[StickySelects.scala 22:54:@5055.4]
  wire  _T_84; // @[StickySelects.scala 22:54:@5056.4]
  wire  _T_85; // @[StickySelects.scala 22:54:@5057.4]
  wire  _T_87; // @[StickySelects.scala 24:52:@5058.4]
  wire  _T_88; // @[StickySelects.scala 24:21:@5059.4]
  reg  _T_91; // @[StickySelects.scala 21:22:@5061.4]
  reg [31:0] _RAND_6;
  wire  _T_96; // @[StickySelects.scala 22:54:@5066.4]
  wire  _T_97; // @[StickySelects.scala 22:54:@5067.4]
  wire  _T_99; // @[StickySelects.scala 24:52:@5068.4]
  wire  _T_100; // @[StickySelects.scala 24:21:@5069.4]
  reg  _T_103; // @[StickySelects.scala 21:22:@5071.4]
  reg [31:0] _RAND_7;
  wire  _T_109; // @[StickySelects.scala 22:54:@5077.4]
  wire  _T_111; // @[StickySelects.scala 24:52:@5078.4]
  wire  _T_112; // @[StickySelects.scala 24:21:@5079.4]
  assign _T_20 = io_ins_1 | io_ins_2; // @[StickySelects.scala 22:54:@5002.4]
  assign _T_21 = _T_20 | io_ins_3; // @[StickySelects.scala 22:54:@5003.4]
  assign _T_22 = _T_21 | io_ins_4; // @[StickySelects.scala 22:54:@5004.4]
  assign _T_23 = _T_22 | io_ins_5; // @[StickySelects.scala 22:54:@5005.4]
  assign _T_24 = _T_23 | io_ins_6; // @[StickySelects.scala 22:54:@5006.4]
  assign _T_25 = _T_24 | io_ins_7; // @[StickySelects.scala 22:54:@5007.4]
  assign _T_27 = io_ins_0 | _T_19; // @[StickySelects.scala 24:52:@5008.4]
  assign _T_28 = _T_25 ? 1'h0 : _T_27; // @[StickySelects.scala 24:21:@5009.4]
  assign _T_32 = io_ins_0 | io_ins_2; // @[StickySelects.scala 22:54:@5012.4]
  assign _T_33 = _T_32 | io_ins_3; // @[StickySelects.scala 22:54:@5013.4]
  assign _T_34 = _T_33 | io_ins_4; // @[StickySelects.scala 22:54:@5014.4]
  assign _T_35 = _T_34 | io_ins_5; // @[StickySelects.scala 22:54:@5015.4]
  assign _T_36 = _T_35 | io_ins_6; // @[StickySelects.scala 22:54:@5016.4]
  assign _T_37 = _T_36 | io_ins_7; // @[StickySelects.scala 22:54:@5017.4]
  assign _T_39 = io_ins_1 | _T_31; // @[StickySelects.scala 24:52:@5018.4]
  assign _T_40 = _T_37 ? 1'h0 : _T_39; // @[StickySelects.scala 24:21:@5019.4]
  assign _T_44 = io_ins_0 | io_ins_1; // @[StickySelects.scala 22:54:@5022.4]
  assign _T_45 = _T_44 | io_ins_3; // @[StickySelects.scala 22:54:@5023.4]
  assign _T_46 = _T_45 | io_ins_4; // @[StickySelects.scala 22:54:@5024.4]
  assign _T_47 = _T_46 | io_ins_5; // @[StickySelects.scala 22:54:@5025.4]
  assign _T_48 = _T_47 | io_ins_6; // @[StickySelects.scala 22:54:@5026.4]
  assign _T_49 = _T_48 | io_ins_7; // @[StickySelects.scala 22:54:@5027.4]
  assign _T_51 = io_ins_2 | _T_43; // @[StickySelects.scala 24:52:@5028.4]
  assign _T_52 = _T_49 ? 1'h0 : _T_51; // @[StickySelects.scala 24:21:@5029.4]
  assign _T_57 = _T_44 | io_ins_2; // @[StickySelects.scala 22:54:@5033.4]
  assign _T_58 = _T_57 | io_ins_4; // @[StickySelects.scala 22:54:@5034.4]
  assign _T_59 = _T_58 | io_ins_5; // @[StickySelects.scala 22:54:@5035.4]
  assign _T_60 = _T_59 | io_ins_6; // @[StickySelects.scala 22:54:@5036.4]
  assign _T_61 = _T_60 | io_ins_7; // @[StickySelects.scala 22:54:@5037.4]
  assign _T_63 = io_ins_3 | _T_55; // @[StickySelects.scala 24:52:@5038.4]
  assign _T_64 = _T_61 ? 1'h0 : _T_63; // @[StickySelects.scala 24:21:@5039.4]
  assign _T_70 = _T_57 | io_ins_3; // @[StickySelects.scala 22:54:@5044.4]
  assign _T_71 = _T_70 | io_ins_5; // @[StickySelects.scala 22:54:@5045.4]
  assign _T_72 = _T_71 | io_ins_6; // @[StickySelects.scala 22:54:@5046.4]
  assign _T_73 = _T_72 | io_ins_7; // @[StickySelects.scala 22:54:@5047.4]
  assign _T_75 = io_ins_4 | _T_67; // @[StickySelects.scala 24:52:@5048.4]
  assign _T_76 = _T_73 ? 1'h0 : _T_75; // @[StickySelects.scala 24:21:@5049.4]
  assign _T_83 = _T_70 | io_ins_4; // @[StickySelects.scala 22:54:@5055.4]
  assign _T_84 = _T_83 | io_ins_6; // @[StickySelects.scala 22:54:@5056.4]
  assign _T_85 = _T_84 | io_ins_7; // @[StickySelects.scala 22:54:@5057.4]
  assign _T_87 = io_ins_5 | _T_79; // @[StickySelects.scala 24:52:@5058.4]
  assign _T_88 = _T_85 ? 1'h0 : _T_87; // @[StickySelects.scala 24:21:@5059.4]
  assign _T_96 = _T_83 | io_ins_5; // @[StickySelects.scala 22:54:@5066.4]
  assign _T_97 = _T_96 | io_ins_7; // @[StickySelects.scala 22:54:@5067.4]
  assign _T_99 = io_ins_6 | _T_91; // @[StickySelects.scala 24:52:@5068.4]
  assign _T_100 = _T_97 ? 1'h0 : _T_99; // @[StickySelects.scala 24:21:@5069.4]
  assign _T_109 = _T_96 | io_ins_6; // @[StickySelects.scala 22:54:@5077.4]
  assign _T_111 = io_ins_7 | _T_103; // @[StickySelects.scala 24:52:@5078.4]
  assign _T_112 = _T_109 ? 1'h0 : _T_111; // @[StickySelects.scala 24:21:@5079.4]
  assign io_outs_0 = _T_25 ? 1'h0 : _T_27; // @[StickySelects.scala 28:52:@5081.4]
  assign io_outs_1 = _T_37 ? 1'h0 : _T_39; // @[StickySelects.scala 28:52:@5082.4]
  assign io_outs_2 = _T_49 ? 1'h0 : _T_51; // @[StickySelects.scala 28:52:@5083.4]
  assign io_outs_3 = _T_61 ? 1'h0 : _T_63; // @[StickySelects.scala 28:52:@5084.4]
  assign io_outs_4 = _T_73 ? 1'h0 : _T_75; // @[StickySelects.scala 28:52:@5085.4]
  assign io_outs_5 = _T_85 ? 1'h0 : _T_87; // @[StickySelects.scala 28:52:@5086.4]
  assign io_outs_6 = _T_97 ? 1'h0 : _T_99; // @[StickySelects.scala 28:52:@5087.4]
  assign io_outs_7 = _T_109 ? 1'h0 : _T_111; // @[StickySelects.scala 28:52:@5088.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_31 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_43 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_55 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_67 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_79 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_91 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_103 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (_T_25) begin
        _T_19 <= 1'h0;
      end else begin
        _T_19 <= _T_27;
      end
    end
    if (reset) begin
      _T_31 <= 1'h0;
    end else begin
      if (_T_37) begin
        _T_31 <= 1'h0;
      end else begin
        _T_31 <= _T_39;
      end
    end
    if (reset) begin
      _T_43 <= 1'h0;
    end else begin
      if (_T_49) begin
        _T_43 <= 1'h0;
      end else begin
        _T_43 <= _T_51;
      end
    end
    if (reset) begin
      _T_55 <= 1'h0;
    end else begin
      if (_T_61) begin
        _T_55 <= 1'h0;
      end else begin
        _T_55 <= _T_63;
      end
    end
    if (reset) begin
      _T_67 <= 1'h0;
    end else begin
      if (_T_73) begin
        _T_67 <= 1'h0;
      end else begin
        _T_67 <= _T_75;
      end
    end
    if (reset) begin
      _T_79 <= 1'h0;
    end else begin
      if (_T_85) begin
        _T_79 <= 1'h0;
      end else begin
        _T_79 <= _T_87;
      end
    end
    if (reset) begin
      _T_91 <= 1'h0;
    end else begin
      if (_T_97) begin
        _T_91 <= 1'h0;
      end else begin
        _T_91 <= _T_99;
      end
    end
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      if (_T_109) begin
        _T_103 <= 1'h0;
      end else begin
        _T_103 <= _T_111;
      end
    end
  end
endmodule
module RetimeWrapper_52( // @[:@5964.2]
  input   clock, // @[:@5965.4]
  input   reset, // @[:@5966.4]
  input   io_flow, // @[:@5967.4]
  input   io_in, // @[:@5967.4]
  output  io_out // @[:@5967.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@5969.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@5969.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@5969.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@5969.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@5969.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@5969.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@5969.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@5982.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@5981.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@5980.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@5979.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@5978.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@5976.4]
endmodule
module x439_lb_0( // @[:@9024.2]
  input        clock, // @[:@9025.4]
  input        reset, // @[:@9026.4]
  input  [2:0] io_rPort_23_banks_0, // @[:@9027.4]
  input        io_rPort_23_ofs_0, // @[:@9027.4]
  input        io_rPort_23_en_0, // @[:@9027.4]
  input        io_rPort_23_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_23_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_22_banks_0, // @[:@9027.4]
  input        io_rPort_22_ofs_0, // @[:@9027.4]
  input        io_rPort_22_en_0, // @[:@9027.4]
  input        io_rPort_22_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_22_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_21_banks_0, // @[:@9027.4]
  input        io_rPort_21_ofs_0, // @[:@9027.4]
  input        io_rPort_21_en_0, // @[:@9027.4]
  input        io_rPort_21_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_21_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_20_banks_0, // @[:@9027.4]
  input        io_rPort_20_ofs_0, // @[:@9027.4]
  input        io_rPort_20_en_0, // @[:@9027.4]
  input        io_rPort_20_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_20_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_19_banks_0, // @[:@9027.4]
  input        io_rPort_19_ofs_0, // @[:@9027.4]
  input        io_rPort_19_en_0, // @[:@9027.4]
  input        io_rPort_19_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_19_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_18_banks_0, // @[:@9027.4]
  input        io_rPort_18_ofs_0, // @[:@9027.4]
  input        io_rPort_18_en_0, // @[:@9027.4]
  input        io_rPort_18_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_18_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_17_banks_0, // @[:@9027.4]
  input        io_rPort_17_ofs_0, // @[:@9027.4]
  input        io_rPort_17_en_0, // @[:@9027.4]
  input        io_rPort_17_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_17_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_16_banks_0, // @[:@9027.4]
  input        io_rPort_16_ofs_0, // @[:@9027.4]
  input        io_rPort_16_en_0, // @[:@9027.4]
  input        io_rPort_16_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_16_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_15_banks_0, // @[:@9027.4]
  input        io_rPort_15_ofs_0, // @[:@9027.4]
  input        io_rPort_15_en_0, // @[:@9027.4]
  input        io_rPort_15_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_15_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_14_banks_0, // @[:@9027.4]
  input        io_rPort_14_ofs_0, // @[:@9027.4]
  input        io_rPort_14_en_0, // @[:@9027.4]
  input        io_rPort_14_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_14_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_13_banks_0, // @[:@9027.4]
  input        io_rPort_13_ofs_0, // @[:@9027.4]
  input        io_rPort_13_en_0, // @[:@9027.4]
  input        io_rPort_13_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_13_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_12_banks_0, // @[:@9027.4]
  input        io_rPort_12_ofs_0, // @[:@9027.4]
  input        io_rPort_12_en_0, // @[:@9027.4]
  input        io_rPort_12_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_12_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_11_banks_0, // @[:@9027.4]
  input        io_rPort_11_ofs_0, // @[:@9027.4]
  input        io_rPort_11_en_0, // @[:@9027.4]
  input        io_rPort_11_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_11_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_10_banks_0, // @[:@9027.4]
  input        io_rPort_10_ofs_0, // @[:@9027.4]
  input        io_rPort_10_en_0, // @[:@9027.4]
  input        io_rPort_10_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_10_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_9_banks_0, // @[:@9027.4]
  input        io_rPort_9_ofs_0, // @[:@9027.4]
  input        io_rPort_9_en_0, // @[:@9027.4]
  input        io_rPort_9_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_9_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_8_banks_0, // @[:@9027.4]
  input        io_rPort_8_ofs_0, // @[:@9027.4]
  input        io_rPort_8_en_0, // @[:@9027.4]
  input        io_rPort_8_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_8_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_7_banks_0, // @[:@9027.4]
  input        io_rPort_7_ofs_0, // @[:@9027.4]
  input        io_rPort_7_en_0, // @[:@9027.4]
  input        io_rPort_7_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_7_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_6_banks_0, // @[:@9027.4]
  input        io_rPort_6_ofs_0, // @[:@9027.4]
  input        io_rPort_6_en_0, // @[:@9027.4]
  input        io_rPort_6_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_6_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_5_banks_0, // @[:@9027.4]
  input        io_rPort_5_ofs_0, // @[:@9027.4]
  input        io_rPort_5_en_0, // @[:@9027.4]
  input        io_rPort_5_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_5_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_4_banks_0, // @[:@9027.4]
  input        io_rPort_4_ofs_0, // @[:@9027.4]
  input        io_rPort_4_en_0, // @[:@9027.4]
  input        io_rPort_4_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_4_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_3_banks_0, // @[:@9027.4]
  input        io_rPort_3_ofs_0, // @[:@9027.4]
  input        io_rPort_3_en_0, // @[:@9027.4]
  input        io_rPort_3_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_3_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_2_banks_0, // @[:@9027.4]
  input        io_rPort_2_ofs_0, // @[:@9027.4]
  input        io_rPort_2_en_0, // @[:@9027.4]
  input        io_rPort_2_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_2_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_1_banks_0, // @[:@9027.4]
  input        io_rPort_1_ofs_0, // @[:@9027.4]
  input        io_rPort_1_en_0, // @[:@9027.4]
  input        io_rPort_1_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_1_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_0_banks_0, // @[:@9027.4]
  input        io_rPort_0_ofs_0, // @[:@9027.4]
  input        io_rPort_0_en_0, // @[:@9027.4]
  input        io_rPort_0_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_0_output_0, // @[:@9027.4]
  input  [2:0] io_wPort_7_banks_0, // @[:@9027.4]
  input        io_wPort_7_ofs_0, // @[:@9027.4]
  input  [7:0] io_wPort_7_data_0, // @[:@9027.4]
  input        io_wPort_7_en_0, // @[:@9027.4]
  input  [2:0] io_wPort_6_banks_0, // @[:@9027.4]
  input        io_wPort_6_ofs_0, // @[:@9027.4]
  input  [7:0] io_wPort_6_data_0, // @[:@9027.4]
  input        io_wPort_6_en_0, // @[:@9027.4]
  input  [2:0] io_wPort_5_banks_0, // @[:@9027.4]
  input        io_wPort_5_ofs_0, // @[:@9027.4]
  input  [7:0] io_wPort_5_data_0, // @[:@9027.4]
  input        io_wPort_5_en_0, // @[:@9027.4]
  input  [2:0] io_wPort_4_banks_0, // @[:@9027.4]
  input        io_wPort_4_ofs_0, // @[:@9027.4]
  input  [7:0] io_wPort_4_data_0, // @[:@9027.4]
  input        io_wPort_4_en_0, // @[:@9027.4]
  input  [2:0] io_wPort_3_banks_0, // @[:@9027.4]
  input        io_wPort_3_ofs_0, // @[:@9027.4]
  input  [7:0] io_wPort_3_data_0, // @[:@9027.4]
  input        io_wPort_3_en_0, // @[:@9027.4]
  input  [2:0] io_wPort_2_banks_0, // @[:@9027.4]
  input        io_wPort_2_ofs_0, // @[:@9027.4]
  input  [7:0] io_wPort_2_data_0, // @[:@9027.4]
  input        io_wPort_2_en_0, // @[:@9027.4]
  input  [2:0] io_wPort_1_banks_0, // @[:@9027.4]
  input        io_wPort_1_ofs_0, // @[:@9027.4]
  input  [7:0] io_wPort_1_data_0, // @[:@9027.4]
  input        io_wPort_1_en_0, // @[:@9027.4]
  input  [2:0] io_wPort_0_banks_0, // @[:@9027.4]
  input        io_wPort_0_ofs_0, // @[:@9027.4]
  input  [7:0] io_wPort_0_data_0, // @[:@9027.4]
  input        io_wPort_0_en_0 // @[:@9027.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@9238.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@9238.4]
  wire  Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9238.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9238.4]
  wire  Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9238.4]
  wire [7:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@9238.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@9238.4]
  wire [7:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@9238.4]
  wire  Mem1D_1_clock; // @[MemPrimitives.scala 64:21:@9254.4]
  wire  Mem1D_1_reset; // @[MemPrimitives.scala 64:21:@9254.4]
  wire  Mem1D_1_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9254.4]
  wire  Mem1D_1_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9254.4]
  wire  Mem1D_1_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9254.4]
  wire [7:0] Mem1D_1_io_w_data_0; // @[MemPrimitives.scala 64:21:@9254.4]
  wire  Mem1D_1_io_w_en_0; // @[MemPrimitives.scala 64:21:@9254.4]
  wire [7:0] Mem1D_1_io_output; // @[MemPrimitives.scala 64:21:@9254.4]
  wire  Mem1D_2_clock; // @[MemPrimitives.scala 64:21:@9270.4]
  wire  Mem1D_2_reset; // @[MemPrimitives.scala 64:21:@9270.4]
  wire  Mem1D_2_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9270.4]
  wire  Mem1D_2_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9270.4]
  wire  Mem1D_2_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9270.4]
  wire [7:0] Mem1D_2_io_w_data_0; // @[MemPrimitives.scala 64:21:@9270.4]
  wire  Mem1D_2_io_w_en_0; // @[MemPrimitives.scala 64:21:@9270.4]
  wire [7:0] Mem1D_2_io_output; // @[MemPrimitives.scala 64:21:@9270.4]
  wire  Mem1D_3_clock; // @[MemPrimitives.scala 64:21:@9286.4]
  wire  Mem1D_3_reset; // @[MemPrimitives.scala 64:21:@9286.4]
  wire  Mem1D_3_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9286.4]
  wire  Mem1D_3_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9286.4]
  wire  Mem1D_3_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9286.4]
  wire [7:0] Mem1D_3_io_w_data_0; // @[MemPrimitives.scala 64:21:@9286.4]
  wire  Mem1D_3_io_w_en_0; // @[MemPrimitives.scala 64:21:@9286.4]
  wire [7:0] Mem1D_3_io_output; // @[MemPrimitives.scala 64:21:@9286.4]
  wire  Mem1D_4_clock; // @[MemPrimitives.scala 64:21:@9302.4]
  wire  Mem1D_4_reset; // @[MemPrimitives.scala 64:21:@9302.4]
  wire  Mem1D_4_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9302.4]
  wire  Mem1D_4_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9302.4]
  wire  Mem1D_4_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9302.4]
  wire [7:0] Mem1D_4_io_w_data_0; // @[MemPrimitives.scala 64:21:@9302.4]
  wire  Mem1D_4_io_w_en_0; // @[MemPrimitives.scala 64:21:@9302.4]
  wire [7:0] Mem1D_4_io_output; // @[MemPrimitives.scala 64:21:@9302.4]
  wire  Mem1D_5_clock; // @[MemPrimitives.scala 64:21:@9318.4]
  wire  Mem1D_5_reset; // @[MemPrimitives.scala 64:21:@9318.4]
  wire  Mem1D_5_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9318.4]
  wire  Mem1D_5_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9318.4]
  wire  Mem1D_5_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9318.4]
  wire [7:0] Mem1D_5_io_w_data_0; // @[MemPrimitives.scala 64:21:@9318.4]
  wire  Mem1D_5_io_w_en_0; // @[MemPrimitives.scala 64:21:@9318.4]
  wire [7:0] Mem1D_5_io_output; // @[MemPrimitives.scala 64:21:@9318.4]
  wire  Mem1D_6_clock; // @[MemPrimitives.scala 64:21:@9334.4]
  wire  Mem1D_6_reset; // @[MemPrimitives.scala 64:21:@9334.4]
  wire  Mem1D_6_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9334.4]
  wire  Mem1D_6_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9334.4]
  wire  Mem1D_6_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9334.4]
  wire [7:0] Mem1D_6_io_w_data_0; // @[MemPrimitives.scala 64:21:@9334.4]
  wire  Mem1D_6_io_w_en_0; // @[MemPrimitives.scala 64:21:@9334.4]
  wire [7:0] Mem1D_6_io_output; // @[MemPrimitives.scala 64:21:@9334.4]
  wire  Mem1D_7_clock; // @[MemPrimitives.scala 64:21:@9350.4]
  wire  Mem1D_7_reset; // @[MemPrimitives.scala 64:21:@9350.4]
  wire  Mem1D_7_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9350.4]
  wire  Mem1D_7_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9350.4]
  wire  Mem1D_7_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9350.4]
  wire [7:0] Mem1D_7_io_w_data_0; // @[MemPrimitives.scala 64:21:@9350.4]
  wire  Mem1D_7_io_w_en_0; // @[MemPrimitives.scala 64:21:@9350.4]
  wire [7:0] Mem1D_7_io_output; // @[MemPrimitives.scala 64:21:@9350.4]
  wire  Mem1D_8_clock; // @[MemPrimitives.scala 64:21:@9366.4]
  wire  Mem1D_8_reset; // @[MemPrimitives.scala 64:21:@9366.4]
  wire  Mem1D_8_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9366.4]
  wire  Mem1D_8_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9366.4]
  wire  Mem1D_8_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9366.4]
  wire [7:0] Mem1D_8_io_w_data_0; // @[MemPrimitives.scala 64:21:@9366.4]
  wire  Mem1D_8_io_w_en_0; // @[MemPrimitives.scala 64:21:@9366.4]
  wire [7:0] Mem1D_8_io_output; // @[MemPrimitives.scala 64:21:@9366.4]
  wire  Mem1D_9_clock; // @[MemPrimitives.scala 64:21:@9382.4]
  wire  Mem1D_9_reset; // @[MemPrimitives.scala 64:21:@9382.4]
  wire  Mem1D_9_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9382.4]
  wire  Mem1D_9_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9382.4]
  wire  Mem1D_9_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9382.4]
  wire [7:0] Mem1D_9_io_w_data_0; // @[MemPrimitives.scala 64:21:@9382.4]
  wire  Mem1D_9_io_w_en_0; // @[MemPrimitives.scala 64:21:@9382.4]
  wire [7:0] Mem1D_9_io_output; // @[MemPrimitives.scala 64:21:@9382.4]
  wire  Mem1D_10_clock; // @[MemPrimitives.scala 64:21:@9398.4]
  wire  Mem1D_10_reset; // @[MemPrimitives.scala 64:21:@9398.4]
  wire  Mem1D_10_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9398.4]
  wire  Mem1D_10_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9398.4]
  wire  Mem1D_10_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9398.4]
  wire [7:0] Mem1D_10_io_w_data_0; // @[MemPrimitives.scala 64:21:@9398.4]
  wire  Mem1D_10_io_w_en_0; // @[MemPrimitives.scala 64:21:@9398.4]
  wire [7:0] Mem1D_10_io_output; // @[MemPrimitives.scala 64:21:@9398.4]
  wire  Mem1D_11_clock; // @[MemPrimitives.scala 64:21:@9414.4]
  wire  Mem1D_11_reset; // @[MemPrimitives.scala 64:21:@9414.4]
  wire  Mem1D_11_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9414.4]
  wire  Mem1D_11_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9414.4]
  wire  Mem1D_11_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9414.4]
  wire [7:0] Mem1D_11_io_w_data_0; // @[MemPrimitives.scala 64:21:@9414.4]
  wire  Mem1D_11_io_w_en_0; // @[MemPrimitives.scala 64:21:@9414.4]
  wire [7:0] Mem1D_11_io_output; // @[MemPrimitives.scala 64:21:@9414.4]
  wire  Mem1D_12_clock; // @[MemPrimitives.scala 64:21:@9430.4]
  wire  Mem1D_12_reset; // @[MemPrimitives.scala 64:21:@9430.4]
  wire  Mem1D_12_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9430.4]
  wire  Mem1D_12_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9430.4]
  wire  Mem1D_12_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9430.4]
  wire [7:0] Mem1D_12_io_w_data_0; // @[MemPrimitives.scala 64:21:@9430.4]
  wire  Mem1D_12_io_w_en_0; // @[MemPrimitives.scala 64:21:@9430.4]
  wire [7:0] Mem1D_12_io_output; // @[MemPrimitives.scala 64:21:@9430.4]
  wire  Mem1D_13_clock; // @[MemPrimitives.scala 64:21:@9446.4]
  wire  Mem1D_13_reset; // @[MemPrimitives.scala 64:21:@9446.4]
  wire  Mem1D_13_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9446.4]
  wire  Mem1D_13_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9446.4]
  wire  Mem1D_13_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9446.4]
  wire [7:0] Mem1D_13_io_w_data_0; // @[MemPrimitives.scala 64:21:@9446.4]
  wire  Mem1D_13_io_w_en_0; // @[MemPrimitives.scala 64:21:@9446.4]
  wire [7:0] Mem1D_13_io_output; // @[MemPrimitives.scala 64:21:@9446.4]
  wire  Mem1D_14_clock; // @[MemPrimitives.scala 64:21:@9462.4]
  wire  Mem1D_14_reset; // @[MemPrimitives.scala 64:21:@9462.4]
  wire  Mem1D_14_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9462.4]
  wire  Mem1D_14_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9462.4]
  wire  Mem1D_14_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9462.4]
  wire [7:0] Mem1D_14_io_w_data_0; // @[MemPrimitives.scala 64:21:@9462.4]
  wire  Mem1D_14_io_w_en_0; // @[MemPrimitives.scala 64:21:@9462.4]
  wire [7:0] Mem1D_14_io_output; // @[MemPrimitives.scala 64:21:@9462.4]
  wire  Mem1D_15_clock; // @[MemPrimitives.scala 64:21:@9478.4]
  wire  Mem1D_15_reset; // @[MemPrimitives.scala 64:21:@9478.4]
  wire  Mem1D_15_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9478.4]
  wire  Mem1D_15_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9478.4]
  wire  Mem1D_15_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9478.4]
  wire [7:0] Mem1D_15_io_w_data_0; // @[MemPrimitives.scala 64:21:@9478.4]
  wire  Mem1D_15_io_w_en_0; // @[MemPrimitives.scala 64:21:@9478.4]
  wire [7:0] Mem1D_15_io_output; // @[MemPrimitives.scala 64:21:@9478.4]
  wire  StickySelects_clock; // @[MemPrimitives.scala 121:29:@9778.4]
  wire  StickySelects_reset; // @[MemPrimitives.scala 121:29:@9778.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 121:29:@9778.4]
  wire  StickySelects_io_ins_1; // @[MemPrimitives.scala 121:29:@9778.4]
  wire  StickySelects_io_ins_2; // @[MemPrimitives.scala 121:29:@9778.4]
  wire  StickySelects_io_ins_3; // @[MemPrimitives.scala 121:29:@9778.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 121:29:@9778.4]
  wire  StickySelects_io_outs_1; // @[MemPrimitives.scala 121:29:@9778.4]
  wire  StickySelects_io_outs_2; // @[MemPrimitives.scala 121:29:@9778.4]
  wire  StickySelects_io_outs_3; // @[MemPrimitives.scala 121:29:@9778.4]
  wire  StickySelects_1_clock; // @[MemPrimitives.scala 121:29:@9818.4]
  wire  StickySelects_1_reset; // @[MemPrimitives.scala 121:29:@9818.4]
  wire  StickySelects_1_io_ins_0; // @[MemPrimitives.scala 121:29:@9818.4]
  wire  StickySelects_1_io_ins_1; // @[MemPrimitives.scala 121:29:@9818.4]
  wire  StickySelects_1_io_ins_2; // @[MemPrimitives.scala 121:29:@9818.4]
  wire  StickySelects_1_io_ins_3; // @[MemPrimitives.scala 121:29:@9818.4]
  wire  StickySelects_1_io_outs_0; // @[MemPrimitives.scala 121:29:@9818.4]
  wire  StickySelects_1_io_outs_1; // @[MemPrimitives.scala 121:29:@9818.4]
  wire  StickySelects_1_io_outs_2; // @[MemPrimitives.scala 121:29:@9818.4]
  wire  StickySelects_1_io_outs_3; // @[MemPrimitives.scala 121:29:@9818.4]
  wire  StickySelects_2_clock; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_reset; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_ins_0; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_ins_1; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_ins_2; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_ins_3; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_ins_4; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_ins_5; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_ins_6; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_ins_7; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_outs_0; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_outs_1; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_outs_2; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_outs_3; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_outs_4; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_outs_5; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_outs_6; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_outs_7; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_3_clock; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_reset; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_ins_0; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_ins_1; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_ins_2; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_ins_3; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_ins_4; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_ins_5; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_ins_6; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_ins_7; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_outs_0; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_outs_1; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_outs_2; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_outs_3; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_outs_4; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_outs_5; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_outs_6; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_outs_7; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_4_clock; // @[MemPrimitives.scala 121:29:@10002.4]
  wire  StickySelects_4_reset; // @[MemPrimitives.scala 121:29:@10002.4]
  wire  StickySelects_4_io_ins_0; // @[MemPrimitives.scala 121:29:@10002.4]
  wire  StickySelects_4_io_ins_1; // @[MemPrimitives.scala 121:29:@10002.4]
  wire  StickySelects_4_io_ins_2; // @[MemPrimitives.scala 121:29:@10002.4]
  wire  StickySelects_4_io_ins_3; // @[MemPrimitives.scala 121:29:@10002.4]
  wire  StickySelects_4_io_outs_0; // @[MemPrimitives.scala 121:29:@10002.4]
  wire  StickySelects_4_io_outs_1; // @[MemPrimitives.scala 121:29:@10002.4]
  wire  StickySelects_4_io_outs_2; // @[MemPrimitives.scala 121:29:@10002.4]
  wire  StickySelects_4_io_outs_3; // @[MemPrimitives.scala 121:29:@10002.4]
  wire  StickySelects_5_clock; // @[MemPrimitives.scala 121:29:@10042.4]
  wire  StickySelects_5_reset; // @[MemPrimitives.scala 121:29:@10042.4]
  wire  StickySelects_5_io_ins_0; // @[MemPrimitives.scala 121:29:@10042.4]
  wire  StickySelects_5_io_ins_1; // @[MemPrimitives.scala 121:29:@10042.4]
  wire  StickySelects_5_io_ins_2; // @[MemPrimitives.scala 121:29:@10042.4]
  wire  StickySelects_5_io_ins_3; // @[MemPrimitives.scala 121:29:@10042.4]
  wire  StickySelects_5_io_outs_0; // @[MemPrimitives.scala 121:29:@10042.4]
  wire  StickySelects_5_io_outs_1; // @[MemPrimitives.scala 121:29:@10042.4]
  wire  StickySelects_5_io_outs_2; // @[MemPrimitives.scala 121:29:@10042.4]
  wire  StickySelects_5_io_outs_3; // @[MemPrimitives.scala 121:29:@10042.4]
  wire  StickySelects_6_clock; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_reset; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_ins_0; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_ins_1; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_ins_2; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_ins_3; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_ins_4; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_ins_5; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_ins_6; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_ins_7; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_outs_0; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_outs_1; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_outs_2; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_outs_3; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_outs_4; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_outs_5; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_outs_6; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_outs_7; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_7_clock; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_reset; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_ins_0; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_ins_1; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_ins_2; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_ins_3; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_ins_4; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_ins_5; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_ins_6; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_ins_7; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_outs_0; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_outs_1; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_outs_2; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_outs_3; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_outs_4; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_outs_5; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_outs_6; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_outs_7; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_8_clock; // @[MemPrimitives.scala 121:29:@10226.4]
  wire  StickySelects_8_reset; // @[MemPrimitives.scala 121:29:@10226.4]
  wire  StickySelects_8_io_ins_0; // @[MemPrimitives.scala 121:29:@10226.4]
  wire  StickySelects_8_io_ins_1; // @[MemPrimitives.scala 121:29:@10226.4]
  wire  StickySelects_8_io_ins_2; // @[MemPrimitives.scala 121:29:@10226.4]
  wire  StickySelects_8_io_ins_3; // @[MemPrimitives.scala 121:29:@10226.4]
  wire  StickySelects_8_io_outs_0; // @[MemPrimitives.scala 121:29:@10226.4]
  wire  StickySelects_8_io_outs_1; // @[MemPrimitives.scala 121:29:@10226.4]
  wire  StickySelects_8_io_outs_2; // @[MemPrimitives.scala 121:29:@10226.4]
  wire  StickySelects_8_io_outs_3; // @[MemPrimitives.scala 121:29:@10226.4]
  wire  StickySelects_9_clock; // @[MemPrimitives.scala 121:29:@10266.4]
  wire  StickySelects_9_reset; // @[MemPrimitives.scala 121:29:@10266.4]
  wire  StickySelects_9_io_ins_0; // @[MemPrimitives.scala 121:29:@10266.4]
  wire  StickySelects_9_io_ins_1; // @[MemPrimitives.scala 121:29:@10266.4]
  wire  StickySelects_9_io_ins_2; // @[MemPrimitives.scala 121:29:@10266.4]
  wire  StickySelects_9_io_ins_3; // @[MemPrimitives.scala 121:29:@10266.4]
  wire  StickySelects_9_io_outs_0; // @[MemPrimitives.scala 121:29:@10266.4]
  wire  StickySelects_9_io_outs_1; // @[MemPrimitives.scala 121:29:@10266.4]
  wire  StickySelects_9_io_outs_2; // @[MemPrimitives.scala 121:29:@10266.4]
  wire  StickySelects_9_io_outs_3; // @[MemPrimitives.scala 121:29:@10266.4]
  wire  StickySelects_10_clock; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_reset; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_ins_0; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_ins_1; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_ins_2; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_ins_3; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_ins_4; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_ins_5; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_ins_6; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_ins_7; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_outs_0; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_outs_1; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_outs_2; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_outs_3; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_outs_4; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_outs_5; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_outs_6; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_outs_7; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_11_clock; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_reset; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_ins_0; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_ins_1; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_ins_2; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_ins_3; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_ins_4; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_ins_5; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_ins_6; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_ins_7; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_outs_0; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_outs_1; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_outs_2; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_outs_3; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_outs_4; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_outs_5; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_outs_6; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_outs_7; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_12_clock; // @[MemPrimitives.scala 121:29:@10450.4]
  wire  StickySelects_12_reset; // @[MemPrimitives.scala 121:29:@10450.4]
  wire  StickySelects_12_io_ins_0; // @[MemPrimitives.scala 121:29:@10450.4]
  wire  StickySelects_12_io_ins_1; // @[MemPrimitives.scala 121:29:@10450.4]
  wire  StickySelects_12_io_ins_2; // @[MemPrimitives.scala 121:29:@10450.4]
  wire  StickySelects_12_io_ins_3; // @[MemPrimitives.scala 121:29:@10450.4]
  wire  StickySelects_12_io_outs_0; // @[MemPrimitives.scala 121:29:@10450.4]
  wire  StickySelects_12_io_outs_1; // @[MemPrimitives.scala 121:29:@10450.4]
  wire  StickySelects_12_io_outs_2; // @[MemPrimitives.scala 121:29:@10450.4]
  wire  StickySelects_12_io_outs_3; // @[MemPrimitives.scala 121:29:@10450.4]
  wire  StickySelects_13_clock; // @[MemPrimitives.scala 121:29:@10490.4]
  wire  StickySelects_13_reset; // @[MemPrimitives.scala 121:29:@10490.4]
  wire  StickySelects_13_io_ins_0; // @[MemPrimitives.scala 121:29:@10490.4]
  wire  StickySelects_13_io_ins_1; // @[MemPrimitives.scala 121:29:@10490.4]
  wire  StickySelects_13_io_ins_2; // @[MemPrimitives.scala 121:29:@10490.4]
  wire  StickySelects_13_io_ins_3; // @[MemPrimitives.scala 121:29:@10490.4]
  wire  StickySelects_13_io_outs_0; // @[MemPrimitives.scala 121:29:@10490.4]
  wire  StickySelects_13_io_outs_1; // @[MemPrimitives.scala 121:29:@10490.4]
  wire  StickySelects_13_io_outs_2; // @[MemPrimitives.scala 121:29:@10490.4]
  wire  StickySelects_13_io_outs_3; // @[MemPrimitives.scala 121:29:@10490.4]
  wire  StickySelects_14_clock; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_reset; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_ins_0; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_ins_1; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_ins_2; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_ins_3; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_ins_4; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_ins_5; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_ins_6; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_ins_7; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_outs_0; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_outs_1; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_outs_2; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_outs_3; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_outs_4; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_outs_5; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_outs_6; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_outs_7; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_15_clock; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_reset; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_ins_0; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_ins_1; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_ins_2; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_ins_3; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_ins_4; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_ins_5; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_ins_6; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_ins_7; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_outs_0; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_outs_1; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_outs_2; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_outs_3; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_outs_4; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_outs_5; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_outs_6; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_outs_7; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@10675.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@10675.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@10675.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@10675.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@10675.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@10683.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@10683.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@10683.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@10683.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@10683.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@10691.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@10691.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@10691.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@10691.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@10691.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@10699.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@10699.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@10699.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@10699.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@10699.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@10723.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@10723.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@10723.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@10723.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@10723.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@10731.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@10731.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@10731.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@10731.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@10731.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@10739.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@10739.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@10739.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@10739.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@10739.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@10747.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@10747.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@10747.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@10747.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@10747.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@10771.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@10771.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@10771.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@10771.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@10771.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@10779.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@10779.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@10779.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@10779.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@10779.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@10787.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@10787.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@10787.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@10787.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@10787.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@10795.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@10795.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@10795.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@10795.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@10795.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@10819.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@10819.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@10819.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@10819.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@10819.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@10827.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@10827.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@10827.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@10827.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@10827.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@10835.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@10835.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@10835.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@10835.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@10835.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@10843.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@10843.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@10843.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@10843.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@10843.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@10867.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@10867.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@10867.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@10867.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@10867.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@10875.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@10875.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@10875.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@10875.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@10875.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@10883.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@10883.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@10883.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@10883.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@10883.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@10891.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@10891.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@10891.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@10891.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@10891.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@10915.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@10915.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@10915.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@10915.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@10915.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@10923.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@10923.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@10923.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@10923.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@10923.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@10931.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@10931.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@10931.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@10931.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@10931.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@10939.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@10939.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@10939.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@10939.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@10939.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@10963.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@10963.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@10963.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@10963.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@10963.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@10971.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@10971.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@10971.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@10971.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@10971.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@10979.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@10979.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@10979.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@10979.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@10979.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@10987.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@10987.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@10987.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@10987.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@10987.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@11011.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@11011.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@11011.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@11011.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@11011.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@11019.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@11019.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@11019.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@11019.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@11019.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@11027.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@11027.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@11027.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@11027.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@11027.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@11035.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@11035.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@11035.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@11035.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@11035.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@11059.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@11059.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@11059.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@11059.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@11059.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@11067.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@11067.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@11067.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@11067.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@11067.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@11075.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@11075.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@11075.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@11075.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@11075.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@11083.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@11083.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@11083.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@11083.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@11083.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@11107.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@11107.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@11107.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@11107.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@11107.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@11115.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@11115.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@11115.4]
  wire  RetimeWrapper_37_io_in; // @[package.scala 93:22:@11115.4]
  wire  RetimeWrapper_37_io_out; // @[package.scala 93:22:@11115.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@11123.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@11123.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@11123.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@11123.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@11123.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@11131.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@11131.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@11131.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@11131.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@11131.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@11155.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@11155.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@11155.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@11155.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@11155.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@11163.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@11163.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@11163.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@11163.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@11163.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@11171.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@11171.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@11171.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@11171.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@11171.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@11179.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@11179.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@11179.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@11179.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@11179.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@11203.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@11203.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@11203.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@11203.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@11203.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@11211.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@11211.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@11211.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@11211.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@11211.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@11219.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@11219.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@11219.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@11219.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@11219.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@11227.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@11227.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@11227.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@11227.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@11227.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@11251.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@11251.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@11251.4]
  wire  RetimeWrapper_48_io_in; // @[package.scala 93:22:@11251.4]
  wire  RetimeWrapper_48_io_out; // @[package.scala 93:22:@11251.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@11259.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@11259.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@11259.4]
  wire  RetimeWrapper_49_io_in; // @[package.scala 93:22:@11259.4]
  wire  RetimeWrapper_49_io_out; // @[package.scala 93:22:@11259.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@11267.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@11267.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@11267.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@11267.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@11267.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@11275.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@11275.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@11275.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@11275.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@11275.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@11299.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@11299.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@11299.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@11299.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@11299.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@11307.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@11307.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@11307.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@11307.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@11307.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@11315.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@11315.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@11315.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@11315.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@11315.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@11323.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@11323.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@11323.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@11323.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@11323.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@11347.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@11347.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@11347.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@11347.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@11347.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@11355.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@11355.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@11355.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@11355.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@11355.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@11363.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@11363.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@11363.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@11363.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@11363.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@11371.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@11371.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@11371.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@11371.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@11371.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@11395.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@11395.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@11395.4]
  wire  RetimeWrapper_60_io_in; // @[package.scala 93:22:@11395.4]
  wire  RetimeWrapper_60_io_out; // @[package.scala 93:22:@11395.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@11403.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@11403.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@11403.4]
  wire  RetimeWrapper_61_io_in; // @[package.scala 93:22:@11403.4]
  wire  RetimeWrapper_61_io_out; // @[package.scala 93:22:@11403.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@11411.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@11411.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@11411.4]
  wire  RetimeWrapper_62_io_in; // @[package.scala 93:22:@11411.4]
  wire  RetimeWrapper_62_io_out; // @[package.scala 93:22:@11411.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@11419.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@11419.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@11419.4]
  wire  RetimeWrapper_63_io_in; // @[package.scala 93:22:@11419.4]
  wire  RetimeWrapper_63_io_out; // @[package.scala 93:22:@11419.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@11443.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@11443.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@11443.4]
  wire  RetimeWrapper_64_io_in; // @[package.scala 93:22:@11443.4]
  wire  RetimeWrapper_64_io_out; // @[package.scala 93:22:@11443.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@11451.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@11451.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@11451.4]
  wire  RetimeWrapper_65_io_in; // @[package.scala 93:22:@11451.4]
  wire  RetimeWrapper_65_io_out; // @[package.scala 93:22:@11451.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@11459.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@11459.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@11459.4]
  wire  RetimeWrapper_66_io_in; // @[package.scala 93:22:@11459.4]
  wire  RetimeWrapper_66_io_out; // @[package.scala 93:22:@11459.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@11467.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@11467.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@11467.4]
  wire  RetimeWrapper_67_io_in; // @[package.scala 93:22:@11467.4]
  wire  RetimeWrapper_67_io_out; // @[package.scala 93:22:@11467.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@11491.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@11491.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@11491.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@11491.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@11491.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@11499.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@11499.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@11499.4]
  wire  RetimeWrapper_69_io_in; // @[package.scala 93:22:@11499.4]
  wire  RetimeWrapper_69_io_out; // @[package.scala 93:22:@11499.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@11507.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@11507.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@11507.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@11507.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@11507.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@11515.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@11515.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@11515.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@11515.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@11515.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@11539.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@11539.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@11539.4]
  wire  RetimeWrapper_72_io_in; // @[package.scala 93:22:@11539.4]
  wire  RetimeWrapper_72_io_out; // @[package.scala 93:22:@11539.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@11547.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@11547.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@11547.4]
  wire  RetimeWrapper_73_io_in; // @[package.scala 93:22:@11547.4]
  wire  RetimeWrapper_73_io_out; // @[package.scala 93:22:@11547.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@11555.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@11555.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@11555.4]
  wire  RetimeWrapper_74_io_in; // @[package.scala 93:22:@11555.4]
  wire  RetimeWrapper_74_io_out; // @[package.scala 93:22:@11555.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@11563.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@11563.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@11563.4]
  wire  RetimeWrapper_75_io_in; // @[package.scala 93:22:@11563.4]
  wire  RetimeWrapper_75_io_out; // @[package.scala 93:22:@11563.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@11587.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@11587.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@11587.4]
  wire  RetimeWrapper_76_io_in; // @[package.scala 93:22:@11587.4]
  wire  RetimeWrapper_76_io_out; // @[package.scala 93:22:@11587.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@11595.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@11595.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@11595.4]
  wire  RetimeWrapper_77_io_in; // @[package.scala 93:22:@11595.4]
  wire  RetimeWrapper_77_io_out; // @[package.scala 93:22:@11595.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@11603.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@11603.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@11603.4]
  wire  RetimeWrapper_78_io_in; // @[package.scala 93:22:@11603.4]
  wire  RetimeWrapper_78_io_out; // @[package.scala 93:22:@11603.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@11611.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@11611.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@11611.4]
  wire  RetimeWrapper_79_io_in; // @[package.scala 93:22:@11611.4]
  wire  RetimeWrapper_79_io_out; // @[package.scala 93:22:@11611.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@11635.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@11635.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@11635.4]
  wire  RetimeWrapper_80_io_in; // @[package.scala 93:22:@11635.4]
  wire  RetimeWrapper_80_io_out; // @[package.scala 93:22:@11635.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@11643.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@11643.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@11643.4]
  wire  RetimeWrapper_81_io_in; // @[package.scala 93:22:@11643.4]
  wire  RetimeWrapper_81_io_out; // @[package.scala 93:22:@11643.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@11651.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@11651.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@11651.4]
  wire  RetimeWrapper_82_io_in; // @[package.scala 93:22:@11651.4]
  wire  RetimeWrapper_82_io_out; // @[package.scala 93:22:@11651.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@11659.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@11659.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@11659.4]
  wire  RetimeWrapper_83_io_in; // @[package.scala 93:22:@11659.4]
  wire  RetimeWrapper_83_io_out; // @[package.scala 93:22:@11659.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@11683.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@11683.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@11683.4]
  wire  RetimeWrapper_84_io_in; // @[package.scala 93:22:@11683.4]
  wire  RetimeWrapper_84_io_out; // @[package.scala 93:22:@11683.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@11691.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@11691.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@11691.4]
  wire  RetimeWrapper_85_io_in; // @[package.scala 93:22:@11691.4]
  wire  RetimeWrapper_85_io_out; // @[package.scala 93:22:@11691.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@11699.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@11699.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@11699.4]
  wire  RetimeWrapper_86_io_in; // @[package.scala 93:22:@11699.4]
  wire  RetimeWrapper_86_io_out; // @[package.scala 93:22:@11699.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@11707.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@11707.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@11707.4]
  wire  RetimeWrapper_87_io_in; // @[package.scala 93:22:@11707.4]
  wire  RetimeWrapper_87_io_out; // @[package.scala 93:22:@11707.4]
  wire  RetimeWrapper_88_clock; // @[package.scala 93:22:@11731.4]
  wire  RetimeWrapper_88_reset; // @[package.scala 93:22:@11731.4]
  wire  RetimeWrapper_88_io_flow; // @[package.scala 93:22:@11731.4]
  wire  RetimeWrapper_88_io_in; // @[package.scala 93:22:@11731.4]
  wire  RetimeWrapper_88_io_out; // @[package.scala 93:22:@11731.4]
  wire  RetimeWrapper_89_clock; // @[package.scala 93:22:@11739.4]
  wire  RetimeWrapper_89_reset; // @[package.scala 93:22:@11739.4]
  wire  RetimeWrapper_89_io_flow; // @[package.scala 93:22:@11739.4]
  wire  RetimeWrapper_89_io_in; // @[package.scala 93:22:@11739.4]
  wire  RetimeWrapper_89_io_out; // @[package.scala 93:22:@11739.4]
  wire  RetimeWrapper_90_clock; // @[package.scala 93:22:@11747.4]
  wire  RetimeWrapper_90_reset; // @[package.scala 93:22:@11747.4]
  wire  RetimeWrapper_90_io_flow; // @[package.scala 93:22:@11747.4]
  wire  RetimeWrapper_90_io_in; // @[package.scala 93:22:@11747.4]
  wire  RetimeWrapper_90_io_out; // @[package.scala 93:22:@11747.4]
  wire  RetimeWrapper_91_clock; // @[package.scala 93:22:@11755.4]
  wire  RetimeWrapper_91_reset; // @[package.scala 93:22:@11755.4]
  wire  RetimeWrapper_91_io_flow; // @[package.scala 93:22:@11755.4]
  wire  RetimeWrapper_91_io_in; // @[package.scala 93:22:@11755.4]
  wire  RetimeWrapper_91_io_out; // @[package.scala 93:22:@11755.4]
  wire  RetimeWrapper_92_clock; // @[package.scala 93:22:@11779.4]
  wire  RetimeWrapper_92_reset; // @[package.scala 93:22:@11779.4]
  wire  RetimeWrapper_92_io_flow; // @[package.scala 93:22:@11779.4]
  wire  RetimeWrapper_92_io_in; // @[package.scala 93:22:@11779.4]
  wire  RetimeWrapper_92_io_out; // @[package.scala 93:22:@11779.4]
  wire  RetimeWrapper_93_clock; // @[package.scala 93:22:@11787.4]
  wire  RetimeWrapper_93_reset; // @[package.scala 93:22:@11787.4]
  wire  RetimeWrapper_93_io_flow; // @[package.scala 93:22:@11787.4]
  wire  RetimeWrapper_93_io_in; // @[package.scala 93:22:@11787.4]
  wire  RetimeWrapper_93_io_out; // @[package.scala 93:22:@11787.4]
  wire  RetimeWrapper_94_clock; // @[package.scala 93:22:@11795.4]
  wire  RetimeWrapper_94_reset; // @[package.scala 93:22:@11795.4]
  wire  RetimeWrapper_94_io_flow; // @[package.scala 93:22:@11795.4]
  wire  RetimeWrapper_94_io_in; // @[package.scala 93:22:@11795.4]
  wire  RetimeWrapper_94_io_out; // @[package.scala 93:22:@11795.4]
  wire  RetimeWrapper_95_clock; // @[package.scala 93:22:@11803.4]
  wire  RetimeWrapper_95_reset; // @[package.scala 93:22:@11803.4]
  wire  RetimeWrapper_95_io_flow; // @[package.scala 93:22:@11803.4]
  wire  RetimeWrapper_95_io_in; // @[package.scala 93:22:@11803.4]
  wire  RetimeWrapper_95_io_out; // @[package.scala 93:22:@11803.4]
  wire  _T_1032; // @[MemPrimitives.scala 82:210:@9494.4]
  wire  _T_1035; // @[MemPrimitives.scala 83:102:@9496.4]
  wire  _T_1037; // @[MemPrimitives.scala 82:210:@9497.4]
  wire  _T_1040; // @[MemPrimitives.scala 83:102:@9499.4]
  wire [9:0] _T_1042; // @[Cat.scala 30:58:@9501.4]
  wire [9:0] _T_1044; // @[Cat.scala 30:58:@9503.4]
  wire [9:0] _T_1045; // @[Mux.scala 31:69:@9504.4]
  wire  _T_1050; // @[MemPrimitives.scala 82:210:@9511.4]
  wire  _T_1053; // @[MemPrimitives.scala 83:102:@9513.4]
  wire  _T_1055; // @[MemPrimitives.scala 82:210:@9514.4]
  wire  _T_1058; // @[MemPrimitives.scala 83:102:@9516.4]
  wire [9:0] _T_1060; // @[Cat.scala 30:58:@9518.4]
  wire [9:0] _T_1062; // @[Cat.scala 30:58:@9520.4]
  wire [9:0] _T_1063; // @[Mux.scala 31:69:@9521.4]
  wire  _T_1068; // @[MemPrimitives.scala 82:210:@9528.4]
  wire  _T_1071; // @[MemPrimitives.scala 83:102:@9530.4]
  wire  _T_1073; // @[MemPrimitives.scala 82:210:@9531.4]
  wire  _T_1076; // @[MemPrimitives.scala 83:102:@9533.4]
  wire [9:0] _T_1078; // @[Cat.scala 30:58:@9535.4]
  wire [9:0] _T_1080; // @[Cat.scala 30:58:@9537.4]
  wire [9:0] _T_1081; // @[Mux.scala 31:69:@9538.4]
  wire  _T_1086; // @[MemPrimitives.scala 82:210:@9545.4]
  wire  _T_1089; // @[MemPrimitives.scala 83:102:@9547.4]
  wire  _T_1091; // @[MemPrimitives.scala 82:210:@9548.4]
  wire  _T_1094; // @[MemPrimitives.scala 83:102:@9550.4]
  wire [9:0] _T_1096; // @[Cat.scala 30:58:@9552.4]
  wire [9:0] _T_1098; // @[Cat.scala 30:58:@9554.4]
  wire [9:0] _T_1099; // @[Mux.scala 31:69:@9555.4]
  wire  _T_1104; // @[MemPrimitives.scala 82:210:@9562.4]
  wire  _T_1107; // @[MemPrimitives.scala 83:102:@9564.4]
  wire  _T_1109; // @[MemPrimitives.scala 82:210:@9565.4]
  wire  _T_1112; // @[MemPrimitives.scala 83:102:@9567.4]
  wire [9:0] _T_1114; // @[Cat.scala 30:58:@9569.4]
  wire [9:0] _T_1116; // @[Cat.scala 30:58:@9571.4]
  wire [9:0] _T_1117; // @[Mux.scala 31:69:@9572.4]
  wire  _T_1122; // @[MemPrimitives.scala 82:210:@9579.4]
  wire  _T_1125; // @[MemPrimitives.scala 83:102:@9581.4]
  wire  _T_1127; // @[MemPrimitives.scala 82:210:@9582.4]
  wire  _T_1130; // @[MemPrimitives.scala 83:102:@9584.4]
  wire [9:0] _T_1132; // @[Cat.scala 30:58:@9586.4]
  wire [9:0] _T_1134; // @[Cat.scala 30:58:@9588.4]
  wire [9:0] _T_1135; // @[Mux.scala 31:69:@9589.4]
  wire  _T_1140; // @[MemPrimitives.scala 82:210:@9596.4]
  wire  _T_1143; // @[MemPrimitives.scala 83:102:@9598.4]
  wire  _T_1145; // @[MemPrimitives.scala 82:210:@9599.4]
  wire  _T_1148; // @[MemPrimitives.scala 83:102:@9601.4]
  wire [9:0] _T_1150; // @[Cat.scala 30:58:@9603.4]
  wire [9:0] _T_1152; // @[Cat.scala 30:58:@9605.4]
  wire [9:0] _T_1153; // @[Mux.scala 31:69:@9606.4]
  wire  _T_1158; // @[MemPrimitives.scala 82:210:@9613.4]
  wire  _T_1161; // @[MemPrimitives.scala 83:102:@9615.4]
  wire  _T_1163; // @[MemPrimitives.scala 82:210:@9616.4]
  wire  _T_1166; // @[MemPrimitives.scala 83:102:@9618.4]
  wire [9:0] _T_1168; // @[Cat.scala 30:58:@9620.4]
  wire [9:0] _T_1170; // @[Cat.scala 30:58:@9622.4]
  wire [9:0] _T_1171; // @[Mux.scala 31:69:@9623.4]
  wire  _T_1176; // @[MemPrimitives.scala 82:210:@9630.4]
  wire  _T_1179; // @[MemPrimitives.scala 83:102:@9632.4]
  wire  _T_1181; // @[MemPrimitives.scala 82:210:@9633.4]
  wire  _T_1184; // @[MemPrimitives.scala 83:102:@9635.4]
  wire [9:0] _T_1186; // @[Cat.scala 30:58:@9637.4]
  wire [9:0] _T_1188; // @[Cat.scala 30:58:@9639.4]
  wire [9:0] _T_1189; // @[Mux.scala 31:69:@9640.4]
  wire  _T_1194; // @[MemPrimitives.scala 82:210:@9647.4]
  wire  _T_1197; // @[MemPrimitives.scala 83:102:@9649.4]
  wire  _T_1199; // @[MemPrimitives.scala 82:210:@9650.4]
  wire  _T_1202; // @[MemPrimitives.scala 83:102:@9652.4]
  wire [9:0] _T_1204; // @[Cat.scala 30:58:@9654.4]
  wire [9:0] _T_1206; // @[Cat.scala 30:58:@9656.4]
  wire [9:0] _T_1207; // @[Mux.scala 31:69:@9657.4]
  wire  _T_1212; // @[MemPrimitives.scala 82:210:@9664.4]
  wire  _T_1215; // @[MemPrimitives.scala 83:102:@9666.4]
  wire  _T_1217; // @[MemPrimitives.scala 82:210:@9667.4]
  wire  _T_1220; // @[MemPrimitives.scala 83:102:@9669.4]
  wire [9:0] _T_1222; // @[Cat.scala 30:58:@9671.4]
  wire [9:0] _T_1224; // @[Cat.scala 30:58:@9673.4]
  wire [9:0] _T_1225; // @[Mux.scala 31:69:@9674.4]
  wire  _T_1230; // @[MemPrimitives.scala 82:210:@9681.4]
  wire  _T_1233; // @[MemPrimitives.scala 83:102:@9683.4]
  wire  _T_1235; // @[MemPrimitives.scala 82:210:@9684.4]
  wire  _T_1238; // @[MemPrimitives.scala 83:102:@9686.4]
  wire [9:0] _T_1240; // @[Cat.scala 30:58:@9688.4]
  wire [9:0] _T_1242; // @[Cat.scala 30:58:@9690.4]
  wire [9:0] _T_1243; // @[Mux.scala 31:69:@9691.4]
  wire  _T_1248; // @[MemPrimitives.scala 82:210:@9698.4]
  wire  _T_1251; // @[MemPrimitives.scala 83:102:@9700.4]
  wire  _T_1253; // @[MemPrimitives.scala 82:210:@9701.4]
  wire  _T_1256; // @[MemPrimitives.scala 83:102:@9703.4]
  wire [9:0] _T_1258; // @[Cat.scala 30:58:@9705.4]
  wire [9:0] _T_1260; // @[Cat.scala 30:58:@9707.4]
  wire [9:0] _T_1261; // @[Mux.scala 31:69:@9708.4]
  wire  _T_1266; // @[MemPrimitives.scala 82:210:@9715.4]
  wire  _T_1269; // @[MemPrimitives.scala 83:102:@9717.4]
  wire  _T_1271; // @[MemPrimitives.scala 82:210:@9718.4]
  wire  _T_1274; // @[MemPrimitives.scala 83:102:@9720.4]
  wire [9:0] _T_1276; // @[Cat.scala 30:58:@9722.4]
  wire [9:0] _T_1278; // @[Cat.scala 30:58:@9724.4]
  wire [9:0] _T_1279; // @[Mux.scala 31:69:@9725.4]
  wire  _T_1284; // @[MemPrimitives.scala 82:210:@9732.4]
  wire  _T_1287; // @[MemPrimitives.scala 83:102:@9734.4]
  wire  _T_1289; // @[MemPrimitives.scala 82:210:@9735.4]
  wire  _T_1292; // @[MemPrimitives.scala 83:102:@9737.4]
  wire [9:0] _T_1294; // @[Cat.scala 30:58:@9739.4]
  wire [9:0] _T_1296; // @[Cat.scala 30:58:@9741.4]
  wire [9:0] _T_1297; // @[Mux.scala 31:69:@9742.4]
  wire  _T_1302; // @[MemPrimitives.scala 82:210:@9749.4]
  wire  _T_1305; // @[MemPrimitives.scala 83:102:@9751.4]
  wire  _T_1307; // @[MemPrimitives.scala 82:210:@9752.4]
  wire  _T_1310; // @[MemPrimitives.scala 83:102:@9754.4]
  wire [9:0] _T_1312; // @[Cat.scala 30:58:@9756.4]
  wire [9:0] _T_1314; // @[Cat.scala 30:58:@9758.4]
  wire [9:0] _T_1315; // @[Mux.scala 31:69:@9759.4]
  wire  _T_1320; // @[MemPrimitives.scala 110:210:@9766.4]
  wire  _T_1325; // @[MemPrimitives.scala 110:210:@9769.4]
  wire  _T_1330; // @[MemPrimitives.scala 110:210:@9772.4]
  wire  _T_1335; // @[MemPrimitives.scala 110:210:@9775.4]
  wire  _T_1339; // @[MemPrimitives.scala 123:41:@9785.4]
  wire  _T_1340; // @[MemPrimitives.scala 123:41:@9786.4]
  wire  _T_1341; // @[MemPrimitives.scala 123:41:@9787.4]
  wire  _T_1342; // @[MemPrimitives.scala 123:41:@9788.4]
  wire [2:0] _T_1344; // @[Cat.scala 30:58:@9790.4]
  wire [2:0] _T_1346; // @[Cat.scala 30:58:@9792.4]
  wire [2:0] _T_1348; // @[Cat.scala 30:58:@9794.4]
  wire [2:0] _T_1350; // @[Cat.scala 30:58:@9796.4]
  wire [2:0] _T_1351; // @[Mux.scala 31:69:@9797.4]
  wire [2:0] _T_1352; // @[Mux.scala 31:69:@9798.4]
  wire [2:0] _T_1353; // @[Mux.scala 31:69:@9799.4]
  wire  _T_1358; // @[MemPrimitives.scala 110:210:@9806.4]
  wire  _T_1363; // @[MemPrimitives.scala 110:210:@9809.4]
  wire  _T_1368; // @[MemPrimitives.scala 110:210:@9812.4]
  wire  _T_1373; // @[MemPrimitives.scala 110:210:@9815.4]
  wire  _T_1377; // @[MemPrimitives.scala 123:41:@9825.4]
  wire  _T_1378; // @[MemPrimitives.scala 123:41:@9826.4]
  wire  _T_1379; // @[MemPrimitives.scala 123:41:@9827.4]
  wire  _T_1380; // @[MemPrimitives.scala 123:41:@9828.4]
  wire [2:0] _T_1382; // @[Cat.scala 30:58:@9830.4]
  wire [2:0] _T_1384; // @[Cat.scala 30:58:@9832.4]
  wire [2:0] _T_1386; // @[Cat.scala 30:58:@9834.4]
  wire [2:0] _T_1388; // @[Cat.scala 30:58:@9836.4]
  wire [2:0] _T_1389; // @[Mux.scala 31:69:@9837.4]
  wire [2:0] _T_1390; // @[Mux.scala 31:69:@9838.4]
  wire [2:0] _T_1391; // @[Mux.scala 31:69:@9839.4]
  wire  _T_1396; // @[MemPrimitives.scala 110:210:@9846.4]
  wire  _T_1401; // @[MemPrimitives.scala 110:210:@9849.4]
  wire  _T_1406; // @[MemPrimitives.scala 110:210:@9852.4]
  wire  _T_1411; // @[MemPrimitives.scala 110:210:@9855.4]
  wire  _T_1416; // @[MemPrimitives.scala 110:210:@9858.4]
  wire  _T_1421; // @[MemPrimitives.scala 110:210:@9861.4]
  wire  _T_1426; // @[MemPrimitives.scala 110:210:@9864.4]
  wire  _T_1431; // @[MemPrimitives.scala 110:210:@9867.4]
  wire  _T_1435; // @[MemPrimitives.scala 123:41:@9881.4]
  wire  _T_1436; // @[MemPrimitives.scala 123:41:@9882.4]
  wire  _T_1437; // @[MemPrimitives.scala 123:41:@9883.4]
  wire  _T_1438; // @[MemPrimitives.scala 123:41:@9884.4]
  wire  _T_1439; // @[MemPrimitives.scala 123:41:@9885.4]
  wire  _T_1440; // @[MemPrimitives.scala 123:41:@9886.4]
  wire  _T_1441; // @[MemPrimitives.scala 123:41:@9887.4]
  wire  _T_1442; // @[MemPrimitives.scala 123:41:@9888.4]
  wire [2:0] _T_1444; // @[Cat.scala 30:58:@9890.4]
  wire [2:0] _T_1446; // @[Cat.scala 30:58:@9892.4]
  wire [2:0] _T_1448; // @[Cat.scala 30:58:@9894.4]
  wire [2:0] _T_1450; // @[Cat.scala 30:58:@9896.4]
  wire [2:0] _T_1452; // @[Cat.scala 30:58:@9898.4]
  wire [2:0] _T_1454; // @[Cat.scala 30:58:@9900.4]
  wire [2:0] _T_1456; // @[Cat.scala 30:58:@9902.4]
  wire [2:0] _T_1458; // @[Cat.scala 30:58:@9904.4]
  wire [2:0] _T_1459; // @[Mux.scala 31:69:@9905.4]
  wire [2:0] _T_1460; // @[Mux.scala 31:69:@9906.4]
  wire [2:0] _T_1461; // @[Mux.scala 31:69:@9907.4]
  wire [2:0] _T_1462; // @[Mux.scala 31:69:@9908.4]
  wire [2:0] _T_1463; // @[Mux.scala 31:69:@9909.4]
  wire [2:0] _T_1464; // @[Mux.scala 31:69:@9910.4]
  wire [2:0] _T_1465; // @[Mux.scala 31:69:@9911.4]
  wire  _T_1470; // @[MemPrimitives.scala 110:210:@9918.4]
  wire  _T_1475; // @[MemPrimitives.scala 110:210:@9921.4]
  wire  _T_1480; // @[MemPrimitives.scala 110:210:@9924.4]
  wire  _T_1485; // @[MemPrimitives.scala 110:210:@9927.4]
  wire  _T_1490; // @[MemPrimitives.scala 110:210:@9930.4]
  wire  _T_1495; // @[MemPrimitives.scala 110:210:@9933.4]
  wire  _T_1500; // @[MemPrimitives.scala 110:210:@9936.4]
  wire  _T_1505; // @[MemPrimitives.scala 110:210:@9939.4]
  wire  _T_1509; // @[MemPrimitives.scala 123:41:@9953.4]
  wire  _T_1510; // @[MemPrimitives.scala 123:41:@9954.4]
  wire  _T_1511; // @[MemPrimitives.scala 123:41:@9955.4]
  wire  _T_1512; // @[MemPrimitives.scala 123:41:@9956.4]
  wire  _T_1513; // @[MemPrimitives.scala 123:41:@9957.4]
  wire  _T_1514; // @[MemPrimitives.scala 123:41:@9958.4]
  wire  _T_1515; // @[MemPrimitives.scala 123:41:@9959.4]
  wire  _T_1516; // @[MemPrimitives.scala 123:41:@9960.4]
  wire [2:0] _T_1518; // @[Cat.scala 30:58:@9962.4]
  wire [2:0] _T_1520; // @[Cat.scala 30:58:@9964.4]
  wire [2:0] _T_1522; // @[Cat.scala 30:58:@9966.4]
  wire [2:0] _T_1524; // @[Cat.scala 30:58:@9968.4]
  wire [2:0] _T_1526; // @[Cat.scala 30:58:@9970.4]
  wire [2:0] _T_1528; // @[Cat.scala 30:58:@9972.4]
  wire [2:0] _T_1530; // @[Cat.scala 30:58:@9974.4]
  wire [2:0] _T_1532; // @[Cat.scala 30:58:@9976.4]
  wire [2:0] _T_1533; // @[Mux.scala 31:69:@9977.4]
  wire [2:0] _T_1534; // @[Mux.scala 31:69:@9978.4]
  wire [2:0] _T_1535; // @[Mux.scala 31:69:@9979.4]
  wire [2:0] _T_1536; // @[Mux.scala 31:69:@9980.4]
  wire [2:0] _T_1537; // @[Mux.scala 31:69:@9981.4]
  wire [2:0] _T_1538; // @[Mux.scala 31:69:@9982.4]
  wire [2:0] _T_1539; // @[Mux.scala 31:69:@9983.4]
  wire  _T_1544; // @[MemPrimitives.scala 110:210:@9990.4]
  wire  _T_1549; // @[MemPrimitives.scala 110:210:@9993.4]
  wire  _T_1554; // @[MemPrimitives.scala 110:210:@9996.4]
  wire  _T_1559; // @[MemPrimitives.scala 110:210:@9999.4]
  wire  _T_1563; // @[MemPrimitives.scala 123:41:@10009.4]
  wire  _T_1564; // @[MemPrimitives.scala 123:41:@10010.4]
  wire  _T_1565; // @[MemPrimitives.scala 123:41:@10011.4]
  wire  _T_1566; // @[MemPrimitives.scala 123:41:@10012.4]
  wire [2:0] _T_1568; // @[Cat.scala 30:58:@10014.4]
  wire [2:0] _T_1570; // @[Cat.scala 30:58:@10016.4]
  wire [2:0] _T_1572; // @[Cat.scala 30:58:@10018.4]
  wire [2:0] _T_1574; // @[Cat.scala 30:58:@10020.4]
  wire [2:0] _T_1575; // @[Mux.scala 31:69:@10021.4]
  wire [2:0] _T_1576; // @[Mux.scala 31:69:@10022.4]
  wire [2:0] _T_1577; // @[Mux.scala 31:69:@10023.4]
  wire  _T_1582; // @[MemPrimitives.scala 110:210:@10030.4]
  wire  _T_1587; // @[MemPrimitives.scala 110:210:@10033.4]
  wire  _T_1592; // @[MemPrimitives.scala 110:210:@10036.4]
  wire  _T_1597; // @[MemPrimitives.scala 110:210:@10039.4]
  wire  _T_1601; // @[MemPrimitives.scala 123:41:@10049.4]
  wire  _T_1602; // @[MemPrimitives.scala 123:41:@10050.4]
  wire  _T_1603; // @[MemPrimitives.scala 123:41:@10051.4]
  wire  _T_1604; // @[MemPrimitives.scala 123:41:@10052.4]
  wire [2:0] _T_1606; // @[Cat.scala 30:58:@10054.4]
  wire [2:0] _T_1608; // @[Cat.scala 30:58:@10056.4]
  wire [2:0] _T_1610; // @[Cat.scala 30:58:@10058.4]
  wire [2:0] _T_1612; // @[Cat.scala 30:58:@10060.4]
  wire [2:0] _T_1613; // @[Mux.scala 31:69:@10061.4]
  wire [2:0] _T_1614; // @[Mux.scala 31:69:@10062.4]
  wire [2:0] _T_1615; // @[Mux.scala 31:69:@10063.4]
  wire  _T_1620; // @[MemPrimitives.scala 110:210:@10070.4]
  wire  _T_1625; // @[MemPrimitives.scala 110:210:@10073.4]
  wire  _T_1630; // @[MemPrimitives.scala 110:210:@10076.4]
  wire  _T_1635; // @[MemPrimitives.scala 110:210:@10079.4]
  wire  _T_1640; // @[MemPrimitives.scala 110:210:@10082.4]
  wire  _T_1645; // @[MemPrimitives.scala 110:210:@10085.4]
  wire  _T_1650; // @[MemPrimitives.scala 110:210:@10088.4]
  wire  _T_1655; // @[MemPrimitives.scala 110:210:@10091.4]
  wire  _T_1659; // @[MemPrimitives.scala 123:41:@10105.4]
  wire  _T_1660; // @[MemPrimitives.scala 123:41:@10106.4]
  wire  _T_1661; // @[MemPrimitives.scala 123:41:@10107.4]
  wire  _T_1662; // @[MemPrimitives.scala 123:41:@10108.4]
  wire  _T_1663; // @[MemPrimitives.scala 123:41:@10109.4]
  wire  _T_1664; // @[MemPrimitives.scala 123:41:@10110.4]
  wire  _T_1665; // @[MemPrimitives.scala 123:41:@10111.4]
  wire  _T_1666; // @[MemPrimitives.scala 123:41:@10112.4]
  wire [2:0] _T_1668; // @[Cat.scala 30:58:@10114.4]
  wire [2:0] _T_1670; // @[Cat.scala 30:58:@10116.4]
  wire [2:0] _T_1672; // @[Cat.scala 30:58:@10118.4]
  wire [2:0] _T_1674; // @[Cat.scala 30:58:@10120.4]
  wire [2:0] _T_1676; // @[Cat.scala 30:58:@10122.4]
  wire [2:0] _T_1678; // @[Cat.scala 30:58:@10124.4]
  wire [2:0] _T_1680; // @[Cat.scala 30:58:@10126.4]
  wire [2:0] _T_1682; // @[Cat.scala 30:58:@10128.4]
  wire [2:0] _T_1683; // @[Mux.scala 31:69:@10129.4]
  wire [2:0] _T_1684; // @[Mux.scala 31:69:@10130.4]
  wire [2:0] _T_1685; // @[Mux.scala 31:69:@10131.4]
  wire [2:0] _T_1686; // @[Mux.scala 31:69:@10132.4]
  wire [2:0] _T_1687; // @[Mux.scala 31:69:@10133.4]
  wire [2:0] _T_1688; // @[Mux.scala 31:69:@10134.4]
  wire [2:0] _T_1689; // @[Mux.scala 31:69:@10135.4]
  wire  _T_1694; // @[MemPrimitives.scala 110:210:@10142.4]
  wire  _T_1699; // @[MemPrimitives.scala 110:210:@10145.4]
  wire  _T_1704; // @[MemPrimitives.scala 110:210:@10148.4]
  wire  _T_1709; // @[MemPrimitives.scala 110:210:@10151.4]
  wire  _T_1714; // @[MemPrimitives.scala 110:210:@10154.4]
  wire  _T_1719; // @[MemPrimitives.scala 110:210:@10157.4]
  wire  _T_1724; // @[MemPrimitives.scala 110:210:@10160.4]
  wire  _T_1729; // @[MemPrimitives.scala 110:210:@10163.4]
  wire  _T_1733; // @[MemPrimitives.scala 123:41:@10177.4]
  wire  _T_1734; // @[MemPrimitives.scala 123:41:@10178.4]
  wire  _T_1735; // @[MemPrimitives.scala 123:41:@10179.4]
  wire  _T_1736; // @[MemPrimitives.scala 123:41:@10180.4]
  wire  _T_1737; // @[MemPrimitives.scala 123:41:@10181.4]
  wire  _T_1738; // @[MemPrimitives.scala 123:41:@10182.4]
  wire  _T_1739; // @[MemPrimitives.scala 123:41:@10183.4]
  wire  _T_1740; // @[MemPrimitives.scala 123:41:@10184.4]
  wire [2:0] _T_1742; // @[Cat.scala 30:58:@10186.4]
  wire [2:0] _T_1744; // @[Cat.scala 30:58:@10188.4]
  wire [2:0] _T_1746; // @[Cat.scala 30:58:@10190.4]
  wire [2:0] _T_1748; // @[Cat.scala 30:58:@10192.4]
  wire [2:0] _T_1750; // @[Cat.scala 30:58:@10194.4]
  wire [2:0] _T_1752; // @[Cat.scala 30:58:@10196.4]
  wire [2:0] _T_1754; // @[Cat.scala 30:58:@10198.4]
  wire [2:0] _T_1756; // @[Cat.scala 30:58:@10200.4]
  wire [2:0] _T_1757; // @[Mux.scala 31:69:@10201.4]
  wire [2:0] _T_1758; // @[Mux.scala 31:69:@10202.4]
  wire [2:0] _T_1759; // @[Mux.scala 31:69:@10203.4]
  wire [2:0] _T_1760; // @[Mux.scala 31:69:@10204.4]
  wire [2:0] _T_1761; // @[Mux.scala 31:69:@10205.4]
  wire [2:0] _T_1762; // @[Mux.scala 31:69:@10206.4]
  wire [2:0] _T_1763; // @[Mux.scala 31:69:@10207.4]
  wire  _T_1768; // @[MemPrimitives.scala 110:210:@10214.4]
  wire  _T_1773; // @[MemPrimitives.scala 110:210:@10217.4]
  wire  _T_1778; // @[MemPrimitives.scala 110:210:@10220.4]
  wire  _T_1783; // @[MemPrimitives.scala 110:210:@10223.4]
  wire  _T_1787; // @[MemPrimitives.scala 123:41:@10233.4]
  wire  _T_1788; // @[MemPrimitives.scala 123:41:@10234.4]
  wire  _T_1789; // @[MemPrimitives.scala 123:41:@10235.4]
  wire  _T_1790; // @[MemPrimitives.scala 123:41:@10236.4]
  wire [2:0] _T_1792; // @[Cat.scala 30:58:@10238.4]
  wire [2:0] _T_1794; // @[Cat.scala 30:58:@10240.4]
  wire [2:0] _T_1796; // @[Cat.scala 30:58:@10242.4]
  wire [2:0] _T_1798; // @[Cat.scala 30:58:@10244.4]
  wire [2:0] _T_1799; // @[Mux.scala 31:69:@10245.4]
  wire [2:0] _T_1800; // @[Mux.scala 31:69:@10246.4]
  wire [2:0] _T_1801; // @[Mux.scala 31:69:@10247.4]
  wire  _T_1806; // @[MemPrimitives.scala 110:210:@10254.4]
  wire  _T_1811; // @[MemPrimitives.scala 110:210:@10257.4]
  wire  _T_1816; // @[MemPrimitives.scala 110:210:@10260.4]
  wire  _T_1821; // @[MemPrimitives.scala 110:210:@10263.4]
  wire  _T_1825; // @[MemPrimitives.scala 123:41:@10273.4]
  wire  _T_1826; // @[MemPrimitives.scala 123:41:@10274.4]
  wire  _T_1827; // @[MemPrimitives.scala 123:41:@10275.4]
  wire  _T_1828; // @[MemPrimitives.scala 123:41:@10276.4]
  wire [2:0] _T_1830; // @[Cat.scala 30:58:@10278.4]
  wire [2:0] _T_1832; // @[Cat.scala 30:58:@10280.4]
  wire [2:0] _T_1834; // @[Cat.scala 30:58:@10282.4]
  wire [2:0] _T_1836; // @[Cat.scala 30:58:@10284.4]
  wire [2:0] _T_1837; // @[Mux.scala 31:69:@10285.4]
  wire [2:0] _T_1838; // @[Mux.scala 31:69:@10286.4]
  wire [2:0] _T_1839; // @[Mux.scala 31:69:@10287.4]
  wire  _T_1844; // @[MemPrimitives.scala 110:210:@10294.4]
  wire  _T_1849; // @[MemPrimitives.scala 110:210:@10297.4]
  wire  _T_1854; // @[MemPrimitives.scala 110:210:@10300.4]
  wire  _T_1859; // @[MemPrimitives.scala 110:210:@10303.4]
  wire  _T_1864; // @[MemPrimitives.scala 110:210:@10306.4]
  wire  _T_1869; // @[MemPrimitives.scala 110:210:@10309.4]
  wire  _T_1874; // @[MemPrimitives.scala 110:210:@10312.4]
  wire  _T_1879; // @[MemPrimitives.scala 110:210:@10315.4]
  wire  _T_1883; // @[MemPrimitives.scala 123:41:@10329.4]
  wire  _T_1884; // @[MemPrimitives.scala 123:41:@10330.4]
  wire  _T_1885; // @[MemPrimitives.scala 123:41:@10331.4]
  wire  _T_1886; // @[MemPrimitives.scala 123:41:@10332.4]
  wire  _T_1887; // @[MemPrimitives.scala 123:41:@10333.4]
  wire  _T_1888; // @[MemPrimitives.scala 123:41:@10334.4]
  wire  _T_1889; // @[MemPrimitives.scala 123:41:@10335.4]
  wire  _T_1890; // @[MemPrimitives.scala 123:41:@10336.4]
  wire [2:0] _T_1892; // @[Cat.scala 30:58:@10338.4]
  wire [2:0] _T_1894; // @[Cat.scala 30:58:@10340.4]
  wire [2:0] _T_1896; // @[Cat.scala 30:58:@10342.4]
  wire [2:0] _T_1898; // @[Cat.scala 30:58:@10344.4]
  wire [2:0] _T_1900; // @[Cat.scala 30:58:@10346.4]
  wire [2:0] _T_1902; // @[Cat.scala 30:58:@10348.4]
  wire [2:0] _T_1904; // @[Cat.scala 30:58:@10350.4]
  wire [2:0] _T_1906; // @[Cat.scala 30:58:@10352.4]
  wire [2:0] _T_1907; // @[Mux.scala 31:69:@10353.4]
  wire [2:0] _T_1908; // @[Mux.scala 31:69:@10354.4]
  wire [2:0] _T_1909; // @[Mux.scala 31:69:@10355.4]
  wire [2:0] _T_1910; // @[Mux.scala 31:69:@10356.4]
  wire [2:0] _T_1911; // @[Mux.scala 31:69:@10357.4]
  wire [2:0] _T_1912; // @[Mux.scala 31:69:@10358.4]
  wire [2:0] _T_1913; // @[Mux.scala 31:69:@10359.4]
  wire  _T_1918; // @[MemPrimitives.scala 110:210:@10366.4]
  wire  _T_1923; // @[MemPrimitives.scala 110:210:@10369.4]
  wire  _T_1928; // @[MemPrimitives.scala 110:210:@10372.4]
  wire  _T_1933; // @[MemPrimitives.scala 110:210:@10375.4]
  wire  _T_1938; // @[MemPrimitives.scala 110:210:@10378.4]
  wire  _T_1943; // @[MemPrimitives.scala 110:210:@10381.4]
  wire  _T_1948; // @[MemPrimitives.scala 110:210:@10384.4]
  wire  _T_1953; // @[MemPrimitives.scala 110:210:@10387.4]
  wire  _T_1957; // @[MemPrimitives.scala 123:41:@10401.4]
  wire  _T_1958; // @[MemPrimitives.scala 123:41:@10402.4]
  wire  _T_1959; // @[MemPrimitives.scala 123:41:@10403.4]
  wire  _T_1960; // @[MemPrimitives.scala 123:41:@10404.4]
  wire  _T_1961; // @[MemPrimitives.scala 123:41:@10405.4]
  wire  _T_1962; // @[MemPrimitives.scala 123:41:@10406.4]
  wire  _T_1963; // @[MemPrimitives.scala 123:41:@10407.4]
  wire  _T_1964; // @[MemPrimitives.scala 123:41:@10408.4]
  wire [2:0] _T_1966; // @[Cat.scala 30:58:@10410.4]
  wire [2:0] _T_1968; // @[Cat.scala 30:58:@10412.4]
  wire [2:0] _T_1970; // @[Cat.scala 30:58:@10414.4]
  wire [2:0] _T_1972; // @[Cat.scala 30:58:@10416.4]
  wire [2:0] _T_1974; // @[Cat.scala 30:58:@10418.4]
  wire [2:0] _T_1976; // @[Cat.scala 30:58:@10420.4]
  wire [2:0] _T_1978; // @[Cat.scala 30:58:@10422.4]
  wire [2:0] _T_1980; // @[Cat.scala 30:58:@10424.4]
  wire [2:0] _T_1981; // @[Mux.scala 31:69:@10425.4]
  wire [2:0] _T_1982; // @[Mux.scala 31:69:@10426.4]
  wire [2:0] _T_1983; // @[Mux.scala 31:69:@10427.4]
  wire [2:0] _T_1984; // @[Mux.scala 31:69:@10428.4]
  wire [2:0] _T_1985; // @[Mux.scala 31:69:@10429.4]
  wire [2:0] _T_1986; // @[Mux.scala 31:69:@10430.4]
  wire [2:0] _T_1987; // @[Mux.scala 31:69:@10431.4]
  wire  _T_1992; // @[MemPrimitives.scala 110:210:@10438.4]
  wire  _T_1997; // @[MemPrimitives.scala 110:210:@10441.4]
  wire  _T_2002; // @[MemPrimitives.scala 110:210:@10444.4]
  wire  _T_2007; // @[MemPrimitives.scala 110:210:@10447.4]
  wire  _T_2011; // @[MemPrimitives.scala 123:41:@10457.4]
  wire  _T_2012; // @[MemPrimitives.scala 123:41:@10458.4]
  wire  _T_2013; // @[MemPrimitives.scala 123:41:@10459.4]
  wire  _T_2014; // @[MemPrimitives.scala 123:41:@10460.4]
  wire [2:0] _T_2016; // @[Cat.scala 30:58:@10462.4]
  wire [2:0] _T_2018; // @[Cat.scala 30:58:@10464.4]
  wire [2:0] _T_2020; // @[Cat.scala 30:58:@10466.4]
  wire [2:0] _T_2022; // @[Cat.scala 30:58:@10468.4]
  wire [2:0] _T_2023; // @[Mux.scala 31:69:@10469.4]
  wire [2:0] _T_2024; // @[Mux.scala 31:69:@10470.4]
  wire [2:0] _T_2025; // @[Mux.scala 31:69:@10471.4]
  wire  _T_2030; // @[MemPrimitives.scala 110:210:@10478.4]
  wire  _T_2035; // @[MemPrimitives.scala 110:210:@10481.4]
  wire  _T_2040; // @[MemPrimitives.scala 110:210:@10484.4]
  wire  _T_2045; // @[MemPrimitives.scala 110:210:@10487.4]
  wire  _T_2049; // @[MemPrimitives.scala 123:41:@10497.4]
  wire  _T_2050; // @[MemPrimitives.scala 123:41:@10498.4]
  wire  _T_2051; // @[MemPrimitives.scala 123:41:@10499.4]
  wire  _T_2052; // @[MemPrimitives.scala 123:41:@10500.4]
  wire [2:0] _T_2054; // @[Cat.scala 30:58:@10502.4]
  wire [2:0] _T_2056; // @[Cat.scala 30:58:@10504.4]
  wire [2:0] _T_2058; // @[Cat.scala 30:58:@10506.4]
  wire [2:0] _T_2060; // @[Cat.scala 30:58:@10508.4]
  wire [2:0] _T_2061; // @[Mux.scala 31:69:@10509.4]
  wire [2:0] _T_2062; // @[Mux.scala 31:69:@10510.4]
  wire [2:0] _T_2063; // @[Mux.scala 31:69:@10511.4]
  wire  _T_2068; // @[MemPrimitives.scala 110:210:@10518.4]
  wire  _T_2073; // @[MemPrimitives.scala 110:210:@10521.4]
  wire  _T_2078; // @[MemPrimitives.scala 110:210:@10524.4]
  wire  _T_2083; // @[MemPrimitives.scala 110:210:@10527.4]
  wire  _T_2088; // @[MemPrimitives.scala 110:210:@10530.4]
  wire  _T_2093; // @[MemPrimitives.scala 110:210:@10533.4]
  wire  _T_2098; // @[MemPrimitives.scala 110:210:@10536.4]
  wire  _T_2103; // @[MemPrimitives.scala 110:210:@10539.4]
  wire  _T_2107; // @[MemPrimitives.scala 123:41:@10553.4]
  wire  _T_2108; // @[MemPrimitives.scala 123:41:@10554.4]
  wire  _T_2109; // @[MemPrimitives.scala 123:41:@10555.4]
  wire  _T_2110; // @[MemPrimitives.scala 123:41:@10556.4]
  wire  _T_2111; // @[MemPrimitives.scala 123:41:@10557.4]
  wire  _T_2112; // @[MemPrimitives.scala 123:41:@10558.4]
  wire  _T_2113; // @[MemPrimitives.scala 123:41:@10559.4]
  wire  _T_2114; // @[MemPrimitives.scala 123:41:@10560.4]
  wire [2:0] _T_2116; // @[Cat.scala 30:58:@10562.4]
  wire [2:0] _T_2118; // @[Cat.scala 30:58:@10564.4]
  wire [2:0] _T_2120; // @[Cat.scala 30:58:@10566.4]
  wire [2:0] _T_2122; // @[Cat.scala 30:58:@10568.4]
  wire [2:0] _T_2124; // @[Cat.scala 30:58:@10570.4]
  wire [2:0] _T_2126; // @[Cat.scala 30:58:@10572.4]
  wire [2:0] _T_2128; // @[Cat.scala 30:58:@10574.4]
  wire [2:0] _T_2130; // @[Cat.scala 30:58:@10576.4]
  wire [2:0] _T_2131; // @[Mux.scala 31:69:@10577.4]
  wire [2:0] _T_2132; // @[Mux.scala 31:69:@10578.4]
  wire [2:0] _T_2133; // @[Mux.scala 31:69:@10579.4]
  wire [2:0] _T_2134; // @[Mux.scala 31:69:@10580.4]
  wire [2:0] _T_2135; // @[Mux.scala 31:69:@10581.4]
  wire [2:0] _T_2136; // @[Mux.scala 31:69:@10582.4]
  wire [2:0] _T_2137; // @[Mux.scala 31:69:@10583.4]
  wire  _T_2142; // @[MemPrimitives.scala 110:210:@10590.4]
  wire  _T_2147; // @[MemPrimitives.scala 110:210:@10593.4]
  wire  _T_2152; // @[MemPrimitives.scala 110:210:@10596.4]
  wire  _T_2157; // @[MemPrimitives.scala 110:210:@10599.4]
  wire  _T_2162; // @[MemPrimitives.scala 110:210:@10602.4]
  wire  _T_2167; // @[MemPrimitives.scala 110:210:@10605.4]
  wire  _T_2172; // @[MemPrimitives.scala 110:210:@10608.4]
  wire  _T_2177; // @[MemPrimitives.scala 110:210:@10611.4]
  wire  _T_2181; // @[MemPrimitives.scala 123:41:@10625.4]
  wire  _T_2182; // @[MemPrimitives.scala 123:41:@10626.4]
  wire  _T_2183; // @[MemPrimitives.scala 123:41:@10627.4]
  wire  _T_2184; // @[MemPrimitives.scala 123:41:@10628.4]
  wire  _T_2185; // @[MemPrimitives.scala 123:41:@10629.4]
  wire  _T_2186; // @[MemPrimitives.scala 123:41:@10630.4]
  wire  _T_2187; // @[MemPrimitives.scala 123:41:@10631.4]
  wire  _T_2188; // @[MemPrimitives.scala 123:41:@10632.4]
  wire [2:0] _T_2190; // @[Cat.scala 30:58:@10634.4]
  wire [2:0] _T_2192; // @[Cat.scala 30:58:@10636.4]
  wire [2:0] _T_2194; // @[Cat.scala 30:58:@10638.4]
  wire [2:0] _T_2196; // @[Cat.scala 30:58:@10640.4]
  wire [2:0] _T_2198; // @[Cat.scala 30:58:@10642.4]
  wire [2:0] _T_2200; // @[Cat.scala 30:58:@10644.4]
  wire [2:0] _T_2202; // @[Cat.scala 30:58:@10646.4]
  wire [2:0] _T_2204; // @[Cat.scala 30:58:@10648.4]
  wire [2:0] _T_2205; // @[Mux.scala 31:69:@10649.4]
  wire [2:0] _T_2206; // @[Mux.scala 31:69:@10650.4]
  wire [2:0] _T_2207; // @[Mux.scala 31:69:@10651.4]
  wire [2:0] _T_2208; // @[Mux.scala 31:69:@10652.4]
  wire [2:0] _T_2209; // @[Mux.scala 31:69:@10653.4]
  wire [2:0] _T_2210; // @[Mux.scala 31:69:@10654.4]
  wire [2:0] _T_2211; // @[Mux.scala 31:69:@10655.4]
  wire  _T_2243; // @[package.scala 96:25:@10696.4 package.scala 96:25:@10697.4]
  wire [7:0] _T_2247; // @[Mux.scala 31:69:@10706.4]
  wire  _T_2240; // @[package.scala 96:25:@10688.4 package.scala 96:25:@10689.4]
  wire [7:0] _T_2248; // @[Mux.scala 31:69:@10707.4]
  wire  _T_2237; // @[package.scala 96:25:@10680.4 package.scala 96:25:@10681.4]
  wire  _T_2278; // @[package.scala 96:25:@10744.4 package.scala 96:25:@10745.4]
  wire [7:0] _T_2282; // @[Mux.scala 31:69:@10754.4]
  wire  _T_2275; // @[package.scala 96:25:@10736.4 package.scala 96:25:@10737.4]
  wire [7:0] _T_2283; // @[Mux.scala 31:69:@10755.4]
  wire  _T_2272; // @[package.scala 96:25:@10728.4 package.scala 96:25:@10729.4]
  wire  _T_2313; // @[package.scala 96:25:@10792.4 package.scala 96:25:@10793.4]
  wire [7:0] _T_2317; // @[Mux.scala 31:69:@10802.4]
  wire  _T_2310; // @[package.scala 96:25:@10784.4 package.scala 96:25:@10785.4]
  wire [7:0] _T_2318; // @[Mux.scala 31:69:@10803.4]
  wire  _T_2307; // @[package.scala 96:25:@10776.4 package.scala 96:25:@10777.4]
  wire  _T_2348; // @[package.scala 96:25:@10840.4 package.scala 96:25:@10841.4]
  wire [7:0] _T_2352; // @[Mux.scala 31:69:@10850.4]
  wire  _T_2345; // @[package.scala 96:25:@10832.4 package.scala 96:25:@10833.4]
  wire [7:0] _T_2353; // @[Mux.scala 31:69:@10851.4]
  wire  _T_2342; // @[package.scala 96:25:@10824.4 package.scala 96:25:@10825.4]
  wire  _T_2383; // @[package.scala 96:25:@10888.4 package.scala 96:25:@10889.4]
  wire [7:0] _T_2387; // @[Mux.scala 31:69:@10898.4]
  wire  _T_2380; // @[package.scala 96:25:@10880.4 package.scala 96:25:@10881.4]
  wire [7:0] _T_2388; // @[Mux.scala 31:69:@10899.4]
  wire  _T_2377; // @[package.scala 96:25:@10872.4 package.scala 96:25:@10873.4]
  wire  _T_2418; // @[package.scala 96:25:@10936.4 package.scala 96:25:@10937.4]
  wire [7:0] _T_2422; // @[Mux.scala 31:69:@10946.4]
  wire  _T_2415; // @[package.scala 96:25:@10928.4 package.scala 96:25:@10929.4]
  wire [7:0] _T_2423; // @[Mux.scala 31:69:@10947.4]
  wire  _T_2412; // @[package.scala 96:25:@10920.4 package.scala 96:25:@10921.4]
  wire  _T_2453; // @[package.scala 96:25:@10984.4 package.scala 96:25:@10985.4]
  wire [7:0] _T_2457; // @[Mux.scala 31:69:@10994.4]
  wire  _T_2450; // @[package.scala 96:25:@10976.4 package.scala 96:25:@10977.4]
  wire [7:0] _T_2458; // @[Mux.scala 31:69:@10995.4]
  wire  _T_2447; // @[package.scala 96:25:@10968.4 package.scala 96:25:@10969.4]
  wire  _T_2488; // @[package.scala 96:25:@11032.4 package.scala 96:25:@11033.4]
  wire [7:0] _T_2492; // @[Mux.scala 31:69:@11042.4]
  wire  _T_2485; // @[package.scala 96:25:@11024.4 package.scala 96:25:@11025.4]
  wire [7:0] _T_2493; // @[Mux.scala 31:69:@11043.4]
  wire  _T_2482; // @[package.scala 96:25:@11016.4 package.scala 96:25:@11017.4]
  wire  _T_2523; // @[package.scala 96:25:@11080.4 package.scala 96:25:@11081.4]
  wire [7:0] _T_2527; // @[Mux.scala 31:69:@11090.4]
  wire  _T_2520; // @[package.scala 96:25:@11072.4 package.scala 96:25:@11073.4]
  wire [7:0] _T_2528; // @[Mux.scala 31:69:@11091.4]
  wire  _T_2517; // @[package.scala 96:25:@11064.4 package.scala 96:25:@11065.4]
  wire  _T_2558; // @[package.scala 96:25:@11128.4 package.scala 96:25:@11129.4]
  wire [7:0] _T_2562; // @[Mux.scala 31:69:@11138.4]
  wire  _T_2555; // @[package.scala 96:25:@11120.4 package.scala 96:25:@11121.4]
  wire [7:0] _T_2563; // @[Mux.scala 31:69:@11139.4]
  wire  _T_2552; // @[package.scala 96:25:@11112.4 package.scala 96:25:@11113.4]
  wire  _T_2593; // @[package.scala 96:25:@11176.4 package.scala 96:25:@11177.4]
  wire [7:0] _T_2597; // @[Mux.scala 31:69:@11186.4]
  wire  _T_2590; // @[package.scala 96:25:@11168.4 package.scala 96:25:@11169.4]
  wire [7:0] _T_2598; // @[Mux.scala 31:69:@11187.4]
  wire  _T_2587; // @[package.scala 96:25:@11160.4 package.scala 96:25:@11161.4]
  wire  _T_2628; // @[package.scala 96:25:@11224.4 package.scala 96:25:@11225.4]
  wire [7:0] _T_2632; // @[Mux.scala 31:69:@11234.4]
  wire  _T_2625; // @[package.scala 96:25:@11216.4 package.scala 96:25:@11217.4]
  wire [7:0] _T_2633; // @[Mux.scala 31:69:@11235.4]
  wire  _T_2622; // @[package.scala 96:25:@11208.4 package.scala 96:25:@11209.4]
  wire  _T_2663; // @[package.scala 96:25:@11272.4 package.scala 96:25:@11273.4]
  wire [7:0] _T_2667; // @[Mux.scala 31:69:@11282.4]
  wire  _T_2660; // @[package.scala 96:25:@11264.4 package.scala 96:25:@11265.4]
  wire [7:0] _T_2668; // @[Mux.scala 31:69:@11283.4]
  wire  _T_2657; // @[package.scala 96:25:@11256.4 package.scala 96:25:@11257.4]
  wire  _T_2698; // @[package.scala 96:25:@11320.4 package.scala 96:25:@11321.4]
  wire [7:0] _T_2702; // @[Mux.scala 31:69:@11330.4]
  wire  _T_2695; // @[package.scala 96:25:@11312.4 package.scala 96:25:@11313.4]
  wire [7:0] _T_2703; // @[Mux.scala 31:69:@11331.4]
  wire  _T_2692; // @[package.scala 96:25:@11304.4 package.scala 96:25:@11305.4]
  wire  _T_2733; // @[package.scala 96:25:@11368.4 package.scala 96:25:@11369.4]
  wire [7:0] _T_2737; // @[Mux.scala 31:69:@11378.4]
  wire  _T_2730; // @[package.scala 96:25:@11360.4 package.scala 96:25:@11361.4]
  wire [7:0] _T_2738; // @[Mux.scala 31:69:@11379.4]
  wire  _T_2727; // @[package.scala 96:25:@11352.4 package.scala 96:25:@11353.4]
  wire  _T_2768; // @[package.scala 96:25:@11416.4 package.scala 96:25:@11417.4]
  wire [7:0] _T_2772; // @[Mux.scala 31:69:@11426.4]
  wire  _T_2765; // @[package.scala 96:25:@11408.4 package.scala 96:25:@11409.4]
  wire [7:0] _T_2773; // @[Mux.scala 31:69:@11427.4]
  wire  _T_2762; // @[package.scala 96:25:@11400.4 package.scala 96:25:@11401.4]
  wire  _T_2803; // @[package.scala 96:25:@11464.4 package.scala 96:25:@11465.4]
  wire [7:0] _T_2807; // @[Mux.scala 31:69:@11474.4]
  wire  _T_2800; // @[package.scala 96:25:@11456.4 package.scala 96:25:@11457.4]
  wire [7:0] _T_2808; // @[Mux.scala 31:69:@11475.4]
  wire  _T_2797; // @[package.scala 96:25:@11448.4 package.scala 96:25:@11449.4]
  wire  _T_2838; // @[package.scala 96:25:@11512.4 package.scala 96:25:@11513.4]
  wire [7:0] _T_2842; // @[Mux.scala 31:69:@11522.4]
  wire  _T_2835; // @[package.scala 96:25:@11504.4 package.scala 96:25:@11505.4]
  wire [7:0] _T_2843; // @[Mux.scala 31:69:@11523.4]
  wire  _T_2832; // @[package.scala 96:25:@11496.4 package.scala 96:25:@11497.4]
  wire  _T_2873; // @[package.scala 96:25:@11560.4 package.scala 96:25:@11561.4]
  wire [7:0] _T_2877; // @[Mux.scala 31:69:@11570.4]
  wire  _T_2870; // @[package.scala 96:25:@11552.4 package.scala 96:25:@11553.4]
  wire [7:0] _T_2878; // @[Mux.scala 31:69:@11571.4]
  wire  _T_2867; // @[package.scala 96:25:@11544.4 package.scala 96:25:@11545.4]
  wire  _T_2908; // @[package.scala 96:25:@11608.4 package.scala 96:25:@11609.4]
  wire [7:0] _T_2912; // @[Mux.scala 31:69:@11618.4]
  wire  _T_2905; // @[package.scala 96:25:@11600.4 package.scala 96:25:@11601.4]
  wire [7:0] _T_2913; // @[Mux.scala 31:69:@11619.4]
  wire  _T_2902; // @[package.scala 96:25:@11592.4 package.scala 96:25:@11593.4]
  wire  _T_2943; // @[package.scala 96:25:@11656.4 package.scala 96:25:@11657.4]
  wire [7:0] _T_2947; // @[Mux.scala 31:69:@11666.4]
  wire  _T_2940; // @[package.scala 96:25:@11648.4 package.scala 96:25:@11649.4]
  wire [7:0] _T_2948; // @[Mux.scala 31:69:@11667.4]
  wire  _T_2937; // @[package.scala 96:25:@11640.4 package.scala 96:25:@11641.4]
  wire  _T_2978; // @[package.scala 96:25:@11704.4 package.scala 96:25:@11705.4]
  wire [7:0] _T_2982; // @[Mux.scala 31:69:@11714.4]
  wire  _T_2975; // @[package.scala 96:25:@11696.4 package.scala 96:25:@11697.4]
  wire [7:0] _T_2983; // @[Mux.scala 31:69:@11715.4]
  wire  _T_2972; // @[package.scala 96:25:@11688.4 package.scala 96:25:@11689.4]
  wire  _T_3013; // @[package.scala 96:25:@11752.4 package.scala 96:25:@11753.4]
  wire [7:0] _T_3017; // @[Mux.scala 31:69:@11762.4]
  wire  _T_3010; // @[package.scala 96:25:@11744.4 package.scala 96:25:@11745.4]
  wire [7:0] _T_3018; // @[Mux.scala 31:69:@11763.4]
  wire  _T_3007; // @[package.scala 96:25:@11736.4 package.scala 96:25:@11737.4]
  wire  _T_3048; // @[package.scala 96:25:@11800.4 package.scala 96:25:@11801.4]
  wire [7:0] _T_3052; // @[Mux.scala 31:69:@11810.4]
  wire  _T_3045; // @[package.scala 96:25:@11792.4 package.scala 96:25:@11793.4]
  wire [7:0] _T_3053; // @[Mux.scala 31:69:@11811.4]
  wire  _T_3042; // @[package.scala 96:25:@11784.4 package.scala 96:25:@11785.4]
  Mem1D_4 Mem1D ( // @[MemPrimitives.scala 64:21:@9238.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  Mem1D_4 Mem1D_1 ( // @[MemPrimitives.scala 64:21:@9254.4]
    .clock(Mem1D_1_clock),
    .reset(Mem1D_1_reset),
    .io_r_ofs_0(Mem1D_1_io_r_ofs_0),
    .io_r_backpressure(Mem1D_1_io_r_backpressure),
    .io_w_ofs_0(Mem1D_1_io_w_ofs_0),
    .io_w_data_0(Mem1D_1_io_w_data_0),
    .io_w_en_0(Mem1D_1_io_w_en_0),
    .io_output(Mem1D_1_io_output)
  );
  Mem1D_4 Mem1D_2 ( // @[MemPrimitives.scala 64:21:@9270.4]
    .clock(Mem1D_2_clock),
    .reset(Mem1D_2_reset),
    .io_r_ofs_0(Mem1D_2_io_r_ofs_0),
    .io_r_backpressure(Mem1D_2_io_r_backpressure),
    .io_w_ofs_0(Mem1D_2_io_w_ofs_0),
    .io_w_data_0(Mem1D_2_io_w_data_0),
    .io_w_en_0(Mem1D_2_io_w_en_0),
    .io_output(Mem1D_2_io_output)
  );
  Mem1D_4 Mem1D_3 ( // @[MemPrimitives.scala 64:21:@9286.4]
    .clock(Mem1D_3_clock),
    .reset(Mem1D_3_reset),
    .io_r_ofs_0(Mem1D_3_io_r_ofs_0),
    .io_r_backpressure(Mem1D_3_io_r_backpressure),
    .io_w_ofs_0(Mem1D_3_io_w_ofs_0),
    .io_w_data_0(Mem1D_3_io_w_data_0),
    .io_w_en_0(Mem1D_3_io_w_en_0),
    .io_output(Mem1D_3_io_output)
  );
  Mem1D_4 Mem1D_4 ( // @[MemPrimitives.scala 64:21:@9302.4]
    .clock(Mem1D_4_clock),
    .reset(Mem1D_4_reset),
    .io_r_ofs_0(Mem1D_4_io_r_ofs_0),
    .io_r_backpressure(Mem1D_4_io_r_backpressure),
    .io_w_ofs_0(Mem1D_4_io_w_ofs_0),
    .io_w_data_0(Mem1D_4_io_w_data_0),
    .io_w_en_0(Mem1D_4_io_w_en_0),
    .io_output(Mem1D_4_io_output)
  );
  Mem1D_4 Mem1D_5 ( // @[MemPrimitives.scala 64:21:@9318.4]
    .clock(Mem1D_5_clock),
    .reset(Mem1D_5_reset),
    .io_r_ofs_0(Mem1D_5_io_r_ofs_0),
    .io_r_backpressure(Mem1D_5_io_r_backpressure),
    .io_w_ofs_0(Mem1D_5_io_w_ofs_0),
    .io_w_data_0(Mem1D_5_io_w_data_0),
    .io_w_en_0(Mem1D_5_io_w_en_0),
    .io_output(Mem1D_5_io_output)
  );
  Mem1D_4 Mem1D_6 ( // @[MemPrimitives.scala 64:21:@9334.4]
    .clock(Mem1D_6_clock),
    .reset(Mem1D_6_reset),
    .io_r_ofs_0(Mem1D_6_io_r_ofs_0),
    .io_r_backpressure(Mem1D_6_io_r_backpressure),
    .io_w_ofs_0(Mem1D_6_io_w_ofs_0),
    .io_w_data_0(Mem1D_6_io_w_data_0),
    .io_w_en_0(Mem1D_6_io_w_en_0),
    .io_output(Mem1D_6_io_output)
  );
  Mem1D_4 Mem1D_7 ( // @[MemPrimitives.scala 64:21:@9350.4]
    .clock(Mem1D_7_clock),
    .reset(Mem1D_7_reset),
    .io_r_ofs_0(Mem1D_7_io_r_ofs_0),
    .io_r_backpressure(Mem1D_7_io_r_backpressure),
    .io_w_ofs_0(Mem1D_7_io_w_ofs_0),
    .io_w_data_0(Mem1D_7_io_w_data_0),
    .io_w_en_0(Mem1D_7_io_w_en_0),
    .io_output(Mem1D_7_io_output)
  );
  Mem1D_4 Mem1D_8 ( // @[MemPrimitives.scala 64:21:@9366.4]
    .clock(Mem1D_8_clock),
    .reset(Mem1D_8_reset),
    .io_r_ofs_0(Mem1D_8_io_r_ofs_0),
    .io_r_backpressure(Mem1D_8_io_r_backpressure),
    .io_w_ofs_0(Mem1D_8_io_w_ofs_0),
    .io_w_data_0(Mem1D_8_io_w_data_0),
    .io_w_en_0(Mem1D_8_io_w_en_0),
    .io_output(Mem1D_8_io_output)
  );
  Mem1D_4 Mem1D_9 ( // @[MemPrimitives.scala 64:21:@9382.4]
    .clock(Mem1D_9_clock),
    .reset(Mem1D_9_reset),
    .io_r_ofs_0(Mem1D_9_io_r_ofs_0),
    .io_r_backpressure(Mem1D_9_io_r_backpressure),
    .io_w_ofs_0(Mem1D_9_io_w_ofs_0),
    .io_w_data_0(Mem1D_9_io_w_data_0),
    .io_w_en_0(Mem1D_9_io_w_en_0),
    .io_output(Mem1D_9_io_output)
  );
  Mem1D_4 Mem1D_10 ( // @[MemPrimitives.scala 64:21:@9398.4]
    .clock(Mem1D_10_clock),
    .reset(Mem1D_10_reset),
    .io_r_ofs_0(Mem1D_10_io_r_ofs_0),
    .io_r_backpressure(Mem1D_10_io_r_backpressure),
    .io_w_ofs_0(Mem1D_10_io_w_ofs_0),
    .io_w_data_0(Mem1D_10_io_w_data_0),
    .io_w_en_0(Mem1D_10_io_w_en_0),
    .io_output(Mem1D_10_io_output)
  );
  Mem1D_4 Mem1D_11 ( // @[MemPrimitives.scala 64:21:@9414.4]
    .clock(Mem1D_11_clock),
    .reset(Mem1D_11_reset),
    .io_r_ofs_0(Mem1D_11_io_r_ofs_0),
    .io_r_backpressure(Mem1D_11_io_r_backpressure),
    .io_w_ofs_0(Mem1D_11_io_w_ofs_0),
    .io_w_data_0(Mem1D_11_io_w_data_0),
    .io_w_en_0(Mem1D_11_io_w_en_0),
    .io_output(Mem1D_11_io_output)
  );
  Mem1D_4 Mem1D_12 ( // @[MemPrimitives.scala 64:21:@9430.4]
    .clock(Mem1D_12_clock),
    .reset(Mem1D_12_reset),
    .io_r_ofs_0(Mem1D_12_io_r_ofs_0),
    .io_r_backpressure(Mem1D_12_io_r_backpressure),
    .io_w_ofs_0(Mem1D_12_io_w_ofs_0),
    .io_w_data_0(Mem1D_12_io_w_data_0),
    .io_w_en_0(Mem1D_12_io_w_en_0),
    .io_output(Mem1D_12_io_output)
  );
  Mem1D_4 Mem1D_13 ( // @[MemPrimitives.scala 64:21:@9446.4]
    .clock(Mem1D_13_clock),
    .reset(Mem1D_13_reset),
    .io_r_ofs_0(Mem1D_13_io_r_ofs_0),
    .io_r_backpressure(Mem1D_13_io_r_backpressure),
    .io_w_ofs_0(Mem1D_13_io_w_ofs_0),
    .io_w_data_0(Mem1D_13_io_w_data_0),
    .io_w_en_0(Mem1D_13_io_w_en_0),
    .io_output(Mem1D_13_io_output)
  );
  Mem1D_4 Mem1D_14 ( // @[MemPrimitives.scala 64:21:@9462.4]
    .clock(Mem1D_14_clock),
    .reset(Mem1D_14_reset),
    .io_r_ofs_0(Mem1D_14_io_r_ofs_0),
    .io_r_backpressure(Mem1D_14_io_r_backpressure),
    .io_w_ofs_0(Mem1D_14_io_w_ofs_0),
    .io_w_data_0(Mem1D_14_io_w_data_0),
    .io_w_en_0(Mem1D_14_io_w_en_0),
    .io_output(Mem1D_14_io_output)
  );
  Mem1D_4 Mem1D_15 ( // @[MemPrimitives.scala 64:21:@9478.4]
    .clock(Mem1D_15_clock),
    .reset(Mem1D_15_reset),
    .io_r_ofs_0(Mem1D_15_io_r_ofs_0),
    .io_r_backpressure(Mem1D_15_io_r_backpressure),
    .io_w_ofs_0(Mem1D_15_io_w_ofs_0),
    .io_w_data_0(Mem1D_15_io_w_data_0),
    .io_w_en_0(Mem1D_15_io_w_en_0),
    .io_output(Mem1D_15_io_output)
  );
  StickySelects StickySelects ( // @[MemPrimitives.scala 121:29:@9778.4]
    .clock(StickySelects_clock),
    .reset(StickySelects_reset),
    .io_ins_0(StickySelects_io_ins_0),
    .io_ins_1(StickySelects_io_ins_1),
    .io_ins_2(StickySelects_io_ins_2),
    .io_ins_3(StickySelects_io_ins_3),
    .io_outs_0(StickySelects_io_outs_0),
    .io_outs_1(StickySelects_io_outs_1),
    .io_outs_2(StickySelects_io_outs_2),
    .io_outs_3(StickySelects_io_outs_3)
  );
  StickySelects StickySelects_1 ( // @[MemPrimitives.scala 121:29:@9818.4]
    .clock(StickySelects_1_clock),
    .reset(StickySelects_1_reset),
    .io_ins_0(StickySelects_1_io_ins_0),
    .io_ins_1(StickySelects_1_io_ins_1),
    .io_ins_2(StickySelects_1_io_ins_2),
    .io_ins_3(StickySelects_1_io_ins_3),
    .io_outs_0(StickySelects_1_io_outs_0),
    .io_outs_1(StickySelects_1_io_outs_1),
    .io_outs_2(StickySelects_1_io_outs_2),
    .io_outs_3(StickySelects_1_io_outs_3)
  );
  StickySelects_2 StickySelects_2 ( // @[MemPrimitives.scala 121:29:@9870.4]
    .clock(StickySelects_2_clock),
    .reset(StickySelects_2_reset),
    .io_ins_0(StickySelects_2_io_ins_0),
    .io_ins_1(StickySelects_2_io_ins_1),
    .io_ins_2(StickySelects_2_io_ins_2),
    .io_ins_3(StickySelects_2_io_ins_3),
    .io_ins_4(StickySelects_2_io_ins_4),
    .io_ins_5(StickySelects_2_io_ins_5),
    .io_ins_6(StickySelects_2_io_ins_6),
    .io_ins_7(StickySelects_2_io_ins_7),
    .io_outs_0(StickySelects_2_io_outs_0),
    .io_outs_1(StickySelects_2_io_outs_1),
    .io_outs_2(StickySelects_2_io_outs_2),
    .io_outs_3(StickySelects_2_io_outs_3),
    .io_outs_4(StickySelects_2_io_outs_4),
    .io_outs_5(StickySelects_2_io_outs_5),
    .io_outs_6(StickySelects_2_io_outs_6),
    .io_outs_7(StickySelects_2_io_outs_7)
  );
  StickySelects_2 StickySelects_3 ( // @[MemPrimitives.scala 121:29:@9942.4]
    .clock(StickySelects_3_clock),
    .reset(StickySelects_3_reset),
    .io_ins_0(StickySelects_3_io_ins_0),
    .io_ins_1(StickySelects_3_io_ins_1),
    .io_ins_2(StickySelects_3_io_ins_2),
    .io_ins_3(StickySelects_3_io_ins_3),
    .io_ins_4(StickySelects_3_io_ins_4),
    .io_ins_5(StickySelects_3_io_ins_5),
    .io_ins_6(StickySelects_3_io_ins_6),
    .io_ins_7(StickySelects_3_io_ins_7),
    .io_outs_0(StickySelects_3_io_outs_0),
    .io_outs_1(StickySelects_3_io_outs_1),
    .io_outs_2(StickySelects_3_io_outs_2),
    .io_outs_3(StickySelects_3_io_outs_3),
    .io_outs_4(StickySelects_3_io_outs_4),
    .io_outs_5(StickySelects_3_io_outs_5),
    .io_outs_6(StickySelects_3_io_outs_6),
    .io_outs_7(StickySelects_3_io_outs_7)
  );
  StickySelects StickySelects_4 ( // @[MemPrimitives.scala 121:29:@10002.4]
    .clock(StickySelects_4_clock),
    .reset(StickySelects_4_reset),
    .io_ins_0(StickySelects_4_io_ins_0),
    .io_ins_1(StickySelects_4_io_ins_1),
    .io_ins_2(StickySelects_4_io_ins_2),
    .io_ins_3(StickySelects_4_io_ins_3),
    .io_outs_0(StickySelects_4_io_outs_0),
    .io_outs_1(StickySelects_4_io_outs_1),
    .io_outs_2(StickySelects_4_io_outs_2),
    .io_outs_3(StickySelects_4_io_outs_3)
  );
  StickySelects StickySelects_5 ( // @[MemPrimitives.scala 121:29:@10042.4]
    .clock(StickySelects_5_clock),
    .reset(StickySelects_5_reset),
    .io_ins_0(StickySelects_5_io_ins_0),
    .io_ins_1(StickySelects_5_io_ins_1),
    .io_ins_2(StickySelects_5_io_ins_2),
    .io_ins_3(StickySelects_5_io_ins_3),
    .io_outs_0(StickySelects_5_io_outs_0),
    .io_outs_1(StickySelects_5_io_outs_1),
    .io_outs_2(StickySelects_5_io_outs_2),
    .io_outs_3(StickySelects_5_io_outs_3)
  );
  StickySelects_2 StickySelects_6 ( // @[MemPrimitives.scala 121:29:@10094.4]
    .clock(StickySelects_6_clock),
    .reset(StickySelects_6_reset),
    .io_ins_0(StickySelects_6_io_ins_0),
    .io_ins_1(StickySelects_6_io_ins_1),
    .io_ins_2(StickySelects_6_io_ins_2),
    .io_ins_3(StickySelects_6_io_ins_3),
    .io_ins_4(StickySelects_6_io_ins_4),
    .io_ins_5(StickySelects_6_io_ins_5),
    .io_ins_6(StickySelects_6_io_ins_6),
    .io_ins_7(StickySelects_6_io_ins_7),
    .io_outs_0(StickySelects_6_io_outs_0),
    .io_outs_1(StickySelects_6_io_outs_1),
    .io_outs_2(StickySelects_6_io_outs_2),
    .io_outs_3(StickySelects_6_io_outs_3),
    .io_outs_4(StickySelects_6_io_outs_4),
    .io_outs_5(StickySelects_6_io_outs_5),
    .io_outs_6(StickySelects_6_io_outs_6),
    .io_outs_7(StickySelects_6_io_outs_7)
  );
  StickySelects_2 StickySelects_7 ( // @[MemPrimitives.scala 121:29:@10166.4]
    .clock(StickySelects_7_clock),
    .reset(StickySelects_7_reset),
    .io_ins_0(StickySelects_7_io_ins_0),
    .io_ins_1(StickySelects_7_io_ins_1),
    .io_ins_2(StickySelects_7_io_ins_2),
    .io_ins_3(StickySelects_7_io_ins_3),
    .io_ins_4(StickySelects_7_io_ins_4),
    .io_ins_5(StickySelects_7_io_ins_5),
    .io_ins_6(StickySelects_7_io_ins_6),
    .io_ins_7(StickySelects_7_io_ins_7),
    .io_outs_0(StickySelects_7_io_outs_0),
    .io_outs_1(StickySelects_7_io_outs_1),
    .io_outs_2(StickySelects_7_io_outs_2),
    .io_outs_3(StickySelects_7_io_outs_3),
    .io_outs_4(StickySelects_7_io_outs_4),
    .io_outs_5(StickySelects_7_io_outs_5),
    .io_outs_6(StickySelects_7_io_outs_6),
    .io_outs_7(StickySelects_7_io_outs_7)
  );
  StickySelects StickySelects_8 ( // @[MemPrimitives.scala 121:29:@10226.4]
    .clock(StickySelects_8_clock),
    .reset(StickySelects_8_reset),
    .io_ins_0(StickySelects_8_io_ins_0),
    .io_ins_1(StickySelects_8_io_ins_1),
    .io_ins_2(StickySelects_8_io_ins_2),
    .io_ins_3(StickySelects_8_io_ins_3),
    .io_outs_0(StickySelects_8_io_outs_0),
    .io_outs_1(StickySelects_8_io_outs_1),
    .io_outs_2(StickySelects_8_io_outs_2),
    .io_outs_3(StickySelects_8_io_outs_3)
  );
  StickySelects StickySelects_9 ( // @[MemPrimitives.scala 121:29:@10266.4]
    .clock(StickySelects_9_clock),
    .reset(StickySelects_9_reset),
    .io_ins_0(StickySelects_9_io_ins_0),
    .io_ins_1(StickySelects_9_io_ins_1),
    .io_ins_2(StickySelects_9_io_ins_2),
    .io_ins_3(StickySelects_9_io_ins_3),
    .io_outs_0(StickySelects_9_io_outs_0),
    .io_outs_1(StickySelects_9_io_outs_1),
    .io_outs_2(StickySelects_9_io_outs_2),
    .io_outs_3(StickySelects_9_io_outs_3)
  );
  StickySelects_2 StickySelects_10 ( // @[MemPrimitives.scala 121:29:@10318.4]
    .clock(StickySelects_10_clock),
    .reset(StickySelects_10_reset),
    .io_ins_0(StickySelects_10_io_ins_0),
    .io_ins_1(StickySelects_10_io_ins_1),
    .io_ins_2(StickySelects_10_io_ins_2),
    .io_ins_3(StickySelects_10_io_ins_3),
    .io_ins_4(StickySelects_10_io_ins_4),
    .io_ins_5(StickySelects_10_io_ins_5),
    .io_ins_6(StickySelects_10_io_ins_6),
    .io_ins_7(StickySelects_10_io_ins_7),
    .io_outs_0(StickySelects_10_io_outs_0),
    .io_outs_1(StickySelects_10_io_outs_1),
    .io_outs_2(StickySelects_10_io_outs_2),
    .io_outs_3(StickySelects_10_io_outs_3),
    .io_outs_4(StickySelects_10_io_outs_4),
    .io_outs_5(StickySelects_10_io_outs_5),
    .io_outs_6(StickySelects_10_io_outs_6),
    .io_outs_7(StickySelects_10_io_outs_7)
  );
  StickySelects_2 StickySelects_11 ( // @[MemPrimitives.scala 121:29:@10390.4]
    .clock(StickySelects_11_clock),
    .reset(StickySelects_11_reset),
    .io_ins_0(StickySelects_11_io_ins_0),
    .io_ins_1(StickySelects_11_io_ins_1),
    .io_ins_2(StickySelects_11_io_ins_2),
    .io_ins_3(StickySelects_11_io_ins_3),
    .io_ins_4(StickySelects_11_io_ins_4),
    .io_ins_5(StickySelects_11_io_ins_5),
    .io_ins_6(StickySelects_11_io_ins_6),
    .io_ins_7(StickySelects_11_io_ins_7),
    .io_outs_0(StickySelects_11_io_outs_0),
    .io_outs_1(StickySelects_11_io_outs_1),
    .io_outs_2(StickySelects_11_io_outs_2),
    .io_outs_3(StickySelects_11_io_outs_3),
    .io_outs_4(StickySelects_11_io_outs_4),
    .io_outs_5(StickySelects_11_io_outs_5),
    .io_outs_6(StickySelects_11_io_outs_6),
    .io_outs_7(StickySelects_11_io_outs_7)
  );
  StickySelects StickySelects_12 ( // @[MemPrimitives.scala 121:29:@10450.4]
    .clock(StickySelects_12_clock),
    .reset(StickySelects_12_reset),
    .io_ins_0(StickySelects_12_io_ins_0),
    .io_ins_1(StickySelects_12_io_ins_1),
    .io_ins_2(StickySelects_12_io_ins_2),
    .io_ins_3(StickySelects_12_io_ins_3),
    .io_outs_0(StickySelects_12_io_outs_0),
    .io_outs_1(StickySelects_12_io_outs_1),
    .io_outs_2(StickySelects_12_io_outs_2),
    .io_outs_3(StickySelects_12_io_outs_3)
  );
  StickySelects StickySelects_13 ( // @[MemPrimitives.scala 121:29:@10490.4]
    .clock(StickySelects_13_clock),
    .reset(StickySelects_13_reset),
    .io_ins_0(StickySelects_13_io_ins_0),
    .io_ins_1(StickySelects_13_io_ins_1),
    .io_ins_2(StickySelects_13_io_ins_2),
    .io_ins_3(StickySelects_13_io_ins_3),
    .io_outs_0(StickySelects_13_io_outs_0),
    .io_outs_1(StickySelects_13_io_outs_1),
    .io_outs_2(StickySelects_13_io_outs_2),
    .io_outs_3(StickySelects_13_io_outs_3)
  );
  StickySelects_2 StickySelects_14 ( // @[MemPrimitives.scala 121:29:@10542.4]
    .clock(StickySelects_14_clock),
    .reset(StickySelects_14_reset),
    .io_ins_0(StickySelects_14_io_ins_0),
    .io_ins_1(StickySelects_14_io_ins_1),
    .io_ins_2(StickySelects_14_io_ins_2),
    .io_ins_3(StickySelects_14_io_ins_3),
    .io_ins_4(StickySelects_14_io_ins_4),
    .io_ins_5(StickySelects_14_io_ins_5),
    .io_ins_6(StickySelects_14_io_ins_6),
    .io_ins_7(StickySelects_14_io_ins_7),
    .io_outs_0(StickySelects_14_io_outs_0),
    .io_outs_1(StickySelects_14_io_outs_1),
    .io_outs_2(StickySelects_14_io_outs_2),
    .io_outs_3(StickySelects_14_io_outs_3),
    .io_outs_4(StickySelects_14_io_outs_4),
    .io_outs_5(StickySelects_14_io_outs_5),
    .io_outs_6(StickySelects_14_io_outs_6),
    .io_outs_7(StickySelects_14_io_outs_7)
  );
  StickySelects_2 StickySelects_15 ( // @[MemPrimitives.scala 121:29:@10614.4]
    .clock(StickySelects_15_clock),
    .reset(StickySelects_15_reset),
    .io_ins_0(StickySelects_15_io_ins_0),
    .io_ins_1(StickySelects_15_io_ins_1),
    .io_ins_2(StickySelects_15_io_ins_2),
    .io_ins_3(StickySelects_15_io_ins_3),
    .io_ins_4(StickySelects_15_io_ins_4),
    .io_ins_5(StickySelects_15_io_ins_5),
    .io_ins_6(StickySelects_15_io_ins_6),
    .io_ins_7(StickySelects_15_io_ins_7),
    .io_outs_0(StickySelects_15_io_outs_0),
    .io_outs_1(StickySelects_15_io_outs_1),
    .io_outs_2(StickySelects_15_io_outs_2),
    .io_outs_3(StickySelects_15_io_outs_3),
    .io_outs_4(StickySelects_15_io_outs_4),
    .io_outs_5(StickySelects_15_io_outs_5),
    .io_outs_6(StickySelects_15_io_outs_6),
    .io_outs_7(StickySelects_15_io_outs_7)
  );
  RetimeWrapper_52 RetimeWrapper ( // @[package.scala 93:22:@10675.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_1 ( // @[package.scala 93:22:@10683.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_2 ( // @[package.scala 93:22:@10691.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_3 ( // @[package.scala 93:22:@10699.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_4 ( // @[package.scala 93:22:@10723.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_5 ( // @[package.scala 93:22:@10731.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_6 ( // @[package.scala 93:22:@10739.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_7 ( // @[package.scala 93:22:@10747.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_8 ( // @[package.scala 93:22:@10771.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_9 ( // @[package.scala 93:22:@10779.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_10 ( // @[package.scala 93:22:@10787.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_11 ( // @[package.scala 93:22:@10795.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_12 ( // @[package.scala 93:22:@10819.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_13 ( // @[package.scala 93:22:@10827.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_14 ( // @[package.scala 93:22:@10835.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_15 ( // @[package.scala 93:22:@10843.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_16 ( // @[package.scala 93:22:@10867.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_17 ( // @[package.scala 93:22:@10875.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_18 ( // @[package.scala 93:22:@10883.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_19 ( // @[package.scala 93:22:@10891.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_20 ( // @[package.scala 93:22:@10915.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_21 ( // @[package.scala 93:22:@10923.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_22 ( // @[package.scala 93:22:@10931.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_23 ( // @[package.scala 93:22:@10939.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_24 ( // @[package.scala 93:22:@10963.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_25 ( // @[package.scala 93:22:@10971.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_26 ( // @[package.scala 93:22:@10979.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_27 ( // @[package.scala 93:22:@10987.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_28 ( // @[package.scala 93:22:@11011.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_29 ( // @[package.scala 93:22:@11019.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_30 ( // @[package.scala 93:22:@11027.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_31 ( // @[package.scala 93:22:@11035.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_32 ( // @[package.scala 93:22:@11059.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_33 ( // @[package.scala 93:22:@11067.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_34 ( // @[package.scala 93:22:@11075.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_35 ( // @[package.scala 93:22:@11083.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_36 ( // @[package.scala 93:22:@11107.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_37 ( // @[package.scala 93:22:@11115.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_38 ( // @[package.scala 93:22:@11123.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_39 ( // @[package.scala 93:22:@11131.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_40 ( // @[package.scala 93:22:@11155.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_41 ( // @[package.scala 93:22:@11163.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_42 ( // @[package.scala 93:22:@11171.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_43 ( // @[package.scala 93:22:@11179.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_44 ( // @[package.scala 93:22:@11203.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_45 ( // @[package.scala 93:22:@11211.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_46 ( // @[package.scala 93:22:@11219.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_47 ( // @[package.scala 93:22:@11227.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_48 ( // @[package.scala 93:22:@11251.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_49 ( // @[package.scala 93:22:@11259.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_50 ( // @[package.scala 93:22:@11267.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_51 ( // @[package.scala 93:22:@11275.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_52 ( // @[package.scala 93:22:@11299.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_53 ( // @[package.scala 93:22:@11307.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_54 ( // @[package.scala 93:22:@11315.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_55 ( // @[package.scala 93:22:@11323.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_56 ( // @[package.scala 93:22:@11347.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_57 ( // @[package.scala 93:22:@11355.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_58 ( // @[package.scala 93:22:@11363.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_59 ( // @[package.scala 93:22:@11371.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_60 ( // @[package.scala 93:22:@11395.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_61 ( // @[package.scala 93:22:@11403.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_62 ( // @[package.scala 93:22:@11411.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_63 ( // @[package.scala 93:22:@11419.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_64 ( // @[package.scala 93:22:@11443.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_65 ( // @[package.scala 93:22:@11451.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_66 ( // @[package.scala 93:22:@11459.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_67 ( // @[package.scala 93:22:@11467.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_68 ( // @[package.scala 93:22:@11491.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_69 ( // @[package.scala 93:22:@11499.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_70 ( // @[package.scala 93:22:@11507.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_71 ( // @[package.scala 93:22:@11515.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_72 ( // @[package.scala 93:22:@11539.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_73 ( // @[package.scala 93:22:@11547.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_74 ( // @[package.scala 93:22:@11555.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_75 ( // @[package.scala 93:22:@11563.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_76 ( // @[package.scala 93:22:@11587.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_77 ( // @[package.scala 93:22:@11595.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_78 ( // @[package.scala 93:22:@11603.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_79 ( // @[package.scala 93:22:@11611.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_80 ( // @[package.scala 93:22:@11635.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_81 ( // @[package.scala 93:22:@11643.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_82 ( // @[package.scala 93:22:@11651.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_83 ( // @[package.scala 93:22:@11659.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_84 ( // @[package.scala 93:22:@11683.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_85 ( // @[package.scala 93:22:@11691.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_86 ( // @[package.scala 93:22:@11699.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_87 ( // @[package.scala 93:22:@11707.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_88 ( // @[package.scala 93:22:@11731.4]
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_89 ( // @[package.scala 93:22:@11739.4]
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_90 ( // @[package.scala 93:22:@11747.4]
    .clock(RetimeWrapper_90_clock),
    .reset(RetimeWrapper_90_reset),
    .io_flow(RetimeWrapper_90_io_flow),
    .io_in(RetimeWrapper_90_io_in),
    .io_out(RetimeWrapper_90_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_91 ( // @[package.scala 93:22:@11755.4]
    .clock(RetimeWrapper_91_clock),
    .reset(RetimeWrapper_91_reset),
    .io_flow(RetimeWrapper_91_io_flow),
    .io_in(RetimeWrapper_91_io_in),
    .io_out(RetimeWrapper_91_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_92 ( // @[package.scala 93:22:@11779.4]
    .clock(RetimeWrapper_92_clock),
    .reset(RetimeWrapper_92_reset),
    .io_flow(RetimeWrapper_92_io_flow),
    .io_in(RetimeWrapper_92_io_in),
    .io_out(RetimeWrapper_92_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_93 ( // @[package.scala 93:22:@11787.4]
    .clock(RetimeWrapper_93_clock),
    .reset(RetimeWrapper_93_reset),
    .io_flow(RetimeWrapper_93_io_flow),
    .io_in(RetimeWrapper_93_io_in),
    .io_out(RetimeWrapper_93_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_94 ( // @[package.scala 93:22:@11795.4]
    .clock(RetimeWrapper_94_clock),
    .reset(RetimeWrapper_94_reset),
    .io_flow(RetimeWrapper_94_io_flow),
    .io_in(RetimeWrapper_94_io_in),
    .io_out(RetimeWrapper_94_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_95 ( // @[package.scala 93:22:@11803.4]
    .clock(RetimeWrapper_95_clock),
    .reset(RetimeWrapper_95_reset),
    .io_flow(RetimeWrapper_95_io_flow),
    .io_in(RetimeWrapper_95_io_in),
    .io_out(RetimeWrapper_95_io_out)
  );
  assign _T_1032 = io_wPort_4_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@9494.4]
  assign _T_1035 = io_wPort_4_en_0 & _T_1032; // @[MemPrimitives.scala 83:102:@9496.4]
  assign _T_1037 = io_wPort_7_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@9497.4]
  assign _T_1040 = io_wPort_7_en_0 & _T_1037; // @[MemPrimitives.scala 83:102:@9499.4]
  assign _T_1042 = {_T_1035,io_wPort_4_data_0,io_wPort_4_ofs_0}; // @[Cat.scala 30:58:@9501.4]
  assign _T_1044 = {_T_1040,io_wPort_7_data_0,io_wPort_7_ofs_0}; // @[Cat.scala 30:58:@9503.4]
  assign _T_1045 = _T_1035 ? _T_1042 : _T_1044; // @[Mux.scala 31:69:@9504.4]
  assign _T_1050 = io_wPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@9511.4]
  assign _T_1053 = io_wPort_0_en_0 & _T_1050; // @[MemPrimitives.scala 83:102:@9513.4]
  assign _T_1055 = io_wPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@9514.4]
  assign _T_1058 = io_wPort_3_en_0 & _T_1055; // @[MemPrimitives.scala 83:102:@9516.4]
  assign _T_1060 = {_T_1053,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9518.4]
  assign _T_1062 = {_T_1058,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@9520.4]
  assign _T_1063 = _T_1053 ? _T_1060 : _T_1062; // @[Mux.scala 31:69:@9521.4]
  assign _T_1068 = io_wPort_5_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@9528.4]
  assign _T_1071 = io_wPort_5_en_0 & _T_1068; // @[MemPrimitives.scala 83:102:@9530.4]
  assign _T_1073 = io_wPort_6_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@9531.4]
  assign _T_1076 = io_wPort_6_en_0 & _T_1073; // @[MemPrimitives.scala 83:102:@9533.4]
  assign _T_1078 = {_T_1071,io_wPort_5_data_0,io_wPort_5_ofs_0}; // @[Cat.scala 30:58:@9535.4]
  assign _T_1080 = {_T_1076,io_wPort_6_data_0,io_wPort_6_ofs_0}; // @[Cat.scala 30:58:@9537.4]
  assign _T_1081 = _T_1071 ? _T_1078 : _T_1080; // @[Mux.scala 31:69:@9538.4]
  assign _T_1086 = io_wPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@9545.4]
  assign _T_1089 = io_wPort_1_en_0 & _T_1086; // @[MemPrimitives.scala 83:102:@9547.4]
  assign _T_1091 = io_wPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@9548.4]
  assign _T_1094 = io_wPort_2_en_0 & _T_1091; // @[MemPrimitives.scala 83:102:@9550.4]
  assign _T_1096 = {_T_1089,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@9552.4]
  assign _T_1098 = {_T_1094,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@9554.4]
  assign _T_1099 = _T_1089 ? _T_1096 : _T_1098; // @[Mux.scala 31:69:@9555.4]
  assign _T_1104 = io_wPort_4_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@9562.4]
  assign _T_1107 = io_wPort_4_en_0 & _T_1104; // @[MemPrimitives.scala 83:102:@9564.4]
  assign _T_1109 = io_wPort_7_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@9565.4]
  assign _T_1112 = io_wPort_7_en_0 & _T_1109; // @[MemPrimitives.scala 83:102:@9567.4]
  assign _T_1114 = {_T_1107,io_wPort_4_data_0,io_wPort_4_ofs_0}; // @[Cat.scala 30:58:@9569.4]
  assign _T_1116 = {_T_1112,io_wPort_7_data_0,io_wPort_7_ofs_0}; // @[Cat.scala 30:58:@9571.4]
  assign _T_1117 = _T_1107 ? _T_1114 : _T_1116; // @[Mux.scala 31:69:@9572.4]
  assign _T_1122 = io_wPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@9579.4]
  assign _T_1125 = io_wPort_0_en_0 & _T_1122; // @[MemPrimitives.scala 83:102:@9581.4]
  assign _T_1127 = io_wPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@9582.4]
  assign _T_1130 = io_wPort_3_en_0 & _T_1127; // @[MemPrimitives.scala 83:102:@9584.4]
  assign _T_1132 = {_T_1125,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9586.4]
  assign _T_1134 = {_T_1130,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@9588.4]
  assign _T_1135 = _T_1125 ? _T_1132 : _T_1134; // @[Mux.scala 31:69:@9589.4]
  assign _T_1140 = io_wPort_5_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@9596.4]
  assign _T_1143 = io_wPort_5_en_0 & _T_1140; // @[MemPrimitives.scala 83:102:@9598.4]
  assign _T_1145 = io_wPort_6_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@9599.4]
  assign _T_1148 = io_wPort_6_en_0 & _T_1145; // @[MemPrimitives.scala 83:102:@9601.4]
  assign _T_1150 = {_T_1143,io_wPort_5_data_0,io_wPort_5_ofs_0}; // @[Cat.scala 30:58:@9603.4]
  assign _T_1152 = {_T_1148,io_wPort_6_data_0,io_wPort_6_ofs_0}; // @[Cat.scala 30:58:@9605.4]
  assign _T_1153 = _T_1143 ? _T_1150 : _T_1152; // @[Mux.scala 31:69:@9606.4]
  assign _T_1158 = io_wPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@9613.4]
  assign _T_1161 = io_wPort_1_en_0 & _T_1158; // @[MemPrimitives.scala 83:102:@9615.4]
  assign _T_1163 = io_wPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@9616.4]
  assign _T_1166 = io_wPort_2_en_0 & _T_1163; // @[MemPrimitives.scala 83:102:@9618.4]
  assign _T_1168 = {_T_1161,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@9620.4]
  assign _T_1170 = {_T_1166,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@9622.4]
  assign _T_1171 = _T_1161 ? _T_1168 : _T_1170; // @[Mux.scala 31:69:@9623.4]
  assign _T_1176 = io_wPort_4_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@9630.4]
  assign _T_1179 = io_wPort_4_en_0 & _T_1176; // @[MemPrimitives.scala 83:102:@9632.4]
  assign _T_1181 = io_wPort_7_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@9633.4]
  assign _T_1184 = io_wPort_7_en_0 & _T_1181; // @[MemPrimitives.scala 83:102:@9635.4]
  assign _T_1186 = {_T_1179,io_wPort_4_data_0,io_wPort_4_ofs_0}; // @[Cat.scala 30:58:@9637.4]
  assign _T_1188 = {_T_1184,io_wPort_7_data_0,io_wPort_7_ofs_0}; // @[Cat.scala 30:58:@9639.4]
  assign _T_1189 = _T_1179 ? _T_1186 : _T_1188; // @[Mux.scala 31:69:@9640.4]
  assign _T_1194 = io_wPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@9647.4]
  assign _T_1197 = io_wPort_0_en_0 & _T_1194; // @[MemPrimitives.scala 83:102:@9649.4]
  assign _T_1199 = io_wPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@9650.4]
  assign _T_1202 = io_wPort_3_en_0 & _T_1199; // @[MemPrimitives.scala 83:102:@9652.4]
  assign _T_1204 = {_T_1197,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9654.4]
  assign _T_1206 = {_T_1202,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@9656.4]
  assign _T_1207 = _T_1197 ? _T_1204 : _T_1206; // @[Mux.scala 31:69:@9657.4]
  assign _T_1212 = io_wPort_5_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@9664.4]
  assign _T_1215 = io_wPort_5_en_0 & _T_1212; // @[MemPrimitives.scala 83:102:@9666.4]
  assign _T_1217 = io_wPort_6_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@9667.4]
  assign _T_1220 = io_wPort_6_en_0 & _T_1217; // @[MemPrimitives.scala 83:102:@9669.4]
  assign _T_1222 = {_T_1215,io_wPort_5_data_0,io_wPort_5_ofs_0}; // @[Cat.scala 30:58:@9671.4]
  assign _T_1224 = {_T_1220,io_wPort_6_data_0,io_wPort_6_ofs_0}; // @[Cat.scala 30:58:@9673.4]
  assign _T_1225 = _T_1215 ? _T_1222 : _T_1224; // @[Mux.scala 31:69:@9674.4]
  assign _T_1230 = io_wPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@9681.4]
  assign _T_1233 = io_wPort_1_en_0 & _T_1230; // @[MemPrimitives.scala 83:102:@9683.4]
  assign _T_1235 = io_wPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@9684.4]
  assign _T_1238 = io_wPort_2_en_0 & _T_1235; // @[MemPrimitives.scala 83:102:@9686.4]
  assign _T_1240 = {_T_1233,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@9688.4]
  assign _T_1242 = {_T_1238,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@9690.4]
  assign _T_1243 = _T_1233 ? _T_1240 : _T_1242; // @[Mux.scala 31:69:@9691.4]
  assign _T_1248 = io_wPort_4_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@9698.4]
  assign _T_1251 = io_wPort_4_en_0 & _T_1248; // @[MemPrimitives.scala 83:102:@9700.4]
  assign _T_1253 = io_wPort_7_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@9701.4]
  assign _T_1256 = io_wPort_7_en_0 & _T_1253; // @[MemPrimitives.scala 83:102:@9703.4]
  assign _T_1258 = {_T_1251,io_wPort_4_data_0,io_wPort_4_ofs_0}; // @[Cat.scala 30:58:@9705.4]
  assign _T_1260 = {_T_1256,io_wPort_7_data_0,io_wPort_7_ofs_0}; // @[Cat.scala 30:58:@9707.4]
  assign _T_1261 = _T_1251 ? _T_1258 : _T_1260; // @[Mux.scala 31:69:@9708.4]
  assign _T_1266 = io_wPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@9715.4]
  assign _T_1269 = io_wPort_0_en_0 & _T_1266; // @[MemPrimitives.scala 83:102:@9717.4]
  assign _T_1271 = io_wPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@9718.4]
  assign _T_1274 = io_wPort_3_en_0 & _T_1271; // @[MemPrimitives.scala 83:102:@9720.4]
  assign _T_1276 = {_T_1269,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9722.4]
  assign _T_1278 = {_T_1274,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@9724.4]
  assign _T_1279 = _T_1269 ? _T_1276 : _T_1278; // @[Mux.scala 31:69:@9725.4]
  assign _T_1284 = io_wPort_5_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@9732.4]
  assign _T_1287 = io_wPort_5_en_0 & _T_1284; // @[MemPrimitives.scala 83:102:@9734.4]
  assign _T_1289 = io_wPort_6_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@9735.4]
  assign _T_1292 = io_wPort_6_en_0 & _T_1289; // @[MemPrimitives.scala 83:102:@9737.4]
  assign _T_1294 = {_T_1287,io_wPort_5_data_0,io_wPort_5_ofs_0}; // @[Cat.scala 30:58:@9739.4]
  assign _T_1296 = {_T_1292,io_wPort_6_data_0,io_wPort_6_ofs_0}; // @[Cat.scala 30:58:@9741.4]
  assign _T_1297 = _T_1287 ? _T_1294 : _T_1296; // @[Mux.scala 31:69:@9742.4]
  assign _T_1302 = io_wPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@9749.4]
  assign _T_1305 = io_wPort_1_en_0 & _T_1302; // @[MemPrimitives.scala 83:102:@9751.4]
  assign _T_1307 = io_wPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@9752.4]
  assign _T_1310 = io_wPort_2_en_0 & _T_1307; // @[MemPrimitives.scala 83:102:@9754.4]
  assign _T_1312 = {_T_1305,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@9756.4]
  assign _T_1314 = {_T_1310,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@9758.4]
  assign _T_1315 = _T_1305 ? _T_1312 : _T_1314; // @[Mux.scala 31:69:@9759.4]
  assign _T_1320 = io_rPort_4_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9766.4]
  assign _T_1325 = io_rPort_12_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9769.4]
  assign _T_1330 = io_rPort_16_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9772.4]
  assign _T_1335 = io_rPort_20_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9775.4]
  assign _T_1339 = StickySelects_io_outs_0; // @[MemPrimitives.scala 123:41:@9785.4]
  assign _T_1340 = StickySelects_io_outs_1; // @[MemPrimitives.scala 123:41:@9786.4]
  assign _T_1341 = StickySelects_io_outs_2; // @[MemPrimitives.scala 123:41:@9787.4]
  assign _T_1342 = StickySelects_io_outs_3; // @[MemPrimitives.scala 123:41:@9788.4]
  assign _T_1344 = {_T_1339,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@9790.4]
  assign _T_1346 = {_T_1340,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@9792.4]
  assign _T_1348 = {_T_1341,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@9794.4]
  assign _T_1350 = {_T_1342,io_rPort_20_backpressure,io_rPort_20_ofs_0}; // @[Cat.scala 30:58:@9796.4]
  assign _T_1351 = _T_1341 ? _T_1348 : _T_1350; // @[Mux.scala 31:69:@9797.4]
  assign _T_1352 = _T_1340 ? _T_1346 : _T_1351; // @[Mux.scala 31:69:@9798.4]
  assign _T_1353 = _T_1339 ? _T_1344 : _T_1352; // @[Mux.scala 31:69:@9799.4]
  assign _T_1358 = io_rPort_5_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9806.4]
  assign _T_1363 = io_rPort_10_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9809.4]
  assign _T_1368 = io_rPort_13_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9812.4]
  assign _T_1373 = io_rPort_23_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9815.4]
  assign _T_1377 = StickySelects_1_io_outs_0; // @[MemPrimitives.scala 123:41:@9825.4]
  assign _T_1378 = StickySelects_1_io_outs_1; // @[MemPrimitives.scala 123:41:@9826.4]
  assign _T_1379 = StickySelects_1_io_outs_2; // @[MemPrimitives.scala 123:41:@9827.4]
  assign _T_1380 = StickySelects_1_io_outs_3; // @[MemPrimitives.scala 123:41:@9828.4]
  assign _T_1382 = {_T_1377,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@9830.4]
  assign _T_1384 = {_T_1378,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@9832.4]
  assign _T_1386 = {_T_1379,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@9834.4]
  assign _T_1388 = {_T_1380,io_rPort_23_backpressure,io_rPort_23_ofs_0}; // @[Cat.scala 30:58:@9836.4]
  assign _T_1389 = _T_1379 ? _T_1386 : _T_1388; // @[Mux.scala 31:69:@9837.4]
  assign _T_1390 = _T_1378 ? _T_1384 : _T_1389; // @[Mux.scala 31:69:@9838.4]
  assign _T_1391 = _T_1377 ? _T_1382 : _T_1390; // @[Mux.scala 31:69:@9839.4]
  assign _T_1396 = io_rPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9846.4]
  assign _T_1401 = io_rPort_7_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9849.4]
  assign _T_1406 = io_rPort_8_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9852.4]
  assign _T_1411 = io_rPort_9_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9855.4]
  assign _T_1416 = io_rPort_14_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9858.4]
  assign _T_1421 = io_rPort_15_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9861.4]
  assign _T_1426 = io_rPort_19_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9864.4]
  assign _T_1431 = io_rPort_22_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9867.4]
  assign _T_1435 = StickySelects_2_io_outs_0; // @[MemPrimitives.scala 123:41:@9881.4]
  assign _T_1436 = StickySelects_2_io_outs_1; // @[MemPrimitives.scala 123:41:@9882.4]
  assign _T_1437 = StickySelects_2_io_outs_2; // @[MemPrimitives.scala 123:41:@9883.4]
  assign _T_1438 = StickySelects_2_io_outs_3; // @[MemPrimitives.scala 123:41:@9884.4]
  assign _T_1439 = StickySelects_2_io_outs_4; // @[MemPrimitives.scala 123:41:@9885.4]
  assign _T_1440 = StickySelects_2_io_outs_5; // @[MemPrimitives.scala 123:41:@9886.4]
  assign _T_1441 = StickySelects_2_io_outs_6; // @[MemPrimitives.scala 123:41:@9887.4]
  assign _T_1442 = StickySelects_2_io_outs_7; // @[MemPrimitives.scala 123:41:@9888.4]
  assign _T_1444 = {_T_1435,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@9890.4]
  assign _T_1446 = {_T_1436,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@9892.4]
  assign _T_1448 = {_T_1437,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@9894.4]
  assign _T_1450 = {_T_1438,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@9896.4]
  assign _T_1452 = {_T_1439,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@9898.4]
  assign _T_1454 = {_T_1440,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@9900.4]
  assign _T_1456 = {_T_1441,io_rPort_19_backpressure,io_rPort_19_ofs_0}; // @[Cat.scala 30:58:@9902.4]
  assign _T_1458 = {_T_1442,io_rPort_22_backpressure,io_rPort_22_ofs_0}; // @[Cat.scala 30:58:@9904.4]
  assign _T_1459 = _T_1441 ? _T_1456 : _T_1458; // @[Mux.scala 31:69:@9905.4]
  assign _T_1460 = _T_1440 ? _T_1454 : _T_1459; // @[Mux.scala 31:69:@9906.4]
  assign _T_1461 = _T_1439 ? _T_1452 : _T_1460; // @[Mux.scala 31:69:@9907.4]
  assign _T_1462 = _T_1438 ? _T_1450 : _T_1461; // @[Mux.scala 31:69:@9908.4]
  assign _T_1463 = _T_1437 ? _T_1448 : _T_1462; // @[Mux.scala 31:69:@9909.4]
  assign _T_1464 = _T_1436 ? _T_1446 : _T_1463; // @[Mux.scala 31:69:@9910.4]
  assign _T_1465 = _T_1435 ? _T_1444 : _T_1464; // @[Mux.scala 31:69:@9911.4]
  assign _T_1470 = io_rPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9918.4]
  assign _T_1475 = io_rPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9921.4]
  assign _T_1480 = io_rPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9924.4]
  assign _T_1485 = io_rPort_6_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9927.4]
  assign _T_1490 = io_rPort_11_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9930.4]
  assign _T_1495 = io_rPort_17_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9933.4]
  assign _T_1500 = io_rPort_18_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9936.4]
  assign _T_1505 = io_rPort_21_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9939.4]
  assign _T_1509 = StickySelects_3_io_outs_0; // @[MemPrimitives.scala 123:41:@9953.4]
  assign _T_1510 = StickySelects_3_io_outs_1; // @[MemPrimitives.scala 123:41:@9954.4]
  assign _T_1511 = StickySelects_3_io_outs_2; // @[MemPrimitives.scala 123:41:@9955.4]
  assign _T_1512 = StickySelects_3_io_outs_3; // @[MemPrimitives.scala 123:41:@9956.4]
  assign _T_1513 = StickySelects_3_io_outs_4; // @[MemPrimitives.scala 123:41:@9957.4]
  assign _T_1514 = StickySelects_3_io_outs_5; // @[MemPrimitives.scala 123:41:@9958.4]
  assign _T_1515 = StickySelects_3_io_outs_6; // @[MemPrimitives.scala 123:41:@9959.4]
  assign _T_1516 = StickySelects_3_io_outs_7; // @[MemPrimitives.scala 123:41:@9960.4]
  assign _T_1518 = {_T_1509,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@9962.4]
  assign _T_1520 = {_T_1510,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@9964.4]
  assign _T_1522 = {_T_1511,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@9966.4]
  assign _T_1524 = {_T_1512,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@9968.4]
  assign _T_1526 = {_T_1513,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@9970.4]
  assign _T_1528 = {_T_1514,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@9972.4]
  assign _T_1530 = {_T_1515,io_rPort_18_backpressure,io_rPort_18_ofs_0}; // @[Cat.scala 30:58:@9974.4]
  assign _T_1532 = {_T_1516,io_rPort_21_backpressure,io_rPort_21_ofs_0}; // @[Cat.scala 30:58:@9976.4]
  assign _T_1533 = _T_1515 ? _T_1530 : _T_1532; // @[Mux.scala 31:69:@9977.4]
  assign _T_1534 = _T_1514 ? _T_1528 : _T_1533; // @[Mux.scala 31:69:@9978.4]
  assign _T_1535 = _T_1513 ? _T_1526 : _T_1534; // @[Mux.scala 31:69:@9979.4]
  assign _T_1536 = _T_1512 ? _T_1524 : _T_1535; // @[Mux.scala 31:69:@9980.4]
  assign _T_1537 = _T_1511 ? _T_1522 : _T_1536; // @[Mux.scala 31:69:@9981.4]
  assign _T_1538 = _T_1510 ? _T_1520 : _T_1537; // @[Mux.scala 31:69:@9982.4]
  assign _T_1539 = _T_1509 ? _T_1518 : _T_1538; // @[Mux.scala 31:69:@9983.4]
  assign _T_1544 = io_rPort_4_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9990.4]
  assign _T_1549 = io_rPort_12_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9993.4]
  assign _T_1554 = io_rPort_16_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9996.4]
  assign _T_1559 = io_rPort_20_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9999.4]
  assign _T_1563 = StickySelects_4_io_outs_0; // @[MemPrimitives.scala 123:41:@10009.4]
  assign _T_1564 = StickySelects_4_io_outs_1; // @[MemPrimitives.scala 123:41:@10010.4]
  assign _T_1565 = StickySelects_4_io_outs_2; // @[MemPrimitives.scala 123:41:@10011.4]
  assign _T_1566 = StickySelects_4_io_outs_3; // @[MemPrimitives.scala 123:41:@10012.4]
  assign _T_1568 = {_T_1563,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@10014.4]
  assign _T_1570 = {_T_1564,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@10016.4]
  assign _T_1572 = {_T_1565,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@10018.4]
  assign _T_1574 = {_T_1566,io_rPort_20_backpressure,io_rPort_20_ofs_0}; // @[Cat.scala 30:58:@10020.4]
  assign _T_1575 = _T_1565 ? _T_1572 : _T_1574; // @[Mux.scala 31:69:@10021.4]
  assign _T_1576 = _T_1564 ? _T_1570 : _T_1575; // @[Mux.scala 31:69:@10022.4]
  assign _T_1577 = _T_1563 ? _T_1568 : _T_1576; // @[Mux.scala 31:69:@10023.4]
  assign _T_1582 = io_rPort_5_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10030.4]
  assign _T_1587 = io_rPort_10_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10033.4]
  assign _T_1592 = io_rPort_13_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10036.4]
  assign _T_1597 = io_rPort_23_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10039.4]
  assign _T_1601 = StickySelects_5_io_outs_0; // @[MemPrimitives.scala 123:41:@10049.4]
  assign _T_1602 = StickySelects_5_io_outs_1; // @[MemPrimitives.scala 123:41:@10050.4]
  assign _T_1603 = StickySelects_5_io_outs_2; // @[MemPrimitives.scala 123:41:@10051.4]
  assign _T_1604 = StickySelects_5_io_outs_3; // @[MemPrimitives.scala 123:41:@10052.4]
  assign _T_1606 = {_T_1601,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@10054.4]
  assign _T_1608 = {_T_1602,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@10056.4]
  assign _T_1610 = {_T_1603,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@10058.4]
  assign _T_1612 = {_T_1604,io_rPort_23_backpressure,io_rPort_23_ofs_0}; // @[Cat.scala 30:58:@10060.4]
  assign _T_1613 = _T_1603 ? _T_1610 : _T_1612; // @[Mux.scala 31:69:@10061.4]
  assign _T_1614 = _T_1602 ? _T_1608 : _T_1613; // @[Mux.scala 31:69:@10062.4]
  assign _T_1615 = _T_1601 ? _T_1606 : _T_1614; // @[Mux.scala 31:69:@10063.4]
  assign _T_1620 = io_rPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10070.4]
  assign _T_1625 = io_rPort_7_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10073.4]
  assign _T_1630 = io_rPort_8_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10076.4]
  assign _T_1635 = io_rPort_9_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10079.4]
  assign _T_1640 = io_rPort_14_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10082.4]
  assign _T_1645 = io_rPort_15_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10085.4]
  assign _T_1650 = io_rPort_19_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10088.4]
  assign _T_1655 = io_rPort_22_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10091.4]
  assign _T_1659 = StickySelects_6_io_outs_0; // @[MemPrimitives.scala 123:41:@10105.4]
  assign _T_1660 = StickySelects_6_io_outs_1; // @[MemPrimitives.scala 123:41:@10106.4]
  assign _T_1661 = StickySelects_6_io_outs_2; // @[MemPrimitives.scala 123:41:@10107.4]
  assign _T_1662 = StickySelects_6_io_outs_3; // @[MemPrimitives.scala 123:41:@10108.4]
  assign _T_1663 = StickySelects_6_io_outs_4; // @[MemPrimitives.scala 123:41:@10109.4]
  assign _T_1664 = StickySelects_6_io_outs_5; // @[MemPrimitives.scala 123:41:@10110.4]
  assign _T_1665 = StickySelects_6_io_outs_6; // @[MemPrimitives.scala 123:41:@10111.4]
  assign _T_1666 = StickySelects_6_io_outs_7; // @[MemPrimitives.scala 123:41:@10112.4]
  assign _T_1668 = {_T_1659,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@10114.4]
  assign _T_1670 = {_T_1660,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@10116.4]
  assign _T_1672 = {_T_1661,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@10118.4]
  assign _T_1674 = {_T_1662,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@10120.4]
  assign _T_1676 = {_T_1663,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@10122.4]
  assign _T_1678 = {_T_1664,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@10124.4]
  assign _T_1680 = {_T_1665,io_rPort_19_backpressure,io_rPort_19_ofs_0}; // @[Cat.scala 30:58:@10126.4]
  assign _T_1682 = {_T_1666,io_rPort_22_backpressure,io_rPort_22_ofs_0}; // @[Cat.scala 30:58:@10128.4]
  assign _T_1683 = _T_1665 ? _T_1680 : _T_1682; // @[Mux.scala 31:69:@10129.4]
  assign _T_1684 = _T_1664 ? _T_1678 : _T_1683; // @[Mux.scala 31:69:@10130.4]
  assign _T_1685 = _T_1663 ? _T_1676 : _T_1684; // @[Mux.scala 31:69:@10131.4]
  assign _T_1686 = _T_1662 ? _T_1674 : _T_1685; // @[Mux.scala 31:69:@10132.4]
  assign _T_1687 = _T_1661 ? _T_1672 : _T_1686; // @[Mux.scala 31:69:@10133.4]
  assign _T_1688 = _T_1660 ? _T_1670 : _T_1687; // @[Mux.scala 31:69:@10134.4]
  assign _T_1689 = _T_1659 ? _T_1668 : _T_1688; // @[Mux.scala 31:69:@10135.4]
  assign _T_1694 = io_rPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10142.4]
  assign _T_1699 = io_rPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10145.4]
  assign _T_1704 = io_rPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10148.4]
  assign _T_1709 = io_rPort_6_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10151.4]
  assign _T_1714 = io_rPort_11_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10154.4]
  assign _T_1719 = io_rPort_17_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10157.4]
  assign _T_1724 = io_rPort_18_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10160.4]
  assign _T_1729 = io_rPort_21_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10163.4]
  assign _T_1733 = StickySelects_7_io_outs_0; // @[MemPrimitives.scala 123:41:@10177.4]
  assign _T_1734 = StickySelects_7_io_outs_1; // @[MemPrimitives.scala 123:41:@10178.4]
  assign _T_1735 = StickySelects_7_io_outs_2; // @[MemPrimitives.scala 123:41:@10179.4]
  assign _T_1736 = StickySelects_7_io_outs_3; // @[MemPrimitives.scala 123:41:@10180.4]
  assign _T_1737 = StickySelects_7_io_outs_4; // @[MemPrimitives.scala 123:41:@10181.4]
  assign _T_1738 = StickySelects_7_io_outs_5; // @[MemPrimitives.scala 123:41:@10182.4]
  assign _T_1739 = StickySelects_7_io_outs_6; // @[MemPrimitives.scala 123:41:@10183.4]
  assign _T_1740 = StickySelects_7_io_outs_7; // @[MemPrimitives.scala 123:41:@10184.4]
  assign _T_1742 = {_T_1733,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@10186.4]
  assign _T_1744 = {_T_1734,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@10188.4]
  assign _T_1746 = {_T_1735,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@10190.4]
  assign _T_1748 = {_T_1736,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@10192.4]
  assign _T_1750 = {_T_1737,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@10194.4]
  assign _T_1752 = {_T_1738,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@10196.4]
  assign _T_1754 = {_T_1739,io_rPort_18_backpressure,io_rPort_18_ofs_0}; // @[Cat.scala 30:58:@10198.4]
  assign _T_1756 = {_T_1740,io_rPort_21_backpressure,io_rPort_21_ofs_0}; // @[Cat.scala 30:58:@10200.4]
  assign _T_1757 = _T_1739 ? _T_1754 : _T_1756; // @[Mux.scala 31:69:@10201.4]
  assign _T_1758 = _T_1738 ? _T_1752 : _T_1757; // @[Mux.scala 31:69:@10202.4]
  assign _T_1759 = _T_1737 ? _T_1750 : _T_1758; // @[Mux.scala 31:69:@10203.4]
  assign _T_1760 = _T_1736 ? _T_1748 : _T_1759; // @[Mux.scala 31:69:@10204.4]
  assign _T_1761 = _T_1735 ? _T_1746 : _T_1760; // @[Mux.scala 31:69:@10205.4]
  assign _T_1762 = _T_1734 ? _T_1744 : _T_1761; // @[Mux.scala 31:69:@10206.4]
  assign _T_1763 = _T_1733 ? _T_1742 : _T_1762; // @[Mux.scala 31:69:@10207.4]
  assign _T_1768 = io_rPort_4_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10214.4]
  assign _T_1773 = io_rPort_12_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10217.4]
  assign _T_1778 = io_rPort_16_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10220.4]
  assign _T_1783 = io_rPort_20_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10223.4]
  assign _T_1787 = StickySelects_8_io_outs_0; // @[MemPrimitives.scala 123:41:@10233.4]
  assign _T_1788 = StickySelects_8_io_outs_1; // @[MemPrimitives.scala 123:41:@10234.4]
  assign _T_1789 = StickySelects_8_io_outs_2; // @[MemPrimitives.scala 123:41:@10235.4]
  assign _T_1790 = StickySelects_8_io_outs_3; // @[MemPrimitives.scala 123:41:@10236.4]
  assign _T_1792 = {_T_1787,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@10238.4]
  assign _T_1794 = {_T_1788,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@10240.4]
  assign _T_1796 = {_T_1789,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@10242.4]
  assign _T_1798 = {_T_1790,io_rPort_20_backpressure,io_rPort_20_ofs_0}; // @[Cat.scala 30:58:@10244.4]
  assign _T_1799 = _T_1789 ? _T_1796 : _T_1798; // @[Mux.scala 31:69:@10245.4]
  assign _T_1800 = _T_1788 ? _T_1794 : _T_1799; // @[Mux.scala 31:69:@10246.4]
  assign _T_1801 = _T_1787 ? _T_1792 : _T_1800; // @[Mux.scala 31:69:@10247.4]
  assign _T_1806 = io_rPort_5_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10254.4]
  assign _T_1811 = io_rPort_10_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10257.4]
  assign _T_1816 = io_rPort_13_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10260.4]
  assign _T_1821 = io_rPort_23_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10263.4]
  assign _T_1825 = StickySelects_9_io_outs_0; // @[MemPrimitives.scala 123:41:@10273.4]
  assign _T_1826 = StickySelects_9_io_outs_1; // @[MemPrimitives.scala 123:41:@10274.4]
  assign _T_1827 = StickySelects_9_io_outs_2; // @[MemPrimitives.scala 123:41:@10275.4]
  assign _T_1828 = StickySelects_9_io_outs_3; // @[MemPrimitives.scala 123:41:@10276.4]
  assign _T_1830 = {_T_1825,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@10278.4]
  assign _T_1832 = {_T_1826,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@10280.4]
  assign _T_1834 = {_T_1827,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@10282.4]
  assign _T_1836 = {_T_1828,io_rPort_23_backpressure,io_rPort_23_ofs_0}; // @[Cat.scala 30:58:@10284.4]
  assign _T_1837 = _T_1827 ? _T_1834 : _T_1836; // @[Mux.scala 31:69:@10285.4]
  assign _T_1838 = _T_1826 ? _T_1832 : _T_1837; // @[Mux.scala 31:69:@10286.4]
  assign _T_1839 = _T_1825 ? _T_1830 : _T_1838; // @[Mux.scala 31:69:@10287.4]
  assign _T_1844 = io_rPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10294.4]
  assign _T_1849 = io_rPort_7_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10297.4]
  assign _T_1854 = io_rPort_8_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10300.4]
  assign _T_1859 = io_rPort_9_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10303.4]
  assign _T_1864 = io_rPort_14_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10306.4]
  assign _T_1869 = io_rPort_15_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10309.4]
  assign _T_1874 = io_rPort_19_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10312.4]
  assign _T_1879 = io_rPort_22_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10315.4]
  assign _T_1883 = StickySelects_10_io_outs_0; // @[MemPrimitives.scala 123:41:@10329.4]
  assign _T_1884 = StickySelects_10_io_outs_1; // @[MemPrimitives.scala 123:41:@10330.4]
  assign _T_1885 = StickySelects_10_io_outs_2; // @[MemPrimitives.scala 123:41:@10331.4]
  assign _T_1886 = StickySelects_10_io_outs_3; // @[MemPrimitives.scala 123:41:@10332.4]
  assign _T_1887 = StickySelects_10_io_outs_4; // @[MemPrimitives.scala 123:41:@10333.4]
  assign _T_1888 = StickySelects_10_io_outs_5; // @[MemPrimitives.scala 123:41:@10334.4]
  assign _T_1889 = StickySelects_10_io_outs_6; // @[MemPrimitives.scala 123:41:@10335.4]
  assign _T_1890 = StickySelects_10_io_outs_7; // @[MemPrimitives.scala 123:41:@10336.4]
  assign _T_1892 = {_T_1883,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@10338.4]
  assign _T_1894 = {_T_1884,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@10340.4]
  assign _T_1896 = {_T_1885,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@10342.4]
  assign _T_1898 = {_T_1886,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@10344.4]
  assign _T_1900 = {_T_1887,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@10346.4]
  assign _T_1902 = {_T_1888,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@10348.4]
  assign _T_1904 = {_T_1889,io_rPort_19_backpressure,io_rPort_19_ofs_0}; // @[Cat.scala 30:58:@10350.4]
  assign _T_1906 = {_T_1890,io_rPort_22_backpressure,io_rPort_22_ofs_0}; // @[Cat.scala 30:58:@10352.4]
  assign _T_1907 = _T_1889 ? _T_1904 : _T_1906; // @[Mux.scala 31:69:@10353.4]
  assign _T_1908 = _T_1888 ? _T_1902 : _T_1907; // @[Mux.scala 31:69:@10354.4]
  assign _T_1909 = _T_1887 ? _T_1900 : _T_1908; // @[Mux.scala 31:69:@10355.4]
  assign _T_1910 = _T_1886 ? _T_1898 : _T_1909; // @[Mux.scala 31:69:@10356.4]
  assign _T_1911 = _T_1885 ? _T_1896 : _T_1910; // @[Mux.scala 31:69:@10357.4]
  assign _T_1912 = _T_1884 ? _T_1894 : _T_1911; // @[Mux.scala 31:69:@10358.4]
  assign _T_1913 = _T_1883 ? _T_1892 : _T_1912; // @[Mux.scala 31:69:@10359.4]
  assign _T_1918 = io_rPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10366.4]
  assign _T_1923 = io_rPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10369.4]
  assign _T_1928 = io_rPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10372.4]
  assign _T_1933 = io_rPort_6_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10375.4]
  assign _T_1938 = io_rPort_11_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10378.4]
  assign _T_1943 = io_rPort_17_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10381.4]
  assign _T_1948 = io_rPort_18_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10384.4]
  assign _T_1953 = io_rPort_21_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10387.4]
  assign _T_1957 = StickySelects_11_io_outs_0; // @[MemPrimitives.scala 123:41:@10401.4]
  assign _T_1958 = StickySelects_11_io_outs_1; // @[MemPrimitives.scala 123:41:@10402.4]
  assign _T_1959 = StickySelects_11_io_outs_2; // @[MemPrimitives.scala 123:41:@10403.4]
  assign _T_1960 = StickySelects_11_io_outs_3; // @[MemPrimitives.scala 123:41:@10404.4]
  assign _T_1961 = StickySelects_11_io_outs_4; // @[MemPrimitives.scala 123:41:@10405.4]
  assign _T_1962 = StickySelects_11_io_outs_5; // @[MemPrimitives.scala 123:41:@10406.4]
  assign _T_1963 = StickySelects_11_io_outs_6; // @[MemPrimitives.scala 123:41:@10407.4]
  assign _T_1964 = StickySelects_11_io_outs_7; // @[MemPrimitives.scala 123:41:@10408.4]
  assign _T_1966 = {_T_1957,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@10410.4]
  assign _T_1968 = {_T_1958,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@10412.4]
  assign _T_1970 = {_T_1959,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@10414.4]
  assign _T_1972 = {_T_1960,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@10416.4]
  assign _T_1974 = {_T_1961,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@10418.4]
  assign _T_1976 = {_T_1962,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@10420.4]
  assign _T_1978 = {_T_1963,io_rPort_18_backpressure,io_rPort_18_ofs_0}; // @[Cat.scala 30:58:@10422.4]
  assign _T_1980 = {_T_1964,io_rPort_21_backpressure,io_rPort_21_ofs_0}; // @[Cat.scala 30:58:@10424.4]
  assign _T_1981 = _T_1963 ? _T_1978 : _T_1980; // @[Mux.scala 31:69:@10425.4]
  assign _T_1982 = _T_1962 ? _T_1976 : _T_1981; // @[Mux.scala 31:69:@10426.4]
  assign _T_1983 = _T_1961 ? _T_1974 : _T_1982; // @[Mux.scala 31:69:@10427.4]
  assign _T_1984 = _T_1960 ? _T_1972 : _T_1983; // @[Mux.scala 31:69:@10428.4]
  assign _T_1985 = _T_1959 ? _T_1970 : _T_1984; // @[Mux.scala 31:69:@10429.4]
  assign _T_1986 = _T_1958 ? _T_1968 : _T_1985; // @[Mux.scala 31:69:@10430.4]
  assign _T_1987 = _T_1957 ? _T_1966 : _T_1986; // @[Mux.scala 31:69:@10431.4]
  assign _T_1992 = io_rPort_4_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10438.4]
  assign _T_1997 = io_rPort_12_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10441.4]
  assign _T_2002 = io_rPort_16_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10444.4]
  assign _T_2007 = io_rPort_20_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10447.4]
  assign _T_2011 = StickySelects_12_io_outs_0; // @[MemPrimitives.scala 123:41:@10457.4]
  assign _T_2012 = StickySelects_12_io_outs_1; // @[MemPrimitives.scala 123:41:@10458.4]
  assign _T_2013 = StickySelects_12_io_outs_2; // @[MemPrimitives.scala 123:41:@10459.4]
  assign _T_2014 = StickySelects_12_io_outs_3; // @[MemPrimitives.scala 123:41:@10460.4]
  assign _T_2016 = {_T_2011,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@10462.4]
  assign _T_2018 = {_T_2012,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@10464.4]
  assign _T_2020 = {_T_2013,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@10466.4]
  assign _T_2022 = {_T_2014,io_rPort_20_backpressure,io_rPort_20_ofs_0}; // @[Cat.scala 30:58:@10468.4]
  assign _T_2023 = _T_2013 ? _T_2020 : _T_2022; // @[Mux.scala 31:69:@10469.4]
  assign _T_2024 = _T_2012 ? _T_2018 : _T_2023; // @[Mux.scala 31:69:@10470.4]
  assign _T_2025 = _T_2011 ? _T_2016 : _T_2024; // @[Mux.scala 31:69:@10471.4]
  assign _T_2030 = io_rPort_5_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10478.4]
  assign _T_2035 = io_rPort_10_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10481.4]
  assign _T_2040 = io_rPort_13_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10484.4]
  assign _T_2045 = io_rPort_23_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10487.4]
  assign _T_2049 = StickySelects_13_io_outs_0; // @[MemPrimitives.scala 123:41:@10497.4]
  assign _T_2050 = StickySelects_13_io_outs_1; // @[MemPrimitives.scala 123:41:@10498.4]
  assign _T_2051 = StickySelects_13_io_outs_2; // @[MemPrimitives.scala 123:41:@10499.4]
  assign _T_2052 = StickySelects_13_io_outs_3; // @[MemPrimitives.scala 123:41:@10500.4]
  assign _T_2054 = {_T_2049,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@10502.4]
  assign _T_2056 = {_T_2050,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@10504.4]
  assign _T_2058 = {_T_2051,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@10506.4]
  assign _T_2060 = {_T_2052,io_rPort_23_backpressure,io_rPort_23_ofs_0}; // @[Cat.scala 30:58:@10508.4]
  assign _T_2061 = _T_2051 ? _T_2058 : _T_2060; // @[Mux.scala 31:69:@10509.4]
  assign _T_2062 = _T_2050 ? _T_2056 : _T_2061; // @[Mux.scala 31:69:@10510.4]
  assign _T_2063 = _T_2049 ? _T_2054 : _T_2062; // @[Mux.scala 31:69:@10511.4]
  assign _T_2068 = io_rPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10518.4]
  assign _T_2073 = io_rPort_7_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10521.4]
  assign _T_2078 = io_rPort_8_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10524.4]
  assign _T_2083 = io_rPort_9_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10527.4]
  assign _T_2088 = io_rPort_14_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10530.4]
  assign _T_2093 = io_rPort_15_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10533.4]
  assign _T_2098 = io_rPort_19_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10536.4]
  assign _T_2103 = io_rPort_22_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10539.4]
  assign _T_2107 = StickySelects_14_io_outs_0; // @[MemPrimitives.scala 123:41:@10553.4]
  assign _T_2108 = StickySelects_14_io_outs_1; // @[MemPrimitives.scala 123:41:@10554.4]
  assign _T_2109 = StickySelects_14_io_outs_2; // @[MemPrimitives.scala 123:41:@10555.4]
  assign _T_2110 = StickySelects_14_io_outs_3; // @[MemPrimitives.scala 123:41:@10556.4]
  assign _T_2111 = StickySelects_14_io_outs_4; // @[MemPrimitives.scala 123:41:@10557.4]
  assign _T_2112 = StickySelects_14_io_outs_5; // @[MemPrimitives.scala 123:41:@10558.4]
  assign _T_2113 = StickySelects_14_io_outs_6; // @[MemPrimitives.scala 123:41:@10559.4]
  assign _T_2114 = StickySelects_14_io_outs_7; // @[MemPrimitives.scala 123:41:@10560.4]
  assign _T_2116 = {_T_2107,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@10562.4]
  assign _T_2118 = {_T_2108,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@10564.4]
  assign _T_2120 = {_T_2109,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@10566.4]
  assign _T_2122 = {_T_2110,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@10568.4]
  assign _T_2124 = {_T_2111,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@10570.4]
  assign _T_2126 = {_T_2112,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@10572.4]
  assign _T_2128 = {_T_2113,io_rPort_19_backpressure,io_rPort_19_ofs_0}; // @[Cat.scala 30:58:@10574.4]
  assign _T_2130 = {_T_2114,io_rPort_22_backpressure,io_rPort_22_ofs_0}; // @[Cat.scala 30:58:@10576.4]
  assign _T_2131 = _T_2113 ? _T_2128 : _T_2130; // @[Mux.scala 31:69:@10577.4]
  assign _T_2132 = _T_2112 ? _T_2126 : _T_2131; // @[Mux.scala 31:69:@10578.4]
  assign _T_2133 = _T_2111 ? _T_2124 : _T_2132; // @[Mux.scala 31:69:@10579.4]
  assign _T_2134 = _T_2110 ? _T_2122 : _T_2133; // @[Mux.scala 31:69:@10580.4]
  assign _T_2135 = _T_2109 ? _T_2120 : _T_2134; // @[Mux.scala 31:69:@10581.4]
  assign _T_2136 = _T_2108 ? _T_2118 : _T_2135; // @[Mux.scala 31:69:@10582.4]
  assign _T_2137 = _T_2107 ? _T_2116 : _T_2136; // @[Mux.scala 31:69:@10583.4]
  assign _T_2142 = io_rPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10590.4]
  assign _T_2147 = io_rPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10593.4]
  assign _T_2152 = io_rPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10596.4]
  assign _T_2157 = io_rPort_6_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10599.4]
  assign _T_2162 = io_rPort_11_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10602.4]
  assign _T_2167 = io_rPort_17_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10605.4]
  assign _T_2172 = io_rPort_18_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10608.4]
  assign _T_2177 = io_rPort_21_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10611.4]
  assign _T_2181 = StickySelects_15_io_outs_0; // @[MemPrimitives.scala 123:41:@10625.4]
  assign _T_2182 = StickySelects_15_io_outs_1; // @[MemPrimitives.scala 123:41:@10626.4]
  assign _T_2183 = StickySelects_15_io_outs_2; // @[MemPrimitives.scala 123:41:@10627.4]
  assign _T_2184 = StickySelects_15_io_outs_3; // @[MemPrimitives.scala 123:41:@10628.4]
  assign _T_2185 = StickySelects_15_io_outs_4; // @[MemPrimitives.scala 123:41:@10629.4]
  assign _T_2186 = StickySelects_15_io_outs_5; // @[MemPrimitives.scala 123:41:@10630.4]
  assign _T_2187 = StickySelects_15_io_outs_6; // @[MemPrimitives.scala 123:41:@10631.4]
  assign _T_2188 = StickySelects_15_io_outs_7; // @[MemPrimitives.scala 123:41:@10632.4]
  assign _T_2190 = {_T_2181,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@10634.4]
  assign _T_2192 = {_T_2182,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@10636.4]
  assign _T_2194 = {_T_2183,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@10638.4]
  assign _T_2196 = {_T_2184,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@10640.4]
  assign _T_2198 = {_T_2185,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@10642.4]
  assign _T_2200 = {_T_2186,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@10644.4]
  assign _T_2202 = {_T_2187,io_rPort_18_backpressure,io_rPort_18_ofs_0}; // @[Cat.scala 30:58:@10646.4]
  assign _T_2204 = {_T_2188,io_rPort_21_backpressure,io_rPort_21_ofs_0}; // @[Cat.scala 30:58:@10648.4]
  assign _T_2205 = _T_2187 ? _T_2202 : _T_2204; // @[Mux.scala 31:69:@10649.4]
  assign _T_2206 = _T_2186 ? _T_2200 : _T_2205; // @[Mux.scala 31:69:@10650.4]
  assign _T_2207 = _T_2185 ? _T_2198 : _T_2206; // @[Mux.scala 31:69:@10651.4]
  assign _T_2208 = _T_2184 ? _T_2196 : _T_2207; // @[Mux.scala 31:69:@10652.4]
  assign _T_2209 = _T_2183 ? _T_2194 : _T_2208; // @[Mux.scala 31:69:@10653.4]
  assign _T_2210 = _T_2182 ? _T_2192 : _T_2209; // @[Mux.scala 31:69:@10654.4]
  assign _T_2211 = _T_2181 ? _T_2190 : _T_2210; // @[Mux.scala 31:69:@10655.4]
  assign _T_2243 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@10696.4 package.scala 96:25:@10697.4]
  assign _T_2247 = _T_2243 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@10706.4]
  assign _T_2240 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@10688.4 package.scala 96:25:@10689.4]
  assign _T_2248 = _T_2240 ? Mem1D_7_io_output : _T_2247; // @[Mux.scala 31:69:@10707.4]
  assign _T_2237 = RetimeWrapper_io_out; // @[package.scala 96:25:@10680.4 package.scala 96:25:@10681.4]
  assign _T_2278 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@10744.4 package.scala 96:25:@10745.4]
  assign _T_2282 = _T_2278 ? Mem1D_10_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@10754.4]
  assign _T_2275 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@10736.4 package.scala 96:25:@10737.4]
  assign _T_2283 = _T_2275 ? Mem1D_6_io_output : _T_2282; // @[Mux.scala 31:69:@10755.4]
  assign _T_2272 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@10728.4 package.scala 96:25:@10729.4]
  assign _T_2313 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@10792.4 package.scala 96:25:@10793.4]
  assign _T_2317 = _T_2313 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@10802.4]
  assign _T_2310 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@10784.4 package.scala 96:25:@10785.4]
  assign _T_2318 = _T_2310 ? Mem1D_7_io_output : _T_2317; // @[Mux.scala 31:69:@10803.4]
  assign _T_2307 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@10776.4 package.scala 96:25:@10777.4]
  assign _T_2348 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@10840.4 package.scala 96:25:@10841.4]
  assign _T_2352 = _T_2348 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@10850.4]
  assign _T_2345 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@10832.4 package.scala 96:25:@10833.4]
  assign _T_2353 = _T_2345 ? Mem1D_7_io_output : _T_2352; // @[Mux.scala 31:69:@10851.4]
  assign _T_2342 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@10824.4 package.scala 96:25:@10825.4]
  assign _T_2383 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@10888.4 package.scala 96:25:@10889.4]
  assign _T_2387 = _T_2383 ? Mem1D_8_io_output : Mem1D_12_io_output; // @[Mux.scala 31:69:@10898.4]
  assign _T_2380 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@10880.4 package.scala 96:25:@10881.4]
  assign _T_2388 = _T_2380 ? Mem1D_4_io_output : _T_2387; // @[Mux.scala 31:69:@10899.4]
  assign _T_2377 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@10872.4 package.scala 96:25:@10873.4]
  assign _T_2418 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@10936.4 package.scala 96:25:@10937.4]
  assign _T_2422 = _T_2418 ? Mem1D_9_io_output : Mem1D_13_io_output; // @[Mux.scala 31:69:@10946.4]
  assign _T_2415 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@10928.4 package.scala 96:25:@10929.4]
  assign _T_2423 = _T_2415 ? Mem1D_5_io_output : _T_2422; // @[Mux.scala 31:69:@10947.4]
  assign _T_2412 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@10920.4 package.scala 96:25:@10921.4]
  assign _T_2453 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@10984.4 package.scala 96:25:@10985.4]
  assign _T_2457 = _T_2453 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@10994.4]
  assign _T_2450 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@10976.4 package.scala 96:25:@10977.4]
  assign _T_2458 = _T_2450 ? Mem1D_7_io_output : _T_2457; // @[Mux.scala 31:69:@10995.4]
  assign _T_2447 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@10968.4 package.scala 96:25:@10969.4]
  assign _T_2488 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@11032.4 package.scala 96:25:@11033.4]
  assign _T_2492 = _T_2488 ? Mem1D_10_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@11042.4]
  assign _T_2485 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@11024.4 package.scala 96:25:@11025.4]
  assign _T_2493 = _T_2485 ? Mem1D_6_io_output : _T_2492; // @[Mux.scala 31:69:@11043.4]
  assign _T_2482 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@11016.4 package.scala 96:25:@11017.4]
  assign _T_2523 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@11080.4 package.scala 96:25:@11081.4]
  assign _T_2527 = _T_2523 ? Mem1D_10_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@11090.4]
  assign _T_2520 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@11072.4 package.scala 96:25:@11073.4]
  assign _T_2528 = _T_2520 ? Mem1D_6_io_output : _T_2527; // @[Mux.scala 31:69:@11091.4]
  assign _T_2517 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@11064.4 package.scala 96:25:@11065.4]
  assign _T_2558 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@11128.4 package.scala 96:25:@11129.4]
  assign _T_2562 = _T_2558 ? Mem1D_10_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@11138.4]
  assign _T_2555 = RetimeWrapper_37_io_out; // @[package.scala 96:25:@11120.4 package.scala 96:25:@11121.4]
  assign _T_2563 = _T_2555 ? Mem1D_6_io_output : _T_2562; // @[Mux.scala 31:69:@11139.4]
  assign _T_2552 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@11112.4 package.scala 96:25:@11113.4]
  assign _T_2593 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@11176.4 package.scala 96:25:@11177.4]
  assign _T_2597 = _T_2593 ? Mem1D_9_io_output : Mem1D_13_io_output; // @[Mux.scala 31:69:@11186.4]
  assign _T_2590 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@11168.4 package.scala 96:25:@11169.4]
  assign _T_2598 = _T_2590 ? Mem1D_5_io_output : _T_2597; // @[Mux.scala 31:69:@11187.4]
  assign _T_2587 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@11160.4 package.scala 96:25:@11161.4]
  assign _T_2628 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@11224.4 package.scala 96:25:@11225.4]
  assign _T_2632 = _T_2628 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@11234.4]
  assign _T_2625 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@11216.4 package.scala 96:25:@11217.4]
  assign _T_2633 = _T_2625 ? Mem1D_7_io_output : _T_2632; // @[Mux.scala 31:69:@11235.4]
  assign _T_2622 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@11208.4 package.scala 96:25:@11209.4]
  assign _T_2663 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@11272.4 package.scala 96:25:@11273.4]
  assign _T_2667 = _T_2663 ? Mem1D_8_io_output : Mem1D_12_io_output; // @[Mux.scala 31:69:@11282.4]
  assign _T_2660 = RetimeWrapper_49_io_out; // @[package.scala 96:25:@11264.4 package.scala 96:25:@11265.4]
  assign _T_2668 = _T_2660 ? Mem1D_4_io_output : _T_2667; // @[Mux.scala 31:69:@11283.4]
  assign _T_2657 = RetimeWrapper_48_io_out; // @[package.scala 96:25:@11256.4 package.scala 96:25:@11257.4]
  assign _T_2698 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@11320.4 package.scala 96:25:@11321.4]
  assign _T_2702 = _T_2698 ? Mem1D_9_io_output : Mem1D_13_io_output; // @[Mux.scala 31:69:@11330.4]
  assign _T_2695 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@11312.4 package.scala 96:25:@11313.4]
  assign _T_2703 = _T_2695 ? Mem1D_5_io_output : _T_2702; // @[Mux.scala 31:69:@11331.4]
  assign _T_2692 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@11304.4 package.scala 96:25:@11305.4]
  assign _T_2733 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@11368.4 package.scala 96:25:@11369.4]
  assign _T_2737 = _T_2733 ? Mem1D_10_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@11378.4]
  assign _T_2730 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@11360.4 package.scala 96:25:@11361.4]
  assign _T_2738 = _T_2730 ? Mem1D_6_io_output : _T_2737; // @[Mux.scala 31:69:@11379.4]
  assign _T_2727 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@11352.4 package.scala 96:25:@11353.4]
  assign _T_2768 = RetimeWrapper_62_io_out; // @[package.scala 96:25:@11416.4 package.scala 96:25:@11417.4]
  assign _T_2772 = _T_2768 ? Mem1D_10_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@11426.4]
  assign _T_2765 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@11408.4 package.scala 96:25:@11409.4]
  assign _T_2773 = _T_2765 ? Mem1D_6_io_output : _T_2772; // @[Mux.scala 31:69:@11427.4]
  assign _T_2762 = RetimeWrapper_60_io_out; // @[package.scala 96:25:@11400.4 package.scala 96:25:@11401.4]
  assign _T_2803 = RetimeWrapper_66_io_out; // @[package.scala 96:25:@11464.4 package.scala 96:25:@11465.4]
  assign _T_2807 = _T_2803 ? Mem1D_8_io_output : Mem1D_12_io_output; // @[Mux.scala 31:69:@11474.4]
  assign _T_2800 = RetimeWrapper_65_io_out; // @[package.scala 96:25:@11456.4 package.scala 96:25:@11457.4]
  assign _T_2808 = _T_2800 ? Mem1D_4_io_output : _T_2807; // @[Mux.scala 31:69:@11475.4]
  assign _T_2797 = RetimeWrapper_64_io_out; // @[package.scala 96:25:@11448.4 package.scala 96:25:@11449.4]
  assign _T_2838 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@11512.4 package.scala 96:25:@11513.4]
  assign _T_2842 = _T_2838 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@11522.4]
  assign _T_2835 = RetimeWrapper_69_io_out; // @[package.scala 96:25:@11504.4 package.scala 96:25:@11505.4]
  assign _T_2843 = _T_2835 ? Mem1D_7_io_output : _T_2842; // @[Mux.scala 31:69:@11523.4]
  assign _T_2832 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@11496.4 package.scala 96:25:@11497.4]
  assign _T_2873 = RetimeWrapper_74_io_out; // @[package.scala 96:25:@11560.4 package.scala 96:25:@11561.4]
  assign _T_2877 = _T_2873 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@11570.4]
  assign _T_2870 = RetimeWrapper_73_io_out; // @[package.scala 96:25:@11552.4 package.scala 96:25:@11553.4]
  assign _T_2878 = _T_2870 ? Mem1D_7_io_output : _T_2877; // @[Mux.scala 31:69:@11571.4]
  assign _T_2867 = RetimeWrapper_72_io_out; // @[package.scala 96:25:@11544.4 package.scala 96:25:@11545.4]
  assign _T_2908 = RetimeWrapper_78_io_out; // @[package.scala 96:25:@11608.4 package.scala 96:25:@11609.4]
  assign _T_2912 = _T_2908 ? Mem1D_10_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@11618.4]
  assign _T_2905 = RetimeWrapper_77_io_out; // @[package.scala 96:25:@11600.4 package.scala 96:25:@11601.4]
  assign _T_2913 = _T_2905 ? Mem1D_6_io_output : _T_2912; // @[Mux.scala 31:69:@11619.4]
  assign _T_2902 = RetimeWrapper_76_io_out; // @[package.scala 96:25:@11592.4 package.scala 96:25:@11593.4]
  assign _T_2943 = RetimeWrapper_82_io_out; // @[package.scala 96:25:@11656.4 package.scala 96:25:@11657.4]
  assign _T_2947 = _T_2943 ? Mem1D_8_io_output : Mem1D_12_io_output; // @[Mux.scala 31:69:@11666.4]
  assign _T_2940 = RetimeWrapper_81_io_out; // @[package.scala 96:25:@11648.4 package.scala 96:25:@11649.4]
  assign _T_2948 = _T_2940 ? Mem1D_4_io_output : _T_2947; // @[Mux.scala 31:69:@11667.4]
  assign _T_2937 = RetimeWrapper_80_io_out; // @[package.scala 96:25:@11640.4 package.scala 96:25:@11641.4]
  assign _T_2978 = RetimeWrapper_86_io_out; // @[package.scala 96:25:@11704.4 package.scala 96:25:@11705.4]
  assign _T_2982 = _T_2978 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@11714.4]
  assign _T_2975 = RetimeWrapper_85_io_out; // @[package.scala 96:25:@11696.4 package.scala 96:25:@11697.4]
  assign _T_2983 = _T_2975 ? Mem1D_7_io_output : _T_2982; // @[Mux.scala 31:69:@11715.4]
  assign _T_2972 = RetimeWrapper_84_io_out; // @[package.scala 96:25:@11688.4 package.scala 96:25:@11689.4]
  assign _T_3013 = RetimeWrapper_90_io_out; // @[package.scala 96:25:@11752.4 package.scala 96:25:@11753.4]
  assign _T_3017 = _T_3013 ? Mem1D_10_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@11762.4]
  assign _T_3010 = RetimeWrapper_89_io_out; // @[package.scala 96:25:@11744.4 package.scala 96:25:@11745.4]
  assign _T_3018 = _T_3010 ? Mem1D_6_io_output : _T_3017; // @[Mux.scala 31:69:@11763.4]
  assign _T_3007 = RetimeWrapper_88_io_out; // @[package.scala 96:25:@11736.4 package.scala 96:25:@11737.4]
  assign _T_3048 = RetimeWrapper_94_io_out; // @[package.scala 96:25:@11800.4 package.scala 96:25:@11801.4]
  assign _T_3052 = _T_3048 ? Mem1D_9_io_output : Mem1D_13_io_output; // @[Mux.scala 31:69:@11810.4]
  assign _T_3045 = RetimeWrapper_93_io_out; // @[package.scala 96:25:@11792.4 package.scala 96:25:@11793.4]
  assign _T_3053 = _T_3045 ? Mem1D_5_io_output : _T_3052; // @[Mux.scala 31:69:@11811.4]
  assign _T_3042 = RetimeWrapper_92_io_out; // @[package.scala 96:25:@11784.4 package.scala 96:25:@11785.4]
  assign io_rPort_23_output_0 = _T_3042 ? Mem1D_1_io_output : _T_3053; // @[MemPrimitives.scala 148:13:@11813.4]
  assign io_rPort_22_output_0 = _T_3007 ? Mem1D_2_io_output : _T_3018; // @[MemPrimitives.scala 148:13:@11765.4]
  assign io_rPort_21_output_0 = _T_2972 ? Mem1D_3_io_output : _T_2983; // @[MemPrimitives.scala 148:13:@11717.4]
  assign io_rPort_20_output_0 = _T_2937 ? Mem1D_io_output : _T_2948; // @[MemPrimitives.scala 148:13:@11669.4]
  assign io_rPort_19_output_0 = _T_2902 ? Mem1D_2_io_output : _T_2913; // @[MemPrimitives.scala 148:13:@11621.4]
  assign io_rPort_18_output_0 = _T_2867 ? Mem1D_3_io_output : _T_2878; // @[MemPrimitives.scala 148:13:@11573.4]
  assign io_rPort_17_output_0 = _T_2832 ? Mem1D_3_io_output : _T_2843; // @[MemPrimitives.scala 148:13:@11525.4]
  assign io_rPort_16_output_0 = _T_2797 ? Mem1D_io_output : _T_2808; // @[MemPrimitives.scala 148:13:@11477.4]
  assign io_rPort_15_output_0 = _T_2762 ? Mem1D_2_io_output : _T_2773; // @[MemPrimitives.scala 148:13:@11429.4]
  assign io_rPort_14_output_0 = _T_2727 ? Mem1D_2_io_output : _T_2738; // @[MemPrimitives.scala 148:13:@11381.4]
  assign io_rPort_13_output_0 = _T_2692 ? Mem1D_1_io_output : _T_2703; // @[MemPrimitives.scala 148:13:@11333.4]
  assign io_rPort_12_output_0 = _T_2657 ? Mem1D_io_output : _T_2668; // @[MemPrimitives.scala 148:13:@11285.4]
  assign io_rPort_11_output_0 = _T_2622 ? Mem1D_3_io_output : _T_2633; // @[MemPrimitives.scala 148:13:@11237.4]
  assign io_rPort_10_output_0 = _T_2587 ? Mem1D_1_io_output : _T_2598; // @[MemPrimitives.scala 148:13:@11189.4]
  assign io_rPort_9_output_0 = _T_2552 ? Mem1D_2_io_output : _T_2563; // @[MemPrimitives.scala 148:13:@11141.4]
  assign io_rPort_8_output_0 = _T_2517 ? Mem1D_2_io_output : _T_2528; // @[MemPrimitives.scala 148:13:@11093.4]
  assign io_rPort_7_output_0 = _T_2482 ? Mem1D_2_io_output : _T_2493; // @[MemPrimitives.scala 148:13:@11045.4]
  assign io_rPort_6_output_0 = _T_2447 ? Mem1D_3_io_output : _T_2458; // @[MemPrimitives.scala 148:13:@10997.4]
  assign io_rPort_5_output_0 = _T_2412 ? Mem1D_1_io_output : _T_2423; // @[MemPrimitives.scala 148:13:@10949.4]
  assign io_rPort_4_output_0 = _T_2377 ? Mem1D_io_output : _T_2388; // @[MemPrimitives.scala 148:13:@10901.4]
  assign io_rPort_3_output_0 = _T_2342 ? Mem1D_3_io_output : _T_2353; // @[MemPrimitives.scala 148:13:@10853.4]
  assign io_rPort_2_output_0 = _T_2307 ? Mem1D_3_io_output : _T_2318; // @[MemPrimitives.scala 148:13:@10805.4]
  assign io_rPort_1_output_0 = _T_2272 ? Mem1D_2_io_output : _T_2283; // @[MemPrimitives.scala 148:13:@10757.4]
  assign io_rPort_0_output_0 = _T_2237 ? Mem1D_3_io_output : _T_2248; // @[MemPrimitives.scala 148:13:@10709.4]
  assign Mem1D_clock = clock; // @[:@9239.4]
  assign Mem1D_reset = reset; // @[:@9240.4]
  assign Mem1D_io_r_ofs_0 = _T_1353[0]; // @[MemPrimitives.scala 127:28:@9803.4]
  assign Mem1D_io_r_backpressure = _T_1353[1]; // @[MemPrimitives.scala 128:32:@9804.4]
  assign Mem1D_io_w_ofs_0 = _T_1045[0]; // @[MemPrimitives.scala 94:28:@9508.4]
  assign Mem1D_io_w_data_0 = _T_1045[8:1]; // @[MemPrimitives.scala 95:29:@9509.4]
  assign Mem1D_io_w_en_0 = _T_1045[9]; // @[MemPrimitives.scala 96:27:@9510.4]
  assign Mem1D_1_clock = clock; // @[:@9255.4]
  assign Mem1D_1_reset = reset; // @[:@9256.4]
  assign Mem1D_1_io_r_ofs_0 = _T_1391[0]; // @[MemPrimitives.scala 127:28:@9843.4]
  assign Mem1D_1_io_r_backpressure = _T_1391[1]; // @[MemPrimitives.scala 128:32:@9844.4]
  assign Mem1D_1_io_w_ofs_0 = _T_1063[0]; // @[MemPrimitives.scala 94:28:@9525.4]
  assign Mem1D_1_io_w_data_0 = _T_1063[8:1]; // @[MemPrimitives.scala 95:29:@9526.4]
  assign Mem1D_1_io_w_en_0 = _T_1063[9]; // @[MemPrimitives.scala 96:27:@9527.4]
  assign Mem1D_2_clock = clock; // @[:@9271.4]
  assign Mem1D_2_reset = reset; // @[:@9272.4]
  assign Mem1D_2_io_r_ofs_0 = _T_1465[0]; // @[MemPrimitives.scala 127:28:@9915.4]
  assign Mem1D_2_io_r_backpressure = _T_1465[1]; // @[MemPrimitives.scala 128:32:@9916.4]
  assign Mem1D_2_io_w_ofs_0 = _T_1081[0]; // @[MemPrimitives.scala 94:28:@9542.4]
  assign Mem1D_2_io_w_data_0 = _T_1081[8:1]; // @[MemPrimitives.scala 95:29:@9543.4]
  assign Mem1D_2_io_w_en_0 = _T_1081[9]; // @[MemPrimitives.scala 96:27:@9544.4]
  assign Mem1D_3_clock = clock; // @[:@9287.4]
  assign Mem1D_3_reset = reset; // @[:@9288.4]
  assign Mem1D_3_io_r_ofs_0 = _T_1539[0]; // @[MemPrimitives.scala 127:28:@9987.4]
  assign Mem1D_3_io_r_backpressure = _T_1539[1]; // @[MemPrimitives.scala 128:32:@9988.4]
  assign Mem1D_3_io_w_ofs_0 = _T_1099[0]; // @[MemPrimitives.scala 94:28:@9559.4]
  assign Mem1D_3_io_w_data_0 = _T_1099[8:1]; // @[MemPrimitives.scala 95:29:@9560.4]
  assign Mem1D_3_io_w_en_0 = _T_1099[9]; // @[MemPrimitives.scala 96:27:@9561.4]
  assign Mem1D_4_clock = clock; // @[:@9303.4]
  assign Mem1D_4_reset = reset; // @[:@9304.4]
  assign Mem1D_4_io_r_ofs_0 = _T_1577[0]; // @[MemPrimitives.scala 127:28:@10027.4]
  assign Mem1D_4_io_r_backpressure = _T_1577[1]; // @[MemPrimitives.scala 128:32:@10028.4]
  assign Mem1D_4_io_w_ofs_0 = _T_1117[0]; // @[MemPrimitives.scala 94:28:@9576.4]
  assign Mem1D_4_io_w_data_0 = _T_1117[8:1]; // @[MemPrimitives.scala 95:29:@9577.4]
  assign Mem1D_4_io_w_en_0 = _T_1117[9]; // @[MemPrimitives.scala 96:27:@9578.4]
  assign Mem1D_5_clock = clock; // @[:@9319.4]
  assign Mem1D_5_reset = reset; // @[:@9320.4]
  assign Mem1D_5_io_r_ofs_0 = _T_1615[0]; // @[MemPrimitives.scala 127:28:@10067.4]
  assign Mem1D_5_io_r_backpressure = _T_1615[1]; // @[MemPrimitives.scala 128:32:@10068.4]
  assign Mem1D_5_io_w_ofs_0 = _T_1135[0]; // @[MemPrimitives.scala 94:28:@9593.4]
  assign Mem1D_5_io_w_data_0 = _T_1135[8:1]; // @[MemPrimitives.scala 95:29:@9594.4]
  assign Mem1D_5_io_w_en_0 = _T_1135[9]; // @[MemPrimitives.scala 96:27:@9595.4]
  assign Mem1D_6_clock = clock; // @[:@9335.4]
  assign Mem1D_6_reset = reset; // @[:@9336.4]
  assign Mem1D_6_io_r_ofs_0 = _T_1689[0]; // @[MemPrimitives.scala 127:28:@10139.4]
  assign Mem1D_6_io_r_backpressure = _T_1689[1]; // @[MemPrimitives.scala 128:32:@10140.4]
  assign Mem1D_6_io_w_ofs_0 = _T_1153[0]; // @[MemPrimitives.scala 94:28:@9610.4]
  assign Mem1D_6_io_w_data_0 = _T_1153[8:1]; // @[MemPrimitives.scala 95:29:@9611.4]
  assign Mem1D_6_io_w_en_0 = _T_1153[9]; // @[MemPrimitives.scala 96:27:@9612.4]
  assign Mem1D_7_clock = clock; // @[:@9351.4]
  assign Mem1D_7_reset = reset; // @[:@9352.4]
  assign Mem1D_7_io_r_ofs_0 = _T_1763[0]; // @[MemPrimitives.scala 127:28:@10211.4]
  assign Mem1D_7_io_r_backpressure = _T_1763[1]; // @[MemPrimitives.scala 128:32:@10212.4]
  assign Mem1D_7_io_w_ofs_0 = _T_1171[0]; // @[MemPrimitives.scala 94:28:@9627.4]
  assign Mem1D_7_io_w_data_0 = _T_1171[8:1]; // @[MemPrimitives.scala 95:29:@9628.4]
  assign Mem1D_7_io_w_en_0 = _T_1171[9]; // @[MemPrimitives.scala 96:27:@9629.4]
  assign Mem1D_8_clock = clock; // @[:@9367.4]
  assign Mem1D_8_reset = reset; // @[:@9368.4]
  assign Mem1D_8_io_r_ofs_0 = _T_1801[0]; // @[MemPrimitives.scala 127:28:@10251.4]
  assign Mem1D_8_io_r_backpressure = _T_1801[1]; // @[MemPrimitives.scala 128:32:@10252.4]
  assign Mem1D_8_io_w_ofs_0 = _T_1189[0]; // @[MemPrimitives.scala 94:28:@9644.4]
  assign Mem1D_8_io_w_data_0 = _T_1189[8:1]; // @[MemPrimitives.scala 95:29:@9645.4]
  assign Mem1D_8_io_w_en_0 = _T_1189[9]; // @[MemPrimitives.scala 96:27:@9646.4]
  assign Mem1D_9_clock = clock; // @[:@9383.4]
  assign Mem1D_9_reset = reset; // @[:@9384.4]
  assign Mem1D_9_io_r_ofs_0 = _T_1839[0]; // @[MemPrimitives.scala 127:28:@10291.4]
  assign Mem1D_9_io_r_backpressure = _T_1839[1]; // @[MemPrimitives.scala 128:32:@10292.4]
  assign Mem1D_9_io_w_ofs_0 = _T_1207[0]; // @[MemPrimitives.scala 94:28:@9661.4]
  assign Mem1D_9_io_w_data_0 = _T_1207[8:1]; // @[MemPrimitives.scala 95:29:@9662.4]
  assign Mem1D_9_io_w_en_0 = _T_1207[9]; // @[MemPrimitives.scala 96:27:@9663.4]
  assign Mem1D_10_clock = clock; // @[:@9399.4]
  assign Mem1D_10_reset = reset; // @[:@9400.4]
  assign Mem1D_10_io_r_ofs_0 = _T_1913[0]; // @[MemPrimitives.scala 127:28:@10363.4]
  assign Mem1D_10_io_r_backpressure = _T_1913[1]; // @[MemPrimitives.scala 128:32:@10364.4]
  assign Mem1D_10_io_w_ofs_0 = _T_1225[0]; // @[MemPrimitives.scala 94:28:@9678.4]
  assign Mem1D_10_io_w_data_0 = _T_1225[8:1]; // @[MemPrimitives.scala 95:29:@9679.4]
  assign Mem1D_10_io_w_en_0 = _T_1225[9]; // @[MemPrimitives.scala 96:27:@9680.4]
  assign Mem1D_11_clock = clock; // @[:@9415.4]
  assign Mem1D_11_reset = reset; // @[:@9416.4]
  assign Mem1D_11_io_r_ofs_0 = _T_1987[0]; // @[MemPrimitives.scala 127:28:@10435.4]
  assign Mem1D_11_io_r_backpressure = _T_1987[1]; // @[MemPrimitives.scala 128:32:@10436.4]
  assign Mem1D_11_io_w_ofs_0 = _T_1243[0]; // @[MemPrimitives.scala 94:28:@9695.4]
  assign Mem1D_11_io_w_data_0 = _T_1243[8:1]; // @[MemPrimitives.scala 95:29:@9696.4]
  assign Mem1D_11_io_w_en_0 = _T_1243[9]; // @[MemPrimitives.scala 96:27:@9697.4]
  assign Mem1D_12_clock = clock; // @[:@9431.4]
  assign Mem1D_12_reset = reset; // @[:@9432.4]
  assign Mem1D_12_io_r_ofs_0 = _T_2025[0]; // @[MemPrimitives.scala 127:28:@10475.4]
  assign Mem1D_12_io_r_backpressure = _T_2025[1]; // @[MemPrimitives.scala 128:32:@10476.4]
  assign Mem1D_12_io_w_ofs_0 = _T_1261[0]; // @[MemPrimitives.scala 94:28:@9712.4]
  assign Mem1D_12_io_w_data_0 = _T_1261[8:1]; // @[MemPrimitives.scala 95:29:@9713.4]
  assign Mem1D_12_io_w_en_0 = _T_1261[9]; // @[MemPrimitives.scala 96:27:@9714.4]
  assign Mem1D_13_clock = clock; // @[:@9447.4]
  assign Mem1D_13_reset = reset; // @[:@9448.4]
  assign Mem1D_13_io_r_ofs_0 = _T_2063[0]; // @[MemPrimitives.scala 127:28:@10515.4]
  assign Mem1D_13_io_r_backpressure = _T_2063[1]; // @[MemPrimitives.scala 128:32:@10516.4]
  assign Mem1D_13_io_w_ofs_0 = _T_1279[0]; // @[MemPrimitives.scala 94:28:@9729.4]
  assign Mem1D_13_io_w_data_0 = _T_1279[8:1]; // @[MemPrimitives.scala 95:29:@9730.4]
  assign Mem1D_13_io_w_en_0 = _T_1279[9]; // @[MemPrimitives.scala 96:27:@9731.4]
  assign Mem1D_14_clock = clock; // @[:@9463.4]
  assign Mem1D_14_reset = reset; // @[:@9464.4]
  assign Mem1D_14_io_r_ofs_0 = _T_2137[0]; // @[MemPrimitives.scala 127:28:@10587.4]
  assign Mem1D_14_io_r_backpressure = _T_2137[1]; // @[MemPrimitives.scala 128:32:@10588.4]
  assign Mem1D_14_io_w_ofs_0 = _T_1297[0]; // @[MemPrimitives.scala 94:28:@9746.4]
  assign Mem1D_14_io_w_data_0 = _T_1297[8:1]; // @[MemPrimitives.scala 95:29:@9747.4]
  assign Mem1D_14_io_w_en_0 = _T_1297[9]; // @[MemPrimitives.scala 96:27:@9748.4]
  assign Mem1D_15_clock = clock; // @[:@9479.4]
  assign Mem1D_15_reset = reset; // @[:@9480.4]
  assign Mem1D_15_io_r_ofs_0 = _T_2211[0]; // @[MemPrimitives.scala 127:28:@10659.4]
  assign Mem1D_15_io_r_backpressure = _T_2211[1]; // @[MemPrimitives.scala 128:32:@10660.4]
  assign Mem1D_15_io_w_ofs_0 = _T_1315[0]; // @[MemPrimitives.scala 94:28:@9763.4]
  assign Mem1D_15_io_w_data_0 = _T_1315[8:1]; // @[MemPrimitives.scala 95:29:@9764.4]
  assign Mem1D_15_io_w_en_0 = _T_1315[9]; // @[MemPrimitives.scala 96:27:@9765.4]
  assign StickySelects_clock = clock; // @[:@9779.4]
  assign StickySelects_reset = reset; // @[:@9780.4]
  assign StickySelects_io_ins_0 = io_rPort_4_en_0 & _T_1320; // @[MemPrimitives.scala 122:60:@9781.4]
  assign StickySelects_io_ins_1 = io_rPort_12_en_0 & _T_1325; // @[MemPrimitives.scala 122:60:@9782.4]
  assign StickySelects_io_ins_2 = io_rPort_16_en_0 & _T_1330; // @[MemPrimitives.scala 122:60:@9783.4]
  assign StickySelects_io_ins_3 = io_rPort_20_en_0 & _T_1335; // @[MemPrimitives.scala 122:60:@9784.4]
  assign StickySelects_1_clock = clock; // @[:@9819.4]
  assign StickySelects_1_reset = reset; // @[:@9820.4]
  assign StickySelects_1_io_ins_0 = io_rPort_5_en_0 & _T_1358; // @[MemPrimitives.scala 122:60:@9821.4]
  assign StickySelects_1_io_ins_1 = io_rPort_10_en_0 & _T_1363; // @[MemPrimitives.scala 122:60:@9822.4]
  assign StickySelects_1_io_ins_2 = io_rPort_13_en_0 & _T_1368; // @[MemPrimitives.scala 122:60:@9823.4]
  assign StickySelects_1_io_ins_3 = io_rPort_23_en_0 & _T_1373; // @[MemPrimitives.scala 122:60:@9824.4]
  assign StickySelects_2_clock = clock; // @[:@9871.4]
  assign StickySelects_2_reset = reset; // @[:@9872.4]
  assign StickySelects_2_io_ins_0 = io_rPort_1_en_0 & _T_1396; // @[MemPrimitives.scala 122:60:@9873.4]
  assign StickySelects_2_io_ins_1 = io_rPort_7_en_0 & _T_1401; // @[MemPrimitives.scala 122:60:@9874.4]
  assign StickySelects_2_io_ins_2 = io_rPort_8_en_0 & _T_1406; // @[MemPrimitives.scala 122:60:@9875.4]
  assign StickySelects_2_io_ins_3 = io_rPort_9_en_0 & _T_1411; // @[MemPrimitives.scala 122:60:@9876.4]
  assign StickySelects_2_io_ins_4 = io_rPort_14_en_0 & _T_1416; // @[MemPrimitives.scala 122:60:@9877.4]
  assign StickySelects_2_io_ins_5 = io_rPort_15_en_0 & _T_1421; // @[MemPrimitives.scala 122:60:@9878.4]
  assign StickySelects_2_io_ins_6 = io_rPort_19_en_0 & _T_1426; // @[MemPrimitives.scala 122:60:@9879.4]
  assign StickySelects_2_io_ins_7 = io_rPort_22_en_0 & _T_1431; // @[MemPrimitives.scala 122:60:@9880.4]
  assign StickySelects_3_clock = clock; // @[:@9943.4]
  assign StickySelects_3_reset = reset; // @[:@9944.4]
  assign StickySelects_3_io_ins_0 = io_rPort_0_en_0 & _T_1470; // @[MemPrimitives.scala 122:60:@9945.4]
  assign StickySelects_3_io_ins_1 = io_rPort_2_en_0 & _T_1475; // @[MemPrimitives.scala 122:60:@9946.4]
  assign StickySelects_3_io_ins_2 = io_rPort_3_en_0 & _T_1480; // @[MemPrimitives.scala 122:60:@9947.4]
  assign StickySelects_3_io_ins_3 = io_rPort_6_en_0 & _T_1485; // @[MemPrimitives.scala 122:60:@9948.4]
  assign StickySelects_3_io_ins_4 = io_rPort_11_en_0 & _T_1490; // @[MemPrimitives.scala 122:60:@9949.4]
  assign StickySelects_3_io_ins_5 = io_rPort_17_en_0 & _T_1495; // @[MemPrimitives.scala 122:60:@9950.4]
  assign StickySelects_3_io_ins_6 = io_rPort_18_en_0 & _T_1500; // @[MemPrimitives.scala 122:60:@9951.4]
  assign StickySelects_3_io_ins_7 = io_rPort_21_en_0 & _T_1505; // @[MemPrimitives.scala 122:60:@9952.4]
  assign StickySelects_4_clock = clock; // @[:@10003.4]
  assign StickySelects_4_reset = reset; // @[:@10004.4]
  assign StickySelects_4_io_ins_0 = io_rPort_4_en_0 & _T_1544; // @[MemPrimitives.scala 122:60:@10005.4]
  assign StickySelects_4_io_ins_1 = io_rPort_12_en_0 & _T_1549; // @[MemPrimitives.scala 122:60:@10006.4]
  assign StickySelects_4_io_ins_2 = io_rPort_16_en_0 & _T_1554; // @[MemPrimitives.scala 122:60:@10007.4]
  assign StickySelects_4_io_ins_3 = io_rPort_20_en_0 & _T_1559; // @[MemPrimitives.scala 122:60:@10008.4]
  assign StickySelects_5_clock = clock; // @[:@10043.4]
  assign StickySelects_5_reset = reset; // @[:@10044.4]
  assign StickySelects_5_io_ins_0 = io_rPort_5_en_0 & _T_1582; // @[MemPrimitives.scala 122:60:@10045.4]
  assign StickySelects_5_io_ins_1 = io_rPort_10_en_0 & _T_1587; // @[MemPrimitives.scala 122:60:@10046.4]
  assign StickySelects_5_io_ins_2 = io_rPort_13_en_0 & _T_1592; // @[MemPrimitives.scala 122:60:@10047.4]
  assign StickySelects_5_io_ins_3 = io_rPort_23_en_0 & _T_1597; // @[MemPrimitives.scala 122:60:@10048.4]
  assign StickySelects_6_clock = clock; // @[:@10095.4]
  assign StickySelects_6_reset = reset; // @[:@10096.4]
  assign StickySelects_6_io_ins_0 = io_rPort_1_en_0 & _T_1620; // @[MemPrimitives.scala 122:60:@10097.4]
  assign StickySelects_6_io_ins_1 = io_rPort_7_en_0 & _T_1625; // @[MemPrimitives.scala 122:60:@10098.4]
  assign StickySelects_6_io_ins_2 = io_rPort_8_en_0 & _T_1630; // @[MemPrimitives.scala 122:60:@10099.4]
  assign StickySelects_6_io_ins_3 = io_rPort_9_en_0 & _T_1635; // @[MemPrimitives.scala 122:60:@10100.4]
  assign StickySelects_6_io_ins_4 = io_rPort_14_en_0 & _T_1640; // @[MemPrimitives.scala 122:60:@10101.4]
  assign StickySelects_6_io_ins_5 = io_rPort_15_en_0 & _T_1645; // @[MemPrimitives.scala 122:60:@10102.4]
  assign StickySelects_6_io_ins_6 = io_rPort_19_en_0 & _T_1650; // @[MemPrimitives.scala 122:60:@10103.4]
  assign StickySelects_6_io_ins_7 = io_rPort_22_en_0 & _T_1655; // @[MemPrimitives.scala 122:60:@10104.4]
  assign StickySelects_7_clock = clock; // @[:@10167.4]
  assign StickySelects_7_reset = reset; // @[:@10168.4]
  assign StickySelects_7_io_ins_0 = io_rPort_0_en_0 & _T_1694; // @[MemPrimitives.scala 122:60:@10169.4]
  assign StickySelects_7_io_ins_1 = io_rPort_2_en_0 & _T_1699; // @[MemPrimitives.scala 122:60:@10170.4]
  assign StickySelects_7_io_ins_2 = io_rPort_3_en_0 & _T_1704; // @[MemPrimitives.scala 122:60:@10171.4]
  assign StickySelects_7_io_ins_3 = io_rPort_6_en_0 & _T_1709; // @[MemPrimitives.scala 122:60:@10172.4]
  assign StickySelects_7_io_ins_4 = io_rPort_11_en_0 & _T_1714; // @[MemPrimitives.scala 122:60:@10173.4]
  assign StickySelects_7_io_ins_5 = io_rPort_17_en_0 & _T_1719; // @[MemPrimitives.scala 122:60:@10174.4]
  assign StickySelects_7_io_ins_6 = io_rPort_18_en_0 & _T_1724; // @[MemPrimitives.scala 122:60:@10175.4]
  assign StickySelects_7_io_ins_7 = io_rPort_21_en_0 & _T_1729; // @[MemPrimitives.scala 122:60:@10176.4]
  assign StickySelects_8_clock = clock; // @[:@10227.4]
  assign StickySelects_8_reset = reset; // @[:@10228.4]
  assign StickySelects_8_io_ins_0 = io_rPort_4_en_0 & _T_1768; // @[MemPrimitives.scala 122:60:@10229.4]
  assign StickySelects_8_io_ins_1 = io_rPort_12_en_0 & _T_1773; // @[MemPrimitives.scala 122:60:@10230.4]
  assign StickySelects_8_io_ins_2 = io_rPort_16_en_0 & _T_1778; // @[MemPrimitives.scala 122:60:@10231.4]
  assign StickySelects_8_io_ins_3 = io_rPort_20_en_0 & _T_1783; // @[MemPrimitives.scala 122:60:@10232.4]
  assign StickySelects_9_clock = clock; // @[:@10267.4]
  assign StickySelects_9_reset = reset; // @[:@10268.4]
  assign StickySelects_9_io_ins_0 = io_rPort_5_en_0 & _T_1806; // @[MemPrimitives.scala 122:60:@10269.4]
  assign StickySelects_9_io_ins_1 = io_rPort_10_en_0 & _T_1811; // @[MemPrimitives.scala 122:60:@10270.4]
  assign StickySelects_9_io_ins_2 = io_rPort_13_en_0 & _T_1816; // @[MemPrimitives.scala 122:60:@10271.4]
  assign StickySelects_9_io_ins_3 = io_rPort_23_en_0 & _T_1821; // @[MemPrimitives.scala 122:60:@10272.4]
  assign StickySelects_10_clock = clock; // @[:@10319.4]
  assign StickySelects_10_reset = reset; // @[:@10320.4]
  assign StickySelects_10_io_ins_0 = io_rPort_1_en_0 & _T_1844; // @[MemPrimitives.scala 122:60:@10321.4]
  assign StickySelects_10_io_ins_1 = io_rPort_7_en_0 & _T_1849; // @[MemPrimitives.scala 122:60:@10322.4]
  assign StickySelects_10_io_ins_2 = io_rPort_8_en_0 & _T_1854; // @[MemPrimitives.scala 122:60:@10323.4]
  assign StickySelects_10_io_ins_3 = io_rPort_9_en_0 & _T_1859; // @[MemPrimitives.scala 122:60:@10324.4]
  assign StickySelects_10_io_ins_4 = io_rPort_14_en_0 & _T_1864; // @[MemPrimitives.scala 122:60:@10325.4]
  assign StickySelects_10_io_ins_5 = io_rPort_15_en_0 & _T_1869; // @[MemPrimitives.scala 122:60:@10326.4]
  assign StickySelects_10_io_ins_6 = io_rPort_19_en_0 & _T_1874; // @[MemPrimitives.scala 122:60:@10327.4]
  assign StickySelects_10_io_ins_7 = io_rPort_22_en_0 & _T_1879; // @[MemPrimitives.scala 122:60:@10328.4]
  assign StickySelects_11_clock = clock; // @[:@10391.4]
  assign StickySelects_11_reset = reset; // @[:@10392.4]
  assign StickySelects_11_io_ins_0 = io_rPort_0_en_0 & _T_1918; // @[MemPrimitives.scala 122:60:@10393.4]
  assign StickySelects_11_io_ins_1 = io_rPort_2_en_0 & _T_1923; // @[MemPrimitives.scala 122:60:@10394.4]
  assign StickySelects_11_io_ins_2 = io_rPort_3_en_0 & _T_1928; // @[MemPrimitives.scala 122:60:@10395.4]
  assign StickySelects_11_io_ins_3 = io_rPort_6_en_0 & _T_1933; // @[MemPrimitives.scala 122:60:@10396.4]
  assign StickySelects_11_io_ins_4 = io_rPort_11_en_0 & _T_1938; // @[MemPrimitives.scala 122:60:@10397.4]
  assign StickySelects_11_io_ins_5 = io_rPort_17_en_0 & _T_1943; // @[MemPrimitives.scala 122:60:@10398.4]
  assign StickySelects_11_io_ins_6 = io_rPort_18_en_0 & _T_1948; // @[MemPrimitives.scala 122:60:@10399.4]
  assign StickySelects_11_io_ins_7 = io_rPort_21_en_0 & _T_1953; // @[MemPrimitives.scala 122:60:@10400.4]
  assign StickySelects_12_clock = clock; // @[:@10451.4]
  assign StickySelects_12_reset = reset; // @[:@10452.4]
  assign StickySelects_12_io_ins_0 = io_rPort_4_en_0 & _T_1992; // @[MemPrimitives.scala 122:60:@10453.4]
  assign StickySelects_12_io_ins_1 = io_rPort_12_en_0 & _T_1997; // @[MemPrimitives.scala 122:60:@10454.4]
  assign StickySelects_12_io_ins_2 = io_rPort_16_en_0 & _T_2002; // @[MemPrimitives.scala 122:60:@10455.4]
  assign StickySelects_12_io_ins_3 = io_rPort_20_en_0 & _T_2007; // @[MemPrimitives.scala 122:60:@10456.4]
  assign StickySelects_13_clock = clock; // @[:@10491.4]
  assign StickySelects_13_reset = reset; // @[:@10492.4]
  assign StickySelects_13_io_ins_0 = io_rPort_5_en_0 & _T_2030; // @[MemPrimitives.scala 122:60:@10493.4]
  assign StickySelects_13_io_ins_1 = io_rPort_10_en_0 & _T_2035; // @[MemPrimitives.scala 122:60:@10494.4]
  assign StickySelects_13_io_ins_2 = io_rPort_13_en_0 & _T_2040; // @[MemPrimitives.scala 122:60:@10495.4]
  assign StickySelects_13_io_ins_3 = io_rPort_23_en_0 & _T_2045; // @[MemPrimitives.scala 122:60:@10496.4]
  assign StickySelects_14_clock = clock; // @[:@10543.4]
  assign StickySelects_14_reset = reset; // @[:@10544.4]
  assign StickySelects_14_io_ins_0 = io_rPort_1_en_0 & _T_2068; // @[MemPrimitives.scala 122:60:@10545.4]
  assign StickySelects_14_io_ins_1 = io_rPort_7_en_0 & _T_2073; // @[MemPrimitives.scala 122:60:@10546.4]
  assign StickySelects_14_io_ins_2 = io_rPort_8_en_0 & _T_2078; // @[MemPrimitives.scala 122:60:@10547.4]
  assign StickySelects_14_io_ins_3 = io_rPort_9_en_0 & _T_2083; // @[MemPrimitives.scala 122:60:@10548.4]
  assign StickySelects_14_io_ins_4 = io_rPort_14_en_0 & _T_2088; // @[MemPrimitives.scala 122:60:@10549.4]
  assign StickySelects_14_io_ins_5 = io_rPort_15_en_0 & _T_2093; // @[MemPrimitives.scala 122:60:@10550.4]
  assign StickySelects_14_io_ins_6 = io_rPort_19_en_0 & _T_2098; // @[MemPrimitives.scala 122:60:@10551.4]
  assign StickySelects_14_io_ins_7 = io_rPort_22_en_0 & _T_2103; // @[MemPrimitives.scala 122:60:@10552.4]
  assign StickySelects_15_clock = clock; // @[:@10615.4]
  assign StickySelects_15_reset = reset; // @[:@10616.4]
  assign StickySelects_15_io_ins_0 = io_rPort_0_en_0 & _T_2142; // @[MemPrimitives.scala 122:60:@10617.4]
  assign StickySelects_15_io_ins_1 = io_rPort_2_en_0 & _T_2147; // @[MemPrimitives.scala 122:60:@10618.4]
  assign StickySelects_15_io_ins_2 = io_rPort_3_en_0 & _T_2152; // @[MemPrimitives.scala 122:60:@10619.4]
  assign StickySelects_15_io_ins_3 = io_rPort_6_en_0 & _T_2157; // @[MemPrimitives.scala 122:60:@10620.4]
  assign StickySelects_15_io_ins_4 = io_rPort_11_en_0 & _T_2162; // @[MemPrimitives.scala 122:60:@10621.4]
  assign StickySelects_15_io_ins_5 = io_rPort_17_en_0 & _T_2167; // @[MemPrimitives.scala 122:60:@10622.4]
  assign StickySelects_15_io_ins_6 = io_rPort_18_en_0 & _T_2172; // @[MemPrimitives.scala 122:60:@10623.4]
  assign StickySelects_15_io_ins_7 = io_rPort_21_en_0 & _T_2177; // @[MemPrimitives.scala 122:60:@10624.4]
  assign RetimeWrapper_clock = clock; // @[:@10676.4]
  assign RetimeWrapper_reset = reset; // @[:@10677.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@10679.4]
  assign RetimeWrapper_io_in = _T_1470 & io_rPort_0_en_0; // @[package.scala 94:16:@10678.4]
  assign RetimeWrapper_1_clock = clock; // @[:@10684.4]
  assign RetimeWrapper_1_reset = reset; // @[:@10685.4]
  assign RetimeWrapper_1_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@10687.4]
  assign RetimeWrapper_1_io_in = _T_1694 & io_rPort_0_en_0; // @[package.scala 94:16:@10686.4]
  assign RetimeWrapper_2_clock = clock; // @[:@10692.4]
  assign RetimeWrapper_2_reset = reset; // @[:@10693.4]
  assign RetimeWrapper_2_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@10695.4]
  assign RetimeWrapper_2_io_in = _T_1918 & io_rPort_0_en_0; // @[package.scala 94:16:@10694.4]
  assign RetimeWrapper_3_clock = clock; // @[:@10700.4]
  assign RetimeWrapper_3_reset = reset; // @[:@10701.4]
  assign RetimeWrapper_3_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@10703.4]
  assign RetimeWrapper_3_io_in = _T_2142 & io_rPort_0_en_0; // @[package.scala 94:16:@10702.4]
  assign RetimeWrapper_4_clock = clock; // @[:@10724.4]
  assign RetimeWrapper_4_reset = reset; // @[:@10725.4]
  assign RetimeWrapper_4_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@10727.4]
  assign RetimeWrapper_4_io_in = _T_1396 & io_rPort_1_en_0; // @[package.scala 94:16:@10726.4]
  assign RetimeWrapper_5_clock = clock; // @[:@10732.4]
  assign RetimeWrapper_5_reset = reset; // @[:@10733.4]
  assign RetimeWrapper_5_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@10735.4]
  assign RetimeWrapper_5_io_in = _T_1620 & io_rPort_1_en_0; // @[package.scala 94:16:@10734.4]
  assign RetimeWrapper_6_clock = clock; // @[:@10740.4]
  assign RetimeWrapper_6_reset = reset; // @[:@10741.4]
  assign RetimeWrapper_6_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@10743.4]
  assign RetimeWrapper_6_io_in = _T_1844 & io_rPort_1_en_0; // @[package.scala 94:16:@10742.4]
  assign RetimeWrapper_7_clock = clock; // @[:@10748.4]
  assign RetimeWrapper_7_reset = reset; // @[:@10749.4]
  assign RetimeWrapper_7_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@10751.4]
  assign RetimeWrapper_7_io_in = _T_2068 & io_rPort_1_en_0; // @[package.scala 94:16:@10750.4]
  assign RetimeWrapper_8_clock = clock; // @[:@10772.4]
  assign RetimeWrapper_8_reset = reset; // @[:@10773.4]
  assign RetimeWrapper_8_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@10775.4]
  assign RetimeWrapper_8_io_in = _T_1475 & io_rPort_2_en_0; // @[package.scala 94:16:@10774.4]
  assign RetimeWrapper_9_clock = clock; // @[:@10780.4]
  assign RetimeWrapper_9_reset = reset; // @[:@10781.4]
  assign RetimeWrapper_9_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@10783.4]
  assign RetimeWrapper_9_io_in = _T_1699 & io_rPort_2_en_0; // @[package.scala 94:16:@10782.4]
  assign RetimeWrapper_10_clock = clock; // @[:@10788.4]
  assign RetimeWrapper_10_reset = reset; // @[:@10789.4]
  assign RetimeWrapper_10_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@10791.4]
  assign RetimeWrapper_10_io_in = _T_1923 & io_rPort_2_en_0; // @[package.scala 94:16:@10790.4]
  assign RetimeWrapper_11_clock = clock; // @[:@10796.4]
  assign RetimeWrapper_11_reset = reset; // @[:@10797.4]
  assign RetimeWrapper_11_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@10799.4]
  assign RetimeWrapper_11_io_in = _T_2147 & io_rPort_2_en_0; // @[package.scala 94:16:@10798.4]
  assign RetimeWrapper_12_clock = clock; // @[:@10820.4]
  assign RetimeWrapper_12_reset = reset; // @[:@10821.4]
  assign RetimeWrapper_12_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@10823.4]
  assign RetimeWrapper_12_io_in = _T_1480 & io_rPort_3_en_0; // @[package.scala 94:16:@10822.4]
  assign RetimeWrapper_13_clock = clock; // @[:@10828.4]
  assign RetimeWrapper_13_reset = reset; // @[:@10829.4]
  assign RetimeWrapper_13_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@10831.4]
  assign RetimeWrapper_13_io_in = _T_1704 & io_rPort_3_en_0; // @[package.scala 94:16:@10830.4]
  assign RetimeWrapper_14_clock = clock; // @[:@10836.4]
  assign RetimeWrapper_14_reset = reset; // @[:@10837.4]
  assign RetimeWrapper_14_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@10839.4]
  assign RetimeWrapper_14_io_in = _T_1928 & io_rPort_3_en_0; // @[package.scala 94:16:@10838.4]
  assign RetimeWrapper_15_clock = clock; // @[:@10844.4]
  assign RetimeWrapper_15_reset = reset; // @[:@10845.4]
  assign RetimeWrapper_15_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@10847.4]
  assign RetimeWrapper_15_io_in = _T_2152 & io_rPort_3_en_0; // @[package.scala 94:16:@10846.4]
  assign RetimeWrapper_16_clock = clock; // @[:@10868.4]
  assign RetimeWrapper_16_reset = reset; // @[:@10869.4]
  assign RetimeWrapper_16_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@10871.4]
  assign RetimeWrapper_16_io_in = _T_1320 & io_rPort_4_en_0; // @[package.scala 94:16:@10870.4]
  assign RetimeWrapper_17_clock = clock; // @[:@10876.4]
  assign RetimeWrapper_17_reset = reset; // @[:@10877.4]
  assign RetimeWrapper_17_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@10879.4]
  assign RetimeWrapper_17_io_in = _T_1544 & io_rPort_4_en_0; // @[package.scala 94:16:@10878.4]
  assign RetimeWrapper_18_clock = clock; // @[:@10884.4]
  assign RetimeWrapper_18_reset = reset; // @[:@10885.4]
  assign RetimeWrapper_18_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@10887.4]
  assign RetimeWrapper_18_io_in = _T_1768 & io_rPort_4_en_0; // @[package.scala 94:16:@10886.4]
  assign RetimeWrapper_19_clock = clock; // @[:@10892.4]
  assign RetimeWrapper_19_reset = reset; // @[:@10893.4]
  assign RetimeWrapper_19_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@10895.4]
  assign RetimeWrapper_19_io_in = _T_1992 & io_rPort_4_en_0; // @[package.scala 94:16:@10894.4]
  assign RetimeWrapper_20_clock = clock; // @[:@10916.4]
  assign RetimeWrapper_20_reset = reset; // @[:@10917.4]
  assign RetimeWrapper_20_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@10919.4]
  assign RetimeWrapper_20_io_in = _T_1358 & io_rPort_5_en_0; // @[package.scala 94:16:@10918.4]
  assign RetimeWrapper_21_clock = clock; // @[:@10924.4]
  assign RetimeWrapper_21_reset = reset; // @[:@10925.4]
  assign RetimeWrapper_21_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@10927.4]
  assign RetimeWrapper_21_io_in = _T_1582 & io_rPort_5_en_0; // @[package.scala 94:16:@10926.4]
  assign RetimeWrapper_22_clock = clock; // @[:@10932.4]
  assign RetimeWrapper_22_reset = reset; // @[:@10933.4]
  assign RetimeWrapper_22_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@10935.4]
  assign RetimeWrapper_22_io_in = _T_1806 & io_rPort_5_en_0; // @[package.scala 94:16:@10934.4]
  assign RetimeWrapper_23_clock = clock; // @[:@10940.4]
  assign RetimeWrapper_23_reset = reset; // @[:@10941.4]
  assign RetimeWrapper_23_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@10943.4]
  assign RetimeWrapper_23_io_in = _T_2030 & io_rPort_5_en_0; // @[package.scala 94:16:@10942.4]
  assign RetimeWrapper_24_clock = clock; // @[:@10964.4]
  assign RetimeWrapper_24_reset = reset; // @[:@10965.4]
  assign RetimeWrapper_24_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@10967.4]
  assign RetimeWrapper_24_io_in = _T_1485 & io_rPort_6_en_0; // @[package.scala 94:16:@10966.4]
  assign RetimeWrapper_25_clock = clock; // @[:@10972.4]
  assign RetimeWrapper_25_reset = reset; // @[:@10973.4]
  assign RetimeWrapper_25_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@10975.4]
  assign RetimeWrapper_25_io_in = _T_1709 & io_rPort_6_en_0; // @[package.scala 94:16:@10974.4]
  assign RetimeWrapper_26_clock = clock; // @[:@10980.4]
  assign RetimeWrapper_26_reset = reset; // @[:@10981.4]
  assign RetimeWrapper_26_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@10983.4]
  assign RetimeWrapper_26_io_in = _T_1933 & io_rPort_6_en_0; // @[package.scala 94:16:@10982.4]
  assign RetimeWrapper_27_clock = clock; // @[:@10988.4]
  assign RetimeWrapper_27_reset = reset; // @[:@10989.4]
  assign RetimeWrapper_27_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@10991.4]
  assign RetimeWrapper_27_io_in = _T_2157 & io_rPort_6_en_0; // @[package.scala 94:16:@10990.4]
  assign RetimeWrapper_28_clock = clock; // @[:@11012.4]
  assign RetimeWrapper_28_reset = reset; // @[:@11013.4]
  assign RetimeWrapper_28_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@11015.4]
  assign RetimeWrapper_28_io_in = _T_1401 & io_rPort_7_en_0; // @[package.scala 94:16:@11014.4]
  assign RetimeWrapper_29_clock = clock; // @[:@11020.4]
  assign RetimeWrapper_29_reset = reset; // @[:@11021.4]
  assign RetimeWrapper_29_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@11023.4]
  assign RetimeWrapper_29_io_in = _T_1625 & io_rPort_7_en_0; // @[package.scala 94:16:@11022.4]
  assign RetimeWrapper_30_clock = clock; // @[:@11028.4]
  assign RetimeWrapper_30_reset = reset; // @[:@11029.4]
  assign RetimeWrapper_30_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@11031.4]
  assign RetimeWrapper_30_io_in = _T_1849 & io_rPort_7_en_0; // @[package.scala 94:16:@11030.4]
  assign RetimeWrapper_31_clock = clock; // @[:@11036.4]
  assign RetimeWrapper_31_reset = reset; // @[:@11037.4]
  assign RetimeWrapper_31_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@11039.4]
  assign RetimeWrapper_31_io_in = _T_2073 & io_rPort_7_en_0; // @[package.scala 94:16:@11038.4]
  assign RetimeWrapper_32_clock = clock; // @[:@11060.4]
  assign RetimeWrapper_32_reset = reset; // @[:@11061.4]
  assign RetimeWrapper_32_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@11063.4]
  assign RetimeWrapper_32_io_in = _T_1406 & io_rPort_8_en_0; // @[package.scala 94:16:@11062.4]
  assign RetimeWrapper_33_clock = clock; // @[:@11068.4]
  assign RetimeWrapper_33_reset = reset; // @[:@11069.4]
  assign RetimeWrapper_33_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@11071.4]
  assign RetimeWrapper_33_io_in = _T_1630 & io_rPort_8_en_0; // @[package.scala 94:16:@11070.4]
  assign RetimeWrapper_34_clock = clock; // @[:@11076.4]
  assign RetimeWrapper_34_reset = reset; // @[:@11077.4]
  assign RetimeWrapper_34_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@11079.4]
  assign RetimeWrapper_34_io_in = _T_1854 & io_rPort_8_en_0; // @[package.scala 94:16:@11078.4]
  assign RetimeWrapper_35_clock = clock; // @[:@11084.4]
  assign RetimeWrapper_35_reset = reset; // @[:@11085.4]
  assign RetimeWrapper_35_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@11087.4]
  assign RetimeWrapper_35_io_in = _T_2078 & io_rPort_8_en_0; // @[package.scala 94:16:@11086.4]
  assign RetimeWrapper_36_clock = clock; // @[:@11108.4]
  assign RetimeWrapper_36_reset = reset; // @[:@11109.4]
  assign RetimeWrapper_36_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@11111.4]
  assign RetimeWrapper_36_io_in = _T_1411 & io_rPort_9_en_0; // @[package.scala 94:16:@11110.4]
  assign RetimeWrapper_37_clock = clock; // @[:@11116.4]
  assign RetimeWrapper_37_reset = reset; // @[:@11117.4]
  assign RetimeWrapper_37_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@11119.4]
  assign RetimeWrapper_37_io_in = _T_1635 & io_rPort_9_en_0; // @[package.scala 94:16:@11118.4]
  assign RetimeWrapper_38_clock = clock; // @[:@11124.4]
  assign RetimeWrapper_38_reset = reset; // @[:@11125.4]
  assign RetimeWrapper_38_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@11127.4]
  assign RetimeWrapper_38_io_in = _T_1859 & io_rPort_9_en_0; // @[package.scala 94:16:@11126.4]
  assign RetimeWrapper_39_clock = clock; // @[:@11132.4]
  assign RetimeWrapper_39_reset = reset; // @[:@11133.4]
  assign RetimeWrapper_39_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@11135.4]
  assign RetimeWrapper_39_io_in = _T_2083 & io_rPort_9_en_0; // @[package.scala 94:16:@11134.4]
  assign RetimeWrapper_40_clock = clock; // @[:@11156.4]
  assign RetimeWrapper_40_reset = reset; // @[:@11157.4]
  assign RetimeWrapper_40_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@11159.4]
  assign RetimeWrapper_40_io_in = _T_1363 & io_rPort_10_en_0; // @[package.scala 94:16:@11158.4]
  assign RetimeWrapper_41_clock = clock; // @[:@11164.4]
  assign RetimeWrapper_41_reset = reset; // @[:@11165.4]
  assign RetimeWrapper_41_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@11167.4]
  assign RetimeWrapper_41_io_in = _T_1587 & io_rPort_10_en_0; // @[package.scala 94:16:@11166.4]
  assign RetimeWrapper_42_clock = clock; // @[:@11172.4]
  assign RetimeWrapper_42_reset = reset; // @[:@11173.4]
  assign RetimeWrapper_42_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@11175.4]
  assign RetimeWrapper_42_io_in = _T_1811 & io_rPort_10_en_0; // @[package.scala 94:16:@11174.4]
  assign RetimeWrapper_43_clock = clock; // @[:@11180.4]
  assign RetimeWrapper_43_reset = reset; // @[:@11181.4]
  assign RetimeWrapper_43_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@11183.4]
  assign RetimeWrapper_43_io_in = _T_2035 & io_rPort_10_en_0; // @[package.scala 94:16:@11182.4]
  assign RetimeWrapper_44_clock = clock; // @[:@11204.4]
  assign RetimeWrapper_44_reset = reset; // @[:@11205.4]
  assign RetimeWrapper_44_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@11207.4]
  assign RetimeWrapper_44_io_in = _T_1490 & io_rPort_11_en_0; // @[package.scala 94:16:@11206.4]
  assign RetimeWrapper_45_clock = clock; // @[:@11212.4]
  assign RetimeWrapper_45_reset = reset; // @[:@11213.4]
  assign RetimeWrapper_45_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@11215.4]
  assign RetimeWrapper_45_io_in = _T_1714 & io_rPort_11_en_0; // @[package.scala 94:16:@11214.4]
  assign RetimeWrapper_46_clock = clock; // @[:@11220.4]
  assign RetimeWrapper_46_reset = reset; // @[:@11221.4]
  assign RetimeWrapper_46_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@11223.4]
  assign RetimeWrapper_46_io_in = _T_1938 & io_rPort_11_en_0; // @[package.scala 94:16:@11222.4]
  assign RetimeWrapper_47_clock = clock; // @[:@11228.4]
  assign RetimeWrapper_47_reset = reset; // @[:@11229.4]
  assign RetimeWrapper_47_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@11231.4]
  assign RetimeWrapper_47_io_in = _T_2162 & io_rPort_11_en_0; // @[package.scala 94:16:@11230.4]
  assign RetimeWrapper_48_clock = clock; // @[:@11252.4]
  assign RetimeWrapper_48_reset = reset; // @[:@11253.4]
  assign RetimeWrapper_48_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@11255.4]
  assign RetimeWrapper_48_io_in = _T_1325 & io_rPort_12_en_0; // @[package.scala 94:16:@11254.4]
  assign RetimeWrapper_49_clock = clock; // @[:@11260.4]
  assign RetimeWrapper_49_reset = reset; // @[:@11261.4]
  assign RetimeWrapper_49_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@11263.4]
  assign RetimeWrapper_49_io_in = _T_1549 & io_rPort_12_en_0; // @[package.scala 94:16:@11262.4]
  assign RetimeWrapper_50_clock = clock; // @[:@11268.4]
  assign RetimeWrapper_50_reset = reset; // @[:@11269.4]
  assign RetimeWrapper_50_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@11271.4]
  assign RetimeWrapper_50_io_in = _T_1773 & io_rPort_12_en_0; // @[package.scala 94:16:@11270.4]
  assign RetimeWrapper_51_clock = clock; // @[:@11276.4]
  assign RetimeWrapper_51_reset = reset; // @[:@11277.4]
  assign RetimeWrapper_51_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@11279.4]
  assign RetimeWrapper_51_io_in = _T_1997 & io_rPort_12_en_0; // @[package.scala 94:16:@11278.4]
  assign RetimeWrapper_52_clock = clock; // @[:@11300.4]
  assign RetimeWrapper_52_reset = reset; // @[:@11301.4]
  assign RetimeWrapper_52_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@11303.4]
  assign RetimeWrapper_52_io_in = _T_1368 & io_rPort_13_en_0; // @[package.scala 94:16:@11302.4]
  assign RetimeWrapper_53_clock = clock; // @[:@11308.4]
  assign RetimeWrapper_53_reset = reset; // @[:@11309.4]
  assign RetimeWrapper_53_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@11311.4]
  assign RetimeWrapper_53_io_in = _T_1592 & io_rPort_13_en_0; // @[package.scala 94:16:@11310.4]
  assign RetimeWrapper_54_clock = clock; // @[:@11316.4]
  assign RetimeWrapper_54_reset = reset; // @[:@11317.4]
  assign RetimeWrapper_54_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@11319.4]
  assign RetimeWrapper_54_io_in = _T_1816 & io_rPort_13_en_0; // @[package.scala 94:16:@11318.4]
  assign RetimeWrapper_55_clock = clock; // @[:@11324.4]
  assign RetimeWrapper_55_reset = reset; // @[:@11325.4]
  assign RetimeWrapper_55_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@11327.4]
  assign RetimeWrapper_55_io_in = _T_2040 & io_rPort_13_en_0; // @[package.scala 94:16:@11326.4]
  assign RetimeWrapper_56_clock = clock; // @[:@11348.4]
  assign RetimeWrapper_56_reset = reset; // @[:@11349.4]
  assign RetimeWrapper_56_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@11351.4]
  assign RetimeWrapper_56_io_in = _T_1416 & io_rPort_14_en_0; // @[package.scala 94:16:@11350.4]
  assign RetimeWrapper_57_clock = clock; // @[:@11356.4]
  assign RetimeWrapper_57_reset = reset; // @[:@11357.4]
  assign RetimeWrapper_57_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@11359.4]
  assign RetimeWrapper_57_io_in = _T_1640 & io_rPort_14_en_0; // @[package.scala 94:16:@11358.4]
  assign RetimeWrapper_58_clock = clock; // @[:@11364.4]
  assign RetimeWrapper_58_reset = reset; // @[:@11365.4]
  assign RetimeWrapper_58_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@11367.4]
  assign RetimeWrapper_58_io_in = _T_1864 & io_rPort_14_en_0; // @[package.scala 94:16:@11366.4]
  assign RetimeWrapper_59_clock = clock; // @[:@11372.4]
  assign RetimeWrapper_59_reset = reset; // @[:@11373.4]
  assign RetimeWrapper_59_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@11375.4]
  assign RetimeWrapper_59_io_in = _T_2088 & io_rPort_14_en_0; // @[package.scala 94:16:@11374.4]
  assign RetimeWrapper_60_clock = clock; // @[:@11396.4]
  assign RetimeWrapper_60_reset = reset; // @[:@11397.4]
  assign RetimeWrapper_60_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@11399.4]
  assign RetimeWrapper_60_io_in = _T_1421 & io_rPort_15_en_0; // @[package.scala 94:16:@11398.4]
  assign RetimeWrapper_61_clock = clock; // @[:@11404.4]
  assign RetimeWrapper_61_reset = reset; // @[:@11405.4]
  assign RetimeWrapper_61_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@11407.4]
  assign RetimeWrapper_61_io_in = _T_1645 & io_rPort_15_en_0; // @[package.scala 94:16:@11406.4]
  assign RetimeWrapper_62_clock = clock; // @[:@11412.4]
  assign RetimeWrapper_62_reset = reset; // @[:@11413.4]
  assign RetimeWrapper_62_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@11415.4]
  assign RetimeWrapper_62_io_in = _T_1869 & io_rPort_15_en_0; // @[package.scala 94:16:@11414.4]
  assign RetimeWrapper_63_clock = clock; // @[:@11420.4]
  assign RetimeWrapper_63_reset = reset; // @[:@11421.4]
  assign RetimeWrapper_63_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@11423.4]
  assign RetimeWrapper_63_io_in = _T_2093 & io_rPort_15_en_0; // @[package.scala 94:16:@11422.4]
  assign RetimeWrapper_64_clock = clock; // @[:@11444.4]
  assign RetimeWrapper_64_reset = reset; // @[:@11445.4]
  assign RetimeWrapper_64_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@11447.4]
  assign RetimeWrapper_64_io_in = _T_1330 & io_rPort_16_en_0; // @[package.scala 94:16:@11446.4]
  assign RetimeWrapper_65_clock = clock; // @[:@11452.4]
  assign RetimeWrapper_65_reset = reset; // @[:@11453.4]
  assign RetimeWrapper_65_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@11455.4]
  assign RetimeWrapper_65_io_in = _T_1554 & io_rPort_16_en_0; // @[package.scala 94:16:@11454.4]
  assign RetimeWrapper_66_clock = clock; // @[:@11460.4]
  assign RetimeWrapper_66_reset = reset; // @[:@11461.4]
  assign RetimeWrapper_66_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@11463.4]
  assign RetimeWrapper_66_io_in = _T_1778 & io_rPort_16_en_0; // @[package.scala 94:16:@11462.4]
  assign RetimeWrapper_67_clock = clock; // @[:@11468.4]
  assign RetimeWrapper_67_reset = reset; // @[:@11469.4]
  assign RetimeWrapper_67_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@11471.4]
  assign RetimeWrapper_67_io_in = _T_2002 & io_rPort_16_en_0; // @[package.scala 94:16:@11470.4]
  assign RetimeWrapper_68_clock = clock; // @[:@11492.4]
  assign RetimeWrapper_68_reset = reset; // @[:@11493.4]
  assign RetimeWrapper_68_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@11495.4]
  assign RetimeWrapper_68_io_in = _T_1495 & io_rPort_17_en_0; // @[package.scala 94:16:@11494.4]
  assign RetimeWrapper_69_clock = clock; // @[:@11500.4]
  assign RetimeWrapper_69_reset = reset; // @[:@11501.4]
  assign RetimeWrapper_69_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@11503.4]
  assign RetimeWrapper_69_io_in = _T_1719 & io_rPort_17_en_0; // @[package.scala 94:16:@11502.4]
  assign RetimeWrapper_70_clock = clock; // @[:@11508.4]
  assign RetimeWrapper_70_reset = reset; // @[:@11509.4]
  assign RetimeWrapper_70_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@11511.4]
  assign RetimeWrapper_70_io_in = _T_1943 & io_rPort_17_en_0; // @[package.scala 94:16:@11510.4]
  assign RetimeWrapper_71_clock = clock; // @[:@11516.4]
  assign RetimeWrapper_71_reset = reset; // @[:@11517.4]
  assign RetimeWrapper_71_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@11519.4]
  assign RetimeWrapper_71_io_in = _T_2167 & io_rPort_17_en_0; // @[package.scala 94:16:@11518.4]
  assign RetimeWrapper_72_clock = clock; // @[:@11540.4]
  assign RetimeWrapper_72_reset = reset; // @[:@11541.4]
  assign RetimeWrapper_72_io_flow = io_rPort_18_backpressure; // @[package.scala 95:18:@11543.4]
  assign RetimeWrapper_72_io_in = _T_1500 & io_rPort_18_en_0; // @[package.scala 94:16:@11542.4]
  assign RetimeWrapper_73_clock = clock; // @[:@11548.4]
  assign RetimeWrapper_73_reset = reset; // @[:@11549.4]
  assign RetimeWrapper_73_io_flow = io_rPort_18_backpressure; // @[package.scala 95:18:@11551.4]
  assign RetimeWrapper_73_io_in = _T_1724 & io_rPort_18_en_0; // @[package.scala 94:16:@11550.4]
  assign RetimeWrapper_74_clock = clock; // @[:@11556.4]
  assign RetimeWrapper_74_reset = reset; // @[:@11557.4]
  assign RetimeWrapper_74_io_flow = io_rPort_18_backpressure; // @[package.scala 95:18:@11559.4]
  assign RetimeWrapper_74_io_in = _T_1948 & io_rPort_18_en_0; // @[package.scala 94:16:@11558.4]
  assign RetimeWrapper_75_clock = clock; // @[:@11564.4]
  assign RetimeWrapper_75_reset = reset; // @[:@11565.4]
  assign RetimeWrapper_75_io_flow = io_rPort_18_backpressure; // @[package.scala 95:18:@11567.4]
  assign RetimeWrapper_75_io_in = _T_2172 & io_rPort_18_en_0; // @[package.scala 94:16:@11566.4]
  assign RetimeWrapper_76_clock = clock; // @[:@11588.4]
  assign RetimeWrapper_76_reset = reset; // @[:@11589.4]
  assign RetimeWrapper_76_io_flow = io_rPort_19_backpressure; // @[package.scala 95:18:@11591.4]
  assign RetimeWrapper_76_io_in = _T_1426 & io_rPort_19_en_0; // @[package.scala 94:16:@11590.4]
  assign RetimeWrapper_77_clock = clock; // @[:@11596.4]
  assign RetimeWrapper_77_reset = reset; // @[:@11597.4]
  assign RetimeWrapper_77_io_flow = io_rPort_19_backpressure; // @[package.scala 95:18:@11599.4]
  assign RetimeWrapper_77_io_in = _T_1650 & io_rPort_19_en_0; // @[package.scala 94:16:@11598.4]
  assign RetimeWrapper_78_clock = clock; // @[:@11604.4]
  assign RetimeWrapper_78_reset = reset; // @[:@11605.4]
  assign RetimeWrapper_78_io_flow = io_rPort_19_backpressure; // @[package.scala 95:18:@11607.4]
  assign RetimeWrapper_78_io_in = _T_1874 & io_rPort_19_en_0; // @[package.scala 94:16:@11606.4]
  assign RetimeWrapper_79_clock = clock; // @[:@11612.4]
  assign RetimeWrapper_79_reset = reset; // @[:@11613.4]
  assign RetimeWrapper_79_io_flow = io_rPort_19_backpressure; // @[package.scala 95:18:@11615.4]
  assign RetimeWrapper_79_io_in = _T_2098 & io_rPort_19_en_0; // @[package.scala 94:16:@11614.4]
  assign RetimeWrapper_80_clock = clock; // @[:@11636.4]
  assign RetimeWrapper_80_reset = reset; // @[:@11637.4]
  assign RetimeWrapper_80_io_flow = io_rPort_20_backpressure; // @[package.scala 95:18:@11639.4]
  assign RetimeWrapper_80_io_in = _T_1335 & io_rPort_20_en_0; // @[package.scala 94:16:@11638.4]
  assign RetimeWrapper_81_clock = clock; // @[:@11644.4]
  assign RetimeWrapper_81_reset = reset; // @[:@11645.4]
  assign RetimeWrapper_81_io_flow = io_rPort_20_backpressure; // @[package.scala 95:18:@11647.4]
  assign RetimeWrapper_81_io_in = _T_1559 & io_rPort_20_en_0; // @[package.scala 94:16:@11646.4]
  assign RetimeWrapper_82_clock = clock; // @[:@11652.4]
  assign RetimeWrapper_82_reset = reset; // @[:@11653.4]
  assign RetimeWrapper_82_io_flow = io_rPort_20_backpressure; // @[package.scala 95:18:@11655.4]
  assign RetimeWrapper_82_io_in = _T_1783 & io_rPort_20_en_0; // @[package.scala 94:16:@11654.4]
  assign RetimeWrapper_83_clock = clock; // @[:@11660.4]
  assign RetimeWrapper_83_reset = reset; // @[:@11661.4]
  assign RetimeWrapper_83_io_flow = io_rPort_20_backpressure; // @[package.scala 95:18:@11663.4]
  assign RetimeWrapper_83_io_in = _T_2007 & io_rPort_20_en_0; // @[package.scala 94:16:@11662.4]
  assign RetimeWrapper_84_clock = clock; // @[:@11684.4]
  assign RetimeWrapper_84_reset = reset; // @[:@11685.4]
  assign RetimeWrapper_84_io_flow = io_rPort_21_backpressure; // @[package.scala 95:18:@11687.4]
  assign RetimeWrapper_84_io_in = _T_1505 & io_rPort_21_en_0; // @[package.scala 94:16:@11686.4]
  assign RetimeWrapper_85_clock = clock; // @[:@11692.4]
  assign RetimeWrapper_85_reset = reset; // @[:@11693.4]
  assign RetimeWrapper_85_io_flow = io_rPort_21_backpressure; // @[package.scala 95:18:@11695.4]
  assign RetimeWrapper_85_io_in = _T_1729 & io_rPort_21_en_0; // @[package.scala 94:16:@11694.4]
  assign RetimeWrapper_86_clock = clock; // @[:@11700.4]
  assign RetimeWrapper_86_reset = reset; // @[:@11701.4]
  assign RetimeWrapper_86_io_flow = io_rPort_21_backpressure; // @[package.scala 95:18:@11703.4]
  assign RetimeWrapper_86_io_in = _T_1953 & io_rPort_21_en_0; // @[package.scala 94:16:@11702.4]
  assign RetimeWrapper_87_clock = clock; // @[:@11708.4]
  assign RetimeWrapper_87_reset = reset; // @[:@11709.4]
  assign RetimeWrapper_87_io_flow = io_rPort_21_backpressure; // @[package.scala 95:18:@11711.4]
  assign RetimeWrapper_87_io_in = _T_2177 & io_rPort_21_en_0; // @[package.scala 94:16:@11710.4]
  assign RetimeWrapper_88_clock = clock; // @[:@11732.4]
  assign RetimeWrapper_88_reset = reset; // @[:@11733.4]
  assign RetimeWrapper_88_io_flow = io_rPort_22_backpressure; // @[package.scala 95:18:@11735.4]
  assign RetimeWrapper_88_io_in = _T_1431 & io_rPort_22_en_0; // @[package.scala 94:16:@11734.4]
  assign RetimeWrapper_89_clock = clock; // @[:@11740.4]
  assign RetimeWrapper_89_reset = reset; // @[:@11741.4]
  assign RetimeWrapper_89_io_flow = io_rPort_22_backpressure; // @[package.scala 95:18:@11743.4]
  assign RetimeWrapper_89_io_in = _T_1655 & io_rPort_22_en_0; // @[package.scala 94:16:@11742.4]
  assign RetimeWrapper_90_clock = clock; // @[:@11748.4]
  assign RetimeWrapper_90_reset = reset; // @[:@11749.4]
  assign RetimeWrapper_90_io_flow = io_rPort_22_backpressure; // @[package.scala 95:18:@11751.4]
  assign RetimeWrapper_90_io_in = _T_1879 & io_rPort_22_en_0; // @[package.scala 94:16:@11750.4]
  assign RetimeWrapper_91_clock = clock; // @[:@11756.4]
  assign RetimeWrapper_91_reset = reset; // @[:@11757.4]
  assign RetimeWrapper_91_io_flow = io_rPort_22_backpressure; // @[package.scala 95:18:@11759.4]
  assign RetimeWrapper_91_io_in = _T_2103 & io_rPort_22_en_0; // @[package.scala 94:16:@11758.4]
  assign RetimeWrapper_92_clock = clock; // @[:@11780.4]
  assign RetimeWrapper_92_reset = reset; // @[:@11781.4]
  assign RetimeWrapper_92_io_flow = io_rPort_23_backpressure; // @[package.scala 95:18:@11783.4]
  assign RetimeWrapper_92_io_in = _T_1373 & io_rPort_23_en_0; // @[package.scala 94:16:@11782.4]
  assign RetimeWrapper_93_clock = clock; // @[:@11788.4]
  assign RetimeWrapper_93_reset = reset; // @[:@11789.4]
  assign RetimeWrapper_93_io_flow = io_rPort_23_backpressure; // @[package.scala 95:18:@11791.4]
  assign RetimeWrapper_93_io_in = _T_1597 & io_rPort_23_en_0; // @[package.scala 94:16:@11790.4]
  assign RetimeWrapper_94_clock = clock; // @[:@11796.4]
  assign RetimeWrapper_94_reset = reset; // @[:@11797.4]
  assign RetimeWrapper_94_io_flow = io_rPort_23_backpressure; // @[package.scala 95:18:@11799.4]
  assign RetimeWrapper_94_io_in = _T_1821 & io_rPort_23_en_0; // @[package.scala 94:16:@11798.4]
  assign RetimeWrapper_95_clock = clock; // @[:@11804.4]
  assign RetimeWrapper_95_reset = reset; // @[:@11805.4]
  assign RetimeWrapper_95_io_flow = io_rPort_23_backpressure; // @[package.scala 95:18:@11807.4]
  assign RetimeWrapper_95_io_in = _T_2045 & io_rPort_23_en_0; // @[package.scala 94:16:@11806.4]
endmodule
module RetimeWrapper_148( // @[:@11827.2]
  input         clock, // @[:@11828.4]
  input         reset, // @[:@11829.4]
  input         io_flow, // @[:@11830.4]
  input  [63:0] io_in, // @[:@11830.4]
  output [63:0] io_out // @[:@11830.4]
);
  wire [63:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@11832.4]
  wire [63:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@11832.4]
  wire [63:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@11832.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@11832.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@11832.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@11832.4]
  RetimeShiftRegister #(.WIDTH(64), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@11832.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@11845.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@11844.4]
  assign sr_init = 64'h0; // @[RetimeShiftRegister.scala 19:16:@11843.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@11842.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@11841.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@11839.4]
endmodule
module SimBlackBoxesfix2fixBox_2( // @[:@11847.2]
  input  [31:0] io_a, // @[:@11850.4]
  output [32:0] io_b // @[:@11850.4]
);
  wire  _T_20; // @[implicits.scala 69:16:@11857.4]
  assign _T_20 = io_a[31]; // @[implicits.scala 69:16:@11857.4]
  assign io_b = {_T_20,io_a}; // @[SimBlackBoxes.scala 99:40:@11862.4]
endmodule
module __2( // @[:@11864.2]
  input  [31:0] io_b, // @[:@11867.4]
  output [32:0] io_result // @[:@11867.4]
);
  wire [31:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@11872.4]
  wire [32:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@11872.4]
  SimBlackBoxesfix2fixBox_2 SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@11872.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@11885.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@11880.4]
endmodule
module RetimeWrapper_149( // @[:@11939.2]
  input         clock, // @[:@11940.4]
  input         reset, // @[:@11941.4]
  input         io_flow, // @[:@11942.4]
  input  [31:0] io_in, // @[:@11942.4]
  output [31:0] io_out // @[:@11942.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@11944.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@11944.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@11944.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@11944.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@11944.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@11944.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@11944.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@11957.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@11956.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@11955.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@11954.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@11953.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@11951.4]
endmodule
module fix2fixBox( // @[:@11959.2]
  input         clock, // @[:@11960.4]
  input         reset, // @[:@11961.4]
  input  [32:0] io_a, // @[:@11962.4]
  input         io_flow, // @[:@11962.4]
  output [31:0] io_b // @[:@11962.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@11972.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@11972.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@11972.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@11972.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@11972.4]
  RetimeWrapper_149 RetimeWrapper ( // @[package.scala 93:22:@11972.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@11979.4]
  assign RetimeWrapper_clock = clock; // @[:@11973.4]
  assign RetimeWrapper_reset = reset; // @[:@11974.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@11976.4]
  assign RetimeWrapper_io_in = io_a[31:0]; // @[package.scala 94:16:@11975.4]
endmodule
module x453_sum( // @[:@11981.2]
  input         clock, // @[:@11982.4]
  input         reset, // @[:@11983.4]
  input  [31:0] io_a, // @[:@11984.4]
  input  [31:0] io_b, // @[:@11984.4]
  input         io_flow, // @[:@11984.4]
  output [31:0] io_result // @[:@11984.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@11992.4]
  wire [32:0] __io_result; // @[Math.scala 709:24:@11992.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@11999.4]
  wire [32:0] __1_io_result; // @[Math.scala 709:24:@11999.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@12017.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@12017.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@12017.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@12017.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@12017.4]
  wire [32:0] a_upcast_number; // @[Math.scala 712:22:@11997.4 Math.scala 713:14:@11998.4]
  wire [32:0] b_upcast_number; // @[Math.scala 712:22:@12004.4 Math.scala 713:14:@12005.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@12006.4]
  __2 _ ( // @[Math.scala 709:24:@11992.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 709:24:@11999.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox fix2fixBox ( // @[Math.scala 141:30:@12017.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@11997.4 Math.scala 713:14:@11998.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@12004.4 Math.scala 713:14:@12005.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@12006.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@12025.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@11995.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@12002.4]
  assign fix2fixBox_clock = clock; // @[:@12018.4]
  assign fix2fixBox_reset = reset; // @[:@12019.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@12020.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@12023.4]
endmodule
module RetimeWrapper_150( // @[:@12039.2]
  input         clock, // @[:@12040.4]
  input         reset, // @[:@12041.4]
  input         io_flow, // @[:@12042.4]
  input  [31:0] io_in, // @[:@12042.4]
  output [31:0] io_out // @[:@12042.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@12044.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@12044.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@12044.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@12044.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@12044.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@12044.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(8)) sr ( // @[RetimeShiftRegister.scala 15:20:@12044.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@12057.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@12056.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@12055.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@12054.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@12053.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@12051.4]
endmodule
module RetimeWrapper_151( // @[:@12071.2]
  input        clock, // @[:@12072.4]
  input        reset, // @[:@12073.4]
  input        io_flow, // @[:@12074.4]
  input  [7:0] io_in, // @[:@12074.4]
  output [7:0] io_out // @[:@12074.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@12076.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@12076.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@12076.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@12076.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@12076.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@12076.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(7)) sr ( // @[RetimeShiftRegister.scala 15:20:@12076.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@12089.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@12088.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@12087.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@12086.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@12085.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@12083.4]
endmodule
module RetimeWrapper_152( // @[:@12103.2]
  input         clock, // @[:@12104.4]
  input         reset, // @[:@12105.4]
  input         io_flow, // @[:@12106.4]
  input  [31:0] io_in, // @[:@12106.4]
  output [31:0] io_out // @[:@12106.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@12108.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@12108.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@12108.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@12108.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@12108.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@12108.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(7)) sr ( // @[RetimeShiftRegister.scala 15:20:@12108.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@12121.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@12120.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@12119.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@12118.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@12117.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@12115.4]
endmodule
module RetimeWrapper_153( // @[:@12135.2]
  input   clock, // @[:@12136.4]
  input   reset, // @[:@12137.4]
  input   io_flow, // @[:@12138.4]
  input   io_in, // @[:@12138.4]
  output  io_out // @[:@12138.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@12140.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@12140.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@12140.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@12140.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@12140.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@12140.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(8)) sr ( // @[RetimeShiftRegister.scala 15:20:@12140.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@12153.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@12152.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@12151.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@12150.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@12149.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@12147.4]
endmodule
module RetimeWrapper_160( // @[:@12655.2]
  input         clock, // @[:@12656.4]
  input         reset, // @[:@12657.4]
  input         io_flow, // @[:@12658.4]
  input  [31:0] io_in, // @[:@12658.4]
  output [31:0] io_out // @[:@12658.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@12660.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@12660.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@12660.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@12660.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@12660.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@12660.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(6)) sr ( // @[RetimeShiftRegister.scala 15:20:@12660.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@12673.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@12672.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@12671.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@12670.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@12669.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@12667.4]
endmodule
module RetimeWrapper_191( // @[:@14979.2]
  input         clock, // @[:@14980.4]
  input         reset, // @[:@14981.4]
  input         io_flow, // @[:@14982.4]
  input  [31:0] io_in, // @[:@14982.4]
  output [31:0] io_out // @[:@14982.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@14984.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@14984.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@14984.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@14984.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@14984.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@14984.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(10)) sr ( // @[RetimeShiftRegister.scala 15:20:@14984.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@14997.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@14996.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@14995.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@14994.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@14993.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@14991.4]
endmodule
module RetimeWrapper_197( // @[:@15319.2]
  input   clock, // @[:@15320.4]
  input   reset, // @[:@15321.4]
  input   io_flow, // @[:@15322.4]
  input   io_in, // @[:@15322.4]
  output  io_out // @[:@15322.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@15324.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@15324.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@15324.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@15324.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@15324.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@15324.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(12)) sr ( // @[RetimeShiftRegister.scala 15:20:@15324.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@15337.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@15336.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@15335.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@15334.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@15333.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@15331.4]
endmodule
module RetimeWrapper_212( // @[:@16095.2]
  input         clock, // @[:@16096.4]
  input         reset, // @[:@16097.4]
  input         io_flow, // @[:@16098.4]
  input  [31:0] io_in, // @[:@16098.4]
  output [31:0] io_out // @[:@16098.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@16100.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@16100.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@16100.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@16100.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@16100.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@16100.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(11)) sr ( // @[RetimeShiftRegister.scala 15:20:@16100.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@16113.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@16112.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@16111.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@16110.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@16109.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@16107.4]
endmodule
module RetimeWrapper_229( // @[:@17527.2]
  input         clock, // @[:@17528.4]
  input         reset, // @[:@17529.4]
  input         io_flow, // @[:@17530.4]
  input  [31:0] io_in, // @[:@17530.4]
  output [31:0] io_out // @[:@17530.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@17532.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@17532.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@17532.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@17532.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@17532.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@17532.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@17532.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@17545.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@17544.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@17543.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@17542.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@17541.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@17539.4]
endmodule
module SimBlackBoxesfix2fixBox_82( // @[:@22215.2]
  input  [7:0] io_a, // @[:@22218.4]
  output [8:0] io_b // @[:@22218.4]
);
  assign io_b = {1'h0,io_a}; // @[SimBlackBoxes.scala 99:40:@22229.4]
endmodule
module __82( // @[:@22231.2]
  input  [7:0] io_b, // @[:@22234.4]
  output [8:0] io_result // @[:@22234.4]
);
  wire [7:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@22239.4]
  wire [8:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@22239.4]
  SimBlackBoxesfix2fixBox_82 SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@22239.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@22252.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@22247.4]
endmodule
module fix2fixBox_40( // @[:@22325.2]
  input        clock, // @[:@22326.4]
  input        reset, // @[:@22327.4]
  input  [8:0] io_a, // @[:@22328.4]
  input        io_flow, // @[:@22328.4]
  output [7:0] io_b // @[:@22328.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@22338.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@22338.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@22338.4]
  wire [7:0] RetimeWrapper_io_in; // @[package.scala 93:22:@22338.4]
  wire [7:0] RetimeWrapper_io_out; // @[package.scala 93:22:@22338.4]
  RetimeWrapper_21 RetimeWrapper ( // @[package.scala 93:22:@22338.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@22345.4]
  assign RetimeWrapper_clock = clock; // @[:@22339.4]
  assign RetimeWrapper_reset = reset; // @[:@22340.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@22342.4]
  assign RetimeWrapper_io_in = io_a[7:0]; // @[package.scala 94:16:@22341.4]
endmodule
module x725_x11( // @[:@22347.2]
  input        clock, // @[:@22348.4]
  input        reset, // @[:@22349.4]
  input  [7:0] io_a, // @[:@22350.4]
  input  [7:0] io_b, // @[:@22350.4]
  input        io_flow, // @[:@22350.4]
  output [7:0] io_result // @[:@22350.4]
);
  wire [7:0] __io_b; // @[Math.scala 709:24:@22358.4]
  wire [8:0] __io_result; // @[Math.scala 709:24:@22358.4]
  wire [7:0] __1_io_b; // @[Math.scala 709:24:@22365.4]
  wire [8:0] __1_io_result; // @[Math.scala 709:24:@22365.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@22375.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@22375.4]
  wire [8:0] fix2fixBox_io_a; // @[Math.scala 141:30:@22375.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@22375.4]
  wire [7:0] fix2fixBox_io_b; // @[Math.scala 141:30:@22375.4]
  wire [8:0] a_upcast_number; // @[Math.scala 712:22:@22363.4 Math.scala 713:14:@22364.4]
  wire [8:0] b_upcast_number; // @[Math.scala 712:22:@22370.4 Math.scala 713:14:@22371.4]
  wire [9:0] _T_21; // @[Math.scala 136:37:@22372.4]
  __82 _ ( // @[Math.scala 709:24:@22358.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __82 __1 ( // @[Math.scala 709:24:@22365.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_40 fix2fixBox ( // @[Math.scala 141:30:@22375.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@22363.4 Math.scala 713:14:@22364.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@22370.4 Math.scala 713:14:@22371.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@22372.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@22383.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@22361.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@22368.4]
  assign fix2fixBox_clock = clock; // @[:@22376.4]
  assign fix2fixBox_reset = reset; // @[:@22377.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@22378.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@22381.4]
endmodule
module fix2fixBox_44( // @[:@22973.2]
  input  [8:0] io_a, // @[:@22976.4]
  output [7:0] io_b // @[:@22976.4]
);
  assign io_b = io_a[7:0]; // @[Converter.scala 95:38:@22986.4]
endmodule
module x729_x11( // @[:@22988.2]
  input  [7:0] io_a, // @[:@22991.4]
  input  [7:0] io_b, // @[:@22991.4]
  output [7:0] io_result // @[:@22991.4]
);
  wire [7:0] __io_b; // @[Math.scala 709:24:@22999.4]
  wire [8:0] __io_result; // @[Math.scala 709:24:@22999.4]
  wire [7:0] __1_io_b; // @[Math.scala 709:24:@23006.4]
  wire [8:0] __1_io_result; // @[Math.scala 709:24:@23006.4]
  wire [8:0] fix2fixBox_io_a; // @[Math.scala 141:30:@23016.4]
  wire [7:0] fix2fixBox_io_b; // @[Math.scala 141:30:@23016.4]
  wire [8:0] a_upcast_number; // @[Math.scala 712:22:@23004.4 Math.scala 713:14:@23005.4]
  wire [8:0] b_upcast_number; // @[Math.scala 712:22:@23011.4 Math.scala 713:14:@23012.4]
  wire [9:0] _T_21; // @[Math.scala 136:37:@23013.4]
  __82 _ ( // @[Math.scala 709:24:@22999.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __82 __1 ( // @[Math.scala 709:24:@23006.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_44 fix2fixBox ( // @[Math.scala 141:30:@23016.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@23004.4 Math.scala 713:14:@23005.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@23011.4 Math.scala 713:14:@23012.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@23013.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@23024.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@23002.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@23009.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@23019.4]
endmodule
module RetimeWrapper_336( // @[:@32371.2]
  input         clock, // @[:@32372.4]
  input         reset, // @[:@32373.4]
  input         io_flow, // @[:@32374.4]
  input  [63:0] io_in, // @[:@32374.4]
  output [63:0] io_out // @[:@32374.4]
);
  wire [63:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@32376.4]
  wire [63:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@32376.4]
  wire [63:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@32376.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@32376.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@32376.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@32376.4]
  RetimeShiftRegister #(.WIDTH(64), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@32376.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@32389.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@32388.4]
  assign sr_init = 64'h0; // @[RetimeShiftRegister.scala 19:16:@32387.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@32386.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@32385.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@32383.4]
endmodule
module x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1( // @[:@32487.2]
  input          clock, // @[:@32488.4]
  input          reset, // @[:@32489.4]
  output         io_in_x426_TREADY, // @[:@32490.4]
  input  [255:0] io_in_x426_TDATA, // @[:@32490.4]
  input  [7:0]   io_in_x426_TID, // @[:@32490.4]
  input  [7:0]   io_in_x426_TDEST, // @[:@32490.4]
  output         io_in_x427_TVALID, // @[:@32490.4]
  input          io_in_x427_TREADY, // @[:@32490.4]
  output [255:0] io_in_x427_TDATA, // @[:@32490.4]
  input          io_sigsIn_backpressure, // @[:@32490.4]
  input          io_sigsIn_datapathEn, // @[:@32490.4]
  input          io_sigsIn_break, // @[:@32490.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_1, // @[:@32490.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_0, // @[:@32490.4]
  input          io_sigsIn_cchainOutputs_0_oobs_0, // @[:@32490.4]
  input          io_sigsIn_cchainOutputs_0_oobs_1, // @[:@32490.4]
  input          io_rr // @[:@32490.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@32504.4]
  wire [31:0] __io_result; // @[Math.scala 709:24:@32504.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@32516.4]
  wire [31:0] __1_io_result; // @[Math.scala 709:24:@32516.4]
  wire  x439_lb_0_clock; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_reset; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [2:0] x439_lb_0_io_rPort_23_banks_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_23_ofs_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_23_en_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_23_backpressure; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [7:0] x439_lb_0_io_rPort_23_output_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [2:0] x439_lb_0_io_rPort_22_banks_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_22_ofs_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_22_en_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_22_backpressure; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [7:0] x439_lb_0_io_rPort_22_output_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [2:0] x439_lb_0_io_rPort_21_banks_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_21_ofs_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_21_en_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_21_backpressure; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [7:0] x439_lb_0_io_rPort_21_output_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [2:0] x439_lb_0_io_rPort_20_banks_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_20_ofs_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_20_en_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_20_backpressure; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [7:0] x439_lb_0_io_rPort_20_output_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [2:0] x439_lb_0_io_rPort_19_banks_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_19_ofs_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_19_en_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_19_backpressure; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [7:0] x439_lb_0_io_rPort_19_output_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [2:0] x439_lb_0_io_rPort_18_banks_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_18_ofs_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_18_en_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_18_backpressure; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [7:0] x439_lb_0_io_rPort_18_output_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [2:0] x439_lb_0_io_rPort_17_banks_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_17_ofs_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_17_en_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_17_backpressure; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [7:0] x439_lb_0_io_rPort_17_output_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [2:0] x439_lb_0_io_rPort_16_banks_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_16_ofs_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_16_en_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_16_backpressure; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [7:0] x439_lb_0_io_rPort_16_output_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [2:0] x439_lb_0_io_rPort_15_banks_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_15_ofs_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_15_en_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_15_backpressure; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [7:0] x439_lb_0_io_rPort_15_output_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [2:0] x439_lb_0_io_rPort_14_banks_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_14_ofs_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_14_en_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_14_backpressure; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [7:0] x439_lb_0_io_rPort_14_output_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [2:0] x439_lb_0_io_rPort_13_banks_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_13_ofs_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_13_en_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_13_backpressure; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [7:0] x439_lb_0_io_rPort_13_output_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [2:0] x439_lb_0_io_rPort_12_banks_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_12_ofs_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_12_en_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_12_backpressure; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [7:0] x439_lb_0_io_rPort_12_output_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [2:0] x439_lb_0_io_rPort_11_banks_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_11_ofs_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_11_en_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_11_backpressure; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [7:0] x439_lb_0_io_rPort_11_output_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [2:0] x439_lb_0_io_rPort_10_banks_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_10_ofs_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_10_en_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_10_backpressure; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [7:0] x439_lb_0_io_rPort_10_output_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [2:0] x439_lb_0_io_rPort_9_banks_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_9_ofs_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_9_en_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_9_backpressure; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [7:0] x439_lb_0_io_rPort_9_output_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [2:0] x439_lb_0_io_rPort_8_banks_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_8_ofs_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_8_en_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_8_backpressure; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [7:0] x439_lb_0_io_rPort_8_output_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [2:0] x439_lb_0_io_rPort_7_banks_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_7_ofs_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_7_en_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_7_backpressure; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [7:0] x439_lb_0_io_rPort_7_output_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [2:0] x439_lb_0_io_rPort_6_banks_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_6_ofs_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_6_en_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_6_backpressure; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [7:0] x439_lb_0_io_rPort_6_output_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [2:0] x439_lb_0_io_rPort_5_banks_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_5_ofs_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_5_en_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_5_backpressure; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [7:0] x439_lb_0_io_rPort_5_output_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [2:0] x439_lb_0_io_rPort_4_banks_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_4_ofs_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_4_en_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_4_backpressure; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [7:0] x439_lb_0_io_rPort_4_output_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [2:0] x439_lb_0_io_rPort_3_banks_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_3_ofs_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_3_en_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_3_backpressure; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [7:0] x439_lb_0_io_rPort_3_output_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [2:0] x439_lb_0_io_rPort_2_banks_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_2_ofs_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_2_en_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_2_backpressure; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [7:0] x439_lb_0_io_rPort_2_output_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [2:0] x439_lb_0_io_rPort_1_banks_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_1_ofs_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_1_en_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_1_backpressure; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [7:0] x439_lb_0_io_rPort_1_output_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [2:0] x439_lb_0_io_rPort_0_banks_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_0_ofs_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_0_en_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_rPort_0_backpressure; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [7:0] x439_lb_0_io_rPort_0_output_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [2:0] x439_lb_0_io_wPort_7_banks_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_wPort_7_ofs_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [7:0] x439_lb_0_io_wPort_7_data_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_wPort_7_en_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [2:0] x439_lb_0_io_wPort_6_banks_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_wPort_6_ofs_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [7:0] x439_lb_0_io_wPort_6_data_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_wPort_6_en_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [2:0] x439_lb_0_io_wPort_5_banks_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_wPort_5_ofs_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [7:0] x439_lb_0_io_wPort_5_data_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_wPort_5_en_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [2:0] x439_lb_0_io_wPort_4_banks_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_wPort_4_ofs_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [7:0] x439_lb_0_io_wPort_4_data_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_wPort_4_en_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [2:0] x439_lb_0_io_wPort_3_banks_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_wPort_3_ofs_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [7:0] x439_lb_0_io_wPort_3_data_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_wPort_3_en_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [2:0] x439_lb_0_io_wPort_2_banks_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_wPort_2_ofs_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [7:0] x439_lb_0_io_wPort_2_data_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_wPort_2_en_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [2:0] x439_lb_0_io_wPort_1_banks_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_wPort_1_ofs_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [7:0] x439_lb_0_io_wPort_1_data_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_wPort_1_en_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [2:0] x439_lb_0_io_wPort_0_banks_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_wPort_0_ofs_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire [7:0] x439_lb_0_io_wPort_0_data_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  x439_lb_0_io_wPort_0_en_0; // @[m_x439_lb_0.scala 57:17:@32526.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@32752.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@32752.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@32752.4]
  wire [63:0] RetimeWrapper_io_in; // @[package.scala 93:22:@32752.4]
  wire [63:0] RetimeWrapper_io_out; // @[package.scala 93:22:@32752.4]
  wire  x453_sum_1_clock; // @[Math.scala 150:24:@32860.4]
  wire  x453_sum_1_reset; // @[Math.scala 150:24:@32860.4]
  wire [31:0] x453_sum_1_io_a; // @[Math.scala 150:24:@32860.4]
  wire [31:0] x453_sum_1_io_b; // @[Math.scala 150:24:@32860.4]
  wire  x453_sum_1_io_flow; // @[Math.scala 150:24:@32860.4]
  wire [31:0] x453_sum_1_io_result; // @[Math.scala 150:24:@32860.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@32870.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@32870.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@32870.4]
  wire [31:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@32870.4]
  wire [31:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@32870.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@32879.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@32879.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@32879.4]
  wire [7:0] RetimeWrapper_2_io_in; // @[package.scala 93:22:@32879.4]
  wire [7:0] RetimeWrapper_2_io_out; // @[package.scala 93:22:@32879.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@32888.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@32888.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@32888.4]
  wire [31:0] RetimeWrapper_3_io_in; // @[package.scala 93:22:@32888.4]
  wire [31:0] RetimeWrapper_3_io_out; // @[package.scala 93:22:@32888.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@32897.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@32897.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@32897.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@32897.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@32897.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@32906.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@32906.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@32906.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@32906.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@32906.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@32919.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@32919.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@32919.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@32919.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@32919.4]
  wire  x459_rdcol_1_clock; // @[Math.scala 150:24:@32942.4]
  wire  x459_rdcol_1_reset; // @[Math.scala 150:24:@32942.4]
  wire [31:0] x459_rdcol_1_io_a; // @[Math.scala 150:24:@32942.4]
  wire [31:0] x459_rdcol_1_io_b; // @[Math.scala 150:24:@32942.4]
  wire  x459_rdcol_1_io_flow; // @[Math.scala 150:24:@32942.4]
  wire [31:0] x459_rdcol_1_io_result; // @[Math.scala 150:24:@32942.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@32963.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@32963.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@32963.4]
  wire [31:0] RetimeWrapper_7_io_in; // @[package.scala 93:22:@32963.4]
  wire [31:0] RetimeWrapper_7_io_out; // @[package.scala 93:22:@32963.4]
  wire  x463_sum_1_clock; // @[Math.scala 150:24:@32972.4]
  wire  x463_sum_1_reset; // @[Math.scala 150:24:@32972.4]
  wire [31:0] x463_sum_1_io_a; // @[Math.scala 150:24:@32972.4]
  wire [31:0] x463_sum_1_io_b; // @[Math.scala 150:24:@32972.4]
  wire  x463_sum_1_io_flow; // @[Math.scala 150:24:@32972.4]
  wire [31:0] x463_sum_1_io_result; // @[Math.scala 150:24:@32972.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@32982.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@32982.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@32982.4]
  wire [7:0] RetimeWrapper_8_io_in; // @[package.scala 93:22:@32982.4]
  wire [7:0] RetimeWrapper_8_io_out; // @[package.scala 93:22:@32982.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@32991.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@32991.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@32991.4]
  wire [31:0] RetimeWrapper_9_io_in; // @[package.scala 93:22:@32991.4]
  wire [31:0] RetimeWrapper_9_io_out; // @[package.scala 93:22:@32991.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@33004.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@33004.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@33004.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@33004.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@33004.4]
  wire  x468_rdcol_1_clock; // @[Math.scala 150:24:@33027.4]
  wire  x468_rdcol_1_reset; // @[Math.scala 150:24:@33027.4]
  wire [31:0] x468_rdcol_1_io_a; // @[Math.scala 150:24:@33027.4]
  wire [31:0] x468_rdcol_1_io_b; // @[Math.scala 150:24:@33027.4]
  wire  x468_rdcol_1_io_flow; // @[Math.scala 150:24:@33027.4]
  wire [31:0] x468_rdcol_1_io_result; // @[Math.scala 150:24:@33027.4]
  wire  x472_sum_1_clock; // @[Math.scala 150:24:@33048.4]
  wire  x472_sum_1_reset; // @[Math.scala 150:24:@33048.4]
  wire [31:0] x472_sum_1_io_a; // @[Math.scala 150:24:@33048.4]
  wire [31:0] x472_sum_1_io_b; // @[Math.scala 150:24:@33048.4]
  wire  x472_sum_1_io_flow; // @[Math.scala 150:24:@33048.4]
  wire [31:0] x472_sum_1_io_result; // @[Math.scala 150:24:@33048.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@33058.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@33058.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@33058.4]
  wire [31:0] RetimeWrapper_11_io_in; // @[package.scala 93:22:@33058.4]
  wire [31:0] RetimeWrapper_11_io_out; // @[package.scala 93:22:@33058.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@33067.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@33067.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@33067.4]
  wire [7:0] RetimeWrapper_12_io_in; // @[package.scala 93:22:@33067.4]
  wire [7:0] RetimeWrapper_12_io_out; // @[package.scala 93:22:@33067.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@33080.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@33080.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@33080.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@33080.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@33080.4]
  wire  x477_rdcol_1_clock; // @[Math.scala 150:24:@33103.4]
  wire  x477_rdcol_1_reset; // @[Math.scala 150:24:@33103.4]
  wire [31:0] x477_rdcol_1_io_a; // @[Math.scala 150:24:@33103.4]
  wire [31:0] x477_rdcol_1_io_b; // @[Math.scala 150:24:@33103.4]
  wire  x477_rdcol_1_io_flow; // @[Math.scala 150:24:@33103.4]
  wire [31:0] x477_rdcol_1_io_result; // @[Math.scala 150:24:@33103.4]
  wire  x481_sum_1_clock; // @[Math.scala 150:24:@33124.4]
  wire  x481_sum_1_reset; // @[Math.scala 150:24:@33124.4]
  wire [31:0] x481_sum_1_io_a; // @[Math.scala 150:24:@33124.4]
  wire [31:0] x481_sum_1_io_b; // @[Math.scala 150:24:@33124.4]
  wire  x481_sum_1_io_flow; // @[Math.scala 150:24:@33124.4]
  wire [31:0] x481_sum_1_io_result; // @[Math.scala 150:24:@33124.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@33134.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@33134.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@33134.4]
  wire [31:0] RetimeWrapper_14_io_in; // @[package.scala 93:22:@33134.4]
  wire [31:0] RetimeWrapper_14_io_out; // @[package.scala 93:22:@33134.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@33143.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@33143.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@33143.4]
  wire [7:0] RetimeWrapper_15_io_in; // @[package.scala 93:22:@33143.4]
  wire [7:0] RetimeWrapper_15_io_out; // @[package.scala 93:22:@33143.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@33156.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@33156.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@33156.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@33156.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@33156.4]
  wire  x486_rdrow_1_clock; // @[Math.scala 150:24:@33179.4]
  wire  x486_rdrow_1_reset; // @[Math.scala 150:24:@33179.4]
  wire [31:0] x486_rdrow_1_io_a; // @[Math.scala 150:24:@33179.4]
  wire [31:0] x486_rdrow_1_io_b; // @[Math.scala 150:24:@33179.4]
  wire  x486_rdrow_1_io_flow; // @[Math.scala 150:24:@33179.4]
  wire [31:0] x486_rdrow_1_io_result; // @[Math.scala 150:24:@33179.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@33260.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@33260.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@33260.4]
  wire [31:0] RetimeWrapper_17_io_in; // @[package.scala 93:22:@33260.4]
  wire [31:0] RetimeWrapper_17_io_out; // @[package.scala 93:22:@33260.4]
  wire  x495_sum_1_clock; // @[Math.scala 150:24:@33269.4]
  wire  x495_sum_1_reset; // @[Math.scala 150:24:@33269.4]
  wire [31:0] x495_sum_1_io_a; // @[Math.scala 150:24:@33269.4]
  wire [31:0] x495_sum_1_io_b; // @[Math.scala 150:24:@33269.4]
  wire  x495_sum_1_io_flow; // @[Math.scala 150:24:@33269.4]
  wire [31:0] x495_sum_1_io_result; // @[Math.scala 150:24:@33269.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@33279.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@33279.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@33279.4]
  wire [31:0] RetimeWrapper_18_io_in; // @[package.scala 93:22:@33279.4]
  wire [31:0] RetimeWrapper_18_io_out; // @[package.scala 93:22:@33279.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@33288.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@33288.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@33288.4]
  wire [7:0] RetimeWrapper_19_io_in; // @[package.scala 93:22:@33288.4]
  wire [7:0] RetimeWrapper_19_io_out; // @[package.scala 93:22:@33288.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@33297.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@33297.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@33297.4]
  wire [31:0] RetimeWrapper_20_io_in; // @[package.scala 93:22:@33297.4]
  wire [31:0] RetimeWrapper_20_io_out; // @[package.scala 93:22:@33297.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@33310.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@33310.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@33310.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@33310.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@33310.4]
  wire  x501_sum_1_clock; // @[Math.scala 150:24:@33333.4]
  wire  x501_sum_1_reset; // @[Math.scala 150:24:@33333.4]
  wire [31:0] x501_sum_1_io_a; // @[Math.scala 150:24:@33333.4]
  wire [31:0] x501_sum_1_io_b; // @[Math.scala 150:24:@33333.4]
  wire  x501_sum_1_io_flow; // @[Math.scala 150:24:@33333.4]
  wire [31:0] x501_sum_1_io_result; // @[Math.scala 150:24:@33333.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@33343.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@33343.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@33343.4]
  wire [7:0] RetimeWrapper_22_io_in; // @[package.scala 93:22:@33343.4]
  wire [7:0] RetimeWrapper_22_io_out; // @[package.scala 93:22:@33343.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@33352.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@33352.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@33352.4]
  wire [31:0] RetimeWrapper_23_io_in; // @[package.scala 93:22:@33352.4]
  wire [31:0] RetimeWrapper_23_io_out; // @[package.scala 93:22:@33352.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@33365.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@33365.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@33365.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@33365.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@33365.4]
  wire  x506_sum_1_clock; // @[Math.scala 150:24:@33388.4]
  wire  x506_sum_1_reset; // @[Math.scala 150:24:@33388.4]
  wire [31:0] x506_sum_1_io_a; // @[Math.scala 150:24:@33388.4]
  wire [31:0] x506_sum_1_io_b; // @[Math.scala 150:24:@33388.4]
  wire  x506_sum_1_io_flow; // @[Math.scala 150:24:@33388.4]
  wire [31:0] x506_sum_1_io_result; // @[Math.scala 150:24:@33388.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@33398.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@33398.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@33398.4]
  wire [7:0] RetimeWrapper_25_io_in; // @[package.scala 93:22:@33398.4]
  wire [7:0] RetimeWrapper_25_io_out; // @[package.scala 93:22:@33398.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@33407.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@33407.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@33407.4]
  wire [31:0] RetimeWrapper_26_io_in; // @[package.scala 93:22:@33407.4]
  wire [31:0] RetimeWrapper_26_io_out; // @[package.scala 93:22:@33407.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@33420.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@33420.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@33420.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@33420.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@33420.4]
  wire  x511_sum_1_clock; // @[Math.scala 150:24:@33443.4]
  wire  x511_sum_1_reset; // @[Math.scala 150:24:@33443.4]
  wire [31:0] x511_sum_1_io_a; // @[Math.scala 150:24:@33443.4]
  wire [31:0] x511_sum_1_io_b; // @[Math.scala 150:24:@33443.4]
  wire  x511_sum_1_io_flow; // @[Math.scala 150:24:@33443.4]
  wire [31:0] x511_sum_1_io_result; // @[Math.scala 150:24:@33443.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@33453.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@33453.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@33453.4]
  wire [31:0] RetimeWrapper_28_io_in; // @[package.scala 93:22:@33453.4]
  wire [31:0] RetimeWrapper_28_io_out; // @[package.scala 93:22:@33453.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@33462.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@33462.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@33462.4]
  wire [7:0] RetimeWrapper_29_io_in; // @[package.scala 93:22:@33462.4]
  wire [7:0] RetimeWrapper_29_io_out; // @[package.scala 93:22:@33462.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@33475.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@33475.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@33475.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@33475.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@33475.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@33496.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@33496.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@33496.4]
  wire [31:0] RetimeWrapper_31_io_in; // @[package.scala 93:22:@33496.4]
  wire [31:0] RetimeWrapper_31_io_out; // @[package.scala 93:22:@33496.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@33523.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@33523.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@33523.4]
  wire [31:0] RetimeWrapper_32_io_in; // @[package.scala 93:22:@33523.4]
  wire [31:0] RetimeWrapper_32_io_out; // @[package.scala 93:22:@33523.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@33565.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@33565.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@33565.4]
  wire [31:0] RetimeWrapper_33_io_in; // @[package.scala 93:22:@33565.4]
  wire [31:0] RetimeWrapper_33_io_out; // @[package.scala 93:22:@33565.4]
  wire  x523_sum_1_clock; // @[Math.scala 150:24:@33574.4]
  wire  x523_sum_1_reset; // @[Math.scala 150:24:@33574.4]
  wire [31:0] x523_sum_1_io_a; // @[Math.scala 150:24:@33574.4]
  wire [31:0] x523_sum_1_io_b; // @[Math.scala 150:24:@33574.4]
  wire  x523_sum_1_io_flow; // @[Math.scala 150:24:@33574.4]
  wire [31:0] x523_sum_1_io_result; // @[Math.scala 150:24:@33574.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@33584.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@33584.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@33584.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@33584.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@33584.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@33593.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@33593.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@33593.4]
  wire [31:0] RetimeWrapper_35_io_in; // @[package.scala 93:22:@33593.4]
  wire [31:0] RetimeWrapper_35_io_out; // @[package.scala 93:22:@33593.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@33602.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@33602.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@33602.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@33602.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@33602.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@33611.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@33611.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@33611.4]
  wire  RetimeWrapper_37_io_in; // @[package.scala 93:22:@33611.4]
  wire  RetimeWrapper_37_io_out; // @[package.scala 93:22:@33611.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@33625.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@33625.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@33625.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@33625.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@33625.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@33646.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@33646.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@33646.4]
  wire [31:0] RetimeWrapper_39_io_in; // @[package.scala 93:22:@33646.4]
  wire [31:0] RetimeWrapper_39_io_out; // @[package.scala 93:22:@33646.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@33668.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@33668.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@33668.4]
  wire [31:0] RetimeWrapper_40_io_in; // @[package.scala 93:22:@33668.4]
  wire [31:0] RetimeWrapper_40_io_out; // @[package.scala 93:22:@33668.4]
  wire  x532_sum_1_clock; // @[Math.scala 150:24:@33677.4]
  wire  x532_sum_1_reset; // @[Math.scala 150:24:@33677.4]
  wire [31:0] x532_sum_1_io_a; // @[Math.scala 150:24:@33677.4]
  wire [31:0] x532_sum_1_io_b; // @[Math.scala 150:24:@33677.4]
  wire  x532_sum_1_io_flow; // @[Math.scala 150:24:@33677.4]
  wire [31:0] x532_sum_1_io_result; // @[Math.scala 150:24:@33677.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@33687.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@33687.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@33687.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@33687.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@33687.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@33701.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@33701.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@33701.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@33701.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@33701.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@33722.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@33722.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@33722.4]
  wire [31:0] RetimeWrapper_43_io_in; // @[package.scala 93:22:@33722.4]
  wire [31:0] RetimeWrapper_43_io_out; // @[package.scala 93:22:@33722.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@33746.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@33746.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@33746.4]
  wire [31:0] RetimeWrapper_44_io_in; // @[package.scala 93:22:@33746.4]
  wire [31:0] RetimeWrapper_44_io_out; // @[package.scala 93:22:@33746.4]
  wire  x540_sum_1_clock; // @[Math.scala 150:24:@33755.4]
  wire  x540_sum_1_reset; // @[Math.scala 150:24:@33755.4]
  wire [31:0] x540_sum_1_io_a; // @[Math.scala 150:24:@33755.4]
  wire [31:0] x540_sum_1_io_b; // @[Math.scala 150:24:@33755.4]
  wire  x540_sum_1_io_flow; // @[Math.scala 150:24:@33755.4]
  wire [31:0] x540_sum_1_io_result; // @[Math.scala 150:24:@33755.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@33765.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@33765.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@33765.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@33765.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@33765.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@33779.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@33779.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@33779.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@33779.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@33779.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@33800.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@33800.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@33800.4]
  wire [31:0] RetimeWrapper_47_io_in; // @[package.scala 93:22:@33800.4]
  wire [31:0] RetimeWrapper_47_io_out; // @[package.scala 93:22:@33800.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@33816.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@33816.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@33816.4]
  wire  RetimeWrapper_48_io_in; // @[package.scala 93:22:@33816.4]
  wire  RetimeWrapper_48_io_out; // @[package.scala 93:22:@33816.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@33831.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@33831.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@33831.4]
  wire [31:0] RetimeWrapper_49_io_in; // @[package.scala 93:22:@33831.4]
  wire [31:0] RetimeWrapper_49_io_out; // @[package.scala 93:22:@33831.4]
  wire  x548_sum_1_clock; // @[Math.scala 150:24:@33840.4]
  wire  x548_sum_1_reset; // @[Math.scala 150:24:@33840.4]
  wire [31:0] x548_sum_1_io_a; // @[Math.scala 150:24:@33840.4]
  wire [31:0] x548_sum_1_io_b; // @[Math.scala 150:24:@33840.4]
  wire  x548_sum_1_io_flow; // @[Math.scala 150:24:@33840.4]
  wire [31:0] x548_sum_1_io_result; // @[Math.scala 150:24:@33840.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@33850.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@33850.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@33850.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@33850.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@33850.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@33864.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@33864.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@33864.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@33864.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@33864.4]
  wire  x553_rdcol_1_clock; // @[Math.scala 150:24:@33887.4]
  wire  x553_rdcol_1_reset; // @[Math.scala 150:24:@33887.4]
  wire [31:0] x553_rdcol_1_io_a; // @[Math.scala 150:24:@33887.4]
  wire [31:0] x553_rdcol_1_io_b; // @[Math.scala 150:24:@33887.4]
  wire  x553_rdcol_1_io_flow; // @[Math.scala 150:24:@33887.4]
  wire [31:0] x553_rdcol_1_io_result; // @[Math.scala 150:24:@33887.4]
  wire  x559_sum_1_clock; // @[Math.scala 150:24:@33919.4]
  wire  x559_sum_1_reset; // @[Math.scala 150:24:@33919.4]
  wire [31:0] x559_sum_1_io_a; // @[Math.scala 150:24:@33919.4]
  wire [31:0] x559_sum_1_io_b; // @[Math.scala 150:24:@33919.4]
  wire  x559_sum_1_io_flow; // @[Math.scala 150:24:@33919.4]
  wire [31:0] x559_sum_1_io_result; // @[Math.scala 150:24:@33919.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@33929.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@33929.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@33929.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@33929.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@33929.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@33943.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@33943.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@33943.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@33943.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@33943.4]
  wire  x565_rdcol_1_clock; // @[Math.scala 150:24:@33966.4]
  wire  x565_rdcol_1_reset; // @[Math.scala 150:24:@33966.4]
  wire [31:0] x565_rdcol_1_io_a; // @[Math.scala 150:24:@33966.4]
  wire [31:0] x565_rdcol_1_io_b; // @[Math.scala 150:24:@33966.4]
  wire  x565_rdcol_1_io_flow; // @[Math.scala 150:24:@33966.4]
  wire [31:0] x565_rdcol_1_io_result; // @[Math.scala 150:24:@33966.4]
  wire  x571_sum_1_clock; // @[Math.scala 150:24:@33998.4]
  wire  x571_sum_1_reset; // @[Math.scala 150:24:@33998.4]
  wire [31:0] x571_sum_1_io_a; // @[Math.scala 150:24:@33998.4]
  wire [31:0] x571_sum_1_io_b; // @[Math.scala 150:24:@33998.4]
  wire  x571_sum_1_io_flow; // @[Math.scala 150:24:@33998.4]
  wire [31:0] x571_sum_1_io_result; // @[Math.scala 150:24:@33998.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@34008.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@34008.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@34008.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@34008.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@34008.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@34022.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@34022.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@34022.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@34022.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@34022.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@34043.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@34043.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@34043.4]
  wire [31:0] RetimeWrapper_56_io_in; // @[package.scala 93:22:@34043.4]
  wire [31:0] RetimeWrapper_56_io_out; // @[package.scala 93:22:@34043.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@34070.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@34070.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@34070.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@34070.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@34070.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@34105.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@34105.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@34105.4]
  wire [31:0] RetimeWrapper_58_io_in; // @[package.scala 93:22:@34105.4]
  wire [31:0] RetimeWrapper_58_io_out; // @[package.scala 93:22:@34105.4]
  wire  x583_sum_1_clock; // @[Math.scala 150:24:@34114.4]
  wire  x583_sum_1_reset; // @[Math.scala 150:24:@34114.4]
  wire [31:0] x583_sum_1_io_a; // @[Math.scala 150:24:@34114.4]
  wire [31:0] x583_sum_1_io_b; // @[Math.scala 150:24:@34114.4]
  wire  x583_sum_1_io_flow; // @[Math.scala 150:24:@34114.4]
  wire [31:0] x583_sum_1_io_result; // @[Math.scala 150:24:@34114.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@34124.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@34124.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@34124.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@34124.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@34124.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@34133.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@34133.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@34133.4]
  wire [31:0] RetimeWrapper_60_io_in; // @[package.scala 93:22:@34133.4]
  wire [31:0] RetimeWrapper_60_io_out; // @[package.scala 93:22:@34133.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@34147.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@34147.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@34147.4]
  wire  RetimeWrapper_61_io_in; // @[package.scala 93:22:@34147.4]
  wire  RetimeWrapper_61_io_out; // @[package.scala 93:22:@34147.4]
  wire  x591_sum_1_clock; // @[Math.scala 150:24:@34176.4]
  wire  x591_sum_1_reset; // @[Math.scala 150:24:@34176.4]
  wire [31:0] x591_sum_1_io_a; // @[Math.scala 150:24:@34176.4]
  wire [31:0] x591_sum_1_io_b; // @[Math.scala 150:24:@34176.4]
  wire  x591_sum_1_io_flow; // @[Math.scala 150:24:@34176.4]
  wire [31:0] x591_sum_1_io_result; // @[Math.scala 150:24:@34176.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@34186.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@34186.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@34186.4]
  wire  RetimeWrapper_62_io_in; // @[package.scala 93:22:@34186.4]
  wire  RetimeWrapper_62_io_out; // @[package.scala 93:22:@34186.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@34200.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@34200.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@34200.4]
  wire  RetimeWrapper_63_io_in; // @[package.scala 93:22:@34200.4]
  wire  RetimeWrapper_63_io_out; // @[package.scala 93:22:@34200.4]
  wire  x598_sum_1_clock; // @[Math.scala 150:24:@34227.4]
  wire  x598_sum_1_reset; // @[Math.scala 150:24:@34227.4]
  wire [31:0] x598_sum_1_io_a; // @[Math.scala 150:24:@34227.4]
  wire [31:0] x598_sum_1_io_b; // @[Math.scala 150:24:@34227.4]
  wire  x598_sum_1_io_flow; // @[Math.scala 150:24:@34227.4]
  wire [31:0] x598_sum_1_io_result; // @[Math.scala 150:24:@34227.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@34237.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@34237.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@34237.4]
  wire  RetimeWrapper_64_io_in; // @[package.scala 93:22:@34237.4]
  wire  RetimeWrapper_64_io_out; // @[package.scala 93:22:@34237.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@34251.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@34251.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@34251.4]
  wire  RetimeWrapper_65_io_in; // @[package.scala 93:22:@34251.4]
  wire  RetimeWrapper_65_io_out; // @[package.scala 93:22:@34251.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@34278.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@34278.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@34278.4]
  wire [31:0] RetimeWrapper_66_io_in; // @[package.scala 93:22:@34278.4]
  wire [31:0] RetimeWrapper_66_io_out; // @[package.scala 93:22:@34278.4]
  wire  x605_sum_1_clock; // @[Math.scala 150:24:@34287.4]
  wire  x605_sum_1_reset; // @[Math.scala 150:24:@34287.4]
  wire [31:0] x605_sum_1_io_a; // @[Math.scala 150:24:@34287.4]
  wire [31:0] x605_sum_1_io_b; // @[Math.scala 150:24:@34287.4]
  wire  x605_sum_1_io_flow; // @[Math.scala 150:24:@34287.4]
  wire [31:0] x605_sum_1_io_result; // @[Math.scala 150:24:@34287.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@34297.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@34297.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@34297.4]
  wire [31:0] RetimeWrapper_67_io_in; // @[package.scala 93:22:@34297.4]
  wire [31:0] RetimeWrapper_67_io_out; // @[package.scala 93:22:@34297.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@34306.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@34306.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@34306.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@34306.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@34306.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@34320.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@34320.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@34320.4]
  wire  RetimeWrapper_69_io_in; // @[package.scala 93:22:@34320.4]
  wire  RetimeWrapper_69_io_out; // @[package.scala 93:22:@34320.4]
  wire  x612_sum_1_clock; // @[Math.scala 150:24:@34347.4]
  wire  x612_sum_1_reset; // @[Math.scala 150:24:@34347.4]
  wire [31:0] x612_sum_1_io_a; // @[Math.scala 150:24:@34347.4]
  wire [31:0] x612_sum_1_io_b; // @[Math.scala 150:24:@34347.4]
  wire  x612_sum_1_io_flow; // @[Math.scala 150:24:@34347.4]
  wire [31:0] x612_sum_1_io_result; // @[Math.scala 150:24:@34347.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@34357.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@34357.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@34357.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@34357.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@34357.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@34371.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@34371.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@34371.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@34371.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@34371.4]
  wire  x619_sum_1_clock; // @[Math.scala 150:24:@34398.4]
  wire  x619_sum_1_reset; // @[Math.scala 150:24:@34398.4]
  wire [31:0] x619_sum_1_io_a; // @[Math.scala 150:24:@34398.4]
  wire [31:0] x619_sum_1_io_b; // @[Math.scala 150:24:@34398.4]
  wire  x619_sum_1_io_flow; // @[Math.scala 150:24:@34398.4]
  wire [31:0] x619_sum_1_io_result; // @[Math.scala 150:24:@34398.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@34408.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@34408.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@34408.4]
  wire  RetimeWrapper_72_io_in; // @[package.scala 93:22:@34408.4]
  wire  RetimeWrapper_72_io_out; // @[package.scala 93:22:@34408.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@34422.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@34422.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@34422.4]
  wire  RetimeWrapper_73_io_in; // @[package.scala 93:22:@34422.4]
  wire  RetimeWrapper_73_io_out; // @[package.scala 93:22:@34422.4]
  wire  x624_rdrow_1_clock; // @[Math.scala 150:24:@34445.4]
  wire  x624_rdrow_1_reset; // @[Math.scala 150:24:@34445.4]
  wire [31:0] x624_rdrow_1_io_a; // @[Math.scala 150:24:@34445.4]
  wire [31:0] x624_rdrow_1_io_b; // @[Math.scala 150:24:@34445.4]
  wire  x624_rdrow_1_io_flow; // @[Math.scala 150:24:@34445.4]
  wire [31:0] x624_rdrow_1_io_result; // @[Math.scala 150:24:@34445.4]
  wire  x631_sum_1_clock; // @[Math.scala 150:24:@34499.4]
  wire  x631_sum_1_reset; // @[Math.scala 150:24:@34499.4]
  wire [31:0] x631_sum_1_io_a; // @[Math.scala 150:24:@34499.4]
  wire [31:0] x631_sum_1_io_b; // @[Math.scala 150:24:@34499.4]
  wire  x631_sum_1_io_flow; // @[Math.scala 150:24:@34499.4]
  wire [31:0] x631_sum_1_io_result; // @[Math.scala 150:24:@34499.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@34509.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@34509.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@34509.4]
  wire  RetimeWrapper_74_io_in; // @[package.scala 93:22:@34509.4]
  wire  RetimeWrapper_74_io_out; // @[package.scala 93:22:@34509.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@34518.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@34518.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@34518.4]
  wire [31:0] RetimeWrapper_75_io_in; // @[package.scala 93:22:@34518.4]
  wire [31:0] RetimeWrapper_75_io_out; // @[package.scala 93:22:@34518.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@34532.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@34532.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@34532.4]
  wire  RetimeWrapper_76_io_in; // @[package.scala 93:22:@34532.4]
  wire  RetimeWrapper_76_io_out; // @[package.scala 93:22:@34532.4]
  wire  x639_sum_1_clock; // @[Math.scala 150:24:@34561.4]
  wire  x639_sum_1_reset; // @[Math.scala 150:24:@34561.4]
  wire [31:0] x639_sum_1_io_a; // @[Math.scala 150:24:@34561.4]
  wire [31:0] x639_sum_1_io_b; // @[Math.scala 150:24:@34561.4]
  wire  x639_sum_1_io_flow; // @[Math.scala 150:24:@34561.4]
  wire [31:0] x639_sum_1_io_result; // @[Math.scala 150:24:@34561.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@34571.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@34571.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@34571.4]
  wire  RetimeWrapper_77_io_in; // @[package.scala 93:22:@34571.4]
  wire  RetimeWrapper_77_io_out; // @[package.scala 93:22:@34571.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@34585.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@34585.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@34585.4]
  wire  RetimeWrapper_78_io_in; // @[package.scala 93:22:@34585.4]
  wire  RetimeWrapper_78_io_out; // @[package.scala 93:22:@34585.4]
  wire  x646_sum_1_clock; // @[Math.scala 150:24:@34612.4]
  wire  x646_sum_1_reset; // @[Math.scala 150:24:@34612.4]
  wire [31:0] x646_sum_1_io_a; // @[Math.scala 150:24:@34612.4]
  wire [31:0] x646_sum_1_io_b; // @[Math.scala 150:24:@34612.4]
  wire  x646_sum_1_io_flow; // @[Math.scala 150:24:@34612.4]
  wire [31:0] x646_sum_1_io_result; // @[Math.scala 150:24:@34612.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@34622.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@34622.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@34622.4]
  wire  RetimeWrapper_79_io_in; // @[package.scala 93:22:@34622.4]
  wire  RetimeWrapper_79_io_out; // @[package.scala 93:22:@34622.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@34636.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@34636.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@34636.4]
  wire  RetimeWrapper_80_io_in; // @[package.scala 93:22:@34636.4]
  wire  RetimeWrapper_80_io_out; // @[package.scala 93:22:@34636.4]
  wire  x653_sum_1_clock; // @[Math.scala 150:24:@34663.4]
  wire  x653_sum_1_reset; // @[Math.scala 150:24:@34663.4]
  wire [31:0] x653_sum_1_io_a; // @[Math.scala 150:24:@34663.4]
  wire [31:0] x653_sum_1_io_b; // @[Math.scala 150:24:@34663.4]
  wire  x653_sum_1_io_flow; // @[Math.scala 150:24:@34663.4]
  wire [31:0] x653_sum_1_io_result; // @[Math.scala 150:24:@34663.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@34673.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@34673.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@34673.4]
  wire  RetimeWrapper_81_io_in; // @[package.scala 93:22:@34673.4]
  wire  RetimeWrapper_81_io_out; // @[package.scala 93:22:@34673.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@34687.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@34687.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@34687.4]
  wire  RetimeWrapper_82_io_in; // @[package.scala 93:22:@34687.4]
  wire  RetimeWrapper_82_io_out; // @[package.scala 93:22:@34687.4]
  wire  x660_sum_1_clock; // @[Math.scala 150:24:@34714.4]
  wire  x660_sum_1_reset; // @[Math.scala 150:24:@34714.4]
  wire [31:0] x660_sum_1_io_a; // @[Math.scala 150:24:@34714.4]
  wire [31:0] x660_sum_1_io_b; // @[Math.scala 150:24:@34714.4]
  wire  x660_sum_1_io_flow; // @[Math.scala 150:24:@34714.4]
  wire [31:0] x660_sum_1_io_result; // @[Math.scala 150:24:@34714.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@34724.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@34724.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@34724.4]
  wire  RetimeWrapper_83_io_in; // @[package.scala 93:22:@34724.4]
  wire  RetimeWrapper_83_io_out; // @[package.scala 93:22:@34724.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@34738.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@34738.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@34738.4]
  wire  RetimeWrapper_84_io_in; // @[package.scala 93:22:@34738.4]
  wire  RetimeWrapper_84_io_out; // @[package.scala 93:22:@34738.4]
  wire  x667_sum_1_clock; // @[Math.scala 150:24:@34765.4]
  wire  x667_sum_1_reset; // @[Math.scala 150:24:@34765.4]
  wire [31:0] x667_sum_1_io_a; // @[Math.scala 150:24:@34765.4]
  wire [31:0] x667_sum_1_io_b; // @[Math.scala 150:24:@34765.4]
  wire  x667_sum_1_io_flow; // @[Math.scala 150:24:@34765.4]
  wire [31:0] x667_sum_1_io_result; // @[Math.scala 150:24:@34765.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@34775.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@34775.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@34775.4]
  wire  RetimeWrapper_85_io_in; // @[package.scala 93:22:@34775.4]
  wire  RetimeWrapper_85_io_out; // @[package.scala 93:22:@34775.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@34789.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@34789.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@34789.4]
  wire  RetimeWrapper_86_io_in; // @[package.scala 93:22:@34789.4]
  wire  RetimeWrapper_86_io_out; // @[package.scala 93:22:@34789.4]
  wire  x672_rdrow_1_clock; // @[Math.scala 150:24:@34812.4]
  wire  x672_rdrow_1_reset; // @[Math.scala 150:24:@34812.4]
  wire [31:0] x672_rdrow_1_io_a; // @[Math.scala 150:24:@34812.4]
  wire [31:0] x672_rdrow_1_io_b; // @[Math.scala 150:24:@34812.4]
  wire  x672_rdrow_1_io_flow; // @[Math.scala 150:24:@34812.4]
  wire [31:0] x672_rdrow_1_io_result; // @[Math.scala 150:24:@34812.4]
  wire  x679_sum_1_clock; // @[Math.scala 150:24:@34866.4]
  wire  x679_sum_1_reset; // @[Math.scala 150:24:@34866.4]
  wire [31:0] x679_sum_1_io_a; // @[Math.scala 150:24:@34866.4]
  wire [31:0] x679_sum_1_io_b; // @[Math.scala 150:24:@34866.4]
  wire  x679_sum_1_io_flow; // @[Math.scala 150:24:@34866.4]
  wire [31:0] x679_sum_1_io_result; // @[Math.scala 150:24:@34866.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@34876.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@34876.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@34876.4]
  wire [31:0] RetimeWrapper_87_io_in; // @[package.scala 93:22:@34876.4]
  wire [31:0] RetimeWrapper_87_io_out; // @[package.scala 93:22:@34876.4]
  wire  RetimeWrapper_88_clock; // @[package.scala 93:22:@34885.4]
  wire  RetimeWrapper_88_reset; // @[package.scala 93:22:@34885.4]
  wire  RetimeWrapper_88_io_flow; // @[package.scala 93:22:@34885.4]
  wire  RetimeWrapper_88_io_in; // @[package.scala 93:22:@34885.4]
  wire  RetimeWrapper_88_io_out; // @[package.scala 93:22:@34885.4]
  wire  RetimeWrapper_89_clock; // @[package.scala 93:22:@34899.4]
  wire  RetimeWrapper_89_reset; // @[package.scala 93:22:@34899.4]
  wire  RetimeWrapper_89_io_flow; // @[package.scala 93:22:@34899.4]
  wire  RetimeWrapper_89_io_in; // @[package.scala 93:22:@34899.4]
  wire  RetimeWrapper_89_io_out; // @[package.scala 93:22:@34899.4]
  wire  x687_sum_1_clock; // @[Math.scala 150:24:@34926.4]
  wire  x687_sum_1_reset; // @[Math.scala 150:24:@34926.4]
  wire [31:0] x687_sum_1_io_a; // @[Math.scala 150:24:@34926.4]
  wire [31:0] x687_sum_1_io_b; // @[Math.scala 150:24:@34926.4]
  wire  x687_sum_1_io_flow; // @[Math.scala 150:24:@34926.4]
  wire [31:0] x687_sum_1_io_result; // @[Math.scala 150:24:@34926.4]
  wire  RetimeWrapper_90_clock; // @[package.scala 93:22:@34936.4]
  wire  RetimeWrapper_90_reset; // @[package.scala 93:22:@34936.4]
  wire  RetimeWrapper_90_io_flow; // @[package.scala 93:22:@34936.4]
  wire  RetimeWrapper_90_io_in; // @[package.scala 93:22:@34936.4]
  wire  RetimeWrapper_90_io_out; // @[package.scala 93:22:@34936.4]
  wire  RetimeWrapper_91_clock; // @[package.scala 93:22:@34950.4]
  wire  RetimeWrapper_91_reset; // @[package.scala 93:22:@34950.4]
  wire  RetimeWrapper_91_io_flow; // @[package.scala 93:22:@34950.4]
  wire  RetimeWrapper_91_io_in; // @[package.scala 93:22:@34950.4]
  wire  RetimeWrapper_91_io_out; // @[package.scala 93:22:@34950.4]
  wire  x694_sum_1_clock; // @[Math.scala 150:24:@34979.4]
  wire  x694_sum_1_reset; // @[Math.scala 150:24:@34979.4]
  wire [31:0] x694_sum_1_io_a; // @[Math.scala 150:24:@34979.4]
  wire [31:0] x694_sum_1_io_b; // @[Math.scala 150:24:@34979.4]
  wire  x694_sum_1_io_flow; // @[Math.scala 150:24:@34979.4]
  wire [31:0] x694_sum_1_io_result; // @[Math.scala 150:24:@34979.4]
  wire  RetimeWrapper_92_clock; // @[package.scala 93:22:@34989.4]
  wire  RetimeWrapper_92_reset; // @[package.scala 93:22:@34989.4]
  wire  RetimeWrapper_92_io_flow; // @[package.scala 93:22:@34989.4]
  wire  RetimeWrapper_92_io_in; // @[package.scala 93:22:@34989.4]
  wire  RetimeWrapper_92_io_out; // @[package.scala 93:22:@34989.4]
  wire  RetimeWrapper_93_clock; // @[package.scala 93:22:@35003.4]
  wire  RetimeWrapper_93_reset; // @[package.scala 93:22:@35003.4]
  wire  RetimeWrapper_93_io_flow; // @[package.scala 93:22:@35003.4]
  wire  RetimeWrapper_93_io_in; // @[package.scala 93:22:@35003.4]
  wire  RetimeWrapper_93_io_out; // @[package.scala 93:22:@35003.4]
  wire  x701_sum_1_clock; // @[Math.scala 150:24:@35030.4]
  wire  x701_sum_1_reset; // @[Math.scala 150:24:@35030.4]
  wire [31:0] x701_sum_1_io_a; // @[Math.scala 150:24:@35030.4]
  wire [31:0] x701_sum_1_io_b; // @[Math.scala 150:24:@35030.4]
  wire  x701_sum_1_io_flow; // @[Math.scala 150:24:@35030.4]
  wire [31:0] x701_sum_1_io_result; // @[Math.scala 150:24:@35030.4]
  wire  RetimeWrapper_94_clock; // @[package.scala 93:22:@35040.4]
  wire  RetimeWrapper_94_reset; // @[package.scala 93:22:@35040.4]
  wire  RetimeWrapper_94_io_flow; // @[package.scala 93:22:@35040.4]
  wire  RetimeWrapper_94_io_in; // @[package.scala 93:22:@35040.4]
  wire  RetimeWrapper_94_io_out; // @[package.scala 93:22:@35040.4]
  wire  RetimeWrapper_95_clock; // @[package.scala 93:22:@35054.4]
  wire  RetimeWrapper_95_reset; // @[package.scala 93:22:@35054.4]
  wire  RetimeWrapper_95_io_flow; // @[package.scala 93:22:@35054.4]
  wire  RetimeWrapper_95_io_in; // @[package.scala 93:22:@35054.4]
  wire  RetimeWrapper_95_io_out; // @[package.scala 93:22:@35054.4]
  wire  x708_sum_1_clock; // @[Math.scala 150:24:@35081.4]
  wire  x708_sum_1_reset; // @[Math.scala 150:24:@35081.4]
  wire [31:0] x708_sum_1_io_a; // @[Math.scala 150:24:@35081.4]
  wire [31:0] x708_sum_1_io_b; // @[Math.scala 150:24:@35081.4]
  wire  x708_sum_1_io_flow; // @[Math.scala 150:24:@35081.4]
  wire [31:0] x708_sum_1_io_result; // @[Math.scala 150:24:@35081.4]
  wire  RetimeWrapper_96_clock; // @[package.scala 93:22:@35091.4]
  wire  RetimeWrapper_96_reset; // @[package.scala 93:22:@35091.4]
  wire  RetimeWrapper_96_io_flow; // @[package.scala 93:22:@35091.4]
  wire  RetimeWrapper_96_io_in; // @[package.scala 93:22:@35091.4]
  wire  RetimeWrapper_96_io_out; // @[package.scala 93:22:@35091.4]
  wire  RetimeWrapper_97_clock; // @[package.scala 93:22:@35105.4]
  wire  RetimeWrapper_97_reset; // @[package.scala 93:22:@35105.4]
  wire  RetimeWrapper_97_io_flow; // @[package.scala 93:22:@35105.4]
  wire  RetimeWrapper_97_io_in; // @[package.scala 93:22:@35105.4]
  wire  RetimeWrapper_97_io_out; // @[package.scala 93:22:@35105.4]
  wire  x715_sum_1_clock; // @[Math.scala 150:24:@35132.4]
  wire  x715_sum_1_reset; // @[Math.scala 150:24:@35132.4]
  wire [31:0] x715_sum_1_io_a; // @[Math.scala 150:24:@35132.4]
  wire [31:0] x715_sum_1_io_b; // @[Math.scala 150:24:@35132.4]
  wire  x715_sum_1_io_flow; // @[Math.scala 150:24:@35132.4]
  wire [31:0] x715_sum_1_io_result; // @[Math.scala 150:24:@35132.4]
  wire  RetimeWrapper_98_clock; // @[package.scala 93:22:@35142.4]
  wire  RetimeWrapper_98_reset; // @[package.scala 93:22:@35142.4]
  wire  RetimeWrapper_98_io_flow; // @[package.scala 93:22:@35142.4]
  wire  RetimeWrapper_98_io_in; // @[package.scala 93:22:@35142.4]
  wire  RetimeWrapper_98_io_out; // @[package.scala 93:22:@35142.4]
  wire  RetimeWrapper_99_clock; // @[package.scala 93:22:@35156.4]
  wire  RetimeWrapper_99_reset; // @[package.scala 93:22:@35156.4]
  wire  RetimeWrapper_99_io_flow; // @[package.scala 93:22:@35156.4]
  wire  RetimeWrapper_99_io_in; // @[package.scala 93:22:@35156.4]
  wire  RetimeWrapper_99_io_out; // @[package.scala 93:22:@35156.4]
  wire  x725_x11_1_clock; // @[Math.scala 150:24:@35202.4]
  wire  x725_x11_1_reset; // @[Math.scala 150:24:@35202.4]
  wire [7:0] x725_x11_1_io_a; // @[Math.scala 150:24:@35202.4]
  wire [7:0] x725_x11_1_io_b; // @[Math.scala 150:24:@35202.4]
  wire  x725_x11_1_io_flow; // @[Math.scala 150:24:@35202.4]
  wire [7:0] x725_x11_1_io_result; // @[Math.scala 150:24:@35202.4]
  wire  x726_x12_1_clock; // @[Math.scala 150:24:@35212.4]
  wire  x726_x12_1_reset; // @[Math.scala 150:24:@35212.4]
  wire [7:0] x726_x12_1_io_a; // @[Math.scala 150:24:@35212.4]
  wire [7:0] x726_x12_1_io_b; // @[Math.scala 150:24:@35212.4]
  wire  x726_x12_1_io_flow; // @[Math.scala 150:24:@35212.4]
  wire [7:0] x726_x12_1_io_result; // @[Math.scala 150:24:@35212.4]
  wire  x727_x11_1_clock; // @[Math.scala 150:24:@35222.4]
  wire  x727_x11_1_reset; // @[Math.scala 150:24:@35222.4]
  wire [7:0] x727_x11_1_io_a; // @[Math.scala 150:24:@35222.4]
  wire [7:0] x727_x11_1_io_b; // @[Math.scala 150:24:@35222.4]
  wire  x727_x11_1_io_flow; // @[Math.scala 150:24:@35222.4]
  wire [7:0] x727_x11_1_io_result; // @[Math.scala 150:24:@35222.4]
  wire  x728_x12_1_clock; // @[Math.scala 150:24:@35232.4]
  wire  x728_x12_1_reset; // @[Math.scala 150:24:@35232.4]
  wire [7:0] x728_x12_1_io_a; // @[Math.scala 150:24:@35232.4]
  wire [7:0] x728_x12_1_io_b; // @[Math.scala 150:24:@35232.4]
  wire  x728_x12_1_io_flow; // @[Math.scala 150:24:@35232.4]
  wire [7:0] x728_x12_1_io_result; // @[Math.scala 150:24:@35232.4]
  wire [7:0] x729_x11_1_io_a; // @[Math.scala 150:24:@35242.4]
  wire [7:0] x729_x11_1_io_b; // @[Math.scala 150:24:@35242.4]
  wire [7:0] x729_x11_1_io_result; // @[Math.scala 150:24:@35242.4]
  wire [7:0] x730_x12_1_io_a; // @[Math.scala 150:24:@35252.4]
  wire [7:0] x730_x12_1_io_b; // @[Math.scala 150:24:@35252.4]
  wire [7:0] x730_x12_1_io_result; // @[Math.scala 150:24:@35252.4]
  wire [7:0] x731_x11_1_io_a; // @[Math.scala 150:24:@35262.4]
  wire [7:0] x731_x11_1_io_b; // @[Math.scala 150:24:@35262.4]
  wire [7:0] x731_x11_1_io_result; // @[Math.scala 150:24:@35262.4]
  wire  RetimeWrapper_100_clock; // @[package.scala 93:22:@35272.4]
  wire  RetimeWrapper_100_reset; // @[package.scala 93:22:@35272.4]
  wire  RetimeWrapper_100_io_flow; // @[package.scala 93:22:@35272.4]
  wire [7:0] RetimeWrapper_100_io_in; // @[package.scala 93:22:@35272.4]
  wire [7:0] RetimeWrapper_100_io_out; // @[package.scala 93:22:@35272.4]
  wire [7:0] x732_sum_1_io_a; // @[Math.scala 150:24:@35281.4]
  wire [7:0] x732_sum_1_io_b; // @[Math.scala 150:24:@35281.4]
  wire [7:0] x732_sum_1_io_result; // @[Math.scala 150:24:@35281.4]
  wire  RetimeWrapper_101_clock; // @[package.scala 93:22:@35295.4]
  wire  RetimeWrapper_101_reset; // @[package.scala 93:22:@35295.4]
  wire  RetimeWrapper_101_io_flow; // @[package.scala 93:22:@35295.4]
  wire [7:0] RetimeWrapper_101_io_in; // @[package.scala 93:22:@35295.4]
  wire [7:0] RetimeWrapper_101_io_out; // @[package.scala 93:22:@35295.4]
  wire  x739_x11_1_clock; // @[Math.scala 150:24:@35330.4]
  wire  x739_x11_1_reset; // @[Math.scala 150:24:@35330.4]
  wire [7:0] x739_x11_1_io_a; // @[Math.scala 150:24:@35330.4]
  wire [7:0] x739_x11_1_io_b; // @[Math.scala 150:24:@35330.4]
  wire  x739_x11_1_io_flow; // @[Math.scala 150:24:@35330.4]
  wire [7:0] x739_x11_1_io_result; // @[Math.scala 150:24:@35330.4]
  wire  x740_x12_1_clock; // @[Math.scala 150:24:@35340.4]
  wire  x740_x12_1_reset; // @[Math.scala 150:24:@35340.4]
  wire [7:0] x740_x12_1_io_a; // @[Math.scala 150:24:@35340.4]
  wire [7:0] x740_x12_1_io_b; // @[Math.scala 150:24:@35340.4]
  wire  x740_x12_1_io_flow; // @[Math.scala 150:24:@35340.4]
  wire [7:0] x740_x12_1_io_result; // @[Math.scala 150:24:@35340.4]
  wire  x741_x11_1_clock; // @[Math.scala 150:24:@35350.4]
  wire  x741_x11_1_reset; // @[Math.scala 150:24:@35350.4]
  wire [7:0] x741_x11_1_io_a; // @[Math.scala 150:24:@35350.4]
  wire [7:0] x741_x11_1_io_b; // @[Math.scala 150:24:@35350.4]
  wire  x741_x11_1_io_flow; // @[Math.scala 150:24:@35350.4]
  wire [7:0] x741_x11_1_io_result; // @[Math.scala 150:24:@35350.4]
  wire  x742_x12_1_clock; // @[Math.scala 150:24:@35360.4]
  wire  x742_x12_1_reset; // @[Math.scala 150:24:@35360.4]
  wire [7:0] x742_x12_1_io_a; // @[Math.scala 150:24:@35360.4]
  wire [7:0] x742_x12_1_io_b; // @[Math.scala 150:24:@35360.4]
  wire  x742_x12_1_io_flow; // @[Math.scala 150:24:@35360.4]
  wire [7:0] x742_x12_1_io_result; // @[Math.scala 150:24:@35360.4]
  wire [7:0] x743_x11_1_io_a; // @[Math.scala 150:24:@35370.4]
  wire [7:0] x743_x11_1_io_b; // @[Math.scala 150:24:@35370.4]
  wire [7:0] x743_x11_1_io_result; // @[Math.scala 150:24:@35370.4]
  wire [7:0] x744_x12_1_io_a; // @[Math.scala 150:24:@35380.4]
  wire [7:0] x744_x12_1_io_b; // @[Math.scala 150:24:@35380.4]
  wire [7:0] x744_x12_1_io_result; // @[Math.scala 150:24:@35380.4]
  wire [7:0] x745_x11_1_io_a; // @[Math.scala 150:24:@35390.4]
  wire [7:0] x745_x11_1_io_b; // @[Math.scala 150:24:@35390.4]
  wire [7:0] x745_x11_1_io_result; // @[Math.scala 150:24:@35390.4]
  wire  RetimeWrapper_102_clock; // @[package.scala 93:22:@35400.4]
  wire  RetimeWrapper_102_reset; // @[package.scala 93:22:@35400.4]
  wire  RetimeWrapper_102_io_flow; // @[package.scala 93:22:@35400.4]
  wire [7:0] RetimeWrapper_102_io_in; // @[package.scala 93:22:@35400.4]
  wire [7:0] RetimeWrapper_102_io_out; // @[package.scala 93:22:@35400.4]
  wire [7:0] x746_sum_1_io_a; // @[Math.scala 150:24:@35411.4]
  wire [7:0] x746_sum_1_io_b; // @[Math.scala 150:24:@35411.4]
  wire [7:0] x746_sum_1_io_result; // @[Math.scala 150:24:@35411.4]
  wire  RetimeWrapper_103_clock; // @[package.scala 93:22:@35425.4]
  wire  RetimeWrapper_103_reset; // @[package.scala 93:22:@35425.4]
  wire  RetimeWrapper_103_io_flow; // @[package.scala 93:22:@35425.4]
  wire [7:0] RetimeWrapper_103_io_in; // @[package.scala 93:22:@35425.4]
  wire [7:0] RetimeWrapper_103_io_out; // @[package.scala 93:22:@35425.4]
  wire  x752_x11_1_clock; // @[Math.scala 150:24:@35455.4]
  wire  x752_x11_1_reset; // @[Math.scala 150:24:@35455.4]
  wire [7:0] x752_x11_1_io_a; // @[Math.scala 150:24:@35455.4]
  wire [7:0] x752_x11_1_io_b; // @[Math.scala 150:24:@35455.4]
  wire  x752_x11_1_io_flow; // @[Math.scala 150:24:@35455.4]
  wire [7:0] x752_x11_1_io_result; // @[Math.scala 150:24:@35455.4]
  wire  x753_x12_1_clock; // @[Math.scala 150:24:@35465.4]
  wire  x753_x12_1_reset; // @[Math.scala 150:24:@35465.4]
  wire [7:0] x753_x12_1_io_a; // @[Math.scala 150:24:@35465.4]
  wire [7:0] x753_x12_1_io_b; // @[Math.scala 150:24:@35465.4]
  wire  x753_x12_1_io_flow; // @[Math.scala 150:24:@35465.4]
  wire [7:0] x753_x12_1_io_result; // @[Math.scala 150:24:@35465.4]
  wire  x754_x11_1_clock; // @[Math.scala 150:24:@35475.4]
  wire  x754_x11_1_reset; // @[Math.scala 150:24:@35475.4]
  wire [7:0] x754_x11_1_io_a; // @[Math.scala 150:24:@35475.4]
  wire [7:0] x754_x11_1_io_b; // @[Math.scala 150:24:@35475.4]
  wire  x754_x11_1_io_flow; // @[Math.scala 150:24:@35475.4]
  wire [7:0] x754_x11_1_io_result; // @[Math.scala 150:24:@35475.4]
  wire  x755_x12_1_clock; // @[Math.scala 150:24:@35485.4]
  wire  x755_x12_1_reset; // @[Math.scala 150:24:@35485.4]
  wire [7:0] x755_x12_1_io_a; // @[Math.scala 150:24:@35485.4]
  wire [7:0] x755_x12_1_io_b; // @[Math.scala 150:24:@35485.4]
  wire  x755_x12_1_io_flow; // @[Math.scala 150:24:@35485.4]
  wire [7:0] x755_x12_1_io_result; // @[Math.scala 150:24:@35485.4]
  wire [7:0] x756_x11_1_io_a; // @[Math.scala 150:24:@35495.4]
  wire [7:0] x756_x11_1_io_b; // @[Math.scala 150:24:@35495.4]
  wire [7:0] x756_x11_1_io_result; // @[Math.scala 150:24:@35495.4]
  wire [7:0] x757_x12_1_io_a; // @[Math.scala 150:24:@35505.4]
  wire [7:0] x757_x12_1_io_b; // @[Math.scala 150:24:@35505.4]
  wire [7:0] x757_x12_1_io_result; // @[Math.scala 150:24:@35505.4]
  wire [7:0] x758_x11_1_io_a; // @[Math.scala 150:24:@35515.4]
  wire [7:0] x758_x11_1_io_b; // @[Math.scala 150:24:@35515.4]
  wire [7:0] x758_x11_1_io_result; // @[Math.scala 150:24:@35515.4]
  wire  RetimeWrapper_104_clock; // @[package.scala 93:22:@35525.4]
  wire  RetimeWrapper_104_reset; // @[package.scala 93:22:@35525.4]
  wire  RetimeWrapper_104_io_flow; // @[package.scala 93:22:@35525.4]
  wire [7:0] RetimeWrapper_104_io_in; // @[package.scala 93:22:@35525.4]
  wire [7:0] RetimeWrapper_104_io_out; // @[package.scala 93:22:@35525.4]
  wire [7:0] x759_sum_1_io_a; // @[Math.scala 150:24:@35534.4]
  wire [7:0] x759_sum_1_io_b; // @[Math.scala 150:24:@35534.4]
  wire [7:0] x759_sum_1_io_result; // @[Math.scala 150:24:@35534.4]
  wire  RetimeWrapper_105_clock; // @[package.scala 93:22:@35548.4]
  wire  RetimeWrapper_105_reset; // @[package.scala 93:22:@35548.4]
  wire  RetimeWrapper_105_io_flow; // @[package.scala 93:22:@35548.4]
  wire [7:0] RetimeWrapper_105_io_in; // @[package.scala 93:22:@35548.4]
  wire [7:0] RetimeWrapper_105_io_out; // @[package.scala 93:22:@35548.4]
  wire  x765_x11_1_clock; // @[Math.scala 150:24:@35578.4]
  wire  x765_x11_1_reset; // @[Math.scala 150:24:@35578.4]
  wire [7:0] x765_x11_1_io_a; // @[Math.scala 150:24:@35578.4]
  wire [7:0] x765_x11_1_io_b; // @[Math.scala 150:24:@35578.4]
  wire  x765_x11_1_io_flow; // @[Math.scala 150:24:@35578.4]
  wire [7:0] x765_x11_1_io_result; // @[Math.scala 150:24:@35578.4]
  wire  x766_x12_1_clock; // @[Math.scala 150:24:@35588.4]
  wire  x766_x12_1_reset; // @[Math.scala 150:24:@35588.4]
  wire [7:0] x766_x12_1_io_a; // @[Math.scala 150:24:@35588.4]
  wire [7:0] x766_x12_1_io_b; // @[Math.scala 150:24:@35588.4]
  wire  x766_x12_1_io_flow; // @[Math.scala 150:24:@35588.4]
  wire [7:0] x766_x12_1_io_result; // @[Math.scala 150:24:@35588.4]
  wire  x767_x11_1_clock; // @[Math.scala 150:24:@35598.4]
  wire  x767_x11_1_reset; // @[Math.scala 150:24:@35598.4]
  wire [7:0] x767_x11_1_io_a; // @[Math.scala 150:24:@35598.4]
  wire [7:0] x767_x11_1_io_b; // @[Math.scala 150:24:@35598.4]
  wire  x767_x11_1_io_flow; // @[Math.scala 150:24:@35598.4]
  wire [7:0] x767_x11_1_io_result; // @[Math.scala 150:24:@35598.4]
  wire  x768_x12_1_clock; // @[Math.scala 150:24:@35608.4]
  wire  x768_x12_1_reset; // @[Math.scala 150:24:@35608.4]
  wire [7:0] x768_x12_1_io_a; // @[Math.scala 150:24:@35608.4]
  wire [7:0] x768_x12_1_io_b; // @[Math.scala 150:24:@35608.4]
  wire  x768_x12_1_io_flow; // @[Math.scala 150:24:@35608.4]
  wire [7:0] x768_x12_1_io_result; // @[Math.scala 150:24:@35608.4]
  wire [7:0] x769_x11_1_io_a; // @[Math.scala 150:24:@35618.4]
  wire [7:0] x769_x11_1_io_b; // @[Math.scala 150:24:@35618.4]
  wire [7:0] x769_x11_1_io_result; // @[Math.scala 150:24:@35618.4]
  wire [7:0] x770_x12_1_io_a; // @[Math.scala 150:24:@35628.4]
  wire [7:0] x770_x12_1_io_b; // @[Math.scala 150:24:@35628.4]
  wire [7:0] x770_x12_1_io_result; // @[Math.scala 150:24:@35628.4]
  wire [7:0] x771_x11_1_io_a; // @[Math.scala 150:24:@35638.4]
  wire [7:0] x771_x11_1_io_b; // @[Math.scala 150:24:@35638.4]
  wire [7:0] x771_x11_1_io_result; // @[Math.scala 150:24:@35638.4]
  wire  RetimeWrapper_106_clock; // @[package.scala 93:22:@35648.4]
  wire  RetimeWrapper_106_reset; // @[package.scala 93:22:@35648.4]
  wire  RetimeWrapper_106_io_flow; // @[package.scala 93:22:@35648.4]
  wire [7:0] RetimeWrapper_106_io_in; // @[package.scala 93:22:@35648.4]
  wire [7:0] RetimeWrapper_106_io_out; // @[package.scala 93:22:@35648.4]
  wire [7:0] x772_sum_1_io_a; // @[Math.scala 150:24:@35657.4]
  wire [7:0] x772_sum_1_io_b; // @[Math.scala 150:24:@35657.4]
  wire [7:0] x772_sum_1_io_result; // @[Math.scala 150:24:@35657.4]
  wire  RetimeWrapper_107_clock; // @[package.scala 93:22:@35671.4]
  wire  RetimeWrapper_107_reset; // @[package.scala 93:22:@35671.4]
  wire  RetimeWrapper_107_io_flow; // @[package.scala 93:22:@35671.4]
  wire [7:0] RetimeWrapper_107_io_in; // @[package.scala 93:22:@35671.4]
  wire [7:0] RetimeWrapper_107_io_out; // @[package.scala 93:22:@35671.4]
  wire  x777_x11_1_clock; // @[Math.scala 150:24:@35696.4]
  wire  x777_x11_1_reset; // @[Math.scala 150:24:@35696.4]
  wire [7:0] x777_x11_1_io_a; // @[Math.scala 150:24:@35696.4]
  wire [7:0] x777_x11_1_io_b; // @[Math.scala 150:24:@35696.4]
  wire  x777_x11_1_io_flow; // @[Math.scala 150:24:@35696.4]
  wire [7:0] x777_x11_1_io_result; // @[Math.scala 150:24:@35696.4]
  wire  x778_x12_1_clock; // @[Math.scala 150:24:@35706.4]
  wire  x778_x12_1_reset; // @[Math.scala 150:24:@35706.4]
  wire [7:0] x778_x12_1_io_a; // @[Math.scala 150:24:@35706.4]
  wire [7:0] x778_x12_1_io_b; // @[Math.scala 150:24:@35706.4]
  wire  x778_x12_1_io_flow; // @[Math.scala 150:24:@35706.4]
  wire [7:0] x778_x12_1_io_result; // @[Math.scala 150:24:@35706.4]
  wire  x779_x11_1_clock; // @[Math.scala 150:24:@35716.4]
  wire  x779_x11_1_reset; // @[Math.scala 150:24:@35716.4]
  wire [7:0] x779_x11_1_io_a; // @[Math.scala 150:24:@35716.4]
  wire [7:0] x779_x11_1_io_b; // @[Math.scala 150:24:@35716.4]
  wire  x779_x11_1_io_flow; // @[Math.scala 150:24:@35716.4]
  wire [7:0] x779_x11_1_io_result; // @[Math.scala 150:24:@35716.4]
  wire  x780_x12_1_clock; // @[Math.scala 150:24:@35726.4]
  wire  x780_x12_1_reset; // @[Math.scala 150:24:@35726.4]
  wire [7:0] x780_x12_1_io_a; // @[Math.scala 150:24:@35726.4]
  wire [7:0] x780_x12_1_io_b; // @[Math.scala 150:24:@35726.4]
  wire  x780_x12_1_io_flow; // @[Math.scala 150:24:@35726.4]
  wire [7:0] x780_x12_1_io_result; // @[Math.scala 150:24:@35726.4]
  wire [7:0] x781_x11_1_io_a; // @[Math.scala 150:24:@35736.4]
  wire [7:0] x781_x11_1_io_b; // @[Math.scala 150:24:@35736.4]
  wire [7:0] x781_x11_1_io_result; // @[Math.scala 150:24:@35736.4]
  wire [7:0] x782_x12_1_io_a; // @[Math.scala 150:24:@35746.4]
  wire [7:0] x782_x12_1_io_b; // @[Math.scala 150:24:@35746.4]
  wire [7:0] x782_x12_1_io_result; // @[Math.scala 150:24:@35746.4]
  wire [7:0] x783_x11_1_io_a; // @[Math.scala 150:24:@35756.4]
  wire [7:0] x783_x11_1_io_b; // @[Math.scala 150:24:@35756.4]
  wire [7:0] x783_x11_1_io_result; // @[Math.scala 150:24:@35756.4]
  wire  RetimeWrapper_108_clock; // @[package.scala 93:22:@35766.4]
  wire  RetimeWrapper_108_reset; // @[package.scala 93:22:@35766.4]
  wire  RetimeWrapper_108_io_flow; // @[package.scala 93:22:@35766.4]
  wire [7:0] RetimeWrapper_108_io_in; // @[package.scala 93:22:@35766.4]
  wire [7:0] RetimeWrapper_108_io_out; // @[package.scala 93:22:@35766.4]
  wire [7:0] x784_sum_1_io_a; // @[Math.scala 150:24:@35775.4]
  wire [7:0] x784_sum_1_io_b; // @[Math.scala 150:24:@35775.4]
  wire [7:0] x784_sum_1_io_result; // @[Math.scala 150:24:@35775.4]
  wire  RetimeWrapper_109_clock; // @[package.scala 93:22:@35789.4]
  wire  RetimeWrapper_109_reset; // @[package.scala 93:22:@35789.4]
  wire  RetimeWrapper_109_io_flow; // @[package.scala 93:22:@35789.4]
  wire [7:0] RetimeWrapper_109_io_in; // @[package.scala 93:22:@35789.4]
  wire [7:0] RetimeWrapper_109_io_out; // @[package.scala 93:22:@35789.4]
  wire  x788_x11_1_clock; // @[Math.scala 150:24:@35809.4]
  wire  x788_x11_1_reset; // @[Math.scala 150:24:@35809.4]
  wire [7:0] x788_x11_1_io_a; // @[Math.scala 150:24:@35809.4]
  wire [7:0] x788_x11_1_io_b; // @[Math.scala 150:24:@35809.4]
  wire  x788_x11_1_io_flow; // @[Math.scala 150:24:@35809.4]
  wire [7:0] x788_x11_1_io_result; // @[Math.scala 150:24:@35809.4]
  wire  x789_x12_1_clock; // @[Math.scala 150:24:@35819.4]
  wire  x789_x12_1_reset; // @[Math.scala 150:24:@35819.4]
  wire [7:0] x789_x12_1_io_a; // @[Math.scala 150:24:@35819.4]
  wire [7:0] x789_x12_1_io_b; // @[Math.scala 150:24:@35819.4]
  wire  x789_x12_1_io_flow; // @[Math.scala 150:24:@35819.4]
  wire [7:0] x789_x12_1_io_result; // @[Math.scala 150:24:@35819.4]
  wire  x790_x11_1_clock; // @[Math.scala 150:24:@35829.4]
  wire  x790_x11_1_reset; // @[Math.scala 150:24:@35829.4]
  wire [7:0] x790_x11_1_io_a; // @[Math.scala 150:24:@35829.4]
  wire [7:0] x790_x11_1_io_b; // @[Math.scala 150:24:@35829.4]
  wire  x790_x11_1_io_flow; // @[Math.scala 150:24:@35829.4]
  wire [7:0] x790_x11_1_io_result; // @[Math.scala 150:24:@35829.4]
  wire  x791_x12_1_clock; // @[Math.scala 150:24:@35841.4]
  wire  x791_x12_1_reset; // @[Math.scala 150:24:@35841.4]
  wire [7:0] x791_x12_1_io_a; // @[Math.scala 150:24:@35841.4]
  wire [7:0] x791_x12_1_io_b; // @[Math.scala 150:24:@35841.4]
  wire  x791_x12_1_io_flow; // @[Math.scala 150:24:@35841.4]
  wire [7:0] x791_x12_1_io_result; // @[Math.scala 150:24:@35841.4]
  wire [7:0] x792_x11_1_io_a; // @[Math.scala 150:24:@35851.4]
  wire [7:0] x792_x11_1_io_b; // @[Math.scala 150:24:@35851.4]
  wire [7:0] x792_x11_1_io_result; // @[Math.scala 150:24:@35851.4]
  wire [7:0] x793_x12_1_io_a; // @[Math.scala 150:24:@35861.4]
  wire [7:0] x793_x12_1_io_b; // @[Math.scala 150:24:@35861.4]
  wire [7:0] x793_x12_1_io_result; // @[Math.scala 150:24:@35861.4]
  wire [7:0] x794_x11_1_io_a; // @[Math.scala 150:24:@35871.4]
  wire [7:0] x794_x11_1_io_b; // @[Math.scala 150:24:@35871.4]
  wire [7:0] x794_x11_1_io_result; // @[Math.scala 150:24:@35871.4]
  wire  RetimeWrapper_110_clock; // @[package.scala 93:22:@35881.4]
  wire  RetimeWrapper_110_reset; // @[package.scala 93:22:@35881.4]
  wire  RetimeWrapper_110_io_flow; // @[package.scala 93:22:@35881.4]
  wire [7:0] RetimeWrapper_110_io_in; // @[package.scala 93:22:@35881.4]
  wire [7:0] RetimeWrapper_110_io_out; // @[package.scala 93:22:@35881.4]
  wire [7:0] x795_sum_1_io_a; // @[Math.scala 150:24:@35890.4]
  wire [7:0] x795_sum_1_io_b; // @[Math.scala 150:24:@35890.4]
  wire [7:0] x795_sum_1_io_result; // @[Math.scala 150:24:@35890.4]
  wire  RetimeWrapper_111_clock; // @[package.scala 93:22:@35904.4]
  wire  RetimeWrapper_111_reset; // @[package.scala 93:22:@35904.4]
  wire  RetimeWrapper_111_io_flow; // @[package.scala 93:22:@35904.4]
  wire [7:0] RetimeWrapper_111_io_in; // @[package.scala 93:22:@35904.4]
  wire [7:0] RetimeWrapper_111_io_out; // @[package.scala 93:22:@35904.4]
  wire  x799_x11_1_clock; // @[Math.scala 150:24:@35924.4]
  wire  x799_x11_1_reset; // @[Math.scala 150:24:@35924.4]
  wire [7:0] x799_x11_1_io_a; // @[Math.scala 150:24:@35924.4]
  wire [7:0] x799_x11_1_io_b; // @[Math.scala 150:24:@35924.4]
  wire  x799_x11_1_io_flow; // @[Math.scala 150:24:@35924.4]
  wire [7:0] x799_x11_1_io_result; // @[Math.scala 150:24:@35924.4]
  wire  x800_x12_1_clock; // @[Math.scala 150:24:@35934.4]
  wire  x800_x12_1_reset; // @[Math.scala 150:24:@35934.4]
  wire [7:0] x800_x12_1_io_a; // @[Math.scala 150:24:@35934.4]
  wire [7:0] x800_x12_1_io_b; // @[Math.scala 150:24:@35934.4]
  wire  x800_x12_1_io_flow; // @[Math.scala 150:24:@35934.4]
  wire [7:0] x800_x12_1_io_result; // @[Math.scala 150:24:@35934.4]
  wire  x801_x11_1_clock; // @[Math.scala 150:24:@35944.4]
  wire  x801_x11_1_reset; // @[Math.scala 150:24:@35944.4]
  wire [7:0] x801_x11_1_io_a; // @[Math.scala 150:24:@35944.4]
  wire [7:0] x801_x11_1_io_b; // @[Math.scala 150:24:@35944.4]
  wire  x801_x11_1_io_flow; // @[Math.scala 150:24:@35944.4]
  wire [7:0] x801_x11_1_io_result; // @[Math.scala 150:24:@35944.4]
  wire  x802_x12_1_clock; // @[Math.scala 150:24:@35954.4]
  wire  x802_x12_1_reset; // @[Math.scala 150:24:@35954.4]
  wire [7:0] x802_x12_1_io_a; // @[Math.scala 150:24:@35954.4]
  wire [7:0] x802_x12_1_io_b; // @[Math.scala 150:24:@35954.4]
  wire  x802_x12_1_io_flow; // @[Math.scala 150:24:@35954.4]
  wire [7:0] x802_x12_1_io_result; // @[Math.scala 150:24:@35954.4]
  wire [7:0] x803_x11_1_io_a; // @[Math.scala 150:24:@35964.4]
  wire [7:0] x803_x11_1_io_b; // @[Math.scala 150:24:@35964.4]
  wire [7:0] x803_x11_1_io_result; // @[Math.scala 150:24:@35964.4]
  wire [7:0] x804_x12_1_io_a; // @[Math.scala 150:24:@35974.4]
  wire [7:0] x804_x12_1_io_b; // @[Math.scala 150:24:@35974.4]
  wire [7:0] x804_x12_1_io_result; // @[Math.scala 150:24:@35974.4]
  wire [7:0] x805_x11_1_io_a; // @[Math.scala 150:24:@35984.4]
  wire [7:0] x805_x11_1_io_b; // @[Math.scala 150:24:@35984.4]
  wire [7:0] x805_x11_1_io_result; // @[Math.scala 150:24:@35984.4]
  wire  RetimeWrapper_112_clock; // @[package.scala 93:22:@35994.4]
  wire  RetimeWrapper_112_reset; // @[package.scala 93:22:@35994.4]
  wire  RetimeWrapper_112_io_flow; // @[package.scala 93:22:@35994.4]
  wire [7:0] RetimeWrapper_112_io_in; // @[package.scala 93:22:@35994.4]
  wire [7:0] RetimeWrapper_112_io_out; // @[package.scala 93:22:@35994.4]
  wire [7:0] x806_sum_1_io_a; // @[Math.scala 150:24:@36003.4]
  wire [7:0] x806_sum_1_io_b; // @[Math.scala 150:24:@36003.4]
  wire [7:0] x806_sum_1_io_result; // @[Math.scala 150:24:@36003.4]
  wire  RetimeWrapper_113_clock; // @[package.scala 93:22:@36017.4]
  wire  RetimeWrapper_113_reset; // @[package.scala 93:22:@36017.4]
  wire  RetimeWrapper_113_io_flow; // @[package.scala 93:22:@36017.4]
  wire [7:0] RetimeWrapper_113_io_in; // @[package.scala 93:22:@36017.4]
  wire [7:0] RetimeWrapper_113_io_out; // @[package.scala 93:22:@36017.4]
  wire  x811_x11_1_clock; // @[Math.scala 150:24:@36042.4]
  wire  x811_x11_1_reset; // @[Math.scala 150:24:@36042.4]
  wire [7:0] x811_x11_1_io_a; // @[Math.scala 150:24:@36042.4]
  wire [7:0] x811_x11_1_io_b; // @[Math.scala 150:24:@36042.4]
  wire  x811_x11_1_io_flow; // @[Math.scala 150:24:@36042.4]
  wire [7:0] x811_x11_1_io_result; // @[Math.scala 150:24:@36042.4]
  wire  x812_x12_1_clock; // @[Math.scala 150:24:@36052.4]
  wire  x812_x12_1_reset; // @[Math.scala 150:24:@36052.4]
  wire [7:0] x812_x12_1_io_a; // @[Math.scala 150:24:@36052.4]
  wire [7:0] x812_x12_1_io_b; // @[Math.scala 150:24:@36052.4]
  wire  x812_x12_1_io_flow; // @[Math.scala 150:24:@36052.4]
  wire [7:0] x812_x12_1_io_result; // @[Math.scala 150:24:@36052.4]
  wire  x813_x11_1_clock; // @[Math.scala 150:24:@36062.4]
  wire  x813_x11_1_reset; // @[Math.scala 150:24:@36062.4]
  wire [7:0] x813_x11_1_io_a; // @[Math.scala 150:24:@36062.4]
  wire [7:0] x813_x11_1_io_b; // @[Math.scala 150:24:@36062.4]
  wire  x813_x11_1_io_flow; // @[Math.scala 150:24:@36062.4]
  wire [7:0] x813_x11_1_io_result; // @[Math.scala 150:24:@36062.4]
  wire  x814_x12_1_clock; // @[Math.scala 150:24:@36072.4]
  wire  x814_x12_1_reset; // @[Math.scala 150:24:@36072.4]
  wire [7:0] x814_x12_1_io_a; // @[Math.scala 150:24:@36072.4]
  wire [7:0] x814_x12_1_io_b; // @[Math.scala 150:24:@36072.4]
  wire  x814_x12_1_io_flow; // @[Math.scala 150:24:@36072.4]
  wire [7:0] x814_x12_1_io_result; // @[Math.scala 150:24:@36072.4]
  wire [7:0] x815_x11_1_io_a; // @[Math.scala 150:24:@36082.4]
  wire [7:0] x815_x11_1_io_b; // @[Math.scala 150:24:@36082.4]
  wire [7:0] x815_x11_1_io_result; // @[Math.scala 150:24:@36082.4]
  wire [7:0] x816_x12_1_io_a; // @[Math.scala 150:24:@36092.4]
  wire [7:0] x816_x12_1_io_b; // @[Math.scala 150:24:@36092.4]
  wire [7:0] x816_x12_1_io_result; // @[Math.scala 150:24:@36092.4]
  wire [7:0] x817_x11_1_io_a; // @[Math.scala 150:24:@36102.4]
  wire [7:0] x817_x11_1_io_b; // @[Math.scala 150:24:@36102.4]
  wire [7:0] x817_x11_1_io_result; // @[Math.scala 150:24:@36102.4]
  wire  RetimeWrapper_114_clock; // @[package.scala 93:22:@36112.4]
  wire  RetimeWrapper_114_reset; // @[package.scala 93:22:@36112.4]
  wire  RetimeWrapper_114_io_flow; // @[package.scala 93:22:@36112.4]
  wire [7:0] RetimeWrapper_114_io_in; // @[package.scala 93:22:@36112.4]
  wire [7:0] RetimeWrapper_114_io_out; // @[package.scala 93:22:@36112.4]
  wire [7:0] x818_sum_1_io_a; // @[Math.scala 150:24:@36121.4]
  wire [7:0] x818_sum_1_io_b; // @[Math.scala 150:24:@36121.4]
  wire [7:0] x818_sum_1_io_result; // @[Math.scala 150:24:@36121.4]
  wire  RetimeWrapper_115_clock; // @[package.scala 93:22:@36135.4]
  wire  RetimeWrapper_115_reset; // @[package.scala 93:22:@36135.4]
  wire  RetimeWrapper_115_io_flow; // @[package.scala 93:22:@36135.4]
  wire [7:0] RetimeWrapper_115_io_in; // @[package.scala 93:22:@36135.4]
  wire [7:0] RetimeWrapper_115_io_out; // @[package.scala 93:22:@36135.4]
  wire  RetimeWrapper_116_clock; // @[package.scala 93:22:@36163.4]
  wire  RetimeWrapper_116_reset; // @[package.scala 93:22:@36163.4]
  wire  RetimeWrapper_116_io_flow; // @[package.scala 93:22:@36163.4]
  wire [63:0] RetimeWrapper_116_io_in; // @[package.scala 93:22:@36163.4]
  wire [63:0] RetimeWrapper_116_io_out; // @[package.scala 93:22:@36163.4]
  wire  RetimeWrapper_117_clock; // @[package.scala 93:22:@36172.4]
  wire  RetimeWrapper_117_reset; // @[package.scala 93:22:@36172.4]
  wire  RetimeWrapper_117_io_flow; // @[package.scala 93:22:@36172.4]
  wire  RetimeWrapper_117_io_in; // @[package.scala 93:22:@36172.4]
  wire  RetimeWrapper_117_io_out; // @[package.scala 93:22:@36172.4]
  wire  RetimeWrapper_118_clock; // @[package.scala 93:22:@36181.4]
  wire  RetimeWrapper_118_reset; // @[package.scala 93:22:@36181.4]
  wire  RetimeWrapper_118_io_flow; // @[package.scala 93:22:@36181.4]
  wire  RetimeWrapper_118_io_in; // @[package.scala 93:22:@36181.4]
  wire  RetimeWrapper_118_io_out; // @[package.scala 93:22:@36181.4]
  wire  RetimeWrapper_119_clock; // @[package.scala 93:22:@36190.4]
  wire  RetimeWrapper_119_reset; // @[package.scala 93:22:@36190.4]
  wire  RetimeWrapper_119_io_flow; // @[package.scala 93:22:@36190.4]
  wire  RetimeWrapper_119_io_in; // @[package.scala 93:22:@36190.4]
  wire  RetimeWrapper_119_io_out; // @[package.scala 93:22:@36190.4]
  wire  b437; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 62:18:@32524.4]
  wire  b438; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 63:18:@32525.4]
  wire  _T_206; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 68:30:@32740.4]
  wire  _T_207; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 68:37:@32741.4]
  wire  _T_211; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 70:76:@32746.4]
  wire  _T_212; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 70:62:@32747.4]
  wire  _T_214; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 70:101:@32748.4]
  wire [63:0] x902_x440_D1_0_number; // @[package.scala 96:25:@32757.4 package.scala 96:25:@32758.4]
  wire [31:0] b435_number; // @[Math.scala 712:22:@32509.4 Math.scala 713:14:@32510.4]
  wire [31:0] _T_254; // @[Math.scala 499:52:@32785.4]
  wire  x444; // @[Math.scala 499:44:@32793.4]
  wire  x445; // @[Math.scala 499:44:@32800.4]
  wire  x446; // @[Math.scala 499:44:@32807.4]
  wire [31:0] _T_301; // @[Mux.scala 19:72:@32819.4]
  wire [31:0] _T_303; // @[Mux.scala 19:72:@32820.4]
  wire [31:0] _T_305; // @[Mux.scala 19:72:@32821.4]
  wire [31:0] _T_307; // @[Mux.scala 19:72:@32823.4]
  wire [31:0] x447_number; // @[Mux.scala 19:72:@32824.4]
  wire [31:0] _T_319; // @[Math.scala 406:49:@32834.4]
  wire [31:0] _T_321; // @[Math.scala 406:56:@32836.4]
  wire [31:0] _T_322; // @[Math.scala 406:56:@32837.4]
  wire  _T_327; // @[FixedPoint.scala 50:25:@32843.4]
  wire [1:0] _T_331; // @[Bitwise.scala 72:12:@32845.4]
  wire [29:0] _T_332; // @[FixedPoint.scala 18:52:@32846.4]
  wire [31:0] b436_number; // @[Math.scala 712:22:@32521.4 Math.scala 713:14:@32522.4]
  wire  _T_337; // @[FixedPoint.scala 50:25:@32852.4]
  wire [1:0] _T_341; // @[Bitwise.scala 72:12:@32854.4]
  wire [29:0] _T_342; // @[FixedPoint.scala 18:52:@32855.4]
  wire  _T_367; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 113:101:@32916.4]
  wire  _T_371; // @[package.scala 96:25:@32924.4 package.scala 96:25:@32925.4]
  wire  _T_373; // @[implicits.scala 55:10:@32926.4]
  wire  _T_374; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 113:118:@32927.4]
  wire  _T_376; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 113:205:@32929.4]
  wire  _T_377; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 113:224:@32930.4]
  wire  x907_b437_D8; // @[package.scala 96:25:@32911.4 package.scala 96:25:@32912.4]
  wire  _T_378; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 113:250:@32931.4]
  wire  x906_b438_D8; // @[package.scala 96:25:@32902.4 package.scala 96:25:@32903.4]
  wire [31:0] x459_rdcol_number; // @[Math.scala 154:22:@32948.4 Math.scala 155:14:@32949.4]
  wire  _T_391; // @[FixedPoint.scala 50:25:@32955.4]
  wire [1:0] _T_395; // @[Bitwise.scala 72:12:@32957.4]
  wire [29:0] _T_396; // @[FixedPoint.scala 18:52:@32958.4]
  wire  _T_419; // @[package.scala 96:25:@33009.4 package.scala 96:25:@33010.4]
  wire  _T_421; // @[implicits.scala 55:10:@33011.4]
  wire  _T_422; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 132:118:@33012.4]
  wire  _T_424; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 132:205:@33014.4]
  wire  _T_425; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 132:224:@33015.4]
  wire  _T_426; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 132:250:@33016.4]
  wire [31:0] x468_rdcol_number; // @[Math.scala 154:22:@33033.4 Math.scala 155:14:@33034.4]
  wire  _T_439; // @[FixedPoint.scala 50:25:@33040.4]
  wire [1:0] _T_443; // @[Bitwise.scala 72:12:@33042.4]
  wire [29:0] _T_444; // @[FixedPoint.scala 18:52:@33043.4]
  wire  _T_464; // @[package.scala 96:25:@33085.4 package.scala 96:25:@33086.4]
  wire  _T_466; // @[implicits.scala 55:10:@33087.4]
  wire  _T_467; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 149:118:@33088.4]
  wire  _T_469; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 149:205:@33090.4]
  wire  _T_470; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 149:224:@33091.4]
  wire  _T_471; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 149:250:@33092.4]
  wire [31:0] x477_rdcol_number; // @[Math.scala 154:22:@33109.4 Math.scala 155:14:@33110.4]
  wire  _T_484; // @[FixedPoint.scala 50:25:@33116.4]
  wire [1:0] _T_488; // @[Bitwise.scala 72:12:@33118.4]
  wire [29:0] _T_489; // @[FixedPoint.scala 18:52:@33119.4]
  wire  _T_509; // @[package.scala 96:25:@33161.4 package.scala 96:25:@33162.4]
  wire  _T_511; // @[implicits.scala 55:10:@33163.4]
  wire  _T_512; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 166:118:@33164.4]
  wire  _T_514; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 166:205:@33166.4]
  wire  _T_515; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 166:224:@33167.4]
  wire  _T_516; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 166:250:@33168.4]
  wire [31:0] x486_rdrow_number; // @[Math.scala 154:22:@33185.4 Math.scala 155:14:@33186.4]
  wire [31:0] _T_531; // @[Math.scala 499:52:@33192.4]
  wire  x488; // @[Math.scala 499:44:@33200.4]
  wire  x489; // @[Math.scala 499:44:@33207.4]
  wire  x490; // @[Math.scala 499:44:@33214.4]
  wire [31:0] _T_578; // @[Mux.scala 19:72:@33226.4]
  wire [31:0] _T_580; // @[Mux.scala 19:72:@33227.4]
  wire [31:0] _T_582; // @[Mux.scala 19:72:@33228.4]
  wire [31:0] _T_584; // @[Mux.scala 19:72:@33230.4]
  wire [31:0] x491_number; // @[Mux.scala 19:72:@33231.4]
  wire [31:0] _T_598; // @[Math.scala 406:49:@33243.4]
  wire [31:0] _T_600; // @[Math.scala 406:56:@33245.4]
  wire [31:0] _T_601; // @[Math.scala 406:56:@33246.4]
  wire  _T_606; // @[FixedPoint.scala 50:25:@33252.4]
  wire [1:0] _T_610; // @[Bitwise.scala 72:12:@33254.4]
  wire [29:0] _T_611; // @[FixedPoint.scala 18:52:@33255.4]
  wire  _T_637; // @[package.scala 96:25:@33315.4 package.scala 96:25:@33316.4]
  wire  _T_639; // @[implicits.scala 55:10:@33317.4]
  wire  _T_640; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 207:166:@33318.4]
  wire  _T_642; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 207:253:@33320.4]
  wire  _T_643; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 207:272:@33321.4]
  wire  _T_644; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 207:298:@33322.4]
  wire  _T_665; // @[package.scala 96:25:@33370.4 package.scala 96:25:@33371.4]
  wire  _T_667; // @[implicits.scala 55:10:@33372.4]
  wire  _T_668; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 220:166:@33373.4]
  wire  _T_670; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 220:253:@33375.4]
  wire  _T_671; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 220:272:@33376.4]
  wire  _T_672; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 220:298:@33377.4]
  wire  _T_693; // @[package.scala 96:25:@33425.4 package.scala 96:25:@33426.4]
  wire  _T_695; // @[implicits.scala 55:10:@33427.4]
  wire  _T_696; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 233:166:@33428.4]
  wire  _T_698; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 233:253:@33430.4]
  wire  _T_699; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 233:272:@33431.4]
  wire  _T_700; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 233:298:@33432.4]
  wire  _T_721; // @[package.scala 96:25:@33480.4 package.scala 96:25:@33481.4]
  wire  _T_723; // @[implicits.scala 55:10:@33482.4]
  wire  _T_724; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 246:166:@33483.4]
  wire  _T_726; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 246:253:@33485.4]
  wire  _T_727; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 246:272:@33486.4]
  wire  _T_728; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 246:298:@33487.4]
  wire [31:0] x925_x486_rdrow_D10_number; // @[package.scala 96:25:@33501.4 package.scala 96:25:@33502.4]
  wire [31:0] _T_740; // @[Math.scala 406:49:@33508.4]
  wire [31:0] _T_742; // @[Math.scala 406:56:@33510.4]
  wire [31:0] _T_743; // @[Math.scala 406:56:@33511.4]
  wire [31:0] x894_number; // @[implicits.scala 133:21:@33512.4]
  wire  x517; // @[Math.scala 465:44:@33520.4]
  wire [31:0] x926_x477_rdcol_D10_number; // @[package.scala 96:25:@33528.4 package.scala 96:25:@33529.4]
  wire [31:0] _T_761; // @[Math.scala 465:37:@33534.4]
  wire  x518; // @[Math.scala 465:44:@33536.4]
  wire  x519; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 259:24:@33539.4]
  wire [31:0] _T_775; // @[Math.scala 406:49:@33548.4]
  wire [31:0] _T_777; // @[Math.scala 406:56:@33550.4]
  wire [31:0] _T_778; // @[Math.scala 406:56:@33551.4]
  wire  _T_783; // @[FixedPoint.scala 50:25:@33557.4]
  wire [1:0] _T_787; // @[Bitwise.scala 72:12:@33559.4]
  wire [29:0] _T_788; // @[FixedPoint.scala 18:52:@33560.4]
  wire  _T_823; // @[package.scala 96:25:@33630.4 package.scala 96:25:@33631.4]
  wire  _T_825; // @[implicits.scala 55:10:@33632.4]
  wire  _T_826; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 282:194:@33633.4]
  wire  x928_x520_D1; // @[package.scala 96:25:@33589.4 package.scala 96:25:@33590.4]
  wire  _T_827; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 282:282:@33634.4]
  wire  x931_b437_D12; // @[package.scala 96:25:@33616.4 package.scala 96:25:@33617.4]
  wire  _T_828; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 282:290:@33635.4]
  wire  x930_b438_D12; // @[package.scala 96:25:@33607.4 package.scala 96:25:@33608.4]
  wire [31:0] x932_x468_rdcol_D10_number; // @[package.scala 96:25:@33651.4 package.scala 96:25:@33652.4]
  wire [31:0] _T_839; // @[Math.scala 465:37:@33657.4]
  wire  x529; // @[Math.scala 465:44:@33659.4]
  wire  x530; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 290:24:@33662.4]
  wire  _T_870; // @[package.scala 96:25:@33706.4 package.scala 96:25:@33707.4]
  wire  _T_872; // @[implicits.scala 55:10:@33708.4]
  wire  _T_873; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 309:194:@33709.4]
  wire  x934_x531_D1; // @[package.scala 96:25:@33692.4 package.scala 96:25:@33693.4]
  wire  _T_874; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 309:282:@33710.4]
  wire  _T_875; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 309:325:@33711.4]
  wire [31:0] x935_x459_rdcol_D10_number; // @[package.scala 96:25:@33727.4 package.scala 96:25:@33728.4]
  wire [31:0] _T_888; // @[Math.scala 465:37:@33735.4]
  wire  x537; // @[Math.scala 465:44:@33737.4]
  wire  x538; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 319:59:@33740.4]
  wire  _T_919; // @[package.scala 96:25:@33784.4 package.scala 96:25:@33785.4]
  wire  _T_921; // @[implicits.scala 55:10:@33786.4]
  wire  _T_922; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 332:194:@33787.4]
  wire  x937_x539_D1; // @[package.scala 96:25:@33770.4 package.scala 96:25:@33771.4]
  wire  _T_923; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 332:282:@33788.4]
  wire  _T_924; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 332:290:@33789.4]
  wire [31:0] x938_b436_D10_number; // @[package.scala 96:25:@33805.4 package.scala 96:25:@33806.4]
  wire [31:0] _T_935; // @[Math.scala 465:37:@33811.4]
  wire  x545; // @[Math.scala 465:44:@33813.4]
  wire  x939_x545_D1; // @[package.scala 96:25:@33821.4 package.scala 96:25:@33822.4]
  wire  x546; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 342:59:@33825.4]
  wire  _T_969; // @[package.scala 96:25:@33869.4 package.scala 96:25:@33870.4]
  wire  _T_971; // @[implicits.scala 55:10:@33871.4]
  wire  _T_972; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 355:194:@33872.4]
  wire  x941_x547_D1; // @[package.scala 96:25:@33855.4 package.scala 96:25:@33856.4]
  wire  _T_973; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 355:282:@33873.4]
  wire  _T_974; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 355:290:@33874.4]
  wire [31:0] x553_rdcol_number; // @[Math.scala 154:22:@33893.4 Math.scala 155:14:@33894.4]
  wire [31:0] _T_989; // @[Math.scala 465:37:@33899.4]
  wire  x554; // @[Math.scala 465:44:@33901.4]
  wire  x555; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 363:59:@33904.4]
  wire  _T_999; // @[FixedPoint.scala 50:25:@33911.4]
  wire [1:0] _T_1003; // @[Bitwise.scala 72:12:@33913.4]
  wire [29:0] _T_1004; // @[FixedPoint.scala 18:52:@33914.4]
  wire  _T_1027; // @[package.scala 96:25:@33948.4 package.scala 96:25:@33949.4]
  wire  _T_1029; // @[implicits.scala 55:10:@33950.4]
  wire  _T_1030; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 376:194:@33951.4]
  wire  x942_x556_D1; // @[package.scala 96:25:@33934.4 package.scala 96:25:@33935.4]
  wire  _T_1031; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 376:282:@33952.4]
  wire  _T_1032; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 376:290:@33953.4]
  wire [31:0] x565_rdcol_number; // @[Math.scala 154:22:@33972.4 Math.scala 155:14:@33973.4]
  wire [31:0] _T_1047; // @[Math.scala 465:37:@33978.4]
  wire  x566; // @[Math.scala 465:44:@33980.4]
  wire  x567; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 384:59:@33983.4]
  wire  _T_1057; // @[FixedPoint.scala 50:25:@33990.4]
  wire [1:0] _T_1061; // @[Bitwise.scala 72:12:@33992.4]
  wire [29:0] _T_1062; // @[FixedPoint.scala 18:52:@33993.4]
  wire  _T_1085; // @[package.scala 96:25:@34027.4 package.scala 96:25:@34028.4]
  wire  _T_1087; // @[implicits.scala 55:10:@34029.4]
  wire  _T_1088; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 397:194:@34030.4]
  wire  x943_x568_D1; // @[package.scala 96:25:@34013.4 package.scala 96:25:@34014.4]
  wire  _T_1089; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 397:282:@34031.4]
  wire  _T_1090; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 397:290:@34032.4]
  wire [31:0] x944_b435_D10_number; // @[package.scala 96:25:@34048.4 package.scala 96:25:@34049.4]
  wire [31:0] _T_1103; // @[Math.scala 406:49:@34055.4]
  wire [31:0] _T_1105; // @[Math.scala 406:56:@34057.4]
  wire [31:0] _T_1106; // @[Math.scala 406:56:@34058.4]
  wire [31:0] x896_number; // @[implicits.scala 133:21:@34059.4]
  wire  x578; // @[Math.scala 465:44:@34067.4]
  wire  x945_x578_D1; // @[package.scala 96:25:@34075.4 package.scala 96:25:@34076.4]
  wire  x579; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 409:24:@34079.4]
  wire [31:0] _T_1130; // @[Math.scala 406:49:@34088.4]
  wire [31:0] _T_1132; // @[Math.scala 406:56:@34090.4]
  wire [31:0] _T_1133; // @[Math.scala 406:56:@34091.4]
  wire  _T_1138; // @[FixedPoint.scala 50:25:@34097.4]
  wire [1:0] _T_1142; // @[Bitwise.scala 72:12:@34099.4]
  wire [29:0] _T_1143; // @[FixedPoint.scala 18:52:@34100.4]
  wire  _T_1172; // @[package.scala 96:25:@34152.4 package.scala 96:25:@34153.4]
  wire  _T_1174; // @[implicits.scala 55:10:@34154.4]
  wire  _T_1175; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 434:194:@34155.4]
  wire  x947_x580_D1; // @[package.scala 96:25:@34129.4 package.scala 96:25:@34130.4]
  wire  _T_1176; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 434:282:@34156.4]
  wire  _T_1177; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 434:290:@34157.4]
  wire  x589; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 438:59:@34168.4]
  wire  _T_1207; // @[package.scala 96:25:@34205.4 package.scala 96:25:@34206.4]
  wire  _T_1209; // @[implicits.scala 55:10:@34207.4]
  wire  _T_1210; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 451:194:@34208.4]
  wire  x949_x590_D1; // @[package.scala 96:25:@34191.4 package.scala 96:25:@34192.4]
  wire  _T_1211; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 451:282:@34209.4]
  wire  _T_1212; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 451:290:@34210.4]
  wire  x596; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 455:59:@34221.4]
  wire  _T_1240; // @[package.scala 96:25:@34256.4 package.scala 96:25:@34257.4]
  wire  _T_1242; // @[implicits.scala 55:10:@34258.4]
  wire  _T_1243; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 466:194:@34259.4]
  wire  x950_x597_D1; // @[package.scala 96:25:@34242.4 package.scala 96:25:@34243.4]
  wire  _T_1244; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 466:282:@34260.4]
  wire  _T_1245; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 466:290:@34261.4]
  wire  x603; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 470:59:@34272.4]
  wire  _T_1279; // @[package.scala 96:25:@34325.4 package.scala 96:25:@34326.4]
  wire  _T_1281; // @[implicits.scala 55:10:@34327.4]
  wire  _T_1282; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 485:194:@34328.4]
  wire  x953_x604_D2; // @[package.scala 96:25:@34311.4 package.scala 96:25:@34312.4]
  wire  _T_1283; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 485:282:@34329.4]
  wire  _T_1284; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 485:290:@34330.4]
  wire  x610; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 489:59:@34341.4]
  wire  _T_1312; // @[package.scala 96:25:@34376.4 package.scala 96:25:@34377.4]
  wire  _T_1314; // @[implicits.scala 55:10:@34378.4]
  wire  _T_1315; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 500:194:@34379.4]
  wire  x954_x611_D1; // @[package.scala 96:25:@34362.4 package.scala 96:25:@34363.4]
  wire  _T_1316; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 500:282:@34380.4]
  wire  _T_1317; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 500:290:@34381.4]
  wire  x617; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 504:59:@34392.4]
  wire  _T_1345; // @[package.scala 96:25:@34427.4 package.scala 96:25:@34428.4]
  wire  _T_1347; // @[implicits.scala 55:10:@34429.4]
  wire  _T_1348; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 515:194:@34430.4]
  wire  x955_x618_D1; // @[package.scala 96:25:@34413.4 package.scala 96:25:@34414.4]
  wire  _T_1349; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 515:282:@34431.4]
  wire  _T_1350; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 515:290:@34432.4]
  wire [31:0] x624_rdrow_number; // @[Math.scala 154:22:@34451.4 Math.scala 155:14:@34452.4]
  wire [31:0] _T_1367; // @[Math.scala 406:49:@34458.4]
  wire [31:0] _T_1369; // @[Math.scala 406:56:@34460.4]
  wire [31:0] _T_1370; // @[Math.scala 406:56:@34461.4]
  wire [31:0] x898_number; // @[implicits.scala 133:21:@34462.4]
  wire  x626; // @[Math.scala 465:44:@34470.4]
  wire  x627; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 525:24:@34473.4]
  wire [31:0] _T_1391; // @[Math.scala 406:49:@34482.4]
  wire [31:0] _T_1393; // @[Math.scala 406:56:@34484.4]
  wire [31:0] _T_1394; // @[Math.scala 406:56:@34485.4]
  wire  _T_1399; // @[FixedPoint.scala 50:25:@34491.4]
  wire [1:0] _T_1403; // @[Bitwise.scala 72:12:@34493.4]
  wire [29:0] _T_1404; // @[FixedPoint.scala 18:52:@34494.4]
  wire  _T_1430; // @[package.scala 96:25:@34537.4 package.scala 96:25:@34538.4]
  wire  _T_1432; // @[implicits.scala 55:10:@34539.4]
  wire  _T_1433; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 542:194:@34540.4]
  wire  x956_x628_D1; // @[package.scala 96:25:@34514.4 package.scala 96:25:@34515.4]
  wire  _T_1434; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 542:282:@34541.4]
  wire  _T_1435; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 542:290:@34542.4]
  wire  x637; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 546:24:@34553.4]
  wire  _T_1465; // @[package.scala 96:25:@34590.4 package.scala 96:25:@34591.4]
  wire  _T_1467; // @[implicits.scala 55:10:@34592.4]
  wire  _T_1468; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 565:194:@34593.4]
  wire  x958_x638_D1; // @[package.scala 96:25:@34576.4 package.scala 96:25:@34577.4]
  wire  _T_1469; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 565:282:@34594.4]
  wire  _T_1470; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 565:290:@34595.4]
  wire  x644; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 569:59:@34606.4]
  wire  _T_1498; // @[package.scala 96:25:@34641.4 package.scala 96:25:@34642.4]
  wire  _T_1500; // @[implicits.scala 55:10:@34643.4]
  wire  _T_1501; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 580:194:@34644.4]
  wire  x959_x645_D1; // @[package.scala 96:25:@34627.4 package.scala 96:25:@34628.4]
  wire  _T_1502; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 580:282:@34645.4]
  wire  _T_1503; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 580:290:@34646.4]
  wire  x651; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 584:59:@34657.4]
  wire  _T_1531; // @[package.scala 96:25:@34692.4 package.scala 96:25:@34693.4]
  wire  _T_1533; // @[implicits.scala 55:10:@34694.4]
  wire  _T_1534; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 595:194:@34695.4]
  wire  x960_x652_D1; // @[package.scala 96:25:@34678.4 package.scala 96:25:@34679.4]
  wire  _T_1535; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 595:282:@34696.4]
  wire  _T_1536; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 595:290:@34697.4]
  wire  x658; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 599:59:@34708.4]
  wire  _T_1564; // @[package.scala 96:25:@34743.4 package.scala 96:25:@34744.4]
  wire  _T_1566; // @[implicits.scala 55:10:@34745.4]
  wire  _T_1567; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 610:194:@34746.4]
  wire  x961_x659_D1; // @[package.scala 96:25:@34729.4 package.scala 96:25:@34730.4]
  wire  _T_1568; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 610:282:@34747.4]
  wire  _T_1569; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 610:290:@34748.4]
  wire  x665; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 614:59:@34759.4]
  wire  _T_1597; // @[package.scala 96:25:@34794.4 package.scala 96:25:@34795.4]
  wire  _T_1599; // @[implicits.scala 55:10:@34796.4]
  wire  _T_1600; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 625:194:@34797.4]
  wire  x962_x666_D1; // @[package.scala 96:25:@34780.4 package.scala 96:25:@34781.4]
  wire  _T_1601; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 625:282:@34798.4]
  wire  _T_1602; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 625:290:@34799.4]
  wire [31:0] x672_rdrow_number; // @[Math.scala 154:22:@34818.4 Math.scala 155:14:@34819.4]
  wire [31:0] _T_1619; // @[Math.scala 406:49:@34825.4]
  wire [31:0] _T_1621; // @[Math.scala 406:56:@34827.4]
  wire [31:0] _T_1622; // @[Math.scala 406:56:@34828.4]
  wire [31:0] x900_number; // @[implicits.scala 133:21:@34829.4]
  wire  x674; // @[Math.scala 465:44:@34837.4]
  wire  x675; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 635:24:@34840.4]
  wire [31:0] _T_1643; // @[Math.scala 406:49:@34849.4]
  wire [31:0] _T_1645; // @[Math.scala 406:56:@34851.4]
  wire [31:0] _T_1646; // @[Math.scala 406:56:@34852.4]
  wire  _T_1651; // @[FixedPoint.scala 50:25:@34858.4]
  wire [1:0] _T_1655; // @[Bitwise.scala 72:12:@34860.4]
  wire [29:0] _T_1656; // @[FixedPoint.scala 18:52:@34861.4]
  wire  _T_1682; // @[package.scala 96:25:@34904.4 package.scala 96:25:@34905.4]
  wire  _T_1684; // @[implicits.scala 55:10:@34906.4]
  wire  _T_1685; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 652:194:@34907.4]
  wire  x964_x676_D1; // @[package.scala 96:25:@34890.4 package.scala 96:25:@34891.4]
  wire  _T_1686; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 652:282:@34908.4]
  wire  _T_1687; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 652:290:@34909.4]
  wire  x685; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 656:24:@34920.4]
  wire  _T_1715; // @[package.scala 96:25:@34955.4 package.scala 96:25:@34956.4]
  wire  _T_1717; // @[implicits.scala 55:10:@34957.4]
  wire  _T_1718; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 667:194:@34958.4]
  wire  x965_x686_D1; // @[package.scala 96:25:@34941.4 package.scala 96:25:@34942.4]
  wire  _T_1719; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 667:282:@34959.4]
  wire  _T_1720; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 667:290:@34960.4]
  wire  x692; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 671:24:@34971.4]
  wire  _T_1750; // @[package.scala 96:25:@35008.4 package.scala 96:25:@35009.4]
  wire  _T_1752; // @[implicits.scala 55:10:@35010.4]
  wire  _T_1753; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 690:194:@35011.4]
  wire  x966_x693_D1; // @[package.scala 96:25:@34994.4 package.scala 96:25:@34995.4]
  wire  _T_1754; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 690:282:@35012.4]
  wire  _T_1755; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 690:290:@35013.4]
  wire  x699; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 694:59:@35024.4]
  wire  _T_1783; // @[package.scala 96:25:@35059.4 package.scala 96:25:@35060.4]
  wire  _T_1785; // @[implicits.scala 55:10:@35061.4]
  wire  _T_1786; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 705:194:@35062.4]
  wire  x967_x700_D1; // @[package.scala 96:25:@35045.4 package.scala 96:25:@35046.4]
  wire  _T_1787; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 705:282:@35063.4]
  wire  _T_1788; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 705:290:@35064.4]
  wire  x706; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 709:59:@35075.4]
  wire  _T_1816; // @[package.scala 96:25:@35110.4 package.scala 96:25:@35111.4]
  wire  _T_1818; // @[implicits.scala 55:10:@35112.4]
  wire  _T_1819; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 720:194:@35113.4]
  wire  x968_x707_D1; // @[package.scala 96:25:@35096.4 package.scala 96:25:@35097.4]
  wire  _T_1820; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 720:282:@35114.4]
  wire  _T_1821; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 720:290:@35115.4]
  wire  x713; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 724:59:@35126.4]
  wire  _T_1849; // @[package.scala 96:25:@35161.4 package.scala 96:25:@35162.4]
  wire  _T_1851; // @[implicits.scala 55:10:@35163.4]
  wire  _T_1852; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 735:194:@35164.4]
  wire  x969_x714_D1; // @[package.scala 96:25:@35147.4 package.scala 96:25:@35148.4]
  wire  _T_1853; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 735:282:@35165.4]
  wire  _T_1854; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 735:290:@35166.4]
  wire [7:0] x535_rd_0_number; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 305:29:@33695.4 sm_x824_inr_Foreach_SAMPLER_BOX.scala 309:442:@33718.4]
  wire [8:0] _GEN_0; // @[Math.scala 450:32:@35178.4]
  wire [8:0] _T_1860; // @[Math.scala 450:32:@35178.4]
  wire [7:0] x587_rd_0_number; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 430:29:@34141.4 sm_x824_inr_Foreach_SAMPLER_BOX.scala 434:407:@34164.4]
  wire [8:0] _GEN_1; // @[Math.scala 450:32:@35183.4]
  wire [8:0] _T_1864; // @[Math.scala 450:32:@35183.4]
  wire [7:0] x594_rd_0_number; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 447:29:@34194.4 sm_x824_inr_Foreach_SAMPLER_BOX.scala 451:407:@34217.4]
  wire [9:0] _GEN_2; // @[Math.scala 450:32:@35188.4]
  wire [9:0] _T_1868; // @[Math.scala 450:32:@35188.4]
  wire [7:0] x601_rd_0_number; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 462:29:@34245.4 sm_x824_inr_Foreach_SAMPLER_BOX.scala 466:407:@34268.4]
  wire [8:0] _GEN_3; // @[Math.scala 450:32:@35193.4]
  wire [8:0] _T_1872; // @[Math.scala 450:32:@35193.4]
  wire [7:0] x642_rd_0_number; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 561:29:@34579.4 sm_x824_inr_Foreach_SAMPLER_BOX.scala 565:407:@34602.4]
  wire [8:0] _GEN_4; // @[Math.scala 450:32:@35198.4]
  wire [8:0] _T_1876; // @[Math.scala 450:32:@35198.4]
  wire [7:0] x732_sum_number; // @[Math.scala 154:22:@35287.4 Math.scala 155:14:@35288.4]
  wire [3:0] _T_1912; // @[FixedPoint.scala 18:52:@35293.4]
  wire [7:0] x543_rd_0_number; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 328:29:@33773.4 sm_x824_inr_Foreach_SAMPLER_BOX.scala 332:407:@33796.4]
  wire [8:0] _GEN_5; // @[Math.scala 450:32:@35306.4]
  wire [8:0] _T_1919; // @[Math.scala 450:32:@35306.4]
  wire [8:0] _GEN_6; // @[Math.scala 450:32:@35311.4]
  wire [8:0] _T_1923; // @[Math.scala 450:32:@35311.4]
  wire [9:0] _GEN_7; // @[Math.scala 450:32:@35316.4]
  wire [9:0] _T_1927; // @[Math.scala 450:32:@35316.4]
  wire [7:0] x608_rd_0_number; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 481:29:@34314.4 sm_x824_inr_Foreach_SAMPLER_BOX.scala 485:407:@34337.4]
  wire [8:0] _GEN_8; // @[Math.scala 450:32:@35321.4]
  wire [8:0] _T_1931; // @[Math.scala 450:32:@35321.4]
  wire [7:0] x649_rd_0_number; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 576:29:@34630.4 sm_x824_inr_Foreach_SAMPLER_BOX.scala 580:407:@34653.4]
  wire [8:0] _GEN_9; // @[Math.scala 450:32:@35326.4]
  wire [8:0] _T_1935; // @[Math.scala 450:32:@35326.4]
  wire [7:0] x746_sum_number; // @[Math.scala 154:22:@35417.4 Math.scala 155:14:@35418.4]
  wire [3:0] _T_1973; // @[FixedPoint.scala 18:52:@35423.4]
  wire [7:0] x551_rd_0_number; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 351:29:@33858.4 sm_x824_inr_Foreach_SAMPLER_BOX.scala 355:407:@33881.4]
  wire [8:0] _GEN_10; // @[Math.scala 450:32:@35436.4]
  wire [8:0] _T_1980; // @[Math.scala 450:32:@35436.4]
  wire [9:0] _GEN_11; // @[Math.scala 450:32:@35441.4]
  wire [9:0] _T_1984; // @[Math.scala 450:32:@35441.4]
  wire [7:0] x615_rd_0_number; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 496:29:@34365.4 sm_x824_inr_Foreach_SAMPLER_BOX.scala 500:407:@34388.4]
  wire [8:0] _GEN_12; // @[Math.scala 450:32:@35446.4]
  wire [8:0] _T_1988; // @[Math.scala 450:32:@35446.4]
  wire [7:0] x656_rd_0_number; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 591:29:@34681.4 sm_x824_inr_Foreach_SAMPLER_BOX.scala 595:407:@34704.4]
  wire [8:0] _GEN_13; // @[Math.scala 450:32:@35451.4]
  wire [8:0] _T_1992; // @[Math.scala 450:32:@35451.4]
  wire [7:0] x759_sum_number; // @[Math.scala 154:22:@35540.4 Math.scala 155:14:@35541.4]
  wire [3:0] _T_2028; // @[FixedPoint.scala 18:52:@35546.4]
  wire [7:0] x563_rd_0_number; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 372:29:@33937.4 sm_x824_inr_Foreach_SAMPLER_BOX.scala 376:407:@33960.4]
  wire [8:0] _GEN_14; // @[Math.scala 450:32:@35559.4]
  wire [8:0] _T_2035; // @[Math.scala 450:32:@35559.4]
  wire [9:0] _GEN_15; // @[Math.scala 450:32:@35564.4]
  wire [9:0] _T_2039; // @[Math.scala 450:32:@35564.4]
  wire [7:0] x622_rd_0_number; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 511:29:@34416.4 sm_x824_inr_Foreach_SAMPLER_BOX.scala 515:407:@34439.4]
  wire [8:0] _GEN_16; // @[Math.scala 450:32:@35569.4]
  wire [8:0] _T_2043; // @[Math.scala 450:32:@35569.4]
  wire [7:0] x663_rd_0_number; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 606:29:@34732.4 sm_x824_inr_Foreach_SAMPLER_BOX.scala 610:407:@34755.4]
  wire [8:0] _GEN_17; // @[Math.scala 450:32:@35574.4]
  wire [8:0] _T_2047; // @[Math.scala 450:32:@35574.4]
  wire [7:0] x772_sum_number; // @[Math.scala 154:22:@35663.4 Math.scala 155:14:@35664.4]
  wire [3:0] _T_2083; // @[FixedPoint.scala 18:52:@35669.4]
  wire [7:0] x635_rd_0_number; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 538:29:@34526.4 sm_x824_inr_Foreach_SAMPLER_BOX.scala 542:407:@34549.4]
  wire [8:0] _GEN_18; // @[Math.scala 450:32:@35682.4]
  wire [8:0] _T_2090; // @[Math.scala 450:32:@35682.4]
  wire [9:0] _GEN_19; // @[Math.scala 450:32:@35687.4]
  wire [9:0] _T_2094; // @[Math.scala 450:32:@35687.4]
  wire [7:0] x690_rd_0_number; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 663:29:@34944.4 sm_x824_inr_Foreach_SAMPLER_BOX.scala 667:407:@34967.4]
  wire [8:0] _GEN_20; // @[Math.scala 450:32:@35692.4]
  wire [8:0] _T_2098; // @[Math.scala 450:32:@35692.4]
  wire [7:0] x784_sum_number; // @[Math.scala 154:22:@35781.4 Math.scala 155:14:@35782.4]
  wire [3:0] _T_2134; // @[FixedPoint.scala 18:52:@35787.4]
  wire [9:0] _GEN_21; // @[Math.scala 450:32:@35800.4]
  wire [9:0] _T_2141; // @[Math.scala 450:32:@35800.4]
  wire [7:0] x697_rd_0_number; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 686:29:@34997.4 sm_x824_inr_Foreach_SAMPLER_BOX.scala 690:407:@35020.4]
  wire [8:0] _GEN_22; // @[Math.scala 450:32:@35805.4]
  wire [8:0] _T_2145; // @[Math.scala 450:32:@35805.4]
  wire [7:0] x795_sum_number; // @[Math.scala 154:22:@35896.4 Math.scala 155:14:@35897.4]
  wire [3:0] _T_2183; // @[FixedPoint.scala 18:52:@35902.4]
  wire [9:0] _GEN_23; // @[Math.scala 450:32:@35915.4]
  wire [9:0] _T_2190; // @[Math.scala 450:32:@35915.4]
  wire [7:0] x704_rd_0_number; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 701:29:@35048.4 sm_x824_inr_Foreach_SAMPLER_BOX.scala 705:407:@35071.4]
  wire [8:0] _GEN_24; // @[Math.scala 450:32:@35920.4]
  wire [8:0] _T_2194; // @[Math.scala 450:32:@35920.4]
  wire [7:0] x806_sum_number; // @[Math.scala 154:22:@36009.4 Math.scala 155:14:@36010.4]
  wire [3:0] _T_2230; // @[FixedPoint.scala 18:52:@36015.4]
  wire [9:0] _GEN_25; // @[Math.scala 450:32:@36028.4]
  wire [9:0] _T_2237; // @[Math.scala 450:32:@36028.4]
  wire [7:0] x670_rd_0_number; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 621:29:@34783.4 sm_x824_inr_Foreach_SAMPLER_BOX.scala 625:407:@34806.4]
  wire [8:0] _GEN_26; // @[Math.scala 450:32:@36033.4]
  wire [8:0] _T_2241; // @[Math.scala 450:32:@36033.4]
  wire [7:0] x711_rd_0_number; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 716:29:@35099.4 sm_x824_inr_Foreach_SAMPLER_BOX.scala 720:407:@35122.4]
  wire [8:0] _GEN_27; // @[Math.scala 450:32:@36038.4]
  wire [8:0] _T_2245; // @[Math.scala 450:32:@36038.4]
  wire [7:0] x818_sum_number; // @[Math.scala 154:22:@36127.4 Math.scala 155:14:@36128.4]
  wire [3:0] _T_2281; // @[FixedPoint.scala 18:52:@36133.4]
  wire [7:0] x807_number; // @[package.scala 96:25:@36022.4 package.scala 96:25:@36023.4]
  wire [7:0] x819_number; // @[package.scala 96:25:@36140.4 package.scala 96:25:@36141.4]
  wire [7:0] x785_number; // @[package.scala 96:25:@35794.4 package.scala 96:25:@35795.4]
  wire [7:0] x796_number; // @[package.scala 96:25:@35909.4 package.scala 96:25:@35910.4]
  wire [31:0] _T_2302; // @[Cat.scala 30:58:@36156.4]
  wire [7:0] x760_number; // @[package.scala 96:25:@35553.4 package.scala 96:25:@35554.4]
  wire [7:0] x773_number; // @[package.scala 96:25:@35676.4 package.scala 96:25:@35677.4]
  wire [7:0] x733_number; // @[package.scala 96:25:@35300.4 package.scala 96:25:@35301.4]
  wire [7:0] x747_number; // @[package.scala 96:25:@35430.4 package.scala 96:25:@35431.4]
  wire [31:0] _T_2305; // @[Cat.scala 30:58:@36159.4]
  wire  _T_2318; // @[package.scala 96:25:@36195.4 package.scala 96:25:@36196.4]
  wire  _T_2320; // @[implicits.scala 55:10:@36197.4]
  wire  x978_b437_D19; // @[package.scala 96:25:@36177.4 package.scala 96:25:@36178.4]
  wire  _T_2321; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 979:116:@36198.4]
  wire  x979_b438_D19; // @[package.scala 96:25:@36186.4 package.scala 96:25:@36187.4]
  wire  _T_2322; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 979:122:@36199.4]
  wire [31:0] x903_x892_D8_number; // @[package.scala 96:25:@32875.4 package.scala 96:25:@32876.4]
  wire [31:0] x905_x453_sum_D7_number; // @[package.scala 96:25:@32893.4 package.scala 96:25:@32894.4]
  wire [31:0] x910_x463_sum_D6_number; // @[package.scala 96:25:@32996.4 package.scala 96:25:@32997.4]
  wire [31:0] x911_x472_sum_D6_number; // @[package.scala 96:25:@33063.4 package.scala 96:25:@33064.4]
  wire [31:0] x913_x481_sum_D6_number; // @[package.scala 96:25:@33139.4 package.scala 96:25:@33140.4]
  wire [31:0] x916_x893_D7_number; // @[package.scala 96:25:@33284.4 package.scala 96:25:@33285.4]
  wire [31:0] x918_x495_sum_D6_number; // @[package.scala 96:25:@33302.4 package.scala 96:25:@33303.4]
  wire [31:0] x920_x501_sum_D6_number; // @[package.scala 96:25:@33357.4 package.scala 96:25:@33358.4]
  wire [31:0] x922_x506_sum_D6_number; // @[package.scala 96:25:@33412.4 package.scala 96:25:@33413.4]
  wire [31:0] x923_x511_sum_D6_number; // @[package.scala 96:25:@33458.4 package.scala 96:25:@33459.4]
  wire [31:0] x523_sum_number; // @[Math.scala 154:22:@33580.4 Math.scala 155:14:@33581.4]
  wire [31:0] x929_x895_D1_number; // @[package.scala 96:25:@33598.4 package.scala 96:25:@33599.4]
  wire [31:0] x532_sum_number; // @[Math.scala 154:22:@33683.4 Math.scala 155:14:@33684.4]
  wire [31:0] x540_sum_number; // @[Math.scala 154:22:@33761.4 Math.scala 155:14:@33762.4]
  wire [31:0] x548_sum_number; // @[Math.scala 154:22:@33846.4 Math.scala 155:14:@33847.4]
  wire [31:0] x559_sum_number; // @[Math.scala 154:22:@33925.4 Math.scala 155:14:@33926.4]
  wire [31:0] x571_sum_number; // @[Math.scala 154:22:@34004.4 Math.scala 155:14:@34005.4]
  wire [31:0] x583_sum_number; // @[Math.scala 154:22:@34120.4 Math.scala 155:14:@34121.4]
  wire [31:0] x948_x897_D2_number; // @[package.scala 96:25:@34138.4 package.scala 96:25:@34139.4]
  wire [31:0] x591_sum_number; // @[Math.scala 154:22:@34182.4 Math.scala 155:14:@34183.4]
  wire [31:0] x598_sum_number; // @[Math.scala 154:22:@34233.4 Math.scala 155:14:@34234.4]
  wire [31:0] x952_x605_sum_D1_number; // @[package.scala 96:25:@34302.4 package.scala 96:25:@34303.4]
  wire [31:0] x612_sum_number; // @[Math.scala 154:22:@34353.4 Math.scala 155:14:@34354.4]
  wire [31:0] x619_sum_number; // @[Math.scala 154:22:@34404.4 Math.scala 155:14:@34405.4]
  wire [31:0] x631_sum_number; // @[Math.scala 154:22:@34505.4 Math.scala 155:14:@34506.4]
  wire [31:0] x957_x899_D1_number; // @[package.scala 96:25:@34523.4 package.scala 96:25:@34524.4]
  wire [31:0] x639_sum_number; // @[Math.scala 154:22:@34567.4 Math.scala 155:14:@34568.4]
  wire [31:0] x646_sum_number; // @[Math.scala 154:22:@34618.4 Math.scala 155:14:@34619.4]
  wire [31:0] x653_sum_number; // @[Math.scala 154:22:@34669.4 Math.scala 155:14:@34670.4]
  wire [31:0] x660_sum_number; // @[Math.scala 154:22:@34720.4 Math.scala 155:14:@34721.4]
  wire [31:0] x667_sum_number; // @[Math.scala 154:22:@34771.4 Math.scala 155:14:@34772.4]
  wire [31:0] x679_sum_number; // @[Math.scala 154:22:@34872.4 Math.scala 155:14:@34873.4]
  wire [31:0] x963_x901_D1_number; // @[package.scala 96:25:@34881.4 package.scala 96:25:@34882.4]
  wire [31:0] x687_sum_number; // @[Math.scala 154:22:@34932.4 Math.scala 155:14:@34933.4]
  wire [31:0] x694_sum_number; // @[Math.scala 154:22:@34985.4 Math.scala 155:14:@34986.4]
  wire [31:0] x701_sum_number; // @[Math.scala 154:22:@35036.4 Math.scala 155:14:@35037.4]
  wire [31:0] x708_sum_number; // @[Math.scala 154:22:@35087.4 Math.scala 155:14:@35088.4]
  wire [31:0] x715_sum_number; // @[Math.scala 154:22:@35138.4 Math.scala 155:14:@35139.4]
  _ _ ( // @[Math.scala 709:24:@32504.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 709:24:@32516.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  x439_lb_0 x439_lb_0 ( // @[m_x439_lb_0.scala 57:17:@32526.4]
    .clock(x439_lb_0_clock),
    .reset(x439_lb_0_reset),
    .io_rPort_23_banks_0(x439_lb_0_io_rPort_23_banks_0),
    .io_rPort_23_ofs_0(x439_lb_0_io_rPort_23_ofs_0),
    .io_rPort_23_en_0(x439_lb_0_io_rPort_23_en_0),
    .io_rPort_23_backpressure(x439_lb_0_io_rPort_23_backpressure),
    .io_rPort_23_output_0(x439_lb_0_io_rPort_23_output_0),
    .io_rPort_22_banks_0(x439_lb_0_io_rPort_22_banks_0),
    .io_rPort_22_ofs_0(x439_lb_0_io_rPort_22_ofs_0),
    .io_rPort_22_en_0(x439_lb_0_io_rPort_22_en_0),
    .io_rPort_22_backpressure(x439_lb_0_io_rPort_22_backpressure),
    .io_rPort_22_output_0(x439_lb_0_io_rPort_22_output_0),
    .io_rPort_21_banks_0(x439_lb_0_io_rPort_21_banks_0),
    .io_rPort_21_ofs_0(x439_lb_0_io_rPort_21_ofs_0),
    .io_rPort_21_en_0(x439_lb_0_io_rPort_21_en_0),
    .io_rPort_21_backpressure(x439_lb_0_io_rPort_21_backpressure),
    .io_rPort_21_output_0(x439_lb_0_io_rPort_21_output_0),
    .io_rPort_20_banks_0(x439_lb_0_io_rPort_20_banks_0),
    .io_rPort_20_ofs_0(x439_lb_0_io_rPort_20_ofs_0),
    .io_rPort_20_en_0(x439_lb_0_io_rPort_20_en_0),
    .io_rPort_20_backpressure(x439_lb_0_io_rPort_20_backpressure),
    .io_rPort_20_output_0(x439_lb_0_io_rPort_20_output_0),
    .io_rPort_19_banks_0(x439_lb_0_io_rPort_19_banks_0),
    .io_rPort_19_ofs_0(x439_lb_0_io_rPort_19_ofs_0),
    .io_rPort_19_en_0(x439_lb_0_io_rPort_19_en_0),
    .io_rPort_19_backpressure(x439_lb_0_io_rPort_19_backpressure),
    .io_rPort_19_output_0(x439_lb_0_io_rPort_19_output_0),
    .io_rPort_18_banks_0(x439_lb_0_io_rPort_18_banks_0),
    .io_rPort_18_ofs_0(x439_lb_0_io_rPort_18_ofs_0),
    .io_rPort_18_en_0(x439_lb_0_io_rPort_18_en_0),
    .io_rPort_18_backpressure(x439_lb_0_io_rPort_18_backpressure),
    .io_rPort_18_output_0(x439_lb_0_io_rPort_18_output_0),
    .io_rPort_17_banks_0(x439_lb_0_io_rPort_17_banks_0),
    .io_rPort_17_ofs_0(x439_lb_0_io_rPort_17_ofs_0),
    .io_rPort_17_en_0(x439_lb_0_io_rPort_17_en_0),
    .io_rPort_17_backpressure(x439_lb_0_io_rPort_17_backpressure),
    .io_rPort_17_output_0(x439_lb_0_io_rPort_17_output_0),
    .io_rPort_16_banks_0(x439_lb_0_io_rPort_16_banks_0),
    .io_rPort_16_ofs_0(x439_lb_0_io_rPort_16_ofs_0),
    .io_rPort_16_en_0(x439_lb_0_io_rPort_16_en_0),
    .io_rPort_16_backpressure(x439_lb_0_io_rPort_16_backpressure),
    .io_rPort_16_output_0(x439_lb_0_io_rPort_16_output_0),
    .io_rPort_15_banks_0(x439_lb_0_io_rPort_15_banks_0),
    .io_rPort_15_ofs_0(x439_lb_0_io_rPort_15_ofs_0),
    .io_rPort_15_en_0(x439_lb_0_io_rPort_15_en_0),
    .io_rPort_15_backpressure(x439_lb_0_io_rPort_15_backpressure),
    .io_rPort_15_output_0(x439_lb_0_io_rPort_15_output_0),
    .io_rPort_14_banks_0(x439_lb_0_io_rPort_14_banks_0),
    .io_rPort_14_ofs_0(x439_lb_0_io_rPort_14_ofs_0),
    .io_rPort_14_en_0(x439_lb_0_io_rPort_14_en_0),
    .io_rPort_14_backpressure(x439_lb_0_io_rPort_14_backpressure),
    .io_rPort_14_output_0(x439_lb_0_io_rPort_14_output_0),
    .io_rPort_13_banks_0(x439_lb_0_io_rPort_13_banks_0),
    .io_rPort_13_ofs_0(x439_lb_0_io_rPort_13_ofs_0),
    .io_rPort_13_en_0(x439_lb_0_io_rPort_13_en_0),
    .io_rPort_13_backpressure(x439_lb_0_io_rPort_13_backpressure),
    .io_rPort_13_output_0(x439_lb_0_io_rPort_13_output_0),
    .io_rPort_12_banks_0(x439_lb_0_io_rPort_12_banks_0),
    .io_rPort_12_ofs_0(x439_lb_0_io_rPort_12_ofs_0),
    .io_rPort_12_en_0(x439_lb_0_io_rPort_12_en_0),
    .io_rPort_12_backpressure(x439_lb_0_io_rPort_12_backpressure),
    .io_rPort_12_output_0(x439_lb_0_io_rPort_12_output_0),
    .io_rPort_11_banks_0(x439_lb_0_io_rPort_11_banks_0),
    .io_rPort_11_ofs_0(x439_lb_0_io_rPort_11_ofs_0),
    .io_rPort_11_en_0(x439_lb_0_io_rPort_11_en_0),
    .io_rPort_11_backpressure(x439_lb_0_io_rPort_11_backpressure),
    .io_rPort_11_output_0(x439_lb_0_io_rPort_11_output_0),
    .io_rPort_10_banks_0(x439_lb_0_io_rPort_10_banks_0),
    .io_rPort_10_ofs_0(x439_lb_0_io_rPort_10_ofs_0),
    .io_rPort_10_en_0(x439_lb_0_io_rPort_10_en_0),
    .io_rPort_10_backpressure(x439_lb_0_io_rPort_10_backpressure),
    .io_rPort_10_output_0(x439_lb_0_io_rPort_10_output_0),
    .io_rPort_9_banks_0(x439_lb_0_io_rPort_9_banks_0),
    .io_rPort_9_ofs_0(x439_lb_0_io_rPort_9_ofs_0),
    .io_rPort_9_en_0(x439_lb_0_io_rPort_9_en_0),
    .io_rPort_9_backpressure(x439_lb_0_io_rPort_9_backpressure),
    .io_rPort_9_output_0(x439_lb_0_io_rPort_9_output_0),
    .io_rPort_8_banks_0(x439_lb_0_io_rPort_8_banks_0),
    .io_rPort_8_ofs_0(x439_lb_0_io_rPort_8_ofs_0),
    .io_rPort_8_en_0(x439_lb_0_io_rPort_8_en_0),
    .io_rPort_8_backpressure(x439_lb_0_io_rPort_8_backpressure),
    .io_rPort_8_output_0(x439_lb_0_io_rPort_8_output_0),
    .io_rPort_7_banks_0(x439_lb_0_io_rPort_7_banks_0),
    .io_rPort_7_ofs_0(x439_lb_0_io_rPort_7_ofs_0),
    .io_rPort_7_en_0(x439_lb_0_io_rPort_7_en_0),
    .io_rPort_7_backpressure(x439_lb_0_io_rPort_7_backpressure),
    .io_rPort_7_output_0(x439_lb_0_io_rPort_7_output_0),
    .io_rPort_6_banks_0(x439_lb_0_io_rPort_6_banks_0),
    .io_rPort_6_ofs_0(x439_lb_0_io_rPort_6_ofs_0),
    .io_rPort_6_en_0(x439_lb_0_io_rPort_6_en_0),
    .io_rPort_6_backpressure(x439_lb_0_io_rPort_6_backpressure),
    .io_rPort_6_output_0(x439_lb_0_io_rPort_6_output_0),
    .io_rPort_5_banks_0(x439_lb_0_io_rPort_5_banks_0),
    .io_rPort_5_ofs_0(x439_lb_0_io_rPort_5_ofs_0),
    .io_rPort_5_en_0(x439_lb_0_io_rPort_5_en_0),
    .io_rPort_5_backpressure(x439_lb_0_io_rPort_5_backpressure),
    .io_rPort_5_output_0(x439_lb_0_io_rPort_5_output_0),
    .io_rPort_4_banks_0(x439_lb_0_io_rPort_4_banks_0),
    .io_rPort_4_ofs_0(x439_lb_0_io_rPort_4_ofs_0),
    .io_rPort_4_en_0(x439_lb_0_io_rPort_4_en_0),
    .io_rPort_4_backpressure(x439_lb_0_io_rPort_4_backpressure),
    .io_rPort_4_output_0(x439_lb_0_io_rPort_4_output_0),
    .io_rPort_3_banks_0(x439_lb_0_io_rPort_3_banks_0),
    .io_rPort_3_ofs_0(x439_lb_0_io_rPort_3_ofs_0),
    .io_rPort_3_en_0(x439_lb_0_io_rPort_3_en_0),
    .io_rPort_3_backpressure(x439_lb_0_io_rPort_3_backpressure),
    .io_rPort_3_output_0(x439_lb_0_io_rPort_3_output_0),
    .io_rPort_2_banks_0(x439_lb_0_io_rPort_2_banks_0),
    .io_rPort_2_ofs_0(x439_lb_0_io_rPort_2_ofs_0),
    .io_rPort_2_en_0(x439_lb_0_io_rPort_2_en_0),
    .io_rPort_2_backpressure(x439_lb_0_io_rPort_2_backpressure),
    .io_rPort_2_output_0(x439_lb_0_io_rPort_2_output_0),
    .io_rPort_1_banks_0(x439_lb_0_io_rPort_1_banks_0),
    .io_rPort_1_ofs_0(x439_lb_0_io_rPort_1_ofs_0),
    .io_rPort_1_en_0(x439_lb_0_io_rPort_1_en_0),
    .io_rPort_1_backpressure(x439_lb_0_io_rPort_1_backpressure),
    .io_rPort_1_output_0(x439_lb_0_io_rPort_1_output_0),
    .io_rPort_0_banks_0(x439_lb_0_io_rPort_0_banks_0),
    .io_rPort_0_ofs_0(x439_lb_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x439_lb_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x439_lb_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x439_lb_0_io_rPort_0_output_0),
    .io_wPort_7_banks_0(x439_lb_0_io_wPort_7_banks_0),
    .io_wPort_7_ofs_0(x439_lb_0_io_wPort_7_ofs_0),
    .io_wPort_7_data_0(x439_lb_0_io_wPort_7_data_0),
    .io_wPort_7_en_0(x439_lb_0_io_wPort_7_en_0),
    .io_wPort_6_banks_0(x439_lb_0_io_wPort_6_banks_0),
    .io_wPort_6_ofs_0(x439_lb_0_io_wPort_6_ofs_0),
    .io_wPort_6_data_0(x439_lb_0_io_wPort_6_data_0),
    .io_wPort_6_en_0(x439_lb_0_io_wPort_6_en_0),
    .io_wPort_5_banks_0(x439_lb_0_io_wPort_5_banks_0),
    .io_wPort_5_ofs_0(x439_lb_0_io_wPort_5_ofs_0),
    .io_wPort_5_data_0(x439_lb_0_io_wPort_5_data_0),
    .io_wPort_5_en_0(x439_lb_0_io_wPort_5_en_0),
    .io_wPort_4_banks_0(x439_lb_0_io_wPort_4_banks_0),
    .io_wPort_4_ofs_0(x439_lb_0_io_wPort_4_ofs_0),
    .io_wPort_4_data_0(x439_lb_0_io_wPort_4_data_0),
    .io_wPort_4_en_0(x439_lb_0_io_wPort_4_en_0),
    .io_wPort_3_banks_0(x439_lb_0_io_wPort_3_banks_0),
    .io_wPort_3_ofs_0(x439_lb_0_io_wPort_3_ofs_0),
    .io_wPort_3_data_0(x439_lb_0_io_wPort_3_data_0),
    .io_wPort_3_en_0(x439_lb_0_io_wPort_3_en_0),
    .io_wPort_2_banks_0(x439_lb_0_io_wPort_2_banks_0),
    .io_wPort_2_ofs_0(x439_lb_0_io_wPort_2_ofs_0),
    .io_wPort_2_data_0(x439_lb_0_io_wPort_2_data_0),
    .io_wPort_2_en_0(x439_lb_0_io_wPort_2_en_0),
    .io_wPort_1_banks_0(x439_lb_0_io_wPort_1_banks_0),
    .io_wPort_1_ofs_0(x439_lb_0_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(x439_lb_0_io_wPort_1_data_0),
    .io_wPort_1_en_0(x439_lb_0_io_wPort_1_en_0),
    .io_wPort_0_banks_0(x439_lb_0_io_wPort_0_banks_0),
    .io_wPort_0_ofs_0(x439_lb_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x439_lb_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x439_lb_0_io_wPort_0_en_0)
  );
  RetimeWrapper_148 RetimeWrapper ( // @[package.scala 93:22:@32752.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x453_sum x453_sum_1 ( // @[Math.scala 150:24:@32860.4]
    .clock(x453_sum_1_clock),
    .reset(x453_sum_1_reset),
    .io_a(x453_sum_1_io_a),
    .io_b(x453_sum_1_io_b),
    .io_flow(x453_sum_1_io_flow),
    .io_result(x453_sum_1_io_result)
  );
  RetimeWrapper_150 RetimeWrapper_1 ( // @[package.scala 93:22:@32870.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_151 RetimeWrapper_2 ( // @[package.scala 93:22:@32879.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_152 RetimeWrapper_3 ( // @[package.scala 93:22:@32888.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_153 RetimeWrapper_4 ( // @[package.scala 93:22:@32897.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_153 RetimeWrapper_5 ( // @[package.scala 93:22:@32906.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_153 RetimeWrapper_6 ( // @[package.scala 93:22:@32919.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  x453_sum x459_rdcol_1 ( // @[Math.scala 150:24:@32942.4]
    .clock(x459_rdcol_1_clock),
    .reset(x459_rdcol_1_reset),
    .io_a(x459_rdcol_1_io_a),
    .io_b(x459_rdcol_1_io_b),
    .io_flow(x459_rdcol_1_io_flow),
    .io_result(x459_rdcol_1_io_result)
  );
  RetimeWrapper_149 RetimeWrapper_7 ( // @[package.scala 93:22:@32963.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  x453_sum x463_sum_1 ( // @[Math.scala 150:24:@32972.4]
    .clock(x463_sum_1_clock),
    .reset(x463_sum_1_reset),
    .io_a(x463_sum_1_io_a),
    .io_b(x463_sum_1_io_b),
    .io_flow(x463_sum_1_io_flow),
    .io_result(x463_sum_1_io_result)
  );
  RetimeWrapper_151 RetimeWrapper_8 ( // @[package.scala 93:22:@32982.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_160 RetimeWrapper_9 ( // @[package.scala 93:22:@32991.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_153 RetimeWrapper_10 ( // @[package.scala 93:22:@33004.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  x453_sum x468_rdcol_1 ( // @[Math.scala 150:24:@33027.4]
    .clock(x468_rdcol_1_clock),
    .reset(x468_rdcol_1_reset),
    .io_a(x468_rdcol_1_io_a),
    .io_b(x468_rdcol_1_io_b),
    .io_flow(x468_rdcol_1_io_flow),
    .io_result(x468_rdcol_1_io_result)
  );
  x453_sum x472_sum_1 ( // @[Math.scala 150:24:@33048.4]
    .clock(x472_sum_1_clock),
    .reset(x472_sum_1_reset),
    .io_a(x472_sum_1_io_a),
    .io_b(x472_sum_1_io_b),
    .io_flow(x472_sum_1_io_flow),
    .io_result(x472_sum_1_io_result)
  );
  RetimeWrapper_160 RetimeWrapper_11 ( // @[package.scala 93:22:@33058.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_151 RetimeWrapper_12 ( // @[package.scala 93:22:@33067.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_153 RetimeWrapper_13 ( // @[package.scala 93:22:@33080.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  x453_sum x477_rdcol_1 ( // @[Math.scala 150:24:@33103.4]
    .clock(x477_rdcol_1_clock),
    .reset(x477_rdcol_1_reset),
    .io_a(x477_rdcol_1_io_a),
    .io_b(x477_rdcol_1_io_b),
    .io_flow(x477_rdcol_1_io_flow),
    .io_result(x477_rdcol_1_io_result)
  );
  x453_sum x481_sum_1 ( // @[Math.scala 150:24:@33124.4]
    .clock(x481_sum_1_clock),
    .reset(x481_sum_1_reset),
    .io_a(x481_sum_1_io_a),
    .io_b(x481_sum_1_io_b),
    .io_flow(x481_sum_1_io_flow),
    .io_result(x481_sum_1_io_result)
  );
  RetimeWrapper_160 RetimeWrapper_14 ( // @[package.scala 93:22:@33134.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_151 RetimeWrapper_15 ( // @[package.scala 93:22:@33143.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_153 RetimeWrapper_16 ( // @[package.scala 93:22:@33156.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  x453_sum x486_rdrow_1 ( // @[Math.scala 150:24:@33179.4]
    .clock(x486_rdrow_1_clock),
    .reset(x486_rdrow_1_reset),
    .io_a(x486_rdrow_1_io_a),
    .io_b(x486_rdrow_1_io_b),
    .io_flow(x486_rdrow_1_io_flow),
    .io_result(x486_rdrow_1_io_result)
  );
  RetimeWrapper_149 RetimeWrapper_17 ( // @[package.scala 93:22:@33260.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  x453_sum x495_sum_1 ( // @[Math.scala 150:24:@33269.4]
    .clock(x495_sum_1_clock),
    .reset(x495_sum_1_reset),
    .io_a(x495_sum_1_io_a),
    .io_b(x495_sum_1_io_b),
    .io_flow(x495_sum_1_io_flow),
    .io_result(x495_sum_1_io_result)
  );
  RetimeWrapper_152 RetimeWrapper_18 ( // @[package.scala 93:22:@33279.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_151 RetimeWrapper_19 ( // @[package.scala 93:22:@33288.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_160 RetimeWrapper_20 ( // @[package.scala 93:22:@33297.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_153 RetimeWrapper_21 ( // @[package.scala 93:22:@33310.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  x453_sum x501_sum_1 ( // @[Math.scala 150:24:@33333.4]
    .clock(x501_sum_1_clock),
    .reset(x501_sum_1_reset),
    .io_a(x501_sum_1_io_a),
    .io_b(x501_sum_1_io_b),
    .io_flow(x501_sum_1_io_flow),
    .io_result(x501_sum_1_io_result)
  );
  RetimeWrapper_151 RetimeWrapper_22 ( // @[package.scala 93:22:@33343.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_160 RetimeWrapper_23 ( // @[package.scala 93:22:@33352.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_153 RetimeWrapper_24 ( // @[package.scala 93:22:@33365.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  x453_sum x506_sum_1 ( // @[Math.scala 150:24:@33388.4]
    .clock(x506_sum_1_clock),
    .reset(x506_sum_1_reset),
    .io_a(x506_sum_1_io_a),
    .io_b(x506_sum_1_io_b),
    .io_flow(x506_sum_1_io_flow),
    .io_result(x506_sum_1_io_result)
  );
  RetimeWrapper_151 RetimeWrapper_25 ( // @[package.scala 93:22:@33398.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_160 RetimeWrapper_26 ( // @[package.scala 93:22:@33407.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_153 RetimeWrapper_27 ( // @[package.scala 93:22:@33420.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  x453_sum x511_sum_1 ( // @[Math.scala 150:24:@33443.4]
    .clock(x511_sum_1_clock),
    .reset(x511_sum_1_reset),
    .io_a(x511_sum_1_io_a),
    .io_b(x511_sum_1_io_b),
    .io_flow(x511_sum_1_io_flow),
    .io_result(x511_sum_1_io_result)
  );
  RetimeWrapper_160 RetimeWrapper_28 ( // @[package.scala 93:22:@33453.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_151 RetimeWrapper_29 ( // @[package.scala 93:22:@33462.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_153 RetimeWrapper_30 ( // @[package.scala 93:22:@33475.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_191 RetimeWrapper_31 ( // @[package.scala 93:22:@33496.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_191 RetimeWrapper_32 ( // @[package.scala 93:22:@33523.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_191 RetimeWrapper_33 ( // @[package.scala 93:22:@33565.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  x453_sum x523_sum_1 ( // @[Math.scala 150:24:@33574.4]
    .clock(x523_sum_1_clock),
    .reset(x523_sum_1_reset),
    .io_a(x523_sum_1_io_a),
    .io_b(x523_sum_1_io_b),
    .io_flow(x523_sum_1_io_flow),
    .io_result(x523_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_34 ( // @[package.scala 93:22:@33584.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_149 RetimeWrapper_35 ( // @[package.scala 93:22:@33593.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_197 RetimeWrapper_36 ( // @[package.scala 93:22:@33602.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_197 RetimeWrapper_37 ( // @[package.scala 93:22:@33611.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_197 RetimeWrapper_38 ( // @[package.scala 93:22:@33625.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_191 RetimeWrapper_39 ( // @[package.scala 93:22:@33646.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_191 RetimeWrapper_40 ( // @[package.scala 93:22:@33668.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  x453_sum x532_sum_1 ( // @[Math.scala 150:24:@33677.4]
    .clock(x532_sum_1_clock),
    .reset(x532_sum_1_reset),
    .io_a(x532_sum_1_io_a),
    .io_b(x532_sum_1_io_b),
    .io_flow(x532_sum_1_io_flow),
    .io_result(x532_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_41 ( // @[package.scala 93:22:@33687.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_197 RetimeWrapper_42 ( // @[package.scala 93:22:@33701.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_191 RetimeWrapper_43 ( // @[package.scala 93:22:@33722.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_191 RetimeWrapper_44 ( // @[package.scala 93:22:@33746.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  x453_sum x540_sum_1 ( // @[Math.scala 150:24:@33755.4]
    .clock(x540_sum_1_clock),
    .reset(x540_sum_1_reset),
    .io_a(x540_sum_1_io_a),
    .io_b(x540_sum_1_io_b),
    .io_flow(x540_sum_1_io_flow),
    .io_result(x540_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_45 ( // @[package.scala 93:22:@33765.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_197 RetimeWrapper_46 ( // @[package.scala 93:22:@33779.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_191 RetimeWrapper_47 ( // @[package.scala 93:22:@33800.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper RetimeWrapper_48 ( // @[package.scala 93:22:@33816.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_212 RetimeWrapper_49 ( // @[package.scala 93:22:@33831.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  x453_sum x548_sum_1 ( // @[Math.scala 150:24:@33840.4]
    .clock(x548_sum_1_clock),
    .reset(x548_sum_1_reset),
    .io_a(x548_sum_1_io_a),
    .io_b(x548_sum_1_io_b),
    .io_flow(x548_sum_1_io_flow),
    .io_result(x548_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_50 ( // @[package.scala 93:22:@33850.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_197 RetimeWrapper_51 ( // @[package.scala 93:22:@33864.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  x453_sum x553_rdcol_1 ( // @[Math.scala 150:24:@33887.4]
    .clock(x553_rdcol_1_clock),
    .reset(x553_rdcol_1_reset),
    .io_a(x553_rdcol_1_io_a),
    .io_b(x553_rdcol_1_io_b),
    .io_flow(x553_rdcol_1_io_flow),
    .io_result(x553_rdcol_1_io_result)
  );
  x453_sum x559_sum_1 ( // @[Math.scala 150:24:@33919.4]
    .clock(x559_sum_1_clock),
    .reset(x559_sum_1_reset),
    .io_a(x559_sum_1_io_a),
    .io_b(x559_sum_1_io_b),
    .io_flow(x559_sum_1_io_flow),
    .io_result(x559_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_52 ( // @[package.scala 93:22:@33929.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_197 RetimeWrapper_53 ( // @[package.scala 93:22:@33943.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  x453_sum x565_rdcol_1 ( // @[Math.scala 150:24:@33966.4]
    .clock(x565_rdcol_1_clock),
    .reset(x565_rdcol_1_reset),
    .io_a(x565_rdcol_1_io_a),
    .io_b(x565_rdcol_1_io_b),
    .io_flow(x565_rdcol_1_io_flow),
    .io_result(x565_rdcol_1_io_result)
  );
  x453_sum x571_sum_1 ( // @[Math.scala 150:24:@33998.4]
    .clock(x571_sum_1_clock),
    .reset(x571_sum_1_reset),
    .io_a(x571_sum_1_io_a),
    .io_b(x571_sum_1_io_b),
    .io_flow(x571_sum_1_io_flow),
    .io_result(x571_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_54 ( // @[package.scala 93:22:@34008.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_197 RetimeWrapper_55 ( // @[package.scala 93:22:@34022.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper_191 RetimeWrapper_56 ( // @[package.scala 93:22:@34043.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper RetimeWrapper_57 ( // @[package.scala 93:22:@34070.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper_149 RetimeWrapper_58 ( // @[package.scala 93:22:@34105.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  x453_sum x583_sum_1 ( // @[Math.scala 150:24:@34114.4]
    .clock(x583_sum_1_clock),
    .reset(x583_sum_1_reset),
    .io_a(x583_sum_1_io_a),
    .io_b(x583_sum_1_io_b),
    .io_flow(x583_sum_1_io_flow),
    .io_result(x583_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_59 ( // @[package.scala 93:22:@34124.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_229 RetimeWrapper_60 ( // @[package.scala 93:22:@34133.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_197 RetimeWrapper_61 ( // @[package.scala 93:22:@34147.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  x453_sum x591_sum_1 ( // @[Math.scala 150:24:@34176.4]
    .clock(x591_sum_1_clock),
    .reset(x591_sum_1_reset),
    .io_a(x591_sum_1_io_a),
    .io_b(x591_sum_1_io_b),
    .io_flow(x591_sum_1_io_flow),
    .io_result(x591_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_62 ( // @[package.scala 93:22:@34186.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_197 RetimeWrapper_63 ( // @[package.scala 93:22:@34200.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  x453_sum x598_sum_1 ( // @[Math.scala 150:24:@34227.4]
    .clock(x598_sum_1_clock),
    .reset(x598_sum_1_reset),
    .io_a(x598_sum_1_io_a),
    .io_b(x598_sum_1_io_b),
    .io_flow(x598_sum_1_io_flow),
    .io_result(x598_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_64 ( // @[package.scala 93:22:@34237.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_197 RetimeWrapper_65 ( // @[package.scala 93:22:@34251.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper_191 RetimeWrapper_66 ( // @[package.scala 93:22:@34278.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  x453_sum x605_sum_1 ( // @[Math.scala 150:24:@34287.4]
    .clock(x605_sum_1_clock),
    .reset(x605_sum_1_reset),
    .io_a(x605_sum_1_io_a),
    .io_b(x605_sum_1_io_b),
    .io_flow(x605_sum_1_io_flow),
    .io_result(x605_sum_1_io_result)
  );
  RetimeWrapper_149 RetimeWrapper_67 ( // @[package.scala 93:22:@34297.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_68 ( // @[package.scala 93:22:@34306.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_197 RetimeWrapper_69 ( // @[package.scala 93:22:@34320.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  x453_sum x612_sum_1 ( // @[Math.scala 150:24:@34347.4]
    .clock(x612_sum_1_clock),
    .reset(x612_sum_1_reset),
    .io_a(x612_sum_1_io_a),
    .io_b(x612_sum_1_io_b),
    .io_flow(x612_sum_1_io_flow),
    .io_result(x612_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_70 ( // @[package.scala 93:22:@34357.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_197 RetimeWrapper_71 ( // @[package.scala 93:22:@34371.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  x453_sum x619_sum_1 ( // @[Math.scala 150:24:@34398.4]
    .clock(x619_sum_1_clock),
    .reset(x619_sum_1_reset),
    .io_a(x619_sum_1_io_a),
    .io_b(x619_sum_1_io_b),
    .io_flow(x619_sum_1_io_flow),
    .io_result(x619_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_72 ( // @[package.scala 93:22:@34408.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  RetimeWrapper_197 RetimeWrapper_73 ( // @[package.scala 93:22:@34422.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  x453_sum x624_rdrow_1 ( // @[Math.scala 150:24:@34445.4]
    .clock(x624_rdrow_1_clock),
    .reset(x624_rdrow_1_reset),
    .io_a(x624_rdrow_1_io_a),
    .io_b(x624_rdrow_1_io_b),
    .io_flow(x624_rdrow_1_io_flow),
    .io_result(x624_rdrow_1_io_result)
  );
  x453_sum x631_sum_1 ( // @[Math.scala 150:24:@34499.4]
    .clock(x631_sum_1_clock),
    .reset(x631_sum_1_reset),
    .io_a(x631_sum_1_io_a),
    .io_b(x631_sum_1_io_b),
    .io_flow(x631_sum_1_io_flow),
    .io_result(x631_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_74 ( // @[package.scala 93:22:@34509.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  RetimeWrapper_149 RetimeWrapper_75 ( // @[package.scala 93:22:@34518.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_197 RetimeWrapper_76 ( // @[package.scala 93:22:@34532.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  x453_sum x639_sum_1 ( // @[Math.scala 150:24:@34561.4]
    .clock(x639_sum_1_clock),
    .reset(x639_sum_1_reset),
    .io_a(x639_sum_1_io_a),
    .io_b(x639_sum_1_io_b),
    .io_flow(x639_sum_1_io_flow),
    .io_result(x639_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_77 ( // @[package.scala 93:22:@34571.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  RetimeWrapper_197 RetimeWrapper_78 ( // @[package.scala 93:22:@34585.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  x453_sum x646_sum_1 ( // @[Math.scala 150:24:@34612.4]
    .clock(x646_sum_1_clock),
    .reset(x646_sum_1_reset),
    .io_a(x646_sum_1_io_a),
    .io_b(x646_sum_1_io_b),
    .io_flow(x646_sum_1_io_flow),
    .io_result(x646_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_79 ( // @[package.scala 93:22:@34622.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper_197 RetimeWrapper_80 ( // @[package.scala 93:22:@34636.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  x453_sum x653_sum_1 ( // @[Math.scala 150:24:@34663.4]
    .clock(x653_sum_1_clock),
    .reset(x653_sum_1_reset),
    .io_a(x653_sum_1_io_a),
    .io_b(x653_sum_1_io_b),
    .io_flow(x653_sum_1_io_flow),
    .io_result(x653_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_81 ( // @[package.scala 93:22:@34673.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_197 RetimeWrapper_82 ( // @[package.scala 93:22:@34687.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  x453_sum x660_sum_1 ( // @[Math.scala 150:24:@34714.4]
    .clock(x660_sum_1_clock),
    .reset(x660_sum_1_reset),
    .io_a(x660_sum_1_io_a),
    .io_b(x660_sum_1_io_b),
    .io_flow(x660_sum_1_io_flow),
    .io_result(x660_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_83 ( // @[package.scala 93:22:@34724.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  RetimeWrapper_197 RetimeWrapper_84 ( // @[package.scala 93:22:@34738.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  x453_sum x667_sum_1 ( // @[Math.scala 150:24:@34765.4]
    .clock(x667_sum_1_clock),
    .reset(x667_sum_1_reset),
    .io_a(x667_sum_1_io_a),
    .io_b(x667_sum_1_io_b),
    .io_flow(x667_sum_1_io_flow),
    .io_result(x667_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_85 ( // @[package.scala 93:22:@34775.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  RetimeWrapper_197 RetimeWrapper_86 ( // @[package.scala 93:22:@34789.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  x453_sum x672_rdrow_1 ( // @[Math.scala 150:24:@34812.4]
    .clock(x672_rdrow_1_clock),
    .reset(x672_rdrow_1_reset),
    .io_a(x672_rdrow_1_io_a),
    .io_b(x672_rdrow_1_io_b),
    .io_flow(x672_rdrow_1_io_flow),
    .io_result(x672_rdrow_1_io_result)
  );
  x453_sum x679_sum_1 ( // @[Math.scala 150:24:@34866.4]
    .clock(x679_sum_1_clock),
    .reset(x679_sum_1_reset),
    .io_a(x679_sum_1_io_a),
    .io_b(x679_sum_1_io_b),
    .io_flow(x679_sum_1_io_flow),
    .io_result(x679_sum_1_io_result)
  );
  RetimeWrapper_149 RetimeWrapper_87 ( // @[package.scala 93:22:@34876.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  RetimeWrapper RetimeWrapper_88 ( // @[package.scala 93:22:@34885.4]
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  RetimeWrapper_197 RetimeWrapper_89 ( // @[package.scala 93:22:@34899.4]
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  x453_sum x687_sum_1 ( // @[Math.scala 150:24:@34926.4]
    .clock(x687_sum_1_clock),
    .reset(x687_sum_1_reset),
    .io_a(x687_sum_1_io_a),
    .io_b(x687_sum_1_io_b),
    .io_flow(x687_sum_1_io_flow),
    .io_result(x687_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_90 ( // @[package.scala 93:22:@34936.4]
    .clock(RetimeWrapper_90_clock),
    .reset(RetimeWrapper_90_reset),
    .io_flow(RetimeWrapper_90_io_flow),
    .io_in(RetimeWrapper_90_io_in),
    .io_out(RetimeWrapper_90_io_out)
  );
  RetimeWrapper_197 RetimeWrapper_91 ( // @[package.scala 93:22:@34950.4]
    .clock(RetimeWrapper_91_clock),
    .reset(RetimeWrapper_91_reset),
    .io_flow(RetimeWrapper_91_io_flow),
    .io_in(RetimeWrapper_91_io_in),
    .io_out(RetimeWrapper_91_io_out)
  );
  x453_sum x694_sum_1 ( // @[Math.scala 150:24:@34979.4]
    .clock(x694_sum_1_clock),
    .reset(x694_sum_1_reset),
    .io_a(x694_sum_1_io_a),
    .io_b(x694_sum_1_io_b),
    .io_flow(x694_sum_1_io_flow),
    .io_result(x694_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_92 ( // @[package.scala 93:22:@34989.4]
    .clock(RetimeWrapper_92_clock),
    .reset(RetimeWrapper_92_reset),
    .io_flow(RetimeWrapper_92_io_flow),
    .io_in(RetimeWrapper_92_io_in),
    .io_out(RetimeWrapper_92_io_out)
  );
  RetimeWrapper_197 RetimeWrapper_93 ( // @[package.scala 93:22:@35003.4]
    .clock(RetimeWrapper_93_clock),
    .reset(RetimeWrapper_93_reset),
    .io_flow(RetimeWrapper_93_io_flow),
    .io_in(RetimeWrapper_93_io_in),
    .io_out(RetimeWrapper_93_io_out)
  );
  x453_sum x701_sum_1 ( // @[Math.scala 150:24:@35030.4]
    .clock(x701_sum_1_clock),
    .reset(x701_sum_1_reset),
    .io_a(x701_sum_1_io_a),
    .io_b(x701_sum_1_io_b),
    .io_flow(x701_sum_1_io_flow),
    .io_result(x701_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_94 ( // @[package.scala 93:22:@35040.4]
    .clock(RetimeWrapper_94_clock),
    .reset(RetimeWrapper_94_reset),
    .io_flow(RetimeWrapper_94_io_flow),
    .io_in(RetimeWrapper_94_io_in),
    .io_out(RetimeWrapper_94_io_out)
  );
  RetimeWrapper_197 RetimeWrapper_95 ( // @[package.scala 93:22:@35054.4]
    .clock(RetimeWrapper_95_clock),
    .reset(RetimeWrapper_95_reset),
    .io_flow(RetimeWrapper_95_io_flow),
    .io_in(RetimeWrapper_95_io_in),
    .io_out(RetimeWrapper_95_io_out)
  );
  x453_sum x708_sum_1 ( // @[Math.scala 150:24:@35081.4]
    .clock(x708_sum_1_clock),
    .reset(x708_sum_1_reset),
    .io_a(x708_sum_1_io_a),
    .io_b(x708_sum_1_io_b),
    .io_flow(x708_sum_1_io_flow),
    .io_result(x708_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_96 ( // @[package.scala 93:22:@35091.4]
    .clock(RetimeWrapper_96_clock),
    .reset(RetimeWrapper_96_reset),
    .io_flow(RetimeWrapper_96_io_flow),
    .io_in(RetimeWrapper_96_io_in),
    .io_out(RetimeWrapper_96_io_out)
  );
  RetimeWrapper_197 RetimeWrapper_97 ( // @[package.scala 93:22:@35105.4]
    .clock(RetimeWrapper_97_clock),
    .reset(RetimeWrapper_97_reset),
    .io_flow(RetimeWrapper_97_io_flow),
    .io_in(RetimeWrapper_97_io_in),
    .io_out(RetimeWrapper_97_io_out)
  );
  x453_sum x715_sum_1 ( // @[Math.scala 150:24:@35132.4]
    .clock(x715_sum_1_clock),
    .reset(x715_sum_1_reset),
    .io_a(x715_sum_1_io_a),
    .io_b(x715_sum_1_io_b),
    .io_flow(x715_sum_1_io_flow),
    .io_result(x715_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_98 ( // @[package.scala 93:22:@35142.4]
    .clock(RetimeWrapper_98_clock),
    .reset(RetimeWrapper_98_reset),
    .io_flow(RetimeWrapper_98_io_flow),
    .io_in(RetimeWrapper_98_io_in),
    .io_out(RetimeWrapper_98_io_out)
  );
  RetimeWrapper_197 RetimeWrapper_99 ( // @[package.scala 93:22:@35156.4]
    .clock(RetimeWrapper_99_clock),
    .reset(RetimeWrapper_99_reset),
    .io_flow(RetimeWrapper_99_io_flow),
    .io_in(RetimeWrapper_99_io_in),
    .io_out(RetimeWrapper_99_io_out)
  );
  x725_x11 x725_x11_1 ( // @[Math.scala 150:24:@35202.4]
    .clock(x725_x11_1_clock),
    .reset(x725_x11_1_reset),
    .io_a(x725_x11_1_io_a),
    .io_b(x725_x11_1_io_b),
    .io_flow(x725_x11_1_io_flow),
    .io_result(x725_x11_1_io_result)
  );
  x725_x11 x726_x12_1 ( // @[Math.scala 150:24:@35212.4]
    .clock(x726_x12_1_clock),
    .reset(x726_x12_1_reset),
    .io_a(x726_x12_1_io_a),
    .io_b(x726_x12_1_io_b),
    .io_flow(x726_x12_1_io_flow),
    .io_result(x726_x12_1_io_result)
  );
  x725_x11 x727_x11_1 ( // @[Math.scala 150:24:@35222.4]
    .clock(x727_x11_1_clock),
    .reset(x727_x11_1_reset),
    .io_a(x727_x11_1_io_a),
    .io_b(x727_x11_1_io_b),
    .io_flow(x727_x11_1_io_flow),
    .io_result(x727_x11_1_io_result)
  );
  x725_x11 x728_x12_1 ( // @[Math.scala 150:24:@35232.4]
    .clock(x728_x12_1_clock),
    .reset(x728_x12_1_reset),
    .io_a(x728_x12_1_io_a),
    .io_b(x728_x12_1_io_b),
    .io_flow(x728_x12_1_io_flow),
    .io_result(x728_x12_1_io_result)
  );
  x729_x11 x729_x11_1 ( // @[Math.scala 150:24:@35242.4]
    .io_a(x729_x11_1_io_a),
    .io_b(x729_x11_1_io_b),
    .io_result(x729_x11_1_io_result)
  );
  x729_x11 x730_x12_1 ( // @[Math.scala 150:24:@35252.4]
    .io_a(x730_x12_1_io_a),
    .io_b(x730_x12_1_io_b),
    .io_result(x730_x12_1_io_result)
  );
  x729_x11 x731_x11_1 ( // @[Math.scala 150:24:@35262.4]
    .io_a(x731_x11_1_io_a),
    .io_b(x731_x11_1_io_b),
    .io_result(x731_x11_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_100 ( // @[package.scala 93:22:@35272.4]
    .clock(RetimeWrapper_100_clock),
    .reset(RetimeWrapper_100_reset),
    .io_flow(RetimeWrapper_100_io_flow),
    .io_in(RetimeWrapper_100_io_in),
    .io_out(RetimeWrapper_100_io_out)
  );
  x729_x11 x732_sum_1 ( // @[Math.scala 150:24:@35281.4]
    .io_a(x732_sum_1_io_a),
    .io_b(x732_sum_1_io_b),
    .io_result(x732_sum_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_101 ( // @[package.scala 93:22:@35295.4]
    .clock(RetimeWrapper_101_clock),
    .reset(RetimeWrapper_101_reset),
    .io_flow(RetimeWrapper_101_io_flow),
    .io_in(RetimeWrapper_101_io_in),
    .io_out(RetimeWrapper_101_io_out)
  );
  x725_x11 x739_x11_1 ( // @[Math.scala 150:24:@35330.4]
    .clock(x739_x11_1_clock),
    .reset(x739_x11_1_reset),
    .io_a(x739_x11_1_io_a),
    .io_b(x739_x11_1_io_b),
    .io_flow(x739_x11_1_io_flow),
    .io_result(x739_x11_1_io_result)
  );
  x725_x11 x740_x12_1 ( // @[Math.scala 150:24:@35340.4]
    .clock(x740_x12_1_clock),
    .reset(x740_x12_1_reset),
    .io_a(x740_x12_1_io_a),
    .io_b(x740_x12_1_io_b),
    .io_flow(x740_x12_1_io_flow),
    .io_result(x740_x12_1_io_result)
  );
  x725_x11 x741_x11_1 ( // @[Math.scala 150:24:@35350.4]
    .clock(x741_x11_1_clock),
    .reset(x741_x11_1_reset),
    .io_a(x741_x11_1_io_a),
    .io_b(x741_x11_1_io_b),
    .io_flow(x741_x11_1_io_flow),
    .io_result(x741_x11_1_io_result)
  );
  x725_x11 x742_x12_1 ( // @[Math.scala 150:24:@35360.4]
    .clock(x742_x12_1_clock),
    .reset(x742_x12_1_reset),
    .io_a(x742_x12_1_io_a),
    .io_b(x742_x12_1_io_b),
    .io_flow(x742_x12_1_io_flow),
    .io_result(x742_x12_1_io_result)
  );
  x729_x11 x743_x11_1 ( // @[Math.scala 150:24:@35370.4]
    .io_a(x743_x11_1_io_a),
    .io_b(x743_x11_1_io_b),
    .io_result(x743_x11_1_io_result)
  );
  x729_x11 x744_x12_1 ( // @[Math.scala 150:24:@35380.4]
    .io_a(x744_x12_1_io_a),
    .io_b(x744_x12_1_io_b),
    .io_result(x744_x12_1_io_result)
  );
  x729_x11 x745_x11_1 ( // @[Math.scala 150:24:@35390.4]
    .io_a(x745_x11_1_io_a),
    .io_b(x745_x11_1_io_b),
    .io_result(x745_x11_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_102 ( // @[package.scala 93:22:@35400.4]
    .clock(RetimeWrapper_102_clock),
    .reset(RetimeWrapper_102_reset),
    .io_flow(RetimeWrapper_102_io_flow),
    .io_in(RetimeWrapper_102_io_in),
    .io_out(RetimeWrapper_102_io_out)
  );
  x729_x11 x746_sum_1 ( // @[Math.scala 150:24:@35411.4]
    .io_a(x746_sum_1_io_a),
    .io_b(x746_sum_1_io_b),
    .io_result(x746_sum_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_103 ( // @[package.scala 93:22:@35425.4]
    .clock(RetimeWrapper_103_clock),
    .reset(RetimeWrapper_103_reset),
    .io_flow(RetimeWrapper_103_io_flow),
    .io_in(RetimeWrapper_103_io_in),
    .io_out(RetimeWrapper_103_io_out)
  );
  x725_x11 x752_x11_1 ( // @[Math.scala 150:24:@35455.4]
    .clock(x752_x11_1_clock),
    .reset(x752_x11_1_reset),
    .io_a(x752_x11_1_io_a),
    .io_b(x752_x11_1_io_b),
    .io_flow(x752_x11_1_io_flow),
    .io_result(x752_x11_1_io_result)
  );
  x725_x11 x753_x12_1 ( // @[Math.scala 150:24:@35465.4]
    .clock(x753_x12_1_clock),
    .reset(x753_x12_1_reset),
    .io_a(x753_x12_1_io_a),
    .io_b(x753_x12_1_io_b),
    .io_flow(x753_x12_1_io_flow),
    .io_result(x753_x12_1_io_result)
  );
  x725_x11 x754_x11_1 ( // @[Math.scala 150:24:@35475.4]
    .clock(x754_x11_1_clock),
    .reset(x754_x11_1_reset),
    .io_a(x754_x11_1_io_a),
    .io_b(x754_x11_1_io_b),
    .io_flow(x754_x11_1_io_flow),
    .io_result(x754_x11_1_io_result)
  );
  x725_x11 x755_x12_1 ( // @[Math.scala 150:24:@35485.4]
    .clock(x755_x12_1_clock),
    .reset(x755_x12_1_reset),
    .io_a(x755_x12_1_io_a),
    .io_b(x755_x12_1_io_b),
    .io_flow(x755_x12_1_io_flow),
    .io_result(x755_x12_1_io_result)
  );
  x729_x11 x756_x11_1 ( // @[Math.scala 150:24:@35495.4]
    .io_a(x756_x11_1_io_a),
    .io_b(x756_x11_1_io_b),
    .io_result(x756_x11_1_io_result)
  );
  x729_x11 x757_x12_1 ( // @[Math.scala 150:24:@35505.4]
    .io_a(x757_x12_1_io_a),
    .io_b(x757_x12_1_io_b),
    .io_result(x757_x12_1_io_result)
  );
  x729_x11 x758_x11_1 ( // @[Math.scala 150:24:@35515.4]
    .io_a(x758_x11_1_io_a),
    .io_b(x758_x11_1_io_b),
    .io_result(x758_x11_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_104 ( // @[package.scala 93:22:@35525.4]
    .clock(RetimeWrapper_104_clock),
    .reset(RetimeWrapper_104_reset),
    .io_flow(RetimeWrapper_104_io_flow),
    .io_in(RetimeWrapper_104_io_in),
    .io_out(RetimeWrapper_104_io_out)
  );
  x729_x11 x759_sum_1 ( // @[Math.scala 150:24:@35534.4]
    .io_a(x759_sum_1_io_a),
    .io_b(x759_sum_1_io_b),
    .io_result(x759_sum_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_105 ( // @[package.scala 93:22:@35548.4]
    .clock(RetimeWrapper_105_clock),
    .reset(RetimeWrapper_105_reset),
    .io_flow(RetimeWrapper_105_io_flow),
    .io_in(RetimeWrapper_105_io_in),
    .io_out(RetimeWrapper_105_io_out)
  );
  x725_x11 x765_x11_1 ( // @[Math.scala 150:24:@35578.4]
    .clock(x765_x11_1_clock),
    .reset(x765_x11_1_reset),
    .io_a(x765_x11_1_io_a),
    .io_b(x765_x11_1_io_b),
    .io_flow(x765_x11_1_io_flow),
    .io_result(x765_x11_1_io_result)
  );
  x725_x11 x766_x12_1 ( // @[Math.scala 150:24:@35588.4]
    .clock(x766_x12_1_clock),
    .reset(x766_x12_1_reset),
    .io_a(x766_x12_1_io_a),
    .io_b(x766_x12_1_io_b),
    .io_flow(x766_x12_1_io_flow),
    .io_result(x766_x12_1_io_result)
  );
  x725_x11 x767_x11_1 ( // @[Math.scala 150:24:@35598.4]
    .clock(x767_x11_1_clock),
    .reset(x767_x11_1_reset),
    .io_a(x767_x11_1_io_a),
    .io_b(x767_x11_1_io_b),
    .io_flow(x767_x11_1_io_flow),
    .io_result(x767_x11_1_io_result)
  );
  x725_x11 x768_x12_1 ( // @[Math.scala 150:24:@35608.4]
    .clock(x768_x12_1_clock),
    .reset(x768_x12_1_reset),
    .io_a(x768_x12_1_io_a),
    .io_b(x768_x12_1_io_b),
    .io_flow(x768_x12_1_io_flow),
    .io_result(x768_x12_1_io_result)
  );
  x729_x11 x769_x11_1 ( // @[Math.scala 150:24:@35618.4]
    .io_a(x769_x11_1_io_a),
    .io_b(x769_x11_1_io_b),
    .io_result(x769_x11_1_io_result)
  );
  x729_x11 x770_x12_1 ( // @[Math.scala 150:24:@35628.4]
    .io_a(x770_x12_1_io_a),
    .io_b(x770_x12_1_io_b),
    .io_result(x770_x12_1_io_result)
  );
  x729_x11 x771_x11_1 ( // @[Math.scala 150:24:@35638.4]
    .io_a(x771_x11_1_io_a),
    .io_b(x771_x11_1_io_b),
    .io_result(x771_x11_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_106 ( // @[package.scala 93:22:@35648.4]
    .clock(RetimeWrapper_106_clock),
    .reset(RetimeWrapper_106_reset),
    .io_flow(RetimeWrapper_106_io_flow),
    .io_in(RetimeWrapper_106_io_in),
    .io_out(RetimeWrapper_106_io_out)
  );
  x729_x11 x772_sum_1 ( // @[Math.scala 150:24:@35657.4]
    .io_a(x772_sum_1_io_a),
    .io_b(x772_sum_1_io_b),
    .io_result(x772_sum_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_107 ( // @[package.scala 93:22:@35671.4]
    .clock(RetimeWrapper_107_clock),
    .reset(RetimeWrapper_107_reset),
    .io_flow(RetimeWrapper_107_io_flow),
    .io_in(RetimeWrapper_107_io_in),
    .io_out(RetimeWrapper_107_io_out)
  );
  x725_x11 x777_x11_1 ( // @[Math.scala 150:24:@35696.4]
    .clock(x777_x11_1_clock),
    .reset(x777_x11_1_reset),
    .io_a(x777_x11_1_io_a),
    .io_b(x777_x11_1_io_b),
    .io_flow(x777_x11_1_io_flow),
    .io_result(x777_x11_1_io_result)
  );
  x725_x11 x778_x12_1 ( // @[Math.scala 150:24:@35706.4]
    .clock(x778_x12_1_clock),
    .reset(x778_x12_1_reset),
    .io_a(x778_x12_1_io_a),
    .io_b(x778_x12_1_io_b),
    .io_flow(x778_x12_1_io_flow),
    .io_result(x778_x12_1_io_result)
  );
  x725_x11 x779_x11_1 ( // @[Math.scala 150:24:@35716.4]
    .clock(x779_x11_1_clock),
    .reset(x779_x11_1_reset),
    .io_a(x779_x11_1_io_a),
    .io_b(x779_x11_1_io_b),
    .io_flow(x779_x11_1_io_flow),
    .io_result(x779_x11_1_io_result)
  );
  x725_x11 x780_x12_1 ( // @[Math.scala 150:24:@35726.4]
    .clock(x780_x12_1_clock),
    .reset(x780_x12_1_reset),
    .io_a(x780_x12_1_io_a),
    .io_b(x780_x12_1_io_b),
    .io_flow(x780_x12_1_io_flow),
    .io_result(x780_x12_1_io_result)
  );
  x729_x11 x781_x11_1 ( // @[Math.scala 150:24:@35736.4]
    .io_a(x781_x11_1_io_a),
    .io_b(x781_x11_1_io_b),
    .io_result(x781_x11_1_io_result)
  );
  x729_x11 x782_x12_1 ( // @[Math.scala 150:24:@35746.4]
    .io_a(x782_x12_1_io_a),
    .io_b(x782_x12_1_io_b),
    .io_result(x782_x12_1_io_result)
  );
  x729_x11 x783_x11_1 ( // @[Math.scala 150:24:@35756.4]
    .io_a(x783_x11_1_io_a),
    .io_b(x783_x11_1_io_b),
    .io_result(x783_x11_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_108 ( // @[package.scala 93:22:@35766.4]
    .clock(RetimeWrapper_108_clock),
    .reset(RetimeWrapper_108_reset),
    .io_flow(RetimeWrapper_108_io_flow),
    .io_in(RetimeWrapper_108_io_in),
    .io_out(RetimeWrapper_108_io_out)
  );
  x729_x11 x784_sum_1 ( // @[Math.scala 150:24:@35775.4]
    .io_a(x784_sum_1_io_a),
    .io_b(x784_sum_1_io_b),
    .io_result(x784_sum_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_109 ( // @[package.scala 93:22:@35789.4]
    .clock(RetimeWrapper_109_clock),
    .reset(RetimeWrapper_109_reset),
    .io_flow(RetimeWrapper_109_io_flow),
    .io_in(RetimeWrapper_109_io_in),
    .io_out(RetimeWrapper_109_io_out)
  );
  x725_x11 x788_x11_1 ( // @[Math.scala 150:24:@35809.4]
    .clock(x788_x11_1_clock),
    .reset(x788_x11_1_reset),
    .io_a(x788_x11_1_io_a),
    .io_b(x788_x11_1_io_b),
    .io_flow(x788_x11_1_io_flow),
    .io_result(x788_x11_1_io_result)
  );
  x725_x11 x789_x12_1 ( // @[Math.scala 150:24:@35819.4]
    .clock(x789_x12_1_clock),
    .reset(x789_x12_1_reset),
    .io_a(x789_x12_1_io_a),
    .io_b(x789_x12_1_io_b),
    .io_flow(x789_x12_1_io_flow),
    .io_result(x789_x12_1_io_result)
  );
  x725_x11 x790_x11_1 ( // @[Math.scala 150:24:@35829.4]
    .clock(x790_x11_1_clock),
    .reset(x790_x11_1_reset),
    .io_a(x790_x11_1_io_a),
    .io_b(x790_x11_1_io_b),
    .io_flow(x790_x11_1_io_flow),
    .io_result(x790_x11_1_io_result)
  );
  x725_x11 x791_x12_1 ( // @[Math.scala 150:24:@35841.4]
    .clock(x791_x12_1_clock),
    .reset(x791_x12_1_reset),
    .io_a(x791_x12_1_io_a),
    .io_b(x791_x12_1_io_b),
    .io_flow(x791_x12_1_io_flow),
    .io_result(x791_x12_1_io_result)
  );
  x729_x11 x792_x11_1 ( // @[Math.scala 150:24:@35851.4]
    .io_a(x792_x11_1_io_a),
    .io_b(x792_x11_1_io_b),
    .io_result(x792_x11_1_io_result)
  );
  x729_x11 x793_x12_1 ( // @[Math.scala 150:24:@35861.4]
    .io_a(x793_x12_1_io_a),
    .io_b(x793_x12_1_io_b),
    .io_result(x793_x12_1_io_result)
  );
  x729_x11 x794_x11_1 ( // @[Math.scala 150:24:@35871.4]
    .io_a(x794_x11_1_io_a),
    .io_b(x794_x11_1_io_b),
    .io_result(x794_x11_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_110 ( // @[package.scala 93:22:@35881.4]
    .clock(RetimeWrapper_110_clock),
    .reset(RetimeWrapper_110_reset),
    .io_flow(RetimeWrapper_110_io_flow),
    .io_in(RetimeWrapper_110_io_in),
    .io_out(RetimeWrapper_110_io_out)
  );
  x729_x11 x795_sum_1 ( // @[Math.scala 150:24:@35890.4]
    .io_a(x795_sum_1_io_a),
    .io_b(x795_sum_1_io_b),
    .io_result(x795_sum_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_111 ( // @[package.scala 93:22:@35904.4]
    .clock(RetimeWrapper_111_clock),
    .reset(RetimeWrapper_111_reset),
    .io_flow(RetimeWrapper_111_io_flow),
    .io_in(RetimeWrapper_111_io_in),
    .io_out(RetimeWrapper_111_io_out)
  );
  x725_x11 x799_x11_1 ( // @[Math.scala 150:24:@35924.4]
    .clock(x799_x11_1_clock),
    .reset(x799_x11_1_reset),
    .io_a(x799_x11_1_io_a),
    .io_b(x799_x11_1_io_b),
    .io_flow(x799_x11_1_io_flow),
    .io_result(x799_x11_1_io_result)
  );
  x725_x11 x800_x12_1 ( // @[Math.scala 150:24:@35934.4]
    .clock(x800_x12_1_clock),
    .reset(x800_x12_1_reset),
    .io_a(x800_x12_1_io_a),
    .io_b(x800_x12_1_io_b),
    .io_flow(x800_x12_1_io_flow),
    .io_result(x800_x12_1_io_result)
  );
  x725_x11 x801_x11_1 ( // @[Math.scala 150:24:@35944.4]
    .clock(x801_x11_1_clock),
    .reset(x801_x11_1_reset),
    .io_a(x801_x11_1_io_a),
    .io_b(x801_x11_1_io_b),
    .io_flow(x801_x11_1_io_flow),
    .io_result(x801_x11_1_io_result)
  );
  x725_x11 x802_x12_1 ( // @[Math.scala 150:24:@35954.4]
    .clock(x802_x12_1_clock),
    .reset(x802_x12_1_reset),
    .io_a(x802_x12_1_io_a),
    .io_b(x802_x12_1_io_b),
    .io_flow(x802_x12_1_io_flow),
    .io_result(x802_x12_1_io_result)
  );
  x729_x11 x803_x11_1 ( // @[Math.scala 150:24:@35964.4]
    .io_a(x803_x11_1_io_a),
    .io_b(x803_x11_1_io_b),
    .io_result(x803_x11_1_io_result)
  );
  x729_x11 x804_x12_1 ( // @[Math.scala 150:24:@35974.4]
    .io_a(x804_x12_1_io_a),
    .io_b(x804_x12_1_io_b),
    .io_result(x804_x12_1_io_result)
  );
  x729_x11 x805_x11_1 ( // @[Math.scala 150:24:@35984.4]
    .io_a(x805_x11_1_io_a),
    .io_b(x805_x11_1_io_b),
    .io_result(x805_x11_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_112 ( // @[package.scala 93:22:@35994.4]
    .clock(RetimeWrapper_112_clock),
    .reset(RetimeWrapper_112_reset),
    .io_flow(RetimeWrapper_112_io_flow),
    .io_in(RetimeWrapper_112_io_in),
    .io_out(RetimeWrapper_112_io_out)
  );
  x729_x11 x806_sum_1 ( // @[Math.scala 150:24:@36003.4]
    .io_a(x806_sum_1_io_a),
    .io_b(x806_sum_1_io_b),
    .io_result(x806_sum_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_113 ( // @[package.scala 93:22:@36017.4]
    .clock(RetimeWrapper_113_clock),
    .reset(RetimeWrapper_113_reset),
    .io_flow(RetimeWrapper_113_io_flow),
    .io_in(RetimeWrapper_113_io_in),
    .io_out(RetimeWrapper_113_io_out)
  );
  x725_x11 x811_x11_1 ( // @[Math.scala 150:24:@36042.4]
    .clock(x811_x11_1_clock),
    .reset(x811_x11_1_reset),
    .io_a(x811_x11_1_io_a),
    .io_b(x811_x11_1_io_b),
    .io_flow(x811_x11_1_io_flow),
    .io_result(x811_x11_1_io_result)
  );
  x725_x11 x812_x12_1 ( // @[Math.scala 150:24:@36052.4]
    .clock(x812_x12_1_clock),
    .reset(x812_x12_1_reset),
    .io_a(x812_x12_1_io_a),
    .io_b(x812_x12_1_io_b),
    .io_flow(x812_x12_1_io_flow),
    .io_result(x812_x12_1_io_result)
  );
  x725_x11 x813_x11_1 ( // @[Math.scala 150:24:@36062.4]
    .clock(x813_x11_1_clock),
    .reset(x813_x11_1_reset),
    .io_a(x813_x11_1_io_a),
    .io_b(x813_x11_1_io_b),
    .io_flow(x813_x11_1_io_flow),
    .io_result(x813_x11_1_io_result)
  );
  x725_x11 x814_x12_1 ( // @[Math.scala 150:24:@36072.4]
    .clock(x814_x12_1_clock),
    .reset(x814_x12_1_reset),
    .io_a(x814_x12_1_io_a),
    .io_b(x814_x12_1_io_b),
    .io_flow(x814_x12_1_io_flow),
    .io_result(x814_x12_1_io_result)
  );
  x729_x11 x815_x11_1 ( // @[Math.scala 150:24:@36082.4]
    .io_a(x815_x11_1_io_a),
    .io_b(x815_x11_1_io_b),
    .io_result(x815_x11_1_io_result)
  );
  x729_x11 x816_x12_1 ( // @[Math.scala 150:24:@36092.4]
    .io_a(x816_x12_1_io_a),
    .io_b(x816_x12_1_io_b),
    .io_result(x816_x12_1_io_result)
  );
  x729_x11 x817_x11_1 ( // @[Math.scala 150:24:@36102.4]
    .io_a(x817_x11_1_io_a),
    .io_b(x817_x11_1_io_b),
    .io_result(x817_x11_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_114 ( // @[package.scala 93:22:@36112.4]
    .clock(RetimeWrapper_114_clock),
    .reset(RetimeWrapper_114_reset),
    .io_flow(RetimeWrapper_114_io_flow),
    .io_in(RetimeWrapper_114_io_in),
    .io_out(RetimeWrapper_114_io_out)
  );
  x729_x11 x818_sum_1 ( // @[Math.scala 150:24:@36121.4]
    .io_a(x818_sum_1_io_a),
    .io_b(x818_sum_1_io_b),
    .io_result(x818_sum_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_115 ( // @[package.scala 93:22:@36135.4]
    .clock(RetimeWrapper_115_clock),
    .reset(RetimeWrapper_115_reset),
    .io_flow(RetimeWrapper_115_io_flow),
    .io_in(RetimeWrapper_115_io_in),
    .io_out(RetimeWrapper_115_io_out)
  );
  RetimeWrapper_336 RetimeWrapper_116 ( // @[package.scala 93:22:@36163.4]
    .clock(RetimeWrapper_116_clock),
    .reset(RetimeWrapper_116_reset),
    .io_flow(RetimeWrapper_116_io_flow),
    .io_in(RetimeWrapper_116_io_in),
    .io_out(RetimeWrapper_116_io_out)
  );
  RetimeWrapper_12 RetimeWrapper_117 ( // @[package.scala 93:22:@36172.4]
    .clock(RetimeWrapper_117_clock),
    .reset(RetimeWrapper_117_reset),
    .io_flow(RetimeWrapper_117_io_flow),
    .io_in(RetimeWrapper_117_io_in),
    .io_out(RetimeWrapper_117_io_out)
  );
  RetimeWrapper_12 RetimeWrapper_118 ( // @[package.scala 93:22:@36181.4]
    .clock(RetimeWrapper_118_clock),
    .reset(RetimeWrapper_118_reset),
    .io_flow(RetimeWrapper_118_io_flow),
    .io_in(RetimeWrapper_118_io_in),
    .io_out(RetimeWrapper_118_io_out)
  );
  RetimeWrapper_12 RetimeWrapper_119 ( // @[package.scala 93:22:@36190.4]
    .clock(RetimeWrapper_119_clock),
    .reset(RetimeWrapper_119_reset),
    .io_flow(RetimeWrapper_119_io_flow),
    .io_in(RetimeWrapper_119_io_in),
    .io_out(RetimeWrapper_119_io_out)
  );
  assign b437 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 62:18:@32524.4]
  assign b438 = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 63:18:@32525.4]
  assign _T_206 = b437 & b438; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 68:30:@32740.4]
  assign _T_207 = _T_206 & io_sigsIn_datapathEn; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 68:37:@32741.4]
  assign _T_211 = io_in_x426_TID == 8'h0; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 70:76:@32746.4]
  assign _T_212 = _T_207 & _T_211; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 70:62:@32747.4]
  assign _T_214 = io_in_x426_TDEST == 8'h0; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 70:101:@32748.4]
  assign x902_x440_D1_0_number = RetimeWrapper_io_out; // @[package.scala 96:25:@32757.4 package.scala 96:25:@32758.4]
  assign b435_number = __io_result; // @[Math.scala 712:22:@32509.4 Math.scala 713:14:@32510.4]
  assign _T_254 = $signed(b435_number); // @[Math.scala 499:52:@32785.4]
  assign x444 = $signed(32'sh1) == $signed(_T_254); // @[Math.scala 499:44:@32793.4]
  assign x445 = $signed(32'sh2) == $signed(_T_254); // @[Math.scala 499:44:@32800.4]
  assign x446 = $signed(32'sh3) == $signed(_T_254); // @[Math.scala 499:44:@32807.4]
  assign _T_301 = x444 ? 32'h1 : 32'h0; // @[Mux.scala 19:72:@32819.4]
  assign _T_303 = x445 ? 32'h2 : 32'h0; // @[Mux.scala 19:72:@32820.4]
  assign _T_305 = x446 ? 32'h3 : 32'h0; // @[Mux.scala 19:72:@32821.4]
  assign _T_307 = _T_301 | _T_303; // @[Mux.scala 19:72:@32823.4]
  assign x447_number = _T_307 | _T_305; // @[Mux.scala 19:72:@32824.4]
  assign _T_319 = $signed(x447_number); // @[Math.scala 406:49:@32834.4]
  assign _T_321 = $signed(_T_319) & $signed(32'sh3); // @[Math.scala 406:56:@32836.4]
  assign _T_322 = $signed(_T_321); // @[Math.scala 406:56:@32837.4]
  assign _T_327 = x447_number[31]; // @[FixedPoint.scala 50:25:@32843.4]
  assign _T_331 = _T_327 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@32845.4]
  assign _T_332 = x447_number[31:2]; // @[FixedPoint.scala 18:52:@32846.4]
  assign b436_number = __1_io_result; // @[Math.scala 712:22:@32521.4 Math.scala 713:14:@32522.4]
  assign _T_337 = b436_number[31]; // @[FixedPoint.scala 50:25:@32852.4]
  assign _T_341 = _T_337 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@32854.4]
  assign _T_342 = b436_number[31:2]; // @[FixedPoint.scala 18:52:@32855.4]
  assign _T_367 = ~ io_sigsIn_break; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 113:101:@32916.4]
  assign _T_371 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@32924.4 package.scala 96:25:@32925.4]
  assign _T_373 = io_rr ? _T_371 : 1'h0; // @[implicits.scala 55:10:@32926.4]
  assign _T_374 = _T_367 & _T_373; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 113:118:@32927.4]
  assign _T_376 = _T_374 & _T_367; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 113:205:@32929.4]
  assign _T_377 = _T_376 & io_sigsIn_backpressure; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 113:224:@32930.4]
  assign x907_b437_D8 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@32911.4 package.scala 96:25:@32912.4]
  assign _T_378 = _T_377 & x907_b437_D8; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 113:250:@32931.4]
  assign x906_b438_D8 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@32902.4 package.scala 96:25:@32903.4]
  assign x459_rdcol_number = x459_rdcol_1_io_result; // @[Math.scala 154:22:@32948.4 Math.scala 155:14:@32949.4]
  assign _T_391 = x459_rdcol_number[31]; // @[FixedPoint.scala 50:25:@32955.4]
  assign _T_395 = _T_391 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@32957.4]
  assign _T_396 = x459_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@32958.4]
  assign _T_419 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@33009.4 package.scala 96:25:@33010.4]
  assign _T_421 = io_rr ? _T_419 : 1'h0; // @[implicits.scala 55:10:@33011.4]
  assign _T_422 = _T_367 & _T_421; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 132:118:@33012.4]
  assign _T_424 = _T_422 & _T_367; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 132:205:@33014.4]
  assign _T_425 = _T_424 & io_sigsIn_backpressure; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 132:224:@33015.4]
  assign _T_426 = _T_425 & x907_b437_D8; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 132:250:@33016.4]
  assign x468_rdcol_number = x468_rdcol_1_io_result; // @[Math.scala 154:22:@33033.4 Math.scala 155:14:@33034.4]
  assign _T_439 = x468_rdcol_number[31]; // @[FixedPoint.scala 50:25:@33040.4]
  assign _T_443 = _T_439 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@33042.4]
  assign _T_444 = x468_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@33043.4]
  assign _T_464 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@33085.4 package.scala 96:25:@33086.4]
  assign _T_466 = io_rr ? _T_464 : 1'h0; // @[implicits.scala 55:10:@33087.4]
  assign _T_467 = _T_367 & _T_466; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 149:118:@33088.4]
  assign _T_469 = _T_467 & _T_367; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 149:205:@33090.4]
  assign _T_470 = _T_469 & io_sigsIn_backpressure; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 149:224:@33091.4]
  assign _T_471 = _T_470 & x907_b437_D8; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 149:250:@33092.4]
  assign x477_rdcol_number = x477_rdcol_1_io_result; // @[Math.scala 154:22:@33109.4 Math.scala 155:14:@33110.4]
  assign _T_484 = x477_rdcol_number[31]; // @[FixedPoint.scala 50:25:@33116.4]
  assign _T_488 = _T_484 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@33118.4]
  assign _T_489 = x477_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@33119.4]
  assign _T_509 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@33161.4 package.scala 96:25:@33162.4]
  assign _T_511 = io_rr ? _T_509 : 1'h0; // @[implicits.scala 55:10:@33163.4]
  assign _T_512 = _T_367 & _T_511; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 166:118:@33164.4]
  assign _T_514 = _T_512 & _T_367; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 166:205:@33166.4]
  assign _T_515 = _T_514 & io_sigsIn_backpressure; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 166:224:@33167.4]
  assign _T_516 = _T_515 & x907_b437_D8; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 166:250:@33168.4]
  assign x486_rdrow_number = x486_rdrow_1_io_result; // @[Math.scala 154:22:@33185.4 Math.scala 155:14:@33186.4]
  assign _T_531 = $signed(x486_rdrow_number); // @[Math.scala 499:52:@33192.4]
  assign x488 = $signed(32'sh1) == $signed(_T_531); // @[Math.scala 499:44:@33200.4]
  assign x489 = $signed(32'sh2) == $signed(_T_531); // @[Math.scala 499:44:@33207.4]
  assign x490 = $signed(32'sh3) == $signed(_T_531); // @[Math.scala 499:44:@33214.4]
  assign _T_578 = x488 ? 32'h1 : 32'h0; // @[Mux.scala 19:72:@33226.4]
  assign _T_580 = x489 ? 32'h2 : 32'h0; // @[Mux.scala 19:72:@33227.4]
  assign _T_582 = x490 ? 32'h3 : 32'h0; // @[Mux.scala 19:72:@33228.4]
  assign _T_584 = _T_578 | _T_580; // @[Mux.scala 19:72:@33230.4]
  assign x491_number = _T_584 | _T_582; // @[Mux.scala 19:72:@33231.4]
  assign _T_598 = $signed(x491_number); // @[Math.scala 406:49:@33243.4]
  assign _T_600 = $signed(_T_598) & $signed(32'sh3); // @[Math.scala 406:56:@33245.4]
  assign _T_601 = $signed(_T_600); // @[Math.scala 406:56:@33246.4]
  assign _T_606 = x491_number[31]; // @[FixedPoint.scala 50:25:@33252.4]
  assign _T_610 = _T_606 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@33254.4]
  assign _T_611 = x491_number[31:2]; // @[FixedPoint.scala 18:52:@33255.4]
  assign _T_637 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@33315.4 package.scala 96:25:@33316.4]
  assign _T_639 = io_rr ? _T_637 : 1'h0; // @[implicits.scala 55:10:@33317.4]
  assign _T_640 = _T_367 & _T_639; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 207:166:@33318.4]
  assign _T_642 = _T_640 & _T_367; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 207:253:@33320.4]
  assign _T_643 = _T_642 & io_sigsIn_backpressure; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 207:272:@33321.4]
  assign _T_644 = _T_643 & x907_b437_D8; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 207:298:@33322.4]
  assign _T_665 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@33370.4 package.scala 96:25:@33371.4]
  assign _T_667 = io_rr ? _T_665 : 1'h0; // @[implicits.scala 55:10:@33372.4]
  assign _T_668 = _T_367 & _T_667; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 220:166:@33373.4]
  assign _T_670 = _T_668 & _T_367; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 220:253:@33375.4]
  assign _T_671 = _T_670 & io_sigsIn_backpressure; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 220:272:@33376.4]
  assign _T_672 = _T_671 & x907_b437_D8; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 220:298:@33377.4]
  assign _T_693 = RetimeWrapper_27_io_out; // @[package.scala 96:25:@33425.4 package.scala 96:25:@33426.4]
  assign _T_695 = io_rr ? _T_693 : 1'h0; // @[implicits.scala 55:10:@33427.4]
  assign _T_696 = _T_367 & _T_695; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 233:166:@33428.4]
  assign _T_698 = _T_696 & _T_367; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 233:253:@33430.4]
  assign _T_699 = _T_698 & io_sigsIn_backpressure; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 233:272:@33431.4]
  assign _T_700 = _T_699 & x907_b437_D8; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 233:298:@33432.4]
  assign _T_721 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@33480.4 package.scala 96:25:@33481.4]
  assign _T_723 = io_rr ? _T_721 : 1'h0; // @[implicits.scala 55:10:@33482.4]
  assign _T_724 = _T_367 & _T_723; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 246:166:@33483.4]
  assign _T_726 = _T_724 & _T_367; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 246:253:@33485.4]
  assign _T_727 = _T_726 & io_sigsIn_backpressure; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 246:272:@33486.4]
  assign _T_728 = _T_727 & x907_b437_D8; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 246:298:@33487.4]
  assign x925_x486_rdrow_D10_number = RetimeWrapper_31_io_out; // @[package.scala 96:25:@33501.4 package.scala 96:25:@33502.4]
  assign _T_740 = $signed(x925_x486_rdrow_D10_number); // @[Math.scala 406:49:@33508.4]
  assign _T_742 = $signed(_T_740) & $signed(32'sh3); // @[Math.scala 406:56:@33510.4]
  assign _T_743 = $signed(_T_742); // @[Math.scala 406:56:@33511.4]
  assign x894_number = $unsigned(_T_743); // @[implicits.scala 133:21:@33512.4]
  assign x517 = $signed(_T_740) < $signed(32'sh0); // @[Math.scala 465:44:@33520.4]
  assign x926_x477_rdcol_D10_number = RetimeWrapper_32_io_out; // @[package.scala 96:25:@33528.4 package.scala 96:25:@33529.4]
  assign _T_761 = $signed(x926_x477_rdcol_D10_number); // @[Math.scala 465:37:@33534.4]
  assign x518 = $signed(_T_761) < $signed(32'sh0); // @[Math.scala 465:44:@33536.4]
  assign x519 = x517 | x518; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 259:24:@33539.4]
  assign _T_775 = $signed(x894_number); // @[Math.scala 406:49:@33548.4]
  assign _T_777 = $signed(_T_775) & $signed(32'sh3); // @[Math.scala 406:56:@33550.4]
  assign _T_778 = $signed(_T_777); // @[Math.scala 406:56:@33551.4]
  assign _T_783 = x894_number[31]; // @[FixedPoint.scala 50:25:@33557.4]
  assign _T_787 = _T_783 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@33559.4]
  assign _T_788 = x894_number[31:2]; // @[FixedPoint.scala 18:52:@33560.4]
  assign _T_823 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@33630.4 package.scala 96:25:@33631.4]
  assign _T_825 = io_rr ? _T_823 : 1'h0; // @[implicits.scala 55:10:@33632.4]
  assign _T_826 = _T_367 & _T_825; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 282:194:@33633.4]
  assign x928_x520_D1 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@33589.4 package.scala 96:25:@33590.4]
  assign _T_827 = _T_826 & x928_x520_D1; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 282:282:@33634.4]
  assign x931_b437_D12 = RetimeWrapper_37_io_out; // @[package.scala 96:25:@33616.4 package.scala 96:25:@33617.4]
  assign _T_828 = _T_827 & x931_b437_D12; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 282:290:@33635.4]
  assign x930_b438_D12 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@33607.4 package.scala 96:25:@33608.4]
  assign x932_x468_rdcol_D10_number = RetimeWrapper_39_io_out; // @[package.scala 96:25:@33651.4 package.scala 96:25:@33652.4]
  assign _T_839 = $signed(x932_x468_rdcol_D10_number); // @[Math.scala 465:37:@33657.4]
  assign x529 = $signed(_T_839) < $signed(32'sh0); // @[Math.scala 465:44:@33659.4]
  assign x530 = x517 | x529; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 290:24:@33662.4]
  assign _T_870 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@33706.4 package.scala 96:25:@33707.4]
  assign _T_872 = io_rr ? _T_870 : 1'h0; // @[implicits.scala 55:10:@33708.4]
  assign _T_873 = _T_367 & _T_872; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 309:194:@33709.4]
  assign x934_x531_D1 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@33692.4 package.scala 96:25:@33693.4]
  assign _T_874 = _T_873 & x934_x531_D1; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 309:282:@33710.4]
  assign _T_875 = _T_874 & x931_b437_D12; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 309:325:@33711.4]
  assign x935_x459_rdcol_D10_number = RetimeWrapper_43_io_out; // @[package.scala 96:25:@33727.4 package.scala 96:25:@33728.4]
  assign _T_888 = $signed(x935_x459_rdcol_D10_number); // @[Math.scala 465:37:@33735.4]
  assign x537 = $signed(_T_888) < $signed(32'sh0); // @[Math.scala 465:44:@33737.4]
  assign x538 = x517 | x537; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 319:59:@33740.4]
  assign _T_919 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@33784.4 package.scala 96:25:@33785.4]
  assign _T_921 = io_rr ? _T_919 : 1'h0; // @[implicits.scala 55:10:@33786.4]
  assign _T_922 = _T_367 & _T_921; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 332:194:@33787.4]
  assign x937_x539_D1 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@33770.4 package.scala 96:25:@33771.4]
  assign _T_923 = _T_922 & x937_x539_D1; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 332:282:@33788.4]
  assign _T_924 = _T_923 & x931_b437_D12; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 332:290:@33789.4]
  assign x938_b436_D10_number = RetimeWrapper_47_io_out; // @[package.scala 96:25:@33805.4 package.scala 96:25:@33806.4]
  assign _T_935 = $signed(x938_b436_D10_number); // @[Math.scala 465:37:@33811.4]
  assign x545 = $signed(_T_935) < $signed(32'sh0); // @[Math.scala 465:44:@33813.4]
  assign x939_x545_D1 = RetimeWrapper_48_io_out; // @[package.scala 96:25:@33821.4 package.scala 96:25:@33822.4]
  assign x546 = x517 | x939_x545_D1; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 342:59:@33825.4]
  assign _T_969 = RetimeWrapper_51_io_out; // @[package.scala 96:25:@33869.4 package.scala 96:25:@33870.4]
  assign _T_971 = io_rr ? _T_969 : 1'h0; // @[implicits.scala 55:10:@33871.4]
  assign _T_972 = _T_367 & _T_971; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 355:194:@33872.4]
  assign x941_x547_D1 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@33855.4 package.scala 96:25:@33856.4]
  assign _T_973 = _T_972 & x941_x547_D1; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 355:282:@33873.4]
  assign _T_974 = _T_973 & x931_b437_D12; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 355:290:@33874.4]
  assign x553_rdcol_number = x553_rdcol_1_io_result; // @[Math.scala 154:22:@33893.4 Math.scala 155:14:@33894.4]
  assign _T_989 = $signed(x553_rdcol_number); // @[Math.scala 465:37:@33899.4]
  assign x554 = $signed(_T_989) < $signed(32'sh0); // @[Math.scala 465:44:@33901.4]
  assign x555 = x517 | x554; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 363:59:@33904.4]
  assign _T_999 = x553_rdcol_number[31]; // @[FixedPoint.scala 50:25:@33911.4]
  assign _T_1003 = _T_999 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@33913.4]
  assign _T_1004 = x553_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@33914.4]
  assign _T_1027 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@33948.4 package.scala 96:25:@33949.4]
  assign _T_1029 = io_rr ? _T_1027 : 1'h0; // @[implicits.scala 55:10:@33950.4]
  assign _T_1030 = _T_367 & _T_1029; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 376:194:@33951.4]
  assign x942_x556_D1 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@33934.4 package.scala 96:25:@33935.4]
  assign _T_1031 = _T_1030 & x942_x556_D1; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 376:282:@33952.4]
  assign _T_1032 = _T_1031 & x931_b437_D12; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 376:290:@33953.4]
  assign x565_rdcol_number = x565_rdcol_1_io_result; // @[Math.scala 154:22:@33972.4 Math.scala 155:14:@33973.4]
  assign _T_1047 = $signed(x565_rdcol_number); // @[Math.scala 465:37:@33978.4]
  assign x566 = $signed(_T_1047) < $signed(32'sh0); // @[Math.scala 465:44:@33980.4]
  assign x567 = x517 | x566; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 384:59:@33983.4]
  assign _T_1057 = x565_rdcol_number[31]; // @[FixedPoint.scala 50:25:@33990.4]
  assign _T_1061 = _T_1057 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@33992.4]
  assign _T_1062 = x565_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@33993.4]
  assign _T_1085 = RetimeWrapper_55_io_out; // @[package.scala 96:25:@34027.4 package.scala 96:25:@34028.4]
  assign _T_1087 = io_rr ? _T_1085 : 1'h0; // @[implicits.scala 55:10:@34029.4]
  assign _T_1088 = _T_367 & _T_1087; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 397:194:@34030.4]
  assign x943_x568_D1 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@34013.4 package.scala 96:25:@34014.4]
  assign _T_1089 = _T_1088 & x943_x568_D1; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 397:282:@34031.4]
  assign _T_1090 = _T_1089 & x931_b437_D12; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 397:290:@34032.4]
  assign x944_b435_D10_number = RetimeWrapper_56_io_out; // @[package.scala 96:25:@34048.4 package.scala 96:25:@34049.4]
  assign _T_1103 = $signed(x944_b435_D10_number); // @[Math.scala 406:49:@34055.4]
  assign _T_1105 = $signed(_T_1103) & $signed(32'sh3); // @[Math.scala 406:56:@34057.4]
  assign _T_1106 = $signed(_T_1105); // @[Math.scala 406:56:@34058.4]
  assign x896_number = $unsigned(_T_1106); // @[implicits.scala 133:21:@34059.4]
  assign x578 = $signed(_T_1103) < $signed(32'sh0); // @[Math.scala 465:44:@34067.4]
  assign x945_x578_D1 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@34075.4 package.scala 96:25:@34076.4]
  assign x579 = x945_x578_D1 | x518; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 409:24:@34079.4]
  assign _T_1130 = $signed(x896_number); // @[Math.scala 406:49:@34088.4]
  assign _T_1132 = $signed(_T_1130) & $signed(32'sh3); // @[Math.scala 406:56:@34090.4]
  assign _T_1133 = $signed(_T_1132); // @[Math.scala 406:56:@34091.4]
  assign _T_1138 = x896_number[31]; // @[FixedPoint.scala 50:25:@34097.4]
  assign _T_1142 = _T_1138 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@34099.4]
  assign _T_1143 = x896_number[31:2]; // @[FixedPoint.scala 18:52:@34100.4]
  assign _T_1172 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@34152.4 package.scala 96:25:@34153.4]
  assign _T_1174 = io_rr ? _T_1172 : 1'h0; // @[implicits.scala 55:10:@34154.4]
  assign _T_1175 = _T_367 & _T_1174; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 434:194:@34155.4]
  assign x947_x580_D1 = RetimeWrapper_59_io_out; // @[package.scala 96:25:@34129.4 package.scala 96:25:@34130.4]
  assign _T_1176 = _T_1175 & x947_x580_D1; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 434:282:@34156.4]
  assign _T_1177 = _T_1176 & x931_b437_D12; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 434:290:@34157.4]
  assign x589 = x945_x578_D1 | x529; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 438:59:@34168.4]
  assign _T_1207 = RetimeWrapper_63_io_out; // @[package.scala 96:25:@34205.4 package.scala 96:25:@34206.4]
  assign _T_1209 = io_rr ? _T_1207 : 1'h0; // @[implicits.scala 55:10:@34207.4]
  assign _T_1210 = _T_367 & _T_1209; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 451:194:@34208.4]
  assign x949_x590_D1 = RetimeWrapper_62_io_out; // @[package.scala 96:25:@34191.4 package.scala 96:25:@34192.4]
  assign _T_1211 = _T_1210 & x949_x590_D1; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 451:282:@34209.4]
  assign _T_1212 = _T_1211 & x931_b437_D12; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 451:290:@34210.4]
  assign x596 = x945_x578_D1 | x537; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 455:59:@34221.4]
  assign _T_1240 = RetimeWrapper_65_io_out; // @[package.scala 96:25:@34256.4 package.scala 96:25:@34257.4]
  assign _T_1242 = io_rr ? _T_1240 : 1'h0; // @[implicits.scala 55:10:@34258.4]
  assign _T_1243 = _T_367 & _T_1242; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 466:194:@34259.4]
  assign x950_x597_D1 = RetimeWrapper_64_io_out; // @[package.scala 96:25:@34242.4 package.scala 96:25:@34243.4]
  assign _T_1244 = _T_1243 & x950_x597_D1; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 466:282:@34260.4]
  assign _T_1245 = _T_1244 & x931_b437_D12; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 466:290:@34261.4]
  assign x603 = x578 | x545; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 470:59:@34272.4]
  assign _T_1279 = RetimeWrapper_69_io_out; // @[package.scala 96:25:@34325.4 package.scala 96:25:@34326.4]
  assign _T_1281 = io_rr ? _T_1279 : 1'h0; // @[implicits.scala 55:10:@34327.4]
  assign _T_1282 = _T_367 & _T_1281; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 485:194:@34328.4]
  assign x953_x604_D2 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@34311.4 package.scala 96:25:@34312.4]
  assign _T_1283 = _T_1282 & x953_x604_D2; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 485:282:@34329.4]
  assign _T_1284 = _T_1283 & x931_b437_D12; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 485:290:@34330.4]
  assign x610 = x945_x578_D1 | x554; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 489:59:@34341.4]
  assign _T_1312 = RetimeWrapper_71_io_out; // @[package.scala 96:25:@34376.4 package.scala 96:25:@34377.4]
  assign _T_1314 = io_rr ? _T_1312 : 1'h0; // @[implicits.scala 55:10:@34378.4]
  assign _T_1315 = _T_367 & _T_1314; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 500:194:@34379.4]
  assign x954_x611_D1 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@34362.4 package.scala 96:25:@34363.4]
  assign _T_1316 = _T_1315 & x954_x611_D1; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 500:282:@34380.4]
  assign _T_1317 = _T_1316 & x931_b437_D12; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 500:290:@34381.4]
  assign x617 = x945_x578_D1 | x566; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 504:59:@34392.4]
  assign _T_1345 = RetimeWrapper_73_io_out; // @[package.scala 96:25:@34427.4 package.scala 96:25:@34428.4]
  assign _T_1347 = io_rr ? _T_1345 : 1'h0; // @[implicits.scala 55:10:@34429.4]
  assign _T_1348 = _T_367 & _T_1347; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 515:194:@34430.4]
  assign x955_x618_D1 = RetimeWrapper_72_io_out; // @[package.scala 96:25:@34413.4 package.scala 96:25:@34414.4]
  assign _T_1349 = _T_1348 & x955_x618_D1; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 515:282:@34431.4]
  assign _T_1350 = _T_1349 & x931_b437_D12; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 515:290:@34432.4]
  assign x624_rdrow_number = x624_rdrow_1_io_result; // @[Math.scala 154:22:@34451.4 Math.scala 155:14:@34452.4]
  assign _T_1367 = $signed(x624_rdrow_number); // @[Math.scala 406:49:@34458.4]
  assign _T_1369 = $signed(_T_1367) & $signed(32'sh3); // @[Math.scala 406:56:@34460.4]
  assign _T_1370 = $signed(_T_1369); // @[Math.scala 406:56:@34461.4]
  assign x898_number = $unsigned(_T_1370); // @[implicits.scala 133:21:@34462.4]
  assign x626 = $signed(_T_1367) < $signed(32'sh0); // @[Math.scala 465:44:@34470.4]
  assign x627 = x626 | x518; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 525:24:@34473.4]
  assign _T_1391 = $signed(x898_number); // @[Math.scala 406:49:@34482.4]
  assign _T_1393 = $signed(_T_1391) & $signed(32'sh3); // @[Math.scala 406:56:@34484.4]
  assign _T_1394 = $signed(_T_1393); // @[Math.scala 406:56:@34485.4]
  assign _T_1399 = x898_number[31]; // @[FixedPoint.scala 50:25:@34491.4]
  assign _T_1403 = _T_1399 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@34493.4]
  assign _T_1404 = x898_number[31:2]; // @[FixedPoint.scala 18:52:@34494.4]
  assign _T_1430 = RetimeWrapper_76_io_out; // @[package.scala 96:25:@34537.4 package.scala 96:25:@34538.4]
  assign _T_1432 = io_rr ? _T_1430 : 1'h0; // @[implicits.scala 55:10:@34539.4]
  assign _T_1433 = _T_367 & _T_1432; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 542:194:@34540.4]
  assign x956_x628_D1 = RetimeWrapper_74_io_out; // @[package.scala 96:25:@34514.4 package.scala 96:25:@34515.4]
  assign _T_1434 = _T_1433 & x956_x628_D1; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 542:282:@34541.4]
  assign _T_1435 = _T_1434 & x931_b437_D12; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 542:290:@34542.4]
  assign x637 = x626 | x529; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 546:24:@34553.4]
  assign _T_1465 = RetimeWrapper_78_io_out; // @[package.scala 96:25:@34590.4 package.scala 96:25:@34591.4]
  assign _T_1467 = io_rr ? _T_1465 : 1'h0; // @[implicits.scala 55:10:@34592.4]
  assign _T_1468 = _T_367 & _T_1467; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 565:194:@34593.4]
  assign x958_x638_D1 = RetimeWrapper_77_io_out; // @[package.scala 96:25:@34576.4 package.scala 96:25:@34577.4]
  assign _T_1469 = _T_1468 & x958_x638_D1; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 565:282:@34594.4]
  assign _T_1470 = _T_1469 & x931_b437_D12; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 565:290:@34595.4]
  assign x644 = x626 | x537; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 569:59:@34606.4]
  assign _T_1498 = RetimeWrapper_80_io_out; // @[package.scala 96:25:@34641.4 package.scala 96:25:@34642.4]
  assign _T_1500 = io_rr ? _T_1498 : 1'h0; // @[implicits.scala 55:10:@34643.4]
  assign _T_1501 = _T_367 & _T_1500; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 580:194:@34644.4]
  assign x959_x645_D1 = RetimeWrapper_79_io_out; // @[package.scala 96:25:@34627.4 package.scala 96:25:@34628.4]
  assign _T_1502 = _T_1501 & x959_x645_D1; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 580:282:@34645.4]
  assign _T_1503 = _T_1502 & x931_b437_D12; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 580:290:@34646.4]
  assign x651 = x626 | x939_x545_D1; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 584:59:@34657.4]
  assign _T_1531 = RetimeWrapper_82_io_out; // @[package.scala 96:25:@34692.4 package.scala 96:25:@34693.4]
  assign _T_1533 = io_rr ? _T_1531 : 1'h0; // @[implicits.scala 55:10:@34694.4]
  assign _T_1534 = _T_367 & _T_1533; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 595:194:@34695.4]
  assign x960_x652_D1 = RetimeWrapper_81_io_out; // @[package.scala 96:25:@34678.4 package.scala 96:25:@34679.4]
  assign _T_1535 = _T_1534 & x960_x652_D1; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 595:282:@34696.4]
  assign _T_1536 = _T_1535 & x931_b437_D12; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 595:290:@34697.4]
  assign x658 = x626 | x554; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 599:59:@34708.4]
  assign _T_1564 = RetimeWrapper_84_io_out; // @[package.scala 96:25:@34743.4 package.scala 96:25:@34744.4]
  assign _T_1566 = io_rr ? _T_1564 : 1'h0; // @[implicits.scala 55:10:@34745.4]
  assign _T_1567 = _T_367 & _T_1566; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 610:194:@34746.4]
  assign x961_x659_D1 = RetimeWrapper_83_io_out; // @[package.scala 96:25:@34729.4 package.scala 96:25:@34730.4]
  assign _T_1568 = _T_1567 & x961_x659_D1; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 610:282:@34747.4]
  assign _T_1569 = _T_1568 & x931_b437_D12; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 610:290:@34748.4]
  assign x665 = x626 | x566; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 614:59:@34759.4]
  assign _T_1597 = RetimeWrapper_86_io_out; // @[package.scala 96:25:@34794.4 package.scala 96:25:@34795.4]
  assign _T_1599 = io_rr ? _T_1597 : 1'h0; // @[implicits.scala 55:10:@34796.4]
  assign _T_1600 = _T_367 & _T_1599; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 625:194:@34797.4]
  assign x962_x666_D1 = RetimeWrapper_85_io_out; // @[package.scala 96:25:@34780.4 package.scala 96:25:@34781.4]
  assign _T_1601 = _T_1600 & x962_x666_D1; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 625:282:@34798.4]
  assign _T_1602 = _T_1601 & x931_b437_D12; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 625:290:@34799.4]
  assign x672_rdrow_number = x672_rdrow_1_io_result; // @[Math.scala 154:22:@34818.4 Math.scala 155:14:@34819.4]
  assign _T_1619 = $signed(x672_rdrow_number); // @[Math.scala 406:49:@34825.4]
  assign _T_1621 = $signed(_T_1619) & $signed(32'sh3); // @[Math.scala 406:56:@34827.4]
  assign _T_1622 = $signed(_T_1621); // @[Math.scala 406:56:@34828.4]
  assign x900_number = $unsigned(_T_1622); // @[implicits.scala 133:21:@34829.4]
  assign x674 = $signed(_T_1619) < $signed(32'sh0); // @[Math.scala 465:44:@34837.4]
  assign x675 = x674 | x518; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 635:24:@34840.4]
  assign _T_1643 = $signed(x900_number); // @[Math.scala 406:49:@34849.4]
  assign _T_1645 = $signed(_T_1643) & $signed(32'sh3); // @[Math.scala 406:56:@34851.4]
  assign _T_1646 = $signed(_T_1645); // @[Math.scala 406:56:@34852.4]
  assign _T_1651 = x900_number[31]; // @[FixedPoint.scala 50:25:@34858.4]
  assign _T_1655 = _T_1651 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@34860.4]
  assign _T_1656 = x900_number[31:2]; // @[FixedPoint.scala 18:52:@34861.4]
  assign _T_1682 = RetimeWrapper_89_io_out; // @[package.scala 96:25:@34904.4 package.scala 96:25:@34905.4]
  assign _T_1684 = io_rr ? _T_1682 : 1'h0; // @[implicits.scala 55:10:@34906.4]
  assign _T_1685 = _T_367 & _T_1684; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 652:194:@34907.4]
  assign x964_x676_D1 = RetimeWrapper_88_io_out; // @[package.scala 96:25:@34890.4 package.scala 96:25:@34891.4]
  assign _T_1686 = _T_1685 & x964_x676_D1; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 652:282:@34908.4]
  assign _T_1687 = _T_1686 & x931_b437_D12; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 652:290:@34909.4]
  assign x685 = x674 | x529; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 656:24:@34920.4]
  assign _T_1715 = RetimeWrapper_91_io_out; // @[package.scala 96:25:@34955.4 package.scala 96:25:@34956.4]
  assign _T_1717 = io_rr ? _T_1715 : 1'h0; // @[implicits.scala 55:10:@34957.4]
  assign _T_1718 = _T_367 & _T_1717; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 667:194:@34958.4]
  assign x965_x686_D1 = RetimeWrapper_90_io_out; // @[package.scala 96:25:@34941.4 package.scala 96:25:@34942.4]
  assign _T_1719 = _T_1718 & x965_x686_D1; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 667:282:@34959.4]
  assign _T_1720 = _T_1719 & x931_b437_D12; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 667:290:@34960.4]
  assign x692 = x674 | x537; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 671:24:@34971.4]
  assign _T_1750 = RetimeWrapper_93_io_out; // @[package.scala 96:25:@35008.4 package.scala 96:25:@35009.4]
  assign _T_1752 = io_rr ? _T_1750 : 1'h0; // @[implicits.scala 55:10:@35010.4]
  assign _T_1753 = _T_367 & _T_1752; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 690:194:@35011.4]
  assign x966_x693_D1 = RetimeWrapper_92_io_out; // @[package.scala 96:25:@34994.4 package.scala 96:25:@34995.4]
  assign _T_1754 = _T_1753 & x966_x693_D1; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 690:282:@35012.4]
  assign _T_1755 = _T_1754 & x931_b437_D12; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 690:290:@35013.4]
  assign x699 = x674 | x939_x545_D1; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 694:59:@35024.4]
  assign _T_1783 = RetimeWrapper_95_io_out; // @[package.scala 96:25:@35059.4 package.scala 96:25:@35060.4]
  assign _T_1785 = io_rr ? _T_1783 : 1'h0; // @[implicits.scala 55:10:@35061.4]
  assign _T_1786 = _T_367 & _T_1785; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 705:194:@35062.4]
  assign x967_x700_D1 = RetimeWrapper_94_io_out; // @[package.scala 96:25:@35045.4 package.scala 96:25:@35046.4]
  assign _T_1787 = _T_1786 & x967_x700_D1; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 705:282:@35063.4]
  assign _T_1788 = _T_1787 & x931_b437_D12; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 705:290:@35064.4]
  assign x706 = x674 | x554; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 709:59:@35075.4]
  assign _T_1816 = RetimeWrapper_97_io_out; // @[package.scala 96:25:@35110.4 package.scala 96:25:@35111.4]
  assign _T_1818 = io_rr ? _T_1816 : 1'h0; // @[implicits.scala 55:10:@35112.4]
  assign _T_1819 = _T_367 & _T_1818; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 720:194:@35113.4]
  assign x968_x707_D1 = RetimeWrapper_96_io_out; // @[package.scala 96:25:@35096.4 package.scala 96:25:@35097.4]
  assign _T_1820 = _T_1819 & x968_x707_D1; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 720:282:@35114.4]
  assign _T_1821 = _T_1820 & x931_b437_D12; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 720:290:@35115.4]
  assign x713 = x674 | x566; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 724:59:@35126.4]
  assign _T_1849 = RetimeWrapper_99_io_out; // @[package.scala 96:25:@35161.4 package.scala 96:25:@35162.4]
  assign _T_1851 = io_rr ? _T_1849 : 1'h0; // @[implicits.scala 55:10:@35163.4]
  assign _T_1852 = _T_367 & _T_1851; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 735:194:@35164.4]
  assign x969_x714_D1 = RetimeWrapper_98_io_out; // @[package.scala 96:25:@35147.4 package.scala 96:25:@35148.4]
  assign _T_1853 = _T_1852 & x969_x714_D1; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 735:282:@35165.4]
  assign _T_1854 = _T_1853 & x931_b437_D12; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 735:290:@35166.4]
  assign x535_rd_0_number = x439_lb_0_io_rPort_14_output_0; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 305:29:@33695.4 sm_x824_inr_Foreach_SAMPLER_BOX.scala 309:442:@33718.4]
  assign _GEN_0 = {{1'd0}, x535_rd_0_number}; // @[Math.scala 450:32:@35178.4]
  assign _T_1860 = _GEN_0 << 1; // @[Math.scala 450:32:@35178.4]
  assign x587_rd_0_number = x439_lb_0_io_rPort_2_output_0; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 430:29:@34141.4 sm_x824_inr_Foreach_SAMPLER_BOX.scala 434:407:@34164.4]
  assign _GEN_1 = {{1'd0}, x587_rd_0_number}; // @[Math.scala 450:32:@35183.4]
  assign _T_1864 = _GEN_1 << 1; // @[Math.scala 450:32:@35183.4]
  assign x594_rd_0_number = x439_lb_0_io_rPort_15_output_0; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 447:29:@34194.4 sm_x824_inr_Foreach_SAMPLER_BOX.scala 451:407:@34217.4]
  assign _GEN_2 = {{2'd0}, x594_rd_0_number}; // @[Math.scala 450:32:@35188.4]
  assign _T_1868 = _GEN_2 << 2; // @[Math.scala 450:32:@35188.4]
  assign x601_rd_0_number = x439_lb_0_io_rPort_10_output_0; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 462:29:@34245.4 sm_x824_inr_Foreach_SAMPLER_BOX.scala 466:407:@34268.4]
  assign _GEN_3 = {{1'd0}, x601_rd_0_number}; // @[Math.scala 450:32:@35193.4]
  assign _T_1872 = _GEN_3 << 1; // @[Math.scala 450:32:@35193.4]
  assign x642_rd_0_number = x439_lb_0_io_rPort_7_output_0; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 561:29:@34579.4 sm_x824_inr_Foreach_SAMPLER_BOX.scala 565:407:@34602.4]
  assign _GEN_4 = {{1'd0}, x642_rd_0_number}; // @[Math.scala 450:32:@35198.4]
  assign _T_1876 = _GEN_4 << 1; // @[Math.scala 450:32:@35198.4]
  assign x732_sum_number = x732_sum_1_io_result; // @[Math.scala 154:22:@35287.4 Math.scala 155:14:@35288.4]
  assign _T_1912 = x732_sum_number[7:4]; // @[FixedPoint.scala 18:52:@35293.4]
  assign x543_rd_0_number = x439_lb_0_io_rPort_23_output_0; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 328:29:@33773.4 sm_x824_inr_Foreach_SAMPLER_BOX.scala 332:407:@33796.4]
  assign _GEN_5 = {{1'd0}, x543_rd_0_number}; // @[Math.scala 450:32:@35306.4]
  assign _T_1919 = _GEN_5 << 1; // @[Math.scala 450:32:@35306.4]
  assign _GEN_6 = {{1'd0}, x594_rd_0_number}; // @[Math.scala 450:32:@35311.4]
  assign _T_1923 = _GEN_6 << 1; // @[Math.scala 450:32:@35311.4]
  assign _GEN_7 = {{2'd0}, x601_rd_0_number}; // @[Math.scala 450:32:@35316.4]
  assign _T_1927 = _GEN_7 << 2; // @[Math.scala 450:32:@35316.4]
  assign x608_rd_0_number = x439_lb_0_io_rPort_16_output_0; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 481:29:@34314.4 sm_x824_inr_Foreach_SAMPLER_BOX.scala 485:407:@34337.4]
  assign _GEN_8 = {{1'd0}, x608_rd_0_number}; // @[Math.scala 450:32:@35321.4]
  assign _T_1931 = _GEN_8 << 1; // @[Math.scala 450:32:@35321.4]
  assign x649_rd_0_number = x439_lb_0_io_rPort_13_output_0; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 576:29:@34630.4 sm_x824_inr_Foreach_SAMPLER_BOX.scala 580:407:@34653.4]
  assign _GEN_9 = {{1'd0}, x649_rd_0_number}; // @[Math.scala 450:32:@35326.4]
  assign _T_1935 = _GEN_9 << 1; // @[Math.scala 450:32:@35326.4]
  assign x746_sum_number = x746_sum_1_io_result; // @[Math.scala 154:22:@35417.4 Math.scala 155:14:@35418.4]
  assign _T_1973 = x746_sum_number[7:4]; // @[FixedPoint.scala 18:52:@35423.4]
  assign x551_rd_0_number = x439_lb_0_io_rPort_4_output_0; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 351:29:@33858.4 sm_x824_inr_Foreach_SAMPLER_BOX.scala 355:407:@33881.4]
  assign _GEN_10 = {{1'd0}, x551_rd_0_number}; // @[Math.scala 450:32:@35436.4]
  assign _T_1980 = _GEN_10 << 1; // @[Math.scala 450:32:@35436.4]
  assign _GEN_11 = {{2'd0}, x608_rd_0_number}; // @[Math.scala 450:32:@35441.4]
  assign _T_1984 = _GEN_11 << 2; // @[Math.scala 450:32:@35441.4]
  assign x615_rd_0_number = x439_lb_0_io_rPort_6_output_0; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 496:29:@34365.4 sm_x824_inr_Foreach_SAMPLER_BOX.scala 500:407:@34388.4]
  assign _GEN_12 = {{1'd0}, x615_rd_0_number}; // @[Math.scala 450:32:@35446.4]
  assign _T_1988 = _GEN_12 << 1; // @[Math.scala 450:32:@35446.4]
  assign x656_rd_0_number = x439_lb_0_io_rPort_20_output_0; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 591:29:@34681.4 sm_x824_inr_Foreach_SAMPLER_BOX.scala 595:407:@34704.4]
  assign _GEN_13 = {{1'd0}, x656_rd_0_number}; // @[Math.scala 450:32:@35451.4]
  assign _T_1992 = _GEN_13 << 1; // @[Math.scala 450:32:@35451.4]
  assign x759_sum_number = x759_sum_1_io_result; // @[Math.scala 154:22:@35540.4 Math.scala 155:14:@35541.4]
  assign _T_2028 = x759_sum_number[7:4]; // @[FixedPoint.scala 18:52:@35546.4]
  assign x563_rd_0_number = x439_lb_0_io_rPort_17_output_0; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 372:29:@33937.4 sm_x824_inr_Foreach_SAMPLER_BOX.scala 376:407:@33960.4]
  assign _GEN_14 = {{1'd0}, x563_rd_0_number}; // @[Math.scala 450:32:@35559.4]
  assign _T_2035 = _GEN_14 << 1; // @[Math.scala 450:32:@35559.4]
  assign _GEN_15 = {{2'd0}, x615_rd_0_number}; // @[Math.scala 450:32:@35564.4]
  assign _T_2039 = _GEN_15 << 2; // @[Math.scala 450:32:@35564.4]
  assign x622_rd_0_number = x439_lb_0_io_rPort_8_output_0; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 511:29:@34416.4 sm_x824_inr_Foreach_SAMPLER_BOX.scala 515:407:@34439.4]
  assign _GEN_16 = {{1'd0}, x622_rd_0_number}; // @[Math.scala 450:32:@35569.4]
  assign _T_2043 = _GEN_16 << 1; // @[Math.scala 450:32:@35569.4]
  assign x663_rd_0_number = x439_lb_0_io_rPort_18_output_0; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 606:29:@34732.4 sm_x824_inr_Foreach_SAMPLER_BOX.scala 610:407:@34755.4]
  assign _GEN_17 = {{1'd0}, x663_rd_0_number}; // @[Math.scala 450:32:@35574.4]
  assign _T_2047 = _GEN_17 << 1; // @[Math.scala 450:32:@35574.4]
  assign x772_sum_number = x772_sum_1_io_result; // @[Math.scala 154:22:@35663.4 Math.scala 155:14:@35664.4]
  assign _T_2083 = x772_sum_number[7:4]; // @[FixedPoint.scala 18:52:@35669.4]
  assign x635_rd_0_number = x439_lb_0_io_rPort_21_output_0; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 538:29:@34526.4 sm_x824_inr_Foreach_SAMPLER_BOX.scala 542:407:@34549.4]
  assign _GEN_18 = {{1'd0}, x635_rd_0_number}; // @[Math.scala 450:32:@35682.4]
  assign _T_2090 = _GEN_18 << 1; // @[Math.scala 450:32:@35682.4]
  assign _GEN_19 = {{2'd0}, x642_rd_0_number}; // @[Math.scala 450:32:@35687.4]
  assign _T_2094 = _GEN_19 << 2; // @[Math.scala 450:32:@35687.4]
  assign x690_rd_0_number = x439_lb_0_io_rPort_19_output_0; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 663:29:@34944.4 sm_x824_inr_Foreach_SAMPLER_BOX.scala 667:407:@34967.4]
  assign _GEN_20 = {{1'd0}, x690_rd_0_number}; // @[Math.scala 450:32:@35692.4]
  assign _T_2098 = _GEN_20 << 1; // @[Math.scala 450:32:@35692.4]
  assign x784_sum_number = x784_sum_1_io_result; // @[Math.scala 154:22:@35781.4 Math.scala 155:14:@35782.4]
  assign _T_2134 = x784_sum_number[7:4]; // @[FixedPoint.scala 18:52:@35787.4]
  assign _GEN_21 = {{2'd0}, x649_rd_0_number}; // @[Math.scala 450:32:@35800.4]
  assign _T_2141 = _GEN_21 << 2; // @[Math.scala 450:32:@35800.4]
  assign x697_rd_0_number = x439_lb_0_io_rPort_5_output_0; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 686:29:@34997.4 sm_x824_inr_Foreach_SAMPLER_BOX.scala 690:407:@35020.4]
  assign _GEN_22 = {{1'd0}, x697_rd_0_number}; // @[Math.scala 450:32:@35805.4]
  assign _T_2145 = _GEN_22 << 1; // @[Math.scala 450:32:@35805.4]
  assign x795_sum_number = x795_sum_1_io_result; // @[Math.scala 154:22:@35896.4 Math.scala 155:14:@35897.4]
  assign _T_2183 = x795_sum_number[7:4]; // @[FixedPoint.scala 18:52:@35902.4]
  assign _GEN_23 = {{2'd0}, x656_rd_0_number}; // @[Math.scala 450:32:@35915.4]
  assign _T_2190 = _GEN_23 << 2; // @[Math.scala 450:32:@35915.4]
  assign x704_rd_0_number = x439_lb_0_io_rPort_12_output_0; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 701:29:@35048.4 sm_x824_inr_Foreach_SAMPLER_BOX.scala 705:407:@35071.4]
  assign _GEN_24 = {{1'd0}, x704_rd_0_number}; // @[Math.scala 450:32:@35920.4]
  assign _T_2194 = _GEN_24 << 1; // @[Math.scala 450:32:@35920.4]
  assign x806_sum_number = x806_sum_1_io_result; // @[Math.scala 154:22:@36009.4 Math.scala 155:14:@36010.4]
  assign _T_2230 = x806_sum_number[7:4]; // @[FixedPoint.scala 18:52:@36015.4]
  assign _GEN_25 = {{2'd0}, x663_rd_0_number}; // @[Math.scala 450:32:@36028.4]
  assign _T_2237 = _GEN_25 << 2; // @[Math.scala 450:32:@36028.4]
  assign x670_rd_0_number = x439_lb_0_io_rPort_1_output_0; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 621:29:@34783.4 sm_x824_inr_Foreach_SAMPLER_BOX.scala 625:407:@34806.4]
  assign _GEN_26 = {{1'd0}, x670_rd_0_number}; // @[Math.scala 450:32:@36033.4]
  assign _T_2241 = _GEN_26 << 1; // @[Math.scala 450:32:@36033.4]
  assign x711_rd_0_number = x439_lb_0_io_rPort_11_output_0; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 716:29:@35099.4 sm_x824_inr_Foreach_SAMPLER_BOX.scala 720:407:@35122.4]
  assign _GEN_27 = {{1'd0}, x711_rd_0_number}; // @[Math.scala 450:32:@36038.4]
  assign _T_2245 = _GEN_27 << 1; // @[Math.scala 450:32:@36038.4]
  assign x818_sum_number = x818_sum_1_io_result; // @[Math.scala 154:22:@36127.4 Math.scala 155:14:@36128.4]
  assign _T_2281 = x818_sum_number[7:4]; // @[FixedPoint.scala 18:52:@36133.4]
  assign x807_number = RetimeWrapper_113_io_out; // @[package.scala 96:25:@36022.4 package.scala 96:25:@36023.4]
  assign x819_number = RetimeWrapper_115_io_out; // @[package.scala 96:25:@36140.4 package.scala 96:25:@36141.4]
  assign x785_number = RetimeWrapper_109_io_out; // @[package.scala 96:25:@35794.4 package.scala 96:25:@35795.4]
  assign x796_number = RetimeWrapper_111_io_out; // @[package.scala 96:25:@35909.4 package.scala 96:25:@35910.4]
  assign _T_2302 = {x785_number,x796_number,x807_number,x819_number}; // @[Cat.scala 30:58:@36156.4]
  assign x760_number = RetimeWrapper_105_io_out; // @[package.scala 96:25:@35553.4 package.scala 96:25:@35554.4]
  assign x773_number = RetimeWrapper_107_io_out; // @[package.scala 96:25:@35676.4 package.scala 96:25:@35677.4]
  assign x733_number = RetimeWrapper_101_io_out; // @[package.scala 96:25:@35300.4 package.scala 96:25:@35301.4]
  assign x747_number = RetimeWrapper_103_io_out; // @[package.scala 96:25:@35430.4 package.scala 96:25:@35431.4]
  assign _T_2305 = {x733_number,x747_number,x760_number,x773_number}; // @[Cat.scala 30:58:@36159.4]
  assign _T_2318 = RetimeWrapper_119_io_out; // @[package.scala 96:25:@36195.4 package.scala 96:25:@36196.4]
  assign _T_2320 = io_rr ? _T_2318 : 1'h0; // @[implicits.scala 55:10:@36197.4]
  assign x978_b437_D19 = RetimeWrapper_117_io_out; // @[package.scala 96:25:@36177.4 package.scala 96:25:@36178.4]
  assign _T_2321 = _T_2320 & x978_b437_D19; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 979:116:@36198.4]
  assign x979_b438_D19 = RetimeWrapper_118_io_out; // @[package.scala 96:25:@36186.4 package.scala 96:25:@36187.4]
  assign _T_2322 = _T_2321 & x979_b438_D19; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 979:122:@36199.4]
  assign x903_x892_D8_number = RetimeWrapper_1_io_out; // @[package.scala 96:25:@32875.4 package.scala 96:25:@32876.4]
  assign x905_x453_sum_D7_number = RetimeWrapper_3_io_out; // @[package.scala 96:25:@32893.4 package.scala 96:25:@32894.4]
  assign x910_x463_sum_D6_number = RetimeWrapper_9_io_out; // @[package.scala 96:25:@32996.4 package.scala 96:25:@32997.4]
  assign x911_x472_sum_D6_number = RetimeWrapper_11_io_out; // @[package.scala 96:25:@33063.4 package.scala 96:25:@33064.4]
  assign x913_x481_sum_D6_number = RetimeWrapper_14_io_out; // @[package.scala 96:25:@33139.4 package.scala 96:25:@33140.4]
  assign x916_x893_D7_number = RetimeWrapper_18_io_out; // @[package.scala 96:25:@33284.4 package.scala 96:25:@33285.4]
  assign x918_x495_sum_D6_number = RetimeWrapper_20_io_out; // @[package.scala 96:25:@33302.4 package.scala 96:25:@33303.4]
  assign x920_x501_sum_D6_number = RetimeWrapper_23_io_out; // @[package.scala 96:25:@33357.4 package.scala 96:25:@33358.4]
  assign x922_x506_sum_D6_number = RetimeWrapper_26_io_out; // @[package.scala 96:25:@33412.4 package.scala 96:25:@33413.4]
  assign x923_x511_sum_D6_number = RetimeWrapper_28_io_out; // @[package.scala 96:25:@33458.4 package.scala 96:25:@33459.4]
  assign x523_sum_number = x523_sum_1_io_result; // @[Math.scala 154:22:@33580.4 Math.scala 155:14:@33581.4]
  assign x929_x895_D1_number = RetimeWrapper_35_io_out; // @[package.scala 96:25:@33598.4 package.scala 96:25:@33599.4]
  assign x532_sum_number = x532_sum_1_io_result; // @[Math.scala 154:22:@33683.4 Math.scala 155:14:@33684.4]
  assign x540_sum_number = x540_sum_1_io_result; // @[Math.scala 154:22:@33761.4 Math.scala 155:14:@33762.4]
  assign x548_sum_number = x548_sum_1_io_result; // @[Math.scala 154:22:@33846.4 Math.scala 155:14:@33847.4]
  assign x559_sum_number = x559_sum_1_io_result; // @[Math.scala 154:22:@33925.4 Math.scala 155:14:@33926.4]
  assign x571_sum_number = x571_sum_1_io_result; // @[Math.scala 154:22:@34004.4 Math.scala 155:14:@34005.4]
  assign x583_sum_number = x583_sum_1_io_result; // @[Math.scala 154:22:@34120.4 Math.scala 155:14:@34121.4]
  assign x948_x897_D2_number = RetimeWrapper_60_io_out; // @[package.scala 96:25:@34138.4 package.scala 96:25:@34139.4]
  assign x591_sum_number = x591_sum_1_io_result; // @[Math.scala 154:22:@34182.4 Math.scala 155:14:@34183.4]
  assign x598_sum_number = x598_sum_1_io_result; // @[Math.scala 154:22:@34233.4 Math.scala 155:14:@34234.4]
  assign x952_x605_sum_D1_number = RetimeWrapper_67_io_out; // @[package.scala 96:25:@34302.4 package.scala 96:25:@34303.4]
  assign x612_sum_number = x612_sum_1_io_result; // @[Math.scala 154:22:@34353.4 Math.scala 155:14:@34354.4]
  assign x619_sum_number = x619_sum_1_io_result; // @[Math.scala 154:22:@34404.4 Math.scala 155:14:@34405.4]
  assign x631_sum_number = x631_sum_1_io_result; // @[Math.scala 154:22:@34505.4 Math.scala 155:14:@34506.4]
  assign x957_x899_D1_number = RetimeWrapper_75_io_out; // @[package.scala 96:25:@34523.4 package.scala 96:25:@34524.4]
  assign x639_sum_number = x639_sum_1_io_result; // @[Math.scala 154:22:@34567.4 Math.scala 155:14:@34568.4]
  assign x646_sum_number = x646_sum_1_io_result; // @[Math.scala 154:22:@34618.4 Math.scala 155:14:@34619.4]
  assign x653_sum_number = x653_sum_1_io_result; // @[Math.scala 154:22:@34669.4 Math.scala 155:14:@34670.4]
  assign x660_sum_number = x660_sum_1_io_result; // @[Math.scala 154:22:@34720.4 Math.scala 155:14:@34721.4]
  assign x667_sum_number = x667_sum_1_io_result; // @[Math.scala 154:22:@34771.4 Math.scala 155:14:@34772.4]
  assign x679_sum_number = x679_sum_1_io_result; // @[Math.scala 154:22:@34872.4 Math.scala 155:14:@34873.4]
  assign x963_x901_D1_number = RetimeWrapper_87_io_out; // @[package.scala 96:25:@34881.4 package.scala 96:25:@34882.4]
  assign x687_sum_number = x687_sum_1_io_result; // @[Math.scala 154:22:@34932.4 Math.scala 155:14:@34933.4]
  assign x694_sum_number = x694_sum_1_io_result; // @[Math.scala 154:22:@34985.4 Math.scala 155:14:@34986.4]
  assign x701_sum_number = x701_sum_1_io_result; // @[Math.scala 154:22:@35036.4 Math.scala 155:14:@35037.4]
  assign x708_sum_number = x708_sum_1_io_result; // @[Math.scala 154:22:@35087.4 Math.scala 155:14:@35088.4]
  assign x715_sum_number = x715_sum_1_io_result; // @[Math.scala 154:22:@35138.4 Math.scala 155:14:@35139.4]
  assign io_in_x426_TREADY = _T_212 & _T_214; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 68:22:@32742.4 sm_x824_inr_Foreach_SAMPLER_BOX.scala 70:22:@32750.4]
  assign io_in_x427_TVALID = _T_2322 & io_sigsIn_backpressure; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 979:22:@36201.4]
  assign io_in_x427_TDATA = {{192'd0}, RetimeWrapper_116_io_out}; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 980:24:@36202.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 710:17:@32507.4]
  assign __1_io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_1); // @[Math.scala 710:17:@32519.4]
  assign x439_lb_0_clock = clock; // @[:@32527.4]
  assign x439_lb_0_reset = reset; // @[:@32528.4]
  assign x439_lb_0_io_rPort_23_banks_0 = x929_x895_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@33791.4]
  assign x439_lb_0_io_rPort_23_ofs_0 = x540_sum_number[0]; // @[MemInterfaceType.scala 107:54:@33793.4]
  assign x439_lb_0_io_rPort_23_en_0 = _T_924 & x930_b438_D12; // @[MemInterfaceType.scala 110:79:@33795.4]
  assign x439_lb_0_io_rPort_23_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@33794.4]
  assign x439_lb_0_io_rPort_22_banks_0 = x929_x895_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@34034.4]
  assign x439_lb_0_io_rPort_22_ofs_0 = x571_sum_number[0]; // @[MemInterfaceType.scala 107:54:@34036.4]
  assign x439_lb_0_io_rPort_22_en_0 = _T_1090 & x930_b438_D12; // @[MemInterfaceType.scala 110:79:@34038.4]
  assign x439_lb_0_io_rPort_22_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34037.4]
  assign x439_lb_0_io_rPort_21_banks_0 = x957_x899_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@34544.4]
  assign x439_lb_0_io_rPort_21_ofs_0 = x631_sum_number[0]; // @[MemInterfaceType.scala 107:54:@34546.4]
  assign x439_lb_0_io_rPort_21_en_0 = _T_1435 & x930_b438_D12; // @[MemInterfaceType.scala 110:79:@34548.4]
  assign x439_lb_0_io_rPort_21_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34547.4]
  assign x439_lb_0_io_rPort_20_banks_0 = x957_x899_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@34699.4]
  assign x439_lb_0_io_rPort_20_ofs_0 = x653_sum_number[0]; // @[MemInterfaceType.scala 107:54:@34701.4]
  assign x439_lb_0_io_rPort_20_en_0 = _T_1536 & x930_b438_D12; // @[MemInterfaceType.scala 110:79:@34703.4]
  assign x439_lb_0_io_rPort_20_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34702.4]
  assign x439_lb_0_io_rPort_19_banks_0 = x963_x901_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@34962.4]
  assign x439_lb_0_io_rPort_19_ofs_0 = x687_sum_number[0]; // @[MemInterfaceType.scala 107:54:@34964.4]
  assign x439_lb_0_io_rPort_19_en_0 = _T_1720 & x930_b438_D12; // @[MemInterfaceType.scala 110:79:@34966.4]
  assign x439_lb_0_io_rPort_19_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34965.4]
  assign x439_lb_0_io_rPort_18_banks_0 = x957_x899_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@34750.4]
  assign x439_lb_0_io_rPort_18_ofs_0 = x660_sum_number[0]; // @[MemInterfaceType.scala 107:54:@34752.4]
  assign x439_lb_0_io_rPort_18_en_0 = _T_1569 & x930_b438_D12; // @[MemInterfaceType.scala 110:79:@34754.4]
  assign x439_lb_0_io_rPort_18_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34753.4]
  assign x439_lb_0_io_rPort_17_banks_0 = x929_x895_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@33955.4]
  assign x439_lb_0_io_rPort_17_ofs_0 = x559_sum_number[0]; // @[MemInterfaceType.scala 107:54:@33957.4]
  assign x439_lb_0_io_rPort_17_en_0 = _T_1032 & x930_b438_D12; // @[MemInterfaceType.scala 110:79:@33959.4]
  assign x439_lb_0_io_rPort_17_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@33958.4]
  assign x439_lb_0_io_rPort_16_banks_0 = x948_x897_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@34332.4]
  assign x439_lb_0_io_rPort_16_ofs_0 = x952_x605_sum_D1_number[0]; // @[MemInterfaceType.scala 107:54:@34334.4]
  assign x439_lb_0_io_rPort_16_en_0 = _T_1284 & x930_b438_D12; // @[MemInterfaceType.scala 110:79:@34336.4]
  assign x439_lb_0_io_rPort_16_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34335.4]
  assign x439_lb_0_io_rPort_15_banks_0 = x948_x897_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@34212.4]
  assign x439_lb_0_io_rPort_15_ofs_0 = x591_sum_number[0]; // @[MemInterfaceType.scala 107:54:@34214.4]
  assign x439_lb_0_io_rPort_15_en_0 = _T_1212 & x930_b438_D12; // @[MemInterfaceType.scala 110:79:@34216.4]
  assign x439_lb_0_io_rPort_15_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34215.4]
  assign x439_lb_0_io_rPort_14_banks_0 = x929_x895_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@33713.4]
  assign x439_lb_0_io_rPort_14_ofs_0 = x532_sum_number[0]; // @[MemInterfaceType.scala 107:54:@33715.4]
  assign x439_lb_0_io_rPort_14_en_0 = _T_875 & x930_b438_D12; // @[MemInterfaceType.scala 110:79:@33717.4]
  assign x439_lb_0_io_rPort_14_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@33716.4]
  assign x439_lb_0_io_rPort_13_banks_0 = x957_x899_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@34648.4]
  assign x439_lb_0_io_rPort_13_ofs_0 = x646_sum_number[0]; // @[MemInterfaceType.scala 107:54:@34650.4]
  assign x439_lb_0_io_rPort_13_en_0 = _T_1503 & x930_b438_D12; // @[MemInterfaceType.scala 110:79:@34652.4]
  assign x439_lb_0_io_rPort_13_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34651.4]
  assign x439_lb_0_io_rPort_12_banks_0 = x963_x901_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@35066.4]
  assign x439_lb_0_io_rPort_12_ofs_0 = x701_sum_number[0]; // @[MemInterfaceType.scala 107:54:@35068.4]
  assign x439_lb_0_io_rPort_12_en_0 = _T_1788 & x930_b438_D12; // @[MemInterfaceType.scala 110:79:@35070.4]
  assign x439_lb_0_io_rPort_12_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@35069.4]
  assign x439_lb_0_io_rPort_11_banks_0 = x963_x901_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@35117.4]
  assign x439_lb_0_io_rPort_11_ofs_0 = x708_sum_number[0]; // @[MemInterfaceType.scala 107:54:@35119.4]
  assign x439_lb_0_io_rPort_11_en_0 = _T_1821 & x930_b438_D12; // @[MemInterfaceType.scala 110:79:@35121.4]
  assign x439_lb_0_io_rPort_11_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@35120.4]
  assign x439_lb_0_io_rPort_10_banks_0 = x948_x897_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@34263.4]
  assign x439_lb_0_io_rPort_10_ofs_0 = x598_sum_number[0]; // @[MemInterfaceType.scala 107:54:@34265.4]
  assign x439_lb_0_io_rPort_10_en_0 = _T_1245 & x930_b438_D12; // @[MemInterfaceType.scala 110:79:@34267.4]
  assign x439_lb_0_io_rPort_10_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34266.4]
  assign x439_lb_0_io_rPort_9_banks_0 = x963_x901_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@35168.4]
  assign x439_lb_0_io_rPort_9_ofs_0 = x715_sum_number[0]; // @[MemInterfaceType.scala 107:54:@35170.4]
  assign x439_lb_0_io_rPort_9_en_0 = _T_1854 & x930_b438_D12; // @[MemInterfaceType.scala 110:79:@35172.4]
  assign x439_lb_0_io_rPort_9_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@35171.4]
  assign x439_lb_0_io_rPort_8_banks_0 = x948_x897_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@34434.4]
  assign x439_lb_0_io_rPort_8_ofs_0 = x619_sum_number[0]; // @[MemInterfaceType.scala 107:54:@34436.4]
  assign x439_lb_0_io_rPort_8_en_0 = _T_1350 & x930_b438_D12; // @[MemInterfaceType.scala 110:79:@34438.4]
  assign x439_lb_0_io_rPort_8_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34437.4]
  assign x439_lb_0_io_rPort_7_banks_0 = x957_x899_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@34597.4]
  assign x439_lb_0_io_rPort_7_ofs_0 = x639_sum_number[0]; // @[MemInterfaceType.scala 107:54:@34599.4]
  assign x439_lb_0_io_rPort_7_en_0 = _T_1470 & x930_b438_D12; // @[MemInterfaceType.scala 110:79:@34601.4]
  assign x439_lb_0_io_rPort_7_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34600.4]
  assign x439_lb_0_io_rPort_6_banks_0 = x948_x897_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@34383.4]
  assign x439_lb_0_io_rPort_6_ofs_0 = x612_sum_number[0]; // @[MemInterfaceType.scala 107:54:@34385.4]
  assign x439_lb_0_io_rPort_6_en_0 = _T_1317 & x930_b438_D12; // @[MemInterfaceType.scala 110:79:@34387.4]
  assign x439_lb_0_io_rPort_6_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34386.4]
  assign x439_lb_0_io_rPort_5_banks_0 = x963_x901_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@35015.4]
  assign x439_lb_0_io_rPort_5_ofs_0 = x694_sum_number[0]; // @[MemInterfaceType.scala 107:54:@35017.4]
  assign x439_lb_0_io_rPort_5_en_0 = _T_1755 & x930_b438_D12; // @[MemInterfaceType.scala 110:79:@35019.4]
  assign x439_lb_0_io_rPort_5_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@35018.4]
  assign x439_lb_0_io_rPort_4_banks_0 = x929_x895_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@33876.4]
  assign x439_lb_0_io_rPort_4_ofs_0 = x548_sum_number[0]; // @[MemInterfaceType.scala 107:54:@33878.4]
  assign x439_lb_0_io_rPort_4_en_0 = _T_974 & x930_b438_D12; // @[MemInterfaceType.scala 110:79:@33880.4]
  assign x439_lb_0_io_rPort_4_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@33879.4]
  assign x439_lb_0_io_rPort_3_banks_0 = x929_x895_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@33637.4]
  assign x439_lb_0_io_rPort_3_ofs_0 = x523_sum_number[0]; // @[MemInterfaceType.scala 107:54:@33639.4]
  assign x439_lb_0_io_rPort_3_en_0 = _T_828 & x930_b438_D12; // @[MemInterfaceType.scala 110:79:@33641.4]
  assign x439_lb_0_io_rPort_3_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@33640.4]
  assign x439_lb_0_io_rPort_2_banks_0 = x948_x897_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@34159.4]
  assign x439_lb_0_io_rPort_2_ofs_0 = x583_sum_number[0]; // @[MemInterfaceType.scala 107:54:@34161.4]
  assign x439_lb_0_io_rPort_2_en_0 = _T_1177 & x930_b438_D12; // @[MemInterfaceType.scala 110:79:@34163.4]
  assign x439_lb_0_io_rPort_2_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34162.4]
  assign x439_lb_0_io_rPort_1_banks_0 = x957_x899_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@34801.4]
  assign x439_lb_0_io_rPort_1_ofs_0 = x667_sum_number[0]; // @[MemInterfaceType.scala 107:54:@34803.4]
  assign x439_lb_0_io_rPort_1_en_0 = _T_1602 & x930_b438_D12; // @[MemInterfaceType.scala 110:79:@34805.4]
  assign x439_lb_0_io_rPort_1_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34804.4]
  assign x439_lb_0_io_rPort_0_banks_0 = x963_x901_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@34911.4]
  assign x439_lb_0_io_rPort_0_ofs_0 = x679_sum_number[0]; // @[MemInterfaceType.scala 107:54:@34913.4]
  assign x439_lb_0_io_rPort_0_en_0 = _T_1687 & x930_b438_D12; // @[MemInterfaceType.scala 110:79:@34915.4]
  assign x439_lb_0_io_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34914.4]
  assign x439_lb_0_io_wPort_7_banks_0 = x903_x892_D8_number[2:0]; // @[MemInterfaceType.scala 88:58:@32933.4]
  assign x439_lb_0_io_wPort_7_ofs_0 = x905_x453_sum_D7_number[0]; // @[MemInterfaceType.scala 89:54:@32935.4]
  assign x439_lb_0_io_wPort_7_data_0 = RetimeWrapper_2_io_out; // @[MemInterfaceType.scala 90:56:@32936.4]
  assign x439_lb_0_io_wPort_7_en_0 = _T_378 & x906_b438_D8; // @[MemInterfaceType.scala 93:57:@32938.4]
  assign x439_lb_0_io_wPort_6_banks_0 = x916_x893_D7_number[2:0]; // @[MemInterfaceType.scala 88:58:@33434.4]
  assign x439_lb_0_io_wPort_6_ofs_0 = x922_x506_sum_D6_number[0]; // @[MemInterfaceType.scala 89:54:@33436.4]
  assign x439_lb_0_io_wPort_6_data_0 = RetimeWrapper_25_io_out; // @[MemInterfaceType.scala 90:56:@33437.4]
  assign x439_lb_0_io_wPort_6_en_0 = _T_700 & x906_b438_D8; // @[MemInterfaceType.scala 93:57:@33439.4]
  assign x439_lb_0_io_wPort_5_banks_0 = x903_x892_D8_number[2:0]; // @[MemInterfaceType.scala 88:58:@33094.4]
  assign x439_lb_0_io_wPort_5_ofs_0 = x911_x472_sum_D6_number[0]; // @[MemInterfaceType.scala 89:54:@33096.4]
  assign x439_lb_0_io_wPort_5_data_0 = RetimeWrapper_12_io_out; // @[MemInterfaceType.scala 90:56:@33097.4]
  assign x439_lb_0_io_wPort_5_en_0 = _T_471 & x906_b438_D8; // @[MemInterfaceType.scala 93:57:@33099.4]
  assign x439_lb_0_io_wPort_4_banks_0 = x916_x893_D7_number[2:0]; // @[MemInterfaceType.scala 88:58:@33324.4]
  assign x439_lb_0_io_wPort_4_ofs_0 = x918_x495_sum_D6_number[0]; // @[MemInterfaceType.scala 89:54:@33326.4]
  assign x439_lb_0_io_wPort_4_data_0 = RetimeWrapper_19_io_out; // @[MemInterfaceType.scala 90:56:@33327.4]
  assign x439_lb_0_io_wPort_4_en_0 = _T_644 & x906_b438_D8; // @[MemInterfaceType.scala 93:57:@33329.4]
  assign x439_lb_0_io_wPort_3_banks_0 = x903_x892_D8_number[2:0]; // @[MemInterfaceType.scala 88:58:@33018.4]
  assign x439_lb_0_io_wPort_3_ofs_0 = x910_x463_sum_D6_number[0]; // @[MemInterfaceType.scala 89:54:@33020.4]
  assign x439_lb_0_io_wPort_3_data_0 = RetimeWrapper_8_io_out; // @[MemInterfaceType.scala 90:56:@33021.4]
  assign x439_lb_0_io_wPort_3_en_0 = _T_426 & x906_b438_D8; // @[MemInterfaceType.scala 93:57:@33023.4]
  assign x439_lb_0_io_wPort_2_banks_0 = x916_x893_D7_number[2:0]; // @[MemInterfaceType.scala 88:58:@33489.4]
  assign x439_lb_0_io_wPort_2_ofs_0 = x923_x511_sum_D6_number[0]; // @[MemInterfaceType.scala 89:54:@33491.4]
  assign x439_lb_0_io_wPort_2_data_0 = RetimeWrapper_29_io_out; // @[MemInterfaceType.scala 90:56:@33492.4]
  assign x439_lb_0_io_wPort_2_en_0 = _T_728 & x906_b438_D8; // @[MemInterfaceType.scala 93:57:@33494.4]
  assign x439_lb_0_io_wPort_1_banks_0 = x903_x892_D8_number[2:0]; // @[MemInterfaceType.scala 88:58:@33170.4]
  assign x439_lb_0_io_wPort_1_ofs_0 = x913_x481_sum_D6_number[0]; // @[MemInterfaceType.scala 89:54:@33172.4]
  assign x439_lb_0_io_wPort_1_data_0 = RetimeWrapper_15_io_out; // @[MemInterfaceType.scala 90:56:@33173.4]
  assign x439_lb_0_io_wPort_1_en_0 = _T_516 & x906_b438_D8; // @[MemInterfaceType.scala 93:57:@33175.4]
  assign x439_lb_0_io_wPort_0_banks_0 = x916_x893_D7_number[2:0]; // @[MemInterfaceType.scala 88:58:@33379.4]
  assign x439_lb_0_io_wPort_0_ofs_0 = x920_x501_sum_D6_number[0]; // @[MemInterfaceType.scala 89:54:@33381.4]
  assign x439_lb_0_io_wPort_0_data_0 = RetimeWrapper_22_io_out; // @[MemInterfaceType.scala 90:56:@33382.4]
  assign x439_lb_0_io_wPort_0_en_0 = _T_672 & x906_b438_D8; // @[MemInterfaceType.scala 93:57:@33384.4]
  assign RetimeWrapper_clock = clock; // @[:@32753.4]
  assign RetimeWrapper_reset = reset; // @[:@32754.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32756.4]
  assign RetimeWrapper_io_in = io_in_x426_TDATA[63:0]; // @[package.scala 94:16:@32755.4]
  assign x453_sum_1_clock = clock; // @[:@32861.4]
  assign x453_sum_1_reset = reset; // @[:@32862.4]
  assign x453_sum_1_io_a = {_T_331,_T_332}; // @[Math.scala 151:17:@32863.4]
  assign x453_sum_1_io_b = {_T_341,_T_342}; // @[Math.scala 152:17:@32864.4]
  assign x453_sum_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@32865.4]
  assign RetimeWrapper_1_clock = clock; // @[:@32871.4]
  assign RetimeWrapper_1_reset = reset; // @[:@32872.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32874.4]
  assign RetimeWrapper_1_io_in = $unsigned(_T_322); // @[package.scala 94:16:@32873.4]
  assign RetimeWrapper_2_clock = clock; // @[:@32880.4]
  assign RetimeWrapper_2_reset = reset; // @[:@32881.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32883.4]
  assign RetimeWrapper_2_io_in = x902_x440_D1_0_number[7:0]; // @[package.scala 94:16:@32882.4]
  assign RetimeWrapper_3_clock = clock; // @[:@32889.4]
  assign RetimeWrapper_3_reset = reset; // @[:@32890.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32892.4]
  assign RetimeWrapper_3_io_in = x453_sum_1_io_result; // @[package.scala 94:16:@32891.4]
  assign RetimeWrapper_4_clock = clock; // @[:@32898.4]
  assign RetimeWrapper_4_reset = reset; // @[:@32899.4]
  assign RetimeWrapper_4_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32901.4]
  assign RetimeWrapper_4_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@32900.4]
  assign RetimeWrapper_5_clock = clock; // @[:@32907.4]
  assign RetimeWrapper_5_reset = reset; // @[:@32908.4]
  assign RetimeWrapper_5_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32910.4]
  assign RetimeWrapper_5_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@32909.4]
  assign RetimeWrapper_6_clock = clock; // @[:@32920.4]
  assign RetimeWrapper_6_reset = reset; // @[:@32921.4]
  assign RetimeWrapper_6_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32923.4]
  assign RetimeWrapper_6_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@32922.4]
  assign x459_rdcol_1_clock = clock; // @[:@32943.4]
  assign x459_rdcol_1_reset = reset; // @[:@32944.4]
  assign x459_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@32945.4]
  assign x459_rdcol_1_io_b = 32'h1; // @[Math.scala 152:17:@32946.4]
  assign x459_rdcol_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@32947.4]
  assign RetimeWrapper_7_clock = clock; // @[:@32964.4]
  assign RetimeWrapper_7_reset = reset; // @[:@32965.4]
  assign RetimeWrapper_7_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32967.4]
  assign RetimeWrapper_7_io_in = {_T_331,_T_332}; // @[package.scala 94:16:@32966.4]
  assign x463_sum_1_clock = clock; // @[:@32973.4]
  assign x463_sum_1_reset = reset; // @[:@32974.4]
  assign x463_sum_1_io_a = RetimeWrapper_7_io_out; // @[Math.scala 151:17:@32975.4]
  assign x463_sum_1_io_b = {_T_395,_T_396}; // @[Math.scala 152:17:@32976.4]
  assign x463_sum_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@32977.4]
  assign RetimeWrapper_8_clock = clock; // @[:@32983.4]
  assign RetimeWrapper_8_reset = reset; // @[:@32984.4]
  assign RetimeWrapper_8_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32986.4]
  assign RetimeWrapper_8_io_in = x902_x440_D1_0_number[15:8]; // @[package.scala 94:16:@32985.4]
  assign RetimeWrapper_9_clock = clock; // @[:@32992.4]
  assign RetimeWrapper_9_reset = reset; // @[:@32993.4]
  assign RetimeWrapper_9_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32995.4]
  assign RetimeWrapper_9_io_in = x463_sum_1_io_result; // @[package.scala 94:16:@32994.4]
  assign RetimeWrapper_10_clock = clock; // @[:@33005.4]
  assign RetimeWrapper_10_reset = reset; // @[:@33006.4]
  assign RetimeWrapper_10_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33008.4]
  assign RetimeWrapper_10_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33007.4]
  assign x468_rdcol_1_clock = clock; // @[:@33028.4]
  assign x468_rdcol_1_reset = reset; // @[:@33029.4]
  assign x468_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@33030.4]
  assign x468_rdcol_1_io_b = 32'h2; // @[Math.scala 152:17:@33031.4]
  assign x468_rdcol_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@33032.4]
  assign x472_sum_1_clock = clock; // @[:@33049.4]
  assign x472_sum_1_reset = reset; // @[:@33050.4]
  assign x472_sum_1_io_a = RetimeWrapper_7_io_out; // @[Math.scala 151:17:@33051.4]
  assign x472_sum_1_io_b = {_T_443,_T_444}; // @[Math.scala 152:17:@33052.4]
  assign x472_sum_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@33053.4]
  assign RetimeWrapper_11_clock = clock; // @[:@33059.4]
  assign RetimeWrapper_11_reset = reset; // @[:@33060.4]
  assign RetimeWrapper_11_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33062.4]
  assign RetimeWrapper_11_io_in = x472_sum_1_io_result; // @[package.scala 94:16:@33061.4]
  assign RetimeWrapper_12_clock = clock; // @[:@33068.4]
  assign RetimeWrapper_12_reset = reset; // @[:@33069.4]
  assign RetimeWrapper_12_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33071.4]
  assign RetimeWrapper_12_io_in = x902_x440_D1_0_number[23:16]; // @[package.scala 94:16:@33070.4]
  assign RetimeWrapper_13_clock = clock; // @[:@33081.4]
  assign RetimeWrapper_13_reset = reset; // @[:@33082.4]
  assign RetimeWrapper_13_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33084.4]
  assign RetimeWrapper_13_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33083.4]
  assign x477_rdcol_1_clock = clock; // @[:@33104.4]
  assign x477_rdcol_1_reset = reset; // @[:@33105.4]
  assign x477_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@33106.4]
  assign x477_rdcol_1_io_b = 32'h3; // @[Math.scala 152:17:@33107.4]
  assign x477_rdcol_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@33108.4]
  assign x481_sum_1_clock = clock; // @[:@33125.4]
  assign x481_sum_1_reset = reset; // @[:@33126.4]
  assign x481_sum_1_io_a = RetimeWrapper_7_io_out; // @[Math.scala 151:17:@33127.4]
  assign x481_sum_1_io_b = {_T_488,_T_489}; // @[Math.scala 152:17:@33128.4]
  assign x481_sum_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@33129.4]
  assign RetimeWrapper_14_clock = clock; // @[:@33135.4]
  assign RetimeWrapper_14_reset = reset; // @[:@33136.4]
  assign RetimeWrapper_14_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33138.4]
  assign RetimeWrapper_14_io_in = x481_sum_1_io_result; // @[package.scala 94:16:@33137.4]
  assign RetimeWrapper_15_clock = clock; // @[:@33144.4]
  assign RetimeWrapper_15_reset = reset; // @[:@33145.4]
  assign RetimeWrapper_15_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33147.4]
  assign RetimeWrapper_15_io_in = x902_x440_D1_0_number[31:24]; // @[package.scala 94:16:@33146.4]
  assign RetimeWrapper_16_clock = clock; // @[:@33157.4]
  assign RetimeWrapper_16_reset = reset; // @[:@33158.4]
  assign RetimeWrapper_16_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33160.4]
  assign RetimeWrapper_16_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33159.4]
  assign x486_rdrow_1_clock = clock; // @[:@33180.4]
  assign x486_rdrow_1_reset = reset; // @[:@33181.4]
  assign x486_rdrow_1_io_a = __io_result; // @[Math.scala 151:17:@33182.4]
  assign x486_rdrow_1_io_b = 32'h1; // @[Math.scala 152:17:@33183.4]
  assign x486_rdrow_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@33184.4]
  assign RetimeWrapper_17_clock = clock; // @[:@33261.4]
  assign RetimeWrapper_17_reset = reset; // @[:@33262.4]
  assign RetimeWrapper_17_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33264.4]
  assign RetimeWrapper_17_io_in = {_T_341,_T_342}; // @[package.scala 94:16:@33263.4]
  assign x495_sum_1_clock = clock; // @[:@33270.4]
  assign x495_sum_1_reset = reset; // @[:@33271.4]
  assign x495_sum_1_io_a = {_T_610,_T_611}; // @[Math.scala 151:17:@33272.4]
  assign x495_sum_1_io_b = RetimeWrapper_17_io_out; // @[Math.scala 152:17:@33273.4]
  assign x495_sum_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@33274.4]
  assign RetimeWrapper_18_clock = clock; // @[:@33280.4]
  assign RetimeWrapper_18_reset = reset; // @[:@33281.4]
  assign RetimeWrapper_18_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33283.4]
  assign RetimeWrapper_18_io_in = $unsigned(_T_601); // @[package.scala 94:16:@33282.4]
  assign RetimeWrapper_19_clock = clock; // @[:@33289.4]
  assign RetimeWrapper_19_reset = reset; // @[:@33290.4]
  assign RetimeWrapper_19_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33292.4]
  assign RetimeWrapper_19_io_in = x902_x440_D1_0_number[39:32]; // @[package.scala 94:16:@33291.4]
  assign RetimeWrapper_20_clock = clock; // @[:@33298.4]
  assign RetimeWrapper_20_reset = reset; // @[:@33299.4]
  assign RetimeWrapper_20_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33301.4]
  assign RetimeWrapper_20_io_in = x495_sum_1_io_result; // @[package.scala 94:16:@33300.4]
  assign RetimeWrapper_21_clock = clock; // @[:@33311.4]
  assign RetimeWrapper_21_reset = reset; // @[:@33312.4]
  assign RetimeWrapper_21_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33314.4]
  assign RetimeWrapper_21_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33313.4]
  assign x501_sum_1_clock = clock; // @[:@33334.4]
  assign x501_sum_1_reset = reset; // @[:@33335.4]
  assign x501_sum_1_io_a = {_T_610,_T_611}; // @[Math.scala 151:17:@33336.4]
  assign x501_sum_1_io_b = {_T_395,_T_396}; // @[Math.scala 152:17:@33337.4]
  assign x501_sum_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@33338.4]
  assign RetimeWrapper_22_clock = clock; // @[:@33344.4]
  assign RetimeWrapper_22_reset = reset; // @[:@33345.4]
  assign RetimeWrapper_22_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33347.4]
  assign RetimeWrapper_22_io_in = x902_x440_D1_0_number[47:40]; // @[package.scala 94:16:@33346.4]
  assign RetimeWrapper_23_clock = clock; // @[:@33353.4]
  assign RetimeWrapper_23_reset = reset; // @[:@33354.4]
  assign RetimeWrapper_23_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33356.4]
  assign RetimeWrapper_23_io_in = x501_sum_1_io_result; // @[package.scala 94:16:@33355.4]
  assign RetimeWrapper_24_clock = clock; // @[:@33366.4]
  assign RetimeWrapper_24_reset = reset; // @[:@33367.4]
  assign RetimeWrapper_24_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33369.4]
  assign RetimeWrapper_24_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33368.4]
  assign x506_sum_1_clock = clock; // @[:@33389.4]
  assign x506_sum_1_reset = reset; // @[:@33390.4]
  assign x506_sum_1_io_a = {_T_610,_T_611}; // @[Math.scala 151:17:@33391.4]
  assign x506_sum_1_io_b = {_T_443,_T_444}; // @[Math.scala 152:17:@33392.4]
  assign x506_sum_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@33393.4]
  assign RetimeWrapper_25_clock = clock; // @[:@33399.4]
  assign RetimeWrapper_25_reset = reset; // @[:@33400.4]
  assign RetimeWrapper_25_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33402.4]
  assign RetimeWrapper_25_io_in = x902_x440_D1_0_number[55:48]; // @[package.scala 94:16:@33401.4]
  assign RetimeWrapper_26_clock = clock; // @[:@33408.4]
  assign RetimeWrapper_26_reset = reset; // @[:@33409.4]
  assign RetimeWrapper_26_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33411.4]
  assign RetimeWrapper_26_io_in = x506_sum_1_io_result; // @[package.scala 94:16:@33410.4]
  assign RetimeWrapper_27_clock = clock; // @[:@33421.4]
  assign RetimeWrapper_27_reset = reset; // @[:@33422.4]
  assign RetimeWrapper_27_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33424.4]
  assign RetimeWrapper_27_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33423.4]
  assign x511_sum_1_clock = clock; // @[:@33444.4]
  assign x511_sum_1_reset = reset; // @[:@33445.4]
  assign x511_sum_1_io_a = {_T_610,_T_611}; // @[Math.scala 151:17:@33446.4]
  assign x511_sum_1_io_b = {_T_488,_T_489}; // @[Math.scala 152:17:@33447.4]
  assign x511_sum_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@33448.4]
  assign RetimeWrapper_28_clock = clock; // @[:@33454.4]
  assign RetimeWrapper_28_reset = reset; // @[:@33455.4]
  assign RetimeWrapper_28_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33457.4]
  assign RetimeWrapper_28_io_in = x511_sum_1_io_result; // @[package.scala 94:16:@33456.4]
  assign RetimeWrapper_29_clock = clock; // @[:@33463.4]
  assign RetimeWrapper_29_reset = reset; // @[:@33464.4]
  assign RetimeWrapper_29_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33466.4]
  assign RetimeWrapper_29_io_in = x902_x440_D1_0_number[63:56]; // @[package.scala 94:16:@33465.4]
  assign RetimeWrapper_30_clock = clock; // @[:@33476.4]
  assign RetimeWrapper_30_reset = reset; // @[:@33477.4]
  assign RetimeWrapper_30_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33479.4]
  assign RetimeWrapper_30_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33478.4]
  assign RetimeWrapper_31_clock = clock; // @[:@33497.4]
  assign RetimeWrapper_31_reset = reset; // @[:@33498.4]
  assign RetimeWrapper_31_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33500.4]
  assign RetimeWrapper_31_io_in = x486_rdrow_1_io_result; // @[package.scala 94:16:@33499.4]
  assign RetimeWrapper_32_clock = clock; // @[:@33524.4]
  assign RetimeWrapper_32_reset = reset; // @[:@33525.4]
  assign RetimeWrapper_32_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33527.4]
  assign RetimeWrapper_32_io_in = x477_rdcol_1_io_result; // @[package.scala 94:16:@33526.4]
  assign RetimeWrapper_33_clock = clock; // @[:@33566.4]
  assign RetimeWrapper_33_reset = reset; // @[:@33567.4]
  assign RetimeWrapper_33_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33569.4]
  assign RetimeWrapper_33_io_in = {_T_488,_T_489}; // @[package.scala 94:16:@33568.4]
  assign x523_sum_1_clock = clock; // @[:@33575.4]
  assign x523_sum_1_reset = reset; // @[:@33576.4]
  assign x523_sum_1_io_a = {_T_787,_T_788}; // @[Math.scala 151:17:@33577.4]
  assign x523_sum_1_io_b = RetimeWrapper_33_io_out; // @[Math.scala 152:17:@33578.4]
  assign x523_sum_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@33579.4]
  assign RetimeWrapper_34_clock = clock; // @[:@33585.4]
  assign RetimeWrapper_34_reset = reset; // @[:@33586.4]
  assign RetimeWrapper_34_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33588.4]
  assign RetimeWrapper_34_io_in = ~ x519; // @[package.scala 94:16:@33587.4]
  assign RetimeWrapper_35_clock = clock; // @[:@33594.4]
  assign RetimeWrapper_35_reset = reset; // @[:@33595.4]
  assign RetimeWrapper_35_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33597.4]
  assign RetimeWrapper_35_io_in = $unsigned(_T_778); // @[package.scala 94:16:@33596.4]
  assign RetimeWrapper_36_clock = clock; // @[:@33603.4]
  assign RetimeWrapper_36_reset = reset; // @[:@33604.4]
  assign RetimeWrapper_36_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33606.4]
  assign RetimeWrapper_36_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@33605.4]
  assign RetimeWrapper_37_clock = clock; // @[:@33612.4]
  assign RetimeWrapper_37_reset = reset; // @[:@33613.4]
  assign RetimeWrapper_37_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33615.4]
  assign RetimeWrapper_37_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@33614.4]
  assign RetimeWrapper_38_clock = clock; // @[:@33626.4]
  assign RetimeWrapper_38_reset = reset; // @[:@33627.4]
  assign RetimeWrapper_38_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33629.4]
  assign RetimeWrapper_38_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33628.4]
  assign RetimeWrapper_39_clock = clock; // @[:@33647.4]
  assign RetimeWrapper_39_reset = reset; // @[:@33648.4]
  assign RetimeWrapper_39_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33650.4]
  assign RetimeWrapper_39_io_in = x468_rdcol_1_io_result; // @[package.scala 94:16:@33649.4]
  assign RetimeWrapper_40_clock = clock; // @[:@33669.4]
  assign RetimeWrapper_40_reset = reset; // @[:@33670.4]
  assign RetimeWrapper_40_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33672.4]
  assign RetimeWrapper_40_io_in = {_T_443,_T_444}; // @[package.scala 94:16:@33671.4]
  assign x532_sum_1_clock = clock; // @[:@33678.4]
  assign x532_sum_1_reset = reset; // @[:@33679.4]
  assign x532_sum_1_io_a = {_T_787,_T_788}; // @[Math.scala 151:17:@33680.4]
  assign x532_sum_1_io_b = RetimeWrapper_40_io_out; // @[Math.scala 152:17:@33681.4]
  assign x532_sum_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@33682.4]
  assign RetimeWrapper_41_clock = clock; // @[:@33688.4]
  assign RetimeWrapper_41_reset = reset; // @[:@33689.4]
  assign RetimeWrapper_41_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33691.4]
  assign RetimeWrapper_41_io_in = ~ x530; // @[package.scala 94:16:@33690.4]
  assign RetimeWrapper_42_clock = clock; // @[:@33702.4]
  assign RetimeWrapper_42_reset = reset; // @[:@33703.4]
  assign RetimeWrapper_42_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33705.4]
  assign RetimeWrapper_42_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33704.4]
  assign RetimeWrapper_43_clock = clock; // @[:@33723.4]
  assign RetimeWrapper_43_reset = reset; // @[:@33724.4]
  assign RetimeWrapper_43_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33726.4]
  assign RetimeWrapper_43_io_in = x459_rdcol_1_io_result; // @[package.scala 94:16:@33725.4]
  assign RetimeWrapper_44_clock = clock; // @[:@33747.4]
  assign RetimeWrapper_44_reset = reset; // @[:@33748.4]
  assign RetimeWrapper_44_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33750.4]
  assign RetimeWrapper_44_io_in = {_T_395,_T_396}; // @[package.scala 94:16:@33749.4]
  assign x540_sum_1_clock = clock; // @[:@33756.4]
  assign x540_sum_1_reset = reset; // @[:@33757.4]
  assign x540_sum_1_io_a = {_T_787,_T_788}; // @[Math.scala 151:17:@33758.4]
  assign x540_sum_1_io_b = RetimeWrapper_44_io_out; // @[Math.scala 152:17:@33759.4]
  assign x540_sum_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@33760.4]
  assign RetimeWrapper_45_clock = clock; // @[:@33766.4]
  assign RetimeWrapper_45_reset = reset; // @[:@33767.4]
  assign RetimeWrapper_45_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33769.4]
  assign RetimeWrapper_45_io_in = ~ x538; // @[package.scala 94:16:@33768.4]
  assign RetimeWrapper_46_clock = clock; // @[:@33780.4]
  assign RetimeWrapper_46_reset = reset; // @[:@33781.4]
  assign RetimeWrapper_46_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33783.4]
  assign RetimeWrapper_46_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33782.4]
  assign RetimeWrapper_47_clock = clock; // @[:@33801.4]
  assign RetimeWrapper_47_reset = reset; // @[:@33802.4]
  assign RetimeWrapper_47_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33804.4]
  assign RetimeWrapper_47_io_in = __1_io_result; // @[package.scala 94:16:@33803.4]
  assign RetimeWrapper_48_clock = clock; // @[:@33817.4]
  assign RetimeWrapper_48_reset = reset; // @[:@33818.4]
  assign RetimeWrapper_48_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33820.4]
  assign RetimeWrapper_48_io_in = $signed(_T_935) < $signed(32'sh0); // @[package.scala 94:16:@33819.4]
  assign RetimeWrapper_49_clock = clock; // @[:@33832.4]
  assign RetimeWrapper_49_reset = reset; // @[:@33833.4]
  assign RetimeWrapper_49_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33835.4]
  assign RetimeWrapper_49_io_in = {_T_341,_T_342}; // @[package.scala 94:16:@33834.4]
  assign x548_sum_1_clock = clock; // @[:@33841.4]
  assign x548_sum_1_reset = reset; // @[:@33842.4]
  assign x548_sum_1_io_a = {_T_787,_T_788}; // @[Math.scala 151:17:@33843.4]
  assign x548_sum_1_io_b = RetimeWrapper_49_io_out; // @[Math.scala 152:17:@33844.4]
  assign x548_sum_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@33845.4]
  assign RetimeWrapper_50_clock = clock; // @[:@33851.4]
  assign RetimeWrapper_50_reset = reset; // @[:@33852.4]
  assign RetimeWrapper_50_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33854.4]
  assign RetimeWrapper_50_io_in = ~ x546; // @[package.scala 94:16:@33853.4]
  assign RetimeWrapper_51_clock = clock; // @[:@33865.4]
  assign RetimeWrapper_51_reset = reset; // @[:@33866.4]
  assign RetimeWrapper_51_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33868.4]
  assign RetimeWrapper_51_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33867.4]
  assign x553_rdcol_1_clock = clock; // @[:@33888.4]
  assign x553_rdcol_1_reset = reset; // @[:@33889.4]
  assign x553_rdcol_1_io_a = RetimeWrapper_47_io_out; // @[Math.scala 151:17:@33890.4]
  assign x553_rdcol_1_io_b = 32'hffffffff; // @[Math.scala 152:17:@33891.4]
  assign x553_rdcol_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@33892.4]
  assign x559_sum_1_clock = clock; // @[:@33920.4]
  assign x559_sum_1_reset = reset; // @[:@33921.4]
  assign x559_sum_1_io_a = {_T_787,_T_788}; // @[Math.scala 151:17:@33922.4]
  assign x559_sum_1_io_b = {_T_1003,_T_1004}; // @[Math.scala 152:17:@33923.4]
  assign x559_sum_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@33924.4]
  assign RetimeWrapper_52_clock = clock; // @[:@33930.4]
  assign RetimeWrapper_52_reset = reset; // @[:@33931.4]
  assign RetimeWrapper_52_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33933.4]
  assign RetimeWrapper_52_io_in = ~ x555; // @[package.scala 94:16:@33932.4]
  assign RetimeWrapper_53_clock = clock; // @[:@33944.4]
  assign RetimeWrapper_53_reset = reset; // @[:@33945.4]
  assign RetimeWrapper_53_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33947.4]
  assign RetimeWrapper_53_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33946.4]
  assign x565_rdcol_1_clock = clock; // @[:@33967.4]
  assign x565_rdcol_1_reset = reset; // @[:@33968.4]
  assign x565_rdcol_1_io_a = RetimeWrapper_47_io_out; // @[Math.scala 151:17:@33969.4]
  assign x565_rdcol_1_io_b = 32'hfffffffe; // @[Math.scala 152:17:@33970.4]
  assign x565_rdcol_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@33971.4]
  assign x571_sum_1_clock = clock; // @[:@33999.4]
  assign x571_sum_1_reset = reset; // @[:@34000.4]
  assign x571_sum_1_io_a = {_T_787,_T_788}; // @[Math.scala 151:17:@34001.4]
  assign x571_sum_1_io_b = {_T_1061,_T_1062}; // @[Math.scala 152:17:@34002.4]
  assign x571_sum_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@34003.4]
  assign RetimeWrapper_54_clock = clock; // @[:@34009.4]
  assign RetimeWrapper_54_reset = reset; // @[:@34010.4]
  assign RetimeWrapper_54_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34012.4]
  assign RetimeWrapper_54_io_in = ~ x567; // @[package.scala 94:16:@34011.4]
  assign RetimeWrapper_55_clock = clock; // @[:@34023.4]
  assign RetimeWrapper_55_reset = reset; // @[:@34024.4]
  assign RetimeWrapper_55_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34026.4]
  assign RetimeWrapper_55_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34025.4]
  assign RetimeWrapper_56_clock = clock; // @[:@34044.4]
  assign RetimeWrapper_56_reset = reset; // @[:@34045.4]
  assign RetimeWrapper_56_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34047.4]
  assign RetimeWrapper_56_io_in = __io_result; // @[package.scala 94:16:@34046.4]
  assign RetimeWrapper_57_clock = clock; // @[:@34071.4]
  assign RetimeWrapper_57_reset = reset; // @[:@34072.4]
  assign RetimeWrapper_57_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34074.4]
  assign RetimeWrapper_57_io_in = $signed(_T_1103) < $signed(32'sh0); // @[package.scala 94:16:@34073.4]
  assign RetimeWrapper_58_clock = clock; // @[:@34106.4]
  assign RetimeWrapper_58_reset = reset; // @[:@34107.4]
  assign RetimeWrapper_58_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34109.4]
  assign RetimeWrapper_58_io_in = {_T_1142,_T_1143}; // @[package.scala 94:16:@34108.4]
  assign x583_sum_1_clock = clock; // @[:@34115.4]
  assign x583_sum_1_reset = reset; // @[:@34116.4]
  assign x583_sum_1_io_a = RetimeWrapper_58_io_out; // @[Math.scala 151:17:@34117.4]
  assign x583_sum_1_io_b = RetimeWrapper_33_io_out; // @[Math.scala 152:17:@34118.4]
  assign x583_sum_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@34119.4]
  assign RetimeWrapper_59_clock = clock; // @[:@34125.4]
  assign RetimeWrapper_59_reset = reset; // @[:@34126.4]
  assign RetimeWrapper_59_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34128.4]
  assign RetimeWrapper_59_io_in = ~ x579; // @[package.scala 94:16:@34127.4]
  assign RetimeWrapper_60_clock = clock; // @[:@34134.4]
  assign RetimeWrapper_60_reset = reset; // @[:@34135.4]
  assign RetimeWrapper_60_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34137.4]
  assign RetimeWrapper_60_io_in = $unsigned(_T_1133); // @[package.scala 94:16:@34136.4]
  assign RetimeWrapper_61_clock = clock; // @[:@34148.4]
  assign RetimeWrapper_61_reset = reset; // @[:@34149.4]
  assign RetimeWrapper_61_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34151.4]
  assign RetimeWrapper_61_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34150.4]
  assign x591_sum_1_clock = clock; // @[:@34177.4]
  assign x591_sum_1_reset = reset; // @[:@34178.4]
  assign x591_sum_1_io_a = RetimeWrapper_58_io_out; // @[Math.scala 151:17:@34179.4]
  assign x591_sum_1_io_b = RetimeWrapper_40_io_out; // @[Math.scala 152:17:@34180.4]
  assign x591_sum_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@34181.4]
  assign RetimeWrapper_62_clock = clock; // @[:@34187.4]
  assign RetimeWrapper_62_reset = reset; // @[:@34188.4]
  assign RetimeWrapper_62_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34190.4]
  assign RetimeWrapper_62_io_in = ~ x589; // @[package.scala 94:16:@34189.4]
  assign RetimeWrapper_63_clock = clock; // @[:@34201.4]
  assign RetimeWrapper_63_reset = reset; // @[:@34202.4]
  assign RetimeWrapper_63_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34204.4]
  assign RetimeWrapper_63_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34203.4]
  assign x598_sum_1_clock = clock; // @[:@34228.4]
  assign x598_sum_1_reset = reset; // @[:@34229.4]
  assign x598_sum_1_io_a = RetimeWrapper_58_io_out; // @[Math.scala 151:17:@34230.4]
  assign x598_sum_1_io_b = RetimeWrapper_44_io_out; // @[Math.scala 152:17:@34231.4]
  assign x598_sum_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@34232.4]
  assign RetimeWrapper_64_clock = clock; // @[:@34238.4]
  assign RetimeWrapper_64_reset = reset; // @[:@34239.4]
  assign RetimeWrapper_64_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34241.4]
  assign RetimeWrapper_64_io_in = ~ x596; // @[package.scala 94:16:@34240.4]
  assign RetimeWrapper_65_clock = clock; // @[:@34252.4]
  assign RetimeWrapper_65_reset = reset; // @[:@34253.4]
  assign RetimeWrapper_65_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34255.4]
  assign RetimeWrapper_65_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34254.4]
  assign RetimeWrapper_66_clock = clock; // @[:@34279.4]
  assign RetimeWrapper_66_reset = reset; // @[:@34280.4]
  assign RetimeWrapper_66_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34282.4]
  assign RetimeWrapper_66_io_in = {_T_341,_T_342}; // @[package.scala 94:16:@34281.4]
  assign x605_sum_1_clock = clock; // @[:@34288.4]
  assign x605_sum_1_reset = reset; // @[:@34289.4]
  assign x605_sum_1_io_a = {_T_1142,_T_1143}; // @[Math.scala 151:17:@34290.4]
  assign x605_sum_1_io_b = RetimeWrapper_66_io_out; // @[Math.scala 152:17:@34291.4]
  assign x605_sum_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@34292.4]
  assign RetimeWrapper_67_clock = clock; // @[:@34298.4]
  assign RetimeWrapper_67_reset = reset; // @[:@34299.4]
  assign RetimeWrapper_67_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34301.4]
  assign RetimeWrapper_67_io_in = x605_sum_1_io_result; // @[package.scala 94:16:@34300.4]
  assign RetimeWrapper_68_clock = clock; // @[:@34307.4]
  assign RetimeWrapper_68_reset = reset; // @[:@34308.4]
  assign RetimeWrapper_68_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34310.4]
  assign RetimeWrapper_68_io_in = ~ x603; // @[package.scala 94:16:@34309.4]
  assign RetimeWrapper_69_clock = clock; // @[:@34321.4]
  assign RetimeWrapper_69_reset = reset; // @[:@34322.4]
  assign RetimeWrapper_69_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34324.4]
  assign RetimeWrapper_69_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34323.4]
  assign x612_sum_1_clock = clock; // @[:@34348.4]
  assign x612_sum_1_reset = reset; // @[:@34349.4]
  assign x612_sum_1_io_a = RetimeWrapper_58_io_out; // @[Math.scala 151:17:@34350.4]
  assign x612_sum_1_io_b = {_T_1003,_T_1004}; // @[Math.scala 152:17:@34351.4]
  assign x612_sum_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@34352.4]
  assign RetimeWrapper_70_clock = clock; // @[:@34358.4]
  assign RetimeWrapper_70_reset = reset; // @[:@34359.4]
  assign RetimeWrapper_70_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34361.4]
  assign RetimeWrapper_70_io_in = ~ x610; // @[package.scala 94:16:@34360.4]
  assign RetimeWrapper_71_clock = clock; // @[:@34372.4]
  assign RetimeWrapper_71_reset = reset; // @[:@34373.4]
  assign RetimeWrapper_71_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34375.4]
  assign RetimeWrapper_71_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34374.4]
  assign x619_sum_1_clock = clock; // @[:@34399.4]
  assign x619_sum_1_reset = reset; // @[:@34400.4]
  assign x619_sum_1_io_a = RetimeWrapper_58_io_out; // @[Math.scala 151:17:@34401.4]
  assign x619_sum_1_io_b = {_T_1061,_T_1062}; // @[Math.scala 152:17:@34402.4]
  assign x619_sum_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@34403.4]
  assign RetimeWrapper_72_clock = clock; // @[:@34409.4]
  assign RetimeWrapper_72_reset = reset; // @[:@34410.4]
  assign RetimeWrapper_72_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34412.4]
  assign RetimeWrapper_72_io_in = ~ x617; // @[package.scala 94:16:@34411.4]
  assign RetimeWrapper_73_clock = clock; // @[:@34423.4]
  assign RetimeWrapper_73_reset = reset; // @[:@34424.4]
  assign RetimeWrapper_73_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34426.4]
  assign RetimeWrapper_73_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34425.4]
  assign x624_rdrow_1_clock = clock; // @[:@34446.4]
  assign x624_rdrow_1_reset = reset; // @[:@34447.4]
  assign x624_rdrow_1_io_a = RetimeWrapper_56_io_out; // @[Math.scala 151:17:@34448.4]
  assign x624_rdrow_1_io_b = 32'hffffffff; // @[Math.scala 152:17:@34449.4]
  assign x624_rdrow_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@34450.4]
  assign x631_sum_1_clock = clock; // @[:@34500.4]
  assign x631_sum_1_reset = reset; // @[:@34501.4]
  assign x631_sum_1_io_a = {_T_1403,_T_1404}; // @[Math.scala 151:17:@34502.4]
  assign x631_sum_1_io_b = RetimeWrapper_33_io_out; // @[Math.scala 152:17:@34503.4]
  assign x631_sum_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@34504.4]
  assign RetimeWrapper_74_clock = clock; // @[:@34510.4]
  assign RetimeWrapper_74_reset = reset; // @[:@34511.4]
  assign RetimeWrapper_74_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34513.4]
  assign RetimeWrapper_74_io_in = ~ x627; // @[package.scala 94:16:@34512.4]
  assign RetimeWrapper_75_clock = clock; // @[:@34519.4]
  assign RetimeWrapper_75_reset = reset; // @[:@34520.4]
  assign RetimeWrapper_75_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34522.4]
  assign RetimeWrapper_75_io_in = $unsigned(_T_1394); // @[package.scala 94:16:@34521.4]
  assign RetimeWrapper_76_clock = clock; // @[:@34533.4]
  assign RetimeWrapper_76_reset = reset; // @[:@34534.4]
  assign RetimeWrapper_76_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34536.4]
  assign RetimeWrapper_76_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34535.4]
  assign x639_sum_1_clock = clock; // @[:@34562.4]
  assign x639_sum_1_reset = reset; // @[:@34563.4]
  assign x639_sum_1_io_a = {_T_1403,_T_1404}; // @[Math.scala 151:17:@34564.4]
  assign x639_sum_1_io_b = RetimeWrapper_40_io_out; // @[Math.scala 152:17:@34565.4]
  assign x639_sum_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@34566.4]
  assign RetimeWrapper_77_clock = clock; // @[:@34572.4]
  assign RetimeWrapper_77_reset = reset; // @[:@34573.4]
  assign RetimeWrapper_77_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34575.4]
  assign RetimeWrapper_77_io_in = ~ x637; // @[package.scala 94:16:@34574.4]
  assign RetimeWrapper_78_clock = clock; // @[:@34586.4]
  assign RetimeWrapper_78_reset = reset; // @[:@34587.4]
  assign RetimeWrapper_78_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34589.4]
  assign RetimeWrapper_78_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34588.4]
  assign x646_sum_1_clock = clock; // @[:@34613.4]
  assign x646_sum_1_reset = reset; // @[:@34614.4]
  assign x646_sum_1_io_a = {_T_1403,_T_1404}; // @[Math.scala 151:17:@34615.4]
  assign x646_sum_1_io_b = RetimeWrapper_44_io_out; // @[Math.scala 152:17:@34616.4]
  assign x646_sum_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@34617.4]
  assign RetimeWrapper_79_clock = clock; // @[:@34623.4]
  assign RetimeWrapper_79_reset = reset; // @[:@34624.4]
  assign RetimeWrapper_79_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34626.4]
  assign RetimeWrapper_79_io_in = ~ x644; // @[package.scala 94:16:@34625.4]
  assign RetimeWrapper_80_clock = clock; // @[:@34637.4]
  assign RetimeWrapper_80_reset = reset; // @[:@34638.4]
  assign RetimeWrapper_80_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34640.4]
  assign RetimeWrapper_80_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34639.4]
  assign x653_sum_1_clock = clock; // @[:@34664.4]
  assign x653_sum_1_reset = reset; // @[:@34665.4]
  assign x653_sum_1_io_a = {_T_1403,_T_1404}; // @[Math.scala 151:17:@34666.4]
  assign x653_sum_1_io_b = RetimeWrapper_49_io_out; // @[Math.scala 152:17:@34667.4]
  assign x653_sum_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@34668.4]
  assign RetimeWrapper_81_clock = clock; // @[:@34674.4]
  assign RetimeWrapper_81_reset = reset; // @[:@34675.4]
  assign RetimeWrapper_81_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34677.4]
  assign RetimeWrapper_81_io_in = ~ x651; // @[package.scala 94:16:@34676.4]
  assign RetimeWrapper_82_clock = clock; // @[:@34688.4]
  assign RetimeWrapper_82_reset = reset; // @[:@34689.4]
  assign RetimeWrapper_82_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34691.4]
  assign RetimeWrapper_82_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34690.4]
  assign x660_sum_1_clock = clock; // @[:@34715.4]
  assign x660_sum_1_reset = reset; // @[:@34716.4]
  assign x660_sum_1_io_a = {_T_1403,_T_1404}; // @[Math.scala 151:17:@34717.4]
  assign x660_sum_1_io_b = {_T_1003,_T_1004}; // @[Math.scala 152:17:@34718.4]
  assign x660_sum_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@34719.4]
  assign RetimeWrapper_83_clock = clock; // @[:@34725.4]
  assign RetimeWrapper_83_reset = reset; // @[:@34726.4]
  assign RetimeWrapper_83_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34728.4]
  assign RetimeWrapper_83_io_in = ~ x658; // @[package.scala 94:16:@34727.4]
  assign RetimeWrapper_84_clock = clock; // @[:@34739.4]
  assign RetimeWrapper_84_reset = reset; // @[:@34740.4]
  assign RetimeWrapper_84_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34742.4]
  assign RetimeWrapper_84_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34741.4]
  assign x667_sum_1_clock = clock; // @[:@34766.4]
  assign x667_sum_1_reset = reset; // @[:@34767.4]
  assign x667_sum_1_io_a = {_T_1403,_T_1404}; // @[Math.scala 151:17:@34768.4]
  assign x667_sum_1_io_b = {_T_1061,_T_1062}; // @[Math.scala 152:17:@34769.4]
  assign x667_sum_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@34770.4]
  assign RetimeWrapper_85_clock = clock; // @[:@34776.4]
  assign RetimeWrapper_85_reset = reset; // @[:@34777.4]
  assign RetimeWrapper_85_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34779.4]
  assign RetimeWrapper_85_io_in = ~ x665; // @[package.scala 94:16:@34778.4]
  assign RetimeWrapper_86_clock = clock; // @[:@34790.4]
  assign RetimeWrapper_86_reset = reset; // @[:@34791.4]
  assign RetimeWrapper_86_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34793.4]
  assign RetimeWrapper_86_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34792.4]
  assign x672_rdrow_1_clock = clock; // @[:@34813.4]
  assign x672_rdrow_1_reset = reset; // @[:@34814.4]
  assign x672_rdrow_1_io_a = RetimeWrapper_56_io_out; // @[Math.scala 151:17:@34815.4]
  assign x672_rdrow_1_io_b = 32'hfffffffe; // @[Math.scala 152:17:@34816.4]
  assign x672_rdrow_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@34817.4]
  assign x679_sum_1_clock = clock; // @[:@34867.4]
  assign x679_sum_1_reset = reset; // @[:@34868.4]
  assign x679_sum_1_io_a = {_T_1655,_T_1656}; // @[Math.scala 151:17:@34869.4]
  assign x679_sum_1_io_b = RetimeWrapper_33_io_out; // @[Math.scala 152:17:@34870.4]
  assign x679_sum_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@34871.4]
  assign RetimeWrapper_87_clock = clock; // @[:@34877.4]
  assign RetimeWrapper_87_reset = reset; // @[:@34878.4]
  assign RetimeWrapper_87_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34880.4]
  assign RetimeWrapper_87_io_in = $unsigned(_T_1646); // @[package.scala 94:16:@34879.4]
  assign RetimeWrapper_88_clock = clock; // @[:@34886.4]
  assign RetimeWrapper_88_reset = reset; // @[:@34887.4]
  assign RetimeWrapper_88_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34889.4]
  assign RetimeWrapper_88_io_in = ~ x675; // @[package.scala 94:16:@34888.4]
  assign RetimeWrapper_89_clock = clock; // @[:@34900.4]
  assign RetimeWrapper_89_reset = reset; // @[:@34901.4]
  assign RetimeWrapper_89_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34903.4]
  assign RetimeWrapper_89_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34902.4]
  assign x687_sum_1_clock = clock; // @[:@34927.4]
  assign x687_sum_1_reset = reset; // @[:@34928.4]
  assign x687_sum_1_io_a = {_T_1655,_T_1656}; // @[Math.scala 151:17:@34929.4]
  assign x687_sum_1_io_b = RetimeWrapper_40_io_out; // @[Math.scala 152:17:@34930.4]
  assign x687_sum_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@34931.4]
  assign RetimeWrapper_90_clock = clock; // @[:@34937.4]
  assign RetimeWrapper_90_reset = reset; // @[:@34938.4]
  assign RetimeWrapper_90_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34940.4]
  assign RetimeWrapper_90_io_in = ~ x685; // @[package.scala 94:16:@34939.4]
  assign RetimeWrapper_91_clock = clock; // @[:@34951.4]
  assign RetimeWrapper_91_reset = reset; // @[:@34952.4]
  assign RetimeWrapper_91_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34954.4]
  assign RetimeWrapper_91_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34953.4]
  assign x694_sum_1_clock = clock; // @[:@34980.4]
  assign x694_sum_1_reset = reset; // @[:@34981.4]
  assign x694_sum_1_io_a = {_T_1655,_T_1656}; // @[Math.scala 151:17:@34982.4]
  assign x694_sum_1_io_b = RetimeWrapper_44_io_out; // @[Math.scala 152:17:@34983.4]
  assign x694_sum_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@34984.4]
  assign RetimeWrapper_92_clock = clock; // @[:@34990.4]
  assign RetimeWrapper_92_reset = reset; // @[:@34991.4]
  assign RetimeWrapper_92_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34993.4]
  assign RetimeWrapper_92_io_in = ~ x692; // @[package.scala 94:16:@34992.4]
  assign RetimeWrapper_93_clock = clock; // @[:@35004.4]
  assign RetimeWrapper_93_reset = reset; // @[:@35005.4]
  assign RetimeWrapper_93_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35007.4]
  assign RetimeWrapper_93_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@35006.4]
  assign x701_sum_1_clock = clock; // @[:@35031.4]
  assign x701_sum_1_reset = reset; // @[:@35032.4]
  assign x701_sum_1_io_a = {_T_1655,_T_1656}; // @[Math.scala 151:17:@35033.4]
  assign x701_sum_1_io_b = RetimeWrapper_49_io_out; // @[Math.scala 152:17:@35034.4]
  assign x701_sum_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@35035.4]
  assign RetimeWrapper_94_clock = clock; // @[:@35041.4]
  assign RetimeWrapper_94_reset = reset; // @[:@35042.4]
  assign RetimeWrapper_94_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35044.4]
  assign RetimeWrapper_94_io_in = ~ x699; // @[package.scala 94:16:@35043.4]
  assign RetimeWrapper_95_clock = clock; // @[:@35055.4]
  assign RetimeWrapper_95_reset = reset; // @[:@35056.4]
  assign RetimeWrapper_95_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35058.4]
  assign RetimeWrapper_95_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@35057.4]
  assign x708_sum_1_clock = clock; // @[:@35082.4]
  assign x708_sum_1_reset = reset; // @[:@35083.4]
  assign x708_sum_1_io_a = {_T_1655,_T_1656}; // @[Math.scala 151:17:@35084.4]
  assign x708_sum_1_io_b = {_T_1003,_T_1004}; // @[Math.scala 152:17:@35085.4]
  assign x708_sum_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@35086.4]
  assign RetimeWrapper_96_clock = clock; // @[:@35092.4]
  assign RetimeWrapper_96_reset = reset; // @[:@35093.4]
  assign RetimeWrapper_96_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35095.4]
  assign RetimeWrapper_96_io_in = ~ x706; // @[package.scala 94:16:@35094.4]
  assign RetimeWrapper_97_clock = clock; // @[:@35106.4]
  assign RetimeWrapper_97_reset = reset; // @[:@35107.4]
  assign RetimeWrapper_97_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35109.4]
  assign RetimeWrapper_97_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@35108.4]
  assign x715_sum_1_clock = clock; // @[:@35133.4]
  assign x715_sum_1_reset = reset; // @[:@35134.4]
  assign x715_sum_1_io_a = {_T_1655,_T_1656}; // @[Math.scala 151:17:@35135.4]
  assign x715_sum_1_io_b = {_T_1061,_T_1062}; // @[Math.scala 152:17:@35136.4]
  assign x715_sum_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@35137.4]
  assign RetimeWrapper_98_clock = clock; // @[:@35143.4]
  assign RetimeWrapper_98_reset = reset; // @[:@35144.4]
  assign RetimeWrapper_98_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35146.4]
  assign RetimeWrapper_98_io_in = ~ x713; // @[package.scala 94:16:@35145.4]
  assign RetimeWrapper_99_clock = clock; // @[:@35157.4]
  assign RetimeWrapper_99_reset = reset; // @[:@35158.4]
  assign RetimeWrapper_99_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35160.4]
  assign RetimeWrapper_99_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@35159.4]
  assign x725_x11_1_clock = clock; // @[:@35203.4]
  assign x725_x11_1_reset = reset; // @[:@35204.4]
  assign x725_x11_1_io_a = x439_lb_0_io_rPort_3_output_0; // @[Math.scala 151:17:@35205.4]
  assign x725_x11_1_io_b = _T_1860[7:0]; // @[Math.scala 152:17:@35206.4]
  assign x725_x11_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@35207.4]
  assign x726_x12_1_clock = clock; // @[:@35213.4]
  assign x726_x12_1_reset = reset; // @[:@35214.4]
  assign x726_x12_1_io_a = x439_lb_0_io_rPort_23_output_0; // @[Math.scala 151:17:@35215.4]
  assign x726_x12_1_io_b = _T_1864[7:0]; // @[Math.scala 152:17:@35216.4]
  assign x726_x12_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@35217.4]
  assign x727_x11_1_clock = clock; // @[:@35223.4]
  assign x727_x11_1_reset = reset; // @[:@35224.4]
  assign x727_x11_1_io_a = _T_1868[7:0]; // @[Math.scala 151:17:@35225.4]
  assign x727_x11_1_io_b = _T_1872[7:0]; // @[Math.scala 152:17:@35226.4]
  assign x727_x11_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@35227.4]
  assign x728_x12_1_clock = clock; // @[:@35233.4]
  assign x728_x12_1_reset = reset; // @[:@35234.4]
  assign x728_x12_1_io_a = x439_lb_0_io_rPort_21_output_0; // @[Math.scala 151:17:@35235.4]
  assign x728_x12_1_io_b = _T_1876[7:0]; // @[Math.scala 152:17:@35236.4]
  assign x728_x12_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@35237.4]
  assign x729_x11_1_io_a = x725_x11_1_io_result; // @[Math.scala 151:17:@35245.4]
  assign x729_x11_1_io_b = x726_x12_1_io_result; // @[Math.scala 152:17:@35246.4]
  assign x730_x12_1_io_a = x727_x11_1_io_result; // @[Math.scala 151:17:@35255.4]
  assign x730_x12_1_io_b = x728_x12_1_io_result; // @[Math.scala 152:17:@35256.4]
  assign x731_x11_1_io_a = x729_x11_1_io_result; // @[Math.scala 151:17:@35265.4]
  assign x731_x11_1_io_b = x730_x12_1_io_result; // @[Math.scala 152:17:@35266.4]
  assign RetimeWrapper_100_clock = clock; // @[:@35273.4]
  assign RetimeWrapper_100_reset = reset; // @[:@35274.4]
  assign RetimeWrapper_100_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35276.4]
  assign RetimeWrapper_100_io_in = x439_lb_0_io_rPort_13_output_0; // @[package.scala 94:16:@35275.4]
  assign x732_sum_1_io_a = x731_x11_1_io_result; // @[Math.scala 151:17:@35284.4]
  assign x732_sum_1_io_b = RetimeWrapper_100_io_out; // @[Math.scala 152:17:@35285.4]
  assign RetimeWrapper_101_clock = clock; // @[:@35296.4]
  assign RetimeWrapper_101_reset = reset; // @[:@35297.4]
  assign RetimeWrapper_101_io_flow = io_in_x427_TREADY; // @[package.scala 95:18:@35299.4]
  assign RetimeWrapper_101_io_in = {4'h0,_T_1912}; // @[package.scala 94:16:@35298.4]
  assign x739_x11_1_clock = clock; // @[:@35331.4]
  assign x739_x11_1_reset = reset; // @[:@35332.4]
  assign x739_x11_1_io_a = x439_lb_0_io_rPort_14_output_0; // @[Math.scala 151:17:@35333.4]
  assign x739_x11_1_io_b = _T_1919[7:0]; // @[Math.scala 152:17:@35334.4]
  assign x739_x11_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@35335.4]
  assign x740_x12_1_clock = clock; // @[:@35341.4]
  assign x740_x12_1_reset = reset; // @[:@35342.4]
  assign x740_x12_1_io_a = x439_lb_0_io_rPort_4_output_0; // @[Math.scala 151:17:@35343.4]
  assign x740_x12_1_io_b = _T_1923[7:0]; // @[Math.scala 152:17:@35344.4]
  assign x740_x12_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@35345.4]
  assign x741_x11_1_clock = clock; // @[:@35351.4]
  assign x741_x11_1_reset = reset; // @[:@35352.4]
  assign x741_x11_1_io_a = _T_1927[7:0]; // @[Math.scala 151:17:@35353.4]
  assign x741_x11_1_io_b = _T_1931[7:0]; // @[Math.scala 152:17:@35354.4]
  assign x741_x11_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@35355.4]
  assign x742_x12_1_clock = clock; // @[:@35361.4]
  assign x742_x12_1_reset = reset; // @[:@35362.4]
  assign x742_x12_1_io_a = x439_lb_0_io_rPort_7_output_0; // @[Math.scala 151:17:@35363.4]
  assign x742_x12_1_io_b = _T_1935[7:0]; // @[Math.scala 152:17:@35364.4]
  assign x742_x12_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@35365.4]
  assign x743_x11_1_io_a = x739_x11_1_io_result; // @[Math.scala 151:17:@35373.4]
  assign x743_x11_1_io_b = x740_x12_1_io_result; // @[Math.scala 152:17:@35374.4]
  assign x744_x12_1_io_a = x741_x11_1_io_result; // @[Math.scala 151:17:@35383.4]
  assign x744_x12_1_io_b = x742_x12_1_io_result; // @[Math.scala 152:17:@35384.4]
  assign x745_x11_1_io_a = x743_x11_1_io_result; // @[Math.scala 151:17:@35393.4]
  assign x745_x11_1_io_b = x744_x12_1_io_result; // @[Math.scala 152:17:@35394.4]
  assign RetimeWrapper_102_clock = clock; // @[:@35401.4]
  assign RetimeWrapper_102_reset = reset; // @[:@35402.4]
  assign RetimeWrapper_102_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35404.4]
  assign RetimeWrapper_102_io_in = x439_lb_0_io_rPort_20_output_0; // @[package.scala 94:16:@35403.4]
  assign x746_sum_1_io_a = x745_x11_1_io_result; // @[Math.scala 151:17:@35414.4]
  assign x746_sum_1_io_b = RetimeWrapper_102_io_out; // @[Math.scala 152:17:@35415.4]
  assign RetimeWrapper_103_clock = clock; // @[:@35426.4]
  assign RetimeWrapper_103_reset = reset; // @[:@35427.4]
  assign RetimeWrapper_103_io_flow = io_in_x427_TREADY; // @[package.scala 95:18:@35429.4]
  assign RetimeWrapper_103_io_in = {4'h0,_T_1973}; // @[package.scala 94:16:@35428.4]
  assign x752_x11_1_clock = clock; // @[:@35456.4]
  assign x752_x11_1_reset = reset; // @[:@35457.4]
  assign x752_x11_1_io_a = x439_lb_0_io_rPort_23_output_0; // @[Math.scala 151:17:@35458.4]
  assign x752_x11_1_io_b = _T_1980[7:0]; // @[Math.scala 152:17:@35459.4]
  assign x752_x11_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@35460.4]
  assign x753_x12_1_clock = clock; // @[:@35466.4]
  assign x753_x12_1_reset = reset; // @[:@35467.4]
  assign x753_x12_1_io_a = x439_lb_0_io_rPort_17_output_0; // @[Math.scala 151:17:@35468.4]
  assign x753_x12_1_io_b = _T_1872[7:0]; // @[Math.scala 152:17:@35469.4]
  assign x753_x12_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@35470.4]
  assign x754_x11_1_clock = clock; // @[:@35476.4]
  assign x754_x11_1_reset = reset; // @[:@35477.4]
  assign x754_x11_1_io_a = _T_1984[7:0]; // @[Math.scala 151:17:@35478.4]
  assign x754_x11_1_io_b = _T_1988[7:0]; // @[Math.scala 152:17:@35479.4]
  assign x754_x11_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@35480.4]
  assign x755_x12_1_clock = clock; // @[:@35486.4]
  assign x755_x12_1_reset = reset; // @[:@35487.4]
  assign x755_x12_1_io_a = x439_lb_0_io_rPort_13_output_0; // @[Math.scala 151:17:@35488.4]
  assign x755_x12_1_io_b = _T_1992[7:0]; // @[Math.scala 152:17:@35489.4]
  assign x755_x12_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@35490.4]
  assign x756_x11_1_io_a = x752_x11_1_io_result; // @[Math.scala 151:17:@35498.4]
  assign x756_x11_1_io_b = x753_x12_1_io_result; // @[Math.scala 152:17:@35499.4]
  assign x757_x12_1_io_a = x754_x11_1_io_result; // @[Math.scala 151:17:@35508.4]
  assign x757_x12_1_io_b = x755_x12_1_io_result; // @[Math.scala 152:17:@35509.4]
  assign x758_x11_1_io_a = x756_x11_1_io_result; // @[Math.scala 151:17:@35518.4]
  assign x758_x11_1_io_b = x757_x12_1_io_result; // @[Math.scala 152:17:@35519.4]
  assign RetimeWrapper_104_clock = clock; // @[:@35526.4]
  assign RetimeWrapper_104_reset = reset; // @[:@35527.4]
  assign RetimeWrapper_104_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35529.4]
  assign RetimeWrapper_104_io_in = x439_lb_0_io_rPort_18_output_0; // @[package.scala 94:16:@35528.4]
  assign x759_sum_1_io_a = x758_x11_1_io_result; // @[Math.scala 151:17:@35537.4]
  assign x759_sum_1_io_b = RetimeWrapper_104_io_out; // @[Math.scala 152:17:@35538.4]
  assign RetimeWrapper_105_clock = clock; // @[:@35549.4]
  assign RetimeWrapper_105_reset = reset; // @[:@35550.4]
  assign RetimeWrapper_105_io_flow = io_in_x427_TREADY; // @[package.scala 95:18:@35552.4]
  assign RetimeWrapper_105_io_in = {4'h0,_T_2028}; // @[package.scala 94:16:@35551.4]
  assign x765_x11_1_clock = clock; // @[:@35579.4]
  assign x765_x11_1_reset = reset; // @[:@35580.4]
  assign x765_x11_1_io_a = x439_lb_0_io_rPort_4_output_0; // @[Math.scala 151:17:@35581.4]
  assign x765_x11_1_io_b = _T_2035[7:0]; // @[Math.scala 152:17:@35582.4]
  assign x765_x11_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@35583.4]
  assign x766_x12_1_clock = clock; // @[:@35589.4]
  assign x766_x12_1_reset = reset; // @[:@35590.4]
  assign x766_x12_1_io_a = x439_lb_0_io_rPort_22_output_0; // @[Math.scala 151:17:@35591.4]
  assign x766_x12_1_io_b = _T_1931[7:0]; // @[Math.scala 152:17:@35592.4]
  assign x766_x12_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@35593.4]
  assign x767_x11_1_clock = clock; // @[:@35599.4]
  assign x767_x11_1_reset = reset; // @[:@35600.4]
  assign x767_x11_1_io_a = _T_2039[7:0]; // @[Math.scala 151:17:@35601.4]
  assign x767_x11_1_io_b = _T_2043[7:0]; // @[Math.scala 152:17:@35602.4]
  assign x767_x11_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@35603.4]
  assign x768_x12_1_clock = clock; // @[:@35609.4]
  assign x768_x12_1_reset = reset; // @[:@35610.4]
  assign x768_x12_1_io_a = x439_lb_0_io_rPort_20_output_0; // @[Math.scala 151:17:@35611.4]
  assign x768_x12_1_io_b = _T_2047[7:0]; // @[Math.scala 152:17:@35612.4]
  assign x768_x12_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@35613.4]
  assign x769_x11_1_io_a = x765_x11_1_io_result; // @[Math.scala 151:17:@35621.4]
  assign x769_x11_1_io_b = x766_x12_1_io_result; // @[Math.scala 152:17:@35622.4]
  assign x770_x12_1_io_a = x767_x11_1_io_result; // @[Math.scala 151:17:@35631.4]
  assign x770_x12_1_io_b = x768_x12_1_io_result; // @[Math.scala 152:17:@35632.4]
  assign x771_x11_1_io_a = x769_x11_1_io_result; // @[Math.scala 151:17:@35641.4]
  assign x771_x11_1_io_b = x770_x12_1_io_result; // @[Math.scala 152:17:@35642.4]
  assign RetimeWrapper_106_clock = clock; // @[:@35649.4]
  assign RetimeWrapper_106_reset = reset; // @[:@35650.4]
  assign RetimeWrapper_106_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35652.4]
  assign RetimeWrapper_106_io_in = x439_lb_0_io_rPort_1_output_0; // @[package.scala 94:16:@35651.4]
  assign x772_sum_1_io_a = x771_x11_1_io_result; // @[Math.scala 151:17:@35660.4]
  assign x772_sum_1_io_b = RetimeWrapper_106_io_out; // @[Math.scala 152:17:@35661.4]
  assign RetimeWrapper_107_clock = clock; // @[:@35672.4]
  assign RetimeWrapper_107_reset = reset; // @[:@35673.4]
  assign RetimeWrapper_107_io_flow = io_in_x427_TREADY; // @[package.scala 95:18:@35675.4]
  assign RetimeWrapper_107_io_in = {4'h0,_T_2083}; // @[package.scala 94:16:@35674.4]
  assign x777_x11_1_clock = clock; // @[:@35697.4]
  assign x777_x11_1_reset = reset; // @[:@35698.4]
  assign x777_x11_1_io_a = x439_lb_0_io_rPort_2_output_0; // @[Math.scala 151:17:@35699.4]
  assign x777_x11_1_io_b = _T_1923[7:0]; // @[Math.scala 152:17:@35700.4]
  assign x777_x11_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@35701.4]
  assign x778_x12_1_clock = clock; // @[:@35707.4]
  assign x778_x12_1_reset = reset; // @[:@35708.4]
  assign x778_x12_1_io_a = x439_lb_0_io_rPort_10_output_0; // @[Math.scala 151:17:@35709.4]
  assign x778_x12_1_io_b = _T_2090[7:0]; // @[Math.scala 152:17:@35710.4]
  assign x778_x12_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@35711.4]
  assign x779_x11_1_clock = clock; // @[:@35717.4]
  assign x779_x11_1_reset = reset; // @[:@35718.4]
  assign x779_x11_1_io_a = _T_2094[7:0]; // @[Math.scala 151:17:@35719.4]
  assign x779_x11_1_io_b = _T_1935[7:0]; // @[Math.scala 152:17:@35720.4]
  assign x779_x11_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@35721.4]
  assign x780_x12_1_clock = clock; // @[:@35727.4]
  assign x780_x12_1_reset = reset; // @[:@35728.4]
  assign x780_x12_1_io_a = x439_lb_0_io_rPort_0_output_0; // @[Math.scala 151:17:@35729.4]
  assign x780_x12_1_io_b = _T_2098[7:0]; // @[Math.scala 152:17:@35730.4]
  assign x780_x12_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@35731.4]
  assign x781_x11_1_io_a = x777_x11_1_io_result; // @[Math.scala 151:17:@35739.4]
  assign x781_x11_1_io_b = x778_x12_1_io_result; // @[Math.scala 152:17:@35740.4]
  assign x782_x12_1_io_a = x779_x11_1_io_result; // @[Math.scala 151:17:@35749.4]
  assign x782_x12_1_io_b = x780_x12_1_io_result; // @[Math.scala 152:17:@35750.4]
  assign x783_x11_1_io_a = x781_x11_1_io_result; // @[Math.scala 151:17:@35759.4]
  assign x783_x11_1_io_b = x782_x12_1_io_result; // @[Math.scala 152:17:@35760.4]
  assign RetimeWrapper_108_clock = clock; // @[:@35767.4]
  assign RetimeWrapper_108_reset = reset; // @[:@35768.4]
  assign RetimeWrapper_108_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35770.4]
  assign RetimeWrapper_108_io_in = x439_lb_0_io_rPort_5_output_0; // @[package.scala 94:16:@35769.4]
  assign x784_sum_1_io_a = x783_x11_1_io_result; // @[Math.scala 151:17:@35778.4]
  assign x784_sum_1_io_b = RetimeWrapper_108_io_out; // @[Math.scala 152:17:@35779.4]
  assign RetimeWrapper_109_clock = clock; // @[:@35790.4]
  assign RetimeWrapper_109_reset = reset; // @[:@35791.4]
  assign RetimeWrapper_109_io_flow = io_in_x427_TREADY; // @[package.scala 95:18:@35793.4]
  assign RetimeWrapper_109_io_in = {4'h0,_T_2134}; // @[package.scala 94:16:@35792.4]
  assign x788_x11_1_clock = clock; // @[:@35810.4]
  assign x788_x11_1_reset = reset; // @[:@35811.4]
  assign x788_x11_1_io_a = x439_lb_0_io_rPort_15_output_0; // @[Math.scala 151:17:@35812.4]
  assign x788_x11_1_io_b = _T_1872[7:0]; // @[Math.scala 152:17:@35813.4]
  assign x788_x11_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@35814.4]
  assign x789_x12_1_clock = clock; // @[:@35820.4]
  assign x789_x12_1_reset = reset; // @[:@35821.4]
  assign x789_x12_1_io_a = x439_lb_0_io_rPort_16_output_0; // @[Math.scala 151:17:@35822.4]
  assign x789_x12_1_io_b = _T_1876[7:0]; // @[Math.scala 152:17:@35823.4]
  assign x789_x12_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@35824.4]
  assign x790_x11_1_clock = clock; // @[:@35830.4]
  assign x790_x11_1_reset = reset; // @[:@35831.4]
  assign x790_x11_1_io_a = _T_2141[7:0]; // @[Math.scala 151:17:@35832.4]
  assign x790_x11_1_io_b = _T_1992[7:0]; // @[Math.scala 152:17:@35833.4]
  assign x790_x11_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@35834.4]
  assign x791_x12_1_clock = clock; // @[:@35842.4]
  assign x791_x12_1_reset = reset; // @[:@35843.4]
  assign x791_x12_1_io_a = x439_lb_0_io_rPort_19_output_0; // @[Math.scala 151:17:@35844.4]
  assign x791_x12_1_io_b = _T_2145[7:0]; // @[Math.scala 152:17:@35845.4]
  assign x791_x12_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@35846.4]
  assign x792_x11_1_io_a = x788_x11_1_io_result; // @[Math.scala 151:17:@35854.4]
  assign x792_x11_1_io_b = x789_x12_1_io_result; // @[Math.scala 152:17:@35855.4]
  assign x793_x12_1_io_a = x790_x11_1_io_result; // @[Math.scala 151:17:@35864.4]
  assign x793_x12_1_io_b = x791_x12_1_io_result; // @[Math.scala 152:17:@35865.4]
  assign x794_x11_1_io_a = x792_x11_1_io_result; // @[Math.scala 151:17:@35874.4]
  assign x794_x11_1_io_b = x793_x12_1_io_result; // @[Math.scala 152:17:@35875.4]
  assign RetimeWrapper_110_clock = clock; // @[:@35882.4]
  assign RetimeWrapper_110_reset = reset; // @[:@35883.4]
  assign RetimeWrapper_110_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35885.4]
  assign RetimeWrapper_110_io_in = x439_lb_0_io_rPort_12_output_0; // @[package.scala 94:16:@35884.4]
  assign x795_sum_1_io_a = x794_x11_1_io_result; // @[Math.scala 151:17:@35893.4]
  assign x795_sum_1_io_b = RetimeWrapper_110_io_out; // @[Math.scala 152:17:@35894.4]
  assign RetimeWrapper_111_clock = clock; // @[:@35905.4]
  assign RetimeWrapper_111_reset = reset; // @[:@35906.4]
  assign RetimeWrapper_111_io_flow = io_in_x427_TREADY; // @[package.scala 95:18:@35908.4]
  assign RetimeWrapper_111_io_in = {4'h0,_T_2183}; // @[package.scala 94:16:@35907.4]
  assign x799_x11_1_clock = clock; // @[:@35925.4]
  assign x799_x11_1_reset = reset; // @[:@35926.4]
  assign x799_x11_1_io_a = x439_lb_0_io_rPort_10_output_0; // @[Math.scala 151:17:@35927.4]
  assign x799_x11_1_io_b = _T_1931[7:0]; // @[Math.scala 152:17:@35928.4]
  assign x799_x11_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@35929.4]
  assign x800_x12_1_clock = clock; // @[:@35935.4]
  assign x800_x12_1_reset = reset; // @[:@35936.4]
  assign x800_x12_1_io_a = x439_lb_0_io_rPort_6_output_0; // @[Math.scala 151:17:@35937.4]
  assign x800_x12_1_io_b = _T_1935[7:0]; // @[Math.scala 152:17:@35938.4]
  assign x800_x12_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@35939.4]
  assign x801_x11_1_clock = clock; // @[:@35945.4]
  assign x801_x11_1_reset = reset; // @[:@35946.4]
  assign x801_x11_1_io_a = _T_2190[7:0]; // @[Math.scala 151:17:@35947.4]
  assign x801_x11_1_io_b = _T_2047[7:0]; // @[Math.scala 152:17:@35948.4]
  assign x801_x11_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@35949.4]
  assign x802_x12_1_clock = clock; // @[:@35955.4]
  assign x802_x12_1_reset = reset; // @[:@35956.4]
  assign x802_x12_1_io_a = x439_lb_0_io_rPort_5_output_0; // @[Math.scala 151:17:@35957.4]
  assign x802_x12_1_io_b = _T_2194[7:0]; // @[Math.scala 152:17:@35958.4]
  assign x802_x12_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@35959.4]
  assign x803_x11_1_io_a = x799_x11_1_io_result; // @[Math.scala 151:17:@35967.4]
  assign x803_x11_1_io_b = x800_x12_1_io_result; // @[Math.scala 152:17:@35968.4]
  assign x804_x12_1_io_a = x801_x11_1_io_result; // @[Math.scala 151:17:@35977.4]
  assign x804_x12_1_io_b = x802_x12_1_io_result; // @[Math.scala 152:17:@35978.4]
  assign x805_x11_1_io_a = x803_x11_1_io_result; // @[Math.scala 151:17:@35987.4]
  assign x805_x11_1_io_b = x804_x12_1_io_result; // @[Math.scala 152:17:@35988.4]
  assign RetimeWrapper_112_clock = clock; // @[:@35995.4]
  assign RetimeWrapper_112_reset = reset; // @[:@35996.4]
  assign RetimeWrapper_112_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35998.4]
  assign RetimeWrapper_112_io_in = x439_lb_0_io_rPort_11_output_0; // @[package.scala 94:16:@35997.4]
  assign x806_sum_1_io_a = x805_x11_1_io_result; // @[Math.scala 151:17:@36006.4]
  assign x806_sum_1_io_b = RetimeWrapper_112_io_out; // @[Math.scala 152:17:@36007.4]
  assign RetimeWrapper_113_clock = clock; // @[:@36018.4]
  assign RetimeWrapper_113_reset = reset; // @[:@36019.4]
  assign RetimeWrapper_113_io_flow = io_in_x427_TREADY; // @[package.scala 95:18:@36021.4]
  assign RetimeWrapper_113_io_in = {4'h0,_T_2230}; // @[package.scala 94:16:@36020.4]
  assign x811_x11_1_clock = clock; // @[:@36043.4]
  assign x811_x11_1_reset = reset; // @[:@36044.4]
  assign x811_x11_1_io_a = x439_lb_0_io_rPort_16_output_0; // @[Math.scala 151:17:@36045.4]
  assign x811_x11_1_io_b = _T_1988[7:0]; // @[Math.scala 152:17:@36046.4]
  assign x811_x11_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@36047.4]
  assign x812_x12_1_clock = clock; // @[:@36053.4]
  assign x812_x12_1_reset = reset; // @[:@36054.4]
  assign x812_x12_1_io_a = x439_lb_0_io_rPort_8_output_0; // @[Math.scala 151:17:@36055.4]
  assign x812_x12_1_io_b = _T_1992[7:0]; // @[Math.scala 152:17:@36056.4]
  assign x812_x12_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@36057.4]
  assign x813_x11_1_clock = clock; // @[:@36063.4]
  assign x813_x11_1_reset = reset; // @[:@36064.4]
  assign x813_x11_1_io_a = _T_2237[7:0]; // @[Math.scala 151:17:@36065.4]
  assign x813_x11_1_io_b = _T_2241[7:0]; // @[Math.scala 152:17:@36066.4]
  assign x813_x11_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@36067.4]
  assign x814_x12_1_clock = clock; // @[:@36073.4]
  assign x814_x12_1_reset = reset; // @[:@36074.4]
  assign x814_x12_1_io_a = x439_lb_0_io_rPort_12_output_0; // @[Math.scala 151:17:@36075.4]
  assign x814_x12_1_io_b = _T_2245[7:0]; // @[Math.scala 152:17:@36076.4]
  assign x814_x12_1_io_flow = io_in_x427_TREADY; // @[Math.scala 153:20:@36077.4]
  assign x815_x11_1_io_a = x811_x11_1_io_result; // @[Math.scala 151:17:@36085.4]
  assign x815_x11_1_io_b = x812_x12_1_io_result; // @[Math.scala 152:17:@36086.4]
  assign x816_x12_1_io_a = x813_x11_1_io_result; // @[Math.scala 151:17:@36095.4]
  assign x816_x12_1_io_b = x814_x12_1_io_result; // @[Math.scala 152:17:@36096.4]
  assign x817_x11_1_io_a = x815_x11_1_io_result; // @[Math.scala 151:17:@36105.4]
  assign x817_x11_1_io_b = x816_x12_1_io_result; // @[Math.scala 152:17:@36106.4]
  assign RetimeWrapper_114_clock = clock; // @[:@36113.4]
  assign RetimeWrapper_114_reset = reset; // @[:@36114.4]
  assign RetimeWrapper_114_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@36116.4]
  assign RetimeWrapper_114_io_in = x439_lb_0_io_rPort_9_output_0; // @[package.scala 94:16:@36115.4]
  assign x818_sum_1_io_a = x817_x11_1_io_result; // @[Math.scala 151:17:@36124.4]
  assign x818_sum_1_io_b = RetimeWrapper_114_io_out; // @[Math.scala 152:17:@36125.4]
  assign RetimeWrapper_115_clock = clock; // @[:@36136.4]
  assign RetimeWrapper_115_reset = reset; // @[:@36137.4]
  assign RetimeWrapper_115_io_flow = io_in_x427_TREADY; // @[package.scala 95:18:@36139.4]
  assign RetimeWrapper_115_io_in = {4'h0,_T_2281}; // @[package.scala 94:16:@36138.4]
  assign RetimeWrapper_116_clock = clock; // @[:@36164.4]
  assign RetimeWrapper_116_reset = reset; // @[:@36165.4]
  assign RetimeWrapper_116_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@36167.4]
  assign RetimeWrapper_116_io_in = {_T_2305,_T_2302}; // @[package.scala 94:16:@36166.4]
  assign RetimeWrapper_117_clock = clock; // @[:@36173.4]
  assign RetimeWrapper_117_reset = reset; // @[:@36174.4]
  assign RetimeWrapper_117_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@36176.4]
  assign RetimeWrapper_117_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@36175.4]
  assign RetimeWrapper_118_clock = clock; // @[:@36182.4]
  assign RetimeWrapper_118_reset = reset; // @[:@36183.4]
  assign RetimeWrapper_118_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@36185.4]
  assign RetimeWrapper_118_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@36184.4]
  assign RetimeWrapper_119_clock = clock; // @[:@36191.4]
  assign RetimeWrapper_119_reset = reset; // @[:@36192.4]
  assign RetimeWrapper_119_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@36194.4]
  assign RetimeWrapper_119_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@36193.4]
endmodule
module x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1( // @[:@36212.2]
  input          clock, // @[:@36213.4]
  input          reset, // @[:@36214.4]
  input          io_in_x426_TVALID, // @[:@36215.4]
  output         io_in_x426_TREADY, // @[:@36215.4]
  input  [255:0] io_in_x426_TDATA, // @[:@36215.4]
  input  [7:0]   io_in_x426_TID, // @[:@36215.4]
  input  [7:0]   io_in_x426_TDEST, // @[:@36215.4]
  output         io_in_x427_TVALID, // @[:@36215.4]
  input          io_in_x427_TREADY, // @[:@36215.4]
  output [255:0] io_in_x427_TDATA, // @[:@36215.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@36215.4]
  input          io_sigsIn_smChildAcks_0, // @[:@36215.4]
  output         io_sigsOut_smDoneIn_0, // @[:@36215.4]
  output         io_sigsOut_smCtrCopyDone_0, // @[:@36215.4]
  input          io_rr // @[:@36215.4]
);
  wire  x434_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@36225.4]
  wire  x434_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@36225.4]
  wire  x434_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@36225.4]
  wire  x434_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@36225.4]
  wire [31:0] x434_ctrchain_io_output_counts_1; // @[SpatialBlocks.scala 37:22:@36225.4]
  wire [31:0] x434_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@36225.4]
  wire  x434_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@36225.4]
  wire  x434_ctrchain_io_output_oobs_1; // @[SpatialBlocks.scala 37:22:@36225.4]
  wire  x434_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@36225.4]
  wire  x824_inr_Foreach_SAMPLER_BOX_sm_clock; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 32:18:@36284.4]
  wire  x824_inr_Foreach_SAMPLER_BOX_sm_reset; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 32:18:@36284.4]
  wire  x824_inr_Foreach_SAMPLER_BOX_sm_io_enable; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 32:18:@36284.4]
  wire  x824_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 32:18:@36284.4]
  wire  x824_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 32:18:@36284.4]
  wire  x824_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 32:18:@36284.4]
  wire  x824_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 32:18:@36284.4]
  wire  x824_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 32:18:@36284.4]
  wire  x824_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 32:18:@36284.4]
  wire  x824_inr_Foreach_SAMPLER_BOX_sm_io_parentAck; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 32:18:@36284.4]
  wire  x824_inr_Foreach_SAMPLER_BOX_sm_io_backpressure; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 32:18:@36284.4]
  wire  x824_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 32:18:@36284.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@36312.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@36312.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@36312.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@36312.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@36312.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@36354.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@36354.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@36354.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@36354.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@36354.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@36362.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@36362.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@36362.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@36362.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@36362.4]
  wire  x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_clock; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 992:24:@36394.4]
  wire  x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_reset; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 992:24:@36394.4]
  wire  x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x426_TREADY; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 992:24:@36394.4]
  wire [255:0] x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x426_TDATA; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 992:24:@36394.4]
  wire [7:0] x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x426_TID; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 992:24:@36394.4]
  wire [7:0] x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x426_TDEST; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 992:24:@36394.4]
  wire  x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x427_TVALID; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 992:24:@36394.4]
  wire  x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x427_TREADY; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 992:24:@36394.4]
  wire [255:0] x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x427_TDATA; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 992:24:@36394.4]
  wire  x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 992:24:@36394.4]
  wire  x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 992:24:@36394.4]
  wire  x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 992:24:@36394.4]
  wire [31:0] x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 992:24:@36394.4]
  wire [31:0] x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 992:24:@36394.4]
  wire  x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 992:24:@36394.4]
  wire  x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 992:24:@36394.4]
  wire  x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_rr; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 992:24:@36394.4]
  wire  _T_239; // @[package.scala 96:25:@36317.4 package.scala 96:25:@36318.4]
  wire  x824_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[sm_x825_outr_UnitPipe.scala 68:66:@36323.4]
  wire  _T_252; // @[package.scala 96:25:@36359.4 package.scala 96:25:@36360.4]
  wire  _T_258; // @[package.scala 96:25:@36367.4 package.scala 96:25:@36368.4]
  wire  _T_261; // @[SpatialBlocks.scala 110:93:@36370.4]
  wire  x824_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn; // @[SpatialBlocks.scala 110:90:@36371.4]
  wire  _T_263; // @[SpatialBlocks.scala 128:36:@36379.4]
  wire  _T_264; // @[SpatialBlocks.scala 128:78:@36380.4]
  wire  _T_269; // @[SpatialBlocks.scala 130:61:@36389.4]
  x434_ctrchain x434_ctrchain ( // @[SpatialBlocks.scala 37:22:@36225.4]
    .clock(x434_ctrchain_clock),
    .reset(x434_ctrchain_reset),
    .io_input_reset(x434_ctrchain_io_input_reset),
    .io_input_enable(x434_ctrchain_io_input_enable),
    .io_output_counts_1(x434_ctrchain_io_output_counts_1),
    .io_output_counts_0(x434_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x434_ctrchain_io_output_oobs_0),
    .io_output_oobs_1(x434_ctrchain_io_output_oobs_1),
    .io_output_done(x434_ctrchain_io_output_done)
  );
  x824_inr_Foreach_SAMPLER_BOX_sm x824_inr_Foreach_SAMPLER_BOX_sm ( // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 32:18:@36284.4]
    .clock(x824_inr_Foreach_SAMPLER_BOX_sm_clock),
    .reset(x824_inr_Foreach_SAMPLER_BOX_sm_reset),
    .io_enable(x824_inr_Foreach_SAMPLER_BOX_sm_io_enable),
    .io_done(x824_inr_Foreach_SAMPLER_BOX_sm_io_done),
    .io_doneLatch(x824_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch),
    .io_ctrDone(x824_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone),
    .io_datapathEn(x824_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn),
    .io_ctrInc(x824_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc),
    .io_ctrRst(x824_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst),
    .io_parentAck(x824_inr_Foreach_SAMPLER_BOX_sm_io_parentAck),
    .io_backpressure(x824_inr_Foreach_SAMPLER_BOX_sm_io_backpressure),
    .io_break(x824_inr_Foreach_SAMPLER_BOX_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@36312.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@36354.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@36362.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1 x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1 ( // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 992:24:@36394.4]
    .clock(x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_clock),
    .reset(x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_reset),
    .io_in_x426_TREADY(x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x426_TREADY),
    .io_in_x426_TDATA(x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x426_TDATA),
    .io_in_x426_TID(x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x426_TID),
    .io_in_x426_TDEST(x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x426_TDEST),
    .io_in_x427_TVALID(x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x427_TVALID),
    .io_in_x427_TREADY(x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x427_TREADY),
    .io_in_x427_TDATA(x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x427_TDATA),
    .io_sigsIn_backpressure(x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_1(x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsIn_cchainOutputs_0_oobs_1(x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1),
    .io_rr(x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_rr)
  );
  assign _T_239 = RetimeWrapper_io_out; // @[package.scala 96:25:@36317.4 package.scala 96:25:@36318.4]
  assign x824_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure = io_in_x426_TVALID | x824_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x825_outr_UnitPipe.scala 68:66:@36323.4]
  assign _T_252 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@36359.4 package.scala 96:25:@36360.4]
  assign _T_258 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@36367.4 package.scala 96:25:@36368.4]
  assign _T_261 = ~ _T_258; // @[SpatialBlocks.scala 110:93:@36370.4]
  assign x824_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn = _T_252 & _T_261; // @[SpatialBlocks.scala 110:90:@36371.4]
  assign _T_263 = x824_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[SpatialBlocks.scala 128:36:@36379.4]
  assign _T_264 = ~ x824_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[SpatialBlocks.scala 128:78:@36380.4]
  assign _T_269 = x824_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[SpatialBlocks.scala 130:61:@36389.4]
  assign io_in_x426_TREADY = x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x426_TREADY; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 48:23:@36451.4]
  assign io_in_x427_TVALID = x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x427_TVALID; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 49:23:@36461.4]
  assign io_in_x427_TDATA = x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x427_TDATA; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 49:23:@36459.4]
  assign io_sigsOut_smDoneIn_0 = x824_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[SpatialBlocks.scala 127:53:@36377.4]
  assign io_sigsOut_smCtrCopyDone_0 = x824_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[SpatialBlocks.scala 139:125:@36393.4]
  assign x434_ctrchain_clock = clock; // @[:@36226.4]
  assign x434_ctrchain_reset = reset; // @[:@36227.4]
  assign x434_ctrchain_io_input_reset = x824_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[SpatialBlocks.scala 130:103:@36392.4]
  assign x434_ctrchain_io_input_enable = _T_269 & x824_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 104:75:@36347.4 SpatialBlocks.scala 130:45:@36391.4]
  assign x824_inr_Foreach_SAMPLER_BOX_sm_clock = clock; // @[:@36285.4]
  assign x824_inr_Foreach_SAMPLER_BOX_sm_reset = reset; // @[:@36286.4]
  assign x824_inr_Foreach_SAMPLER_BOX_sm_io_enable = x824_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn & x824_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 112:18:@36374.4]
  assign x824_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone = io_rr ? _T_239 : 1'h0; // @[sm_x825_outr_UnitPipe.scala 66:50:@36320.4]
  assign x824_inr_Foreach_SAMPLER_BOX_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 114:21:@36376.4]
  assign x824_inr_Foreach_SAMPLER_BOX_sm_io_backpressure = io_in_x427_TREADY | x824_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[SpatialBlocks.scala 105:24:@36348.4]
  assign x824_inr_Foreach_SAMPLER_BOX_sm_io_break = 1'h0; // @[sm_x825_outr_UnitPipe.scala 70:48:@36326.4]
  assign RetimeWrapper_clock = clock; // @[:@36313.4]
  assign RetimeWrapper_reset = reset; // @[:@36314.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@36316.4]
  assign RetimeWrapper_io_in = x434_ctrchain_io_output_done; // @[package.scala 94:16:@36315.4]
  assign RetimeWrapper_1_clock = clock; // @[:@36355.4]
  assign RetimeWrapper_1_reset = reset; // @[:@36356.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@36358.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@36357.4]
  assign RetimeWrapper_2_clock = clock; // @[:@36363.4]
  assign RetimeWrapper_2_reset = reset; // @[:@36364.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@36366.4]
  assign RetimeWrapper_2_io_in = x824_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[package.scala 94:16:@36365.4]
  assign x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_clock = clock; // @[:@36395.4]
  assign x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_reset = reset; // @[:@36396.4]
  assign x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x426_TDATA = io_in_x426_TDATA; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 48:23:@36450.4]
  assign x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x426_TID = io_in_x426_TID; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 48:23:@36446.4]
  assign x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x426_TDEST = io_in_x426_TDEST; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 48:23:@36445.4]
  assign x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x427_TREADY = io_in_x427_TREADY; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 49:23:@36460.4]
  assign x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure = io_in_x427_TREADY | x824_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 996:22:@36478.4]
  assign x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn = _T_263 & _T_264; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 996:22:@36476.4]
  assign x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break = x824_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 996:22:@36474.4]
  assign x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1 = x434_ctrchain_io_output_counts_1; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 996:22:@36469.4]
  assign x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = x434_ctrchain_io_output_counts_0; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 996:22:@36468.4]
  assign x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x434_ctrchain_io_output_oobs_0; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 996:22:@36466.4]
  assign x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1 = x434_ctrchain_io_output_oobs_1; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 996:22:@36467.4]
  assign x824_inr_Foreach_SAMPLER_BOX_kernelx824_inr_Foreach_SAMPLER_BOX_concrete1_io_rr = io_rr; // @[sm_x824_inr_Foreach_SAMPLER_BOX.scala 995:18:@36462.4]
endmodule
module RootController_kernelRootController_concrete1( // @[:@36491.2]
  input          clock, // @[:@36492.4]
  input          reset, // @[:@36493.4]
  input          io_in_x426_TVALID, // @[:@36494.4]
  output         io_in_x426_TREADY, // @[:@36494.4]
  input  [255:0] io_in_x426_TDATA, // @[:@36494.4]
  input  [7:0]   io_in_x426_TID, // @[:@36494.4]
  input  [7:0]   io_in_x426_TDEST, // @[:@36494.4]
  output         io_in_x427_TVALID, // @[:@36494.4]
  input          io_in_x427_TREADY, // @[:@36494.4]
  output [255:0] io_in_x427_TDATA, // @[:@36494.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@36494.4]
  input          io_sigsIn_smChildAcks_0, // @[:@36494.4]
  output         io_sigsOut_smDoneIn_0, // @[:@36494.4]
  input          io_rr // @[:@36494.4]
);
  wire  x825_outr_UnitPipe_sm_clock; // @[sm_x825_outr_UnitPipe.scala 32:18:@36635.4]
  wire  x825_outr_UnitPipe_sm_reset; // @[sm_x825_outr_UnitPipe.scala 32:18:@36635.4]
  wire  x825_outr_UnitPipe_sm_io_enable; // @[sm_x825_outr_UnitPipe.scala 32:18:@36635.4]
  wire  x825_outr_UnitPipe_sm_io_done; // @[sm_x825_outr_UnitPipe.scala 32:18:@36635.4]
  wire  x825_outr_UnitPipe_sm_io_parentAck; // @[sm_x825_outr_UnitPipe.scala 32:18:@36635.4]
  wire  x825_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x825_outr_UnitPipe.scala 32:18:@36635.4]
  wire  x825_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x825_outr_UnitPipe.scala 32:18:@36635.4]
  wire  x825_outr_UnitPipe_sm_io_childAck_0; // @[sm_x825_outr_UnitPipe.scala 32:18:@36635.4]
  wire  x825_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x825_outr_UnitPipe.scala 32:18:@36635.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@36687.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@36687.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@36687.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@36687.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@36687.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@36695.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@36695.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@36695.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@36695.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@36695.4]
  wire  x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_clock; // @[sm_x825_outr_UnitPipe.scala 75:24:@36722.4]
  wire  x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_reset; // @[sm_x825_outr_UnitPipe.scala 75:24:@36722.4]
  wire  x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_io_in_x426_TVALID; // @[sm_x825_outr_UnitPipe.scala 75:24:@36722.4]
  wire  x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_io_in_x426_TREADY; // @[sm_x825_outr_UnitPipe.scala 75:24:@36722.4]
  wire [255:0] x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_io_in_x426_TDATA; // @[sm_x825_outr_UnitPipe.scala 75:24:@36722.4]
  wire [7:0] x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_io_in_x426_TID; // @[sm_x825_outr_UnitPipe.scala 75:24:@36722.4]
  wire [7:0] x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_io_in_x426_TDEST; // @[sm_x825_outr_UnitPipe.scala 75:24:@36722.4]
  wire  x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_io_in_x427_TVALID; // @[sm_x825_outr_UnitPipe.scala 75:24:@36722.4]
  wire  x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_io_in_x427_TREADY; // @[sm_x825_outr_UnitPipe.scala 75:24:@36722.4]
  wire [255:0] x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_io_in_x427_TDATA; // @[sm_x825_outr_UnitPipe.scala 75:24:@36722.4]
  wire  x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x825_outr_UnitPipe.scala 75:24:@36722.4]
  wire  x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x825_outr_UnitPipe.scala 75:24:@36722.4]
  wire  x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x825_outr_UnitPipe.scala 75:24:@36722.4]
  wire  x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x825_outr_UnitPipe.scala 75:24:@36722.4]
  wire  x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_io_rr; // @[sm_x825_outr_UnitPipe.scala 75:24:@36722.4]
  wire  _T_246; // @[package.scala 96:25:@36692.4 package.scala 96:25:@36693.4]
  wire  _T_252; // @[package.scala 96:25:@36700.4 package.scala 96:25:@36701.4]
  wire  _T_255; // @[SpatialBlocks.scala 110:93:@36703.4]
  x825_outr_UnitPipe_sm x825_outr_UnitPipe_sm ( // @[sm_x825_outr_UnitPipe.scala 32:18:@36635.4]
    .clock(x825_outr_UnitPipe_sm_clock),
    .reset(x825_outr_UnitPipe_sm_reset),
    .io_enable(x825_outr_UnitPipe_sm_io_enable),
    .io_done(x825_outr_UnitPipe_sm_io_done),
    .io_parentAck(x825_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x825_outr_UnitPipe_sm_io_doneIn_0),
    .io_enableOut_0(x825_outr_UnitPipe_sm_io_enableOut_0),
    .io_childAck_0(x825_outr_UnitPipe_sm_io_childAck_0),
    .io_ctrCopyDone_0(x825_outr_UnitPipe_sm_io_ctrCopyDone_0)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@36687.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@36695.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1 x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1 ( // @[sm_x825_outr_UnitPipe.scala 75:24:@36722.4]
    .clock(x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_clock),
    .reset(x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_reset),
    .io_in_x426_TVALID(x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_io_in_x426_TVALID),
    .io_in_x426_TREADY(x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_io_in_x426_TREADY),
    .io_in_x426_TDATA(x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_io_in_x426_TDATA),
    .io_in_x426_TID(x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_io_in_x426_TID),
    .io_in_x426_TDEST(x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_io_in_x426_TDEST),
    .io_in_x427_TVALID(x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_io_in_x427_TVALID),
    .io_in_x427_TREADY(x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_io_in_x427_TREADY),
    .io_in_x427_TDATA(x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_io_in_x427_TDATA),
    .io_sigsIn_smEnableOuts_0(x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smCtrCopyDone_0(x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_rr(x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_246 = RetimeWrapper_io_out; // @[package.scala 96:25:@36692.4 package.scala 96:25:@36693.4]
  assign _T_252 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@36700.4 package.scala 96:25:@36701.4]
  assign _T_255 = ~ _T_252; // @[SpatialBlocks.scala 110:93:@36703.4]
  assign io_in_x426_TREADY = x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_io_in_x426_TREADY; // @[sm_x825_outr_UnitPipe.scala 48:23:@36777.4]
  assign io_in_x427_TVALID = x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_io_in_x427_TVALID; // @[sm_x825_outr_UnitPipe.scala 49:23:@36787.4]
  assign io_in_x427_TDATA = x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_io_in_x427_TDATA; // @[sm_x825_outr_UnitPipe.scala 49:23:@36785.4]
  assign io_sigsOut_smDoneIn_0 = x825_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 127:53:@36710.4]
  assign x825_outr_UnitPipe_sm_clock = clock; // @[:@36636.4]
  assign x825_outr_UnitPipe_sm_reset = reset; // @[:@36637.4]
  assign x825_outr_UnitPipe_sm_io_enable = _T_246 & _T_255; // @[SpatialBlocks.scala 112:18:@36707.4]
  assign x825_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 114:21:@36709.4]
  assign x825_outr_UnitPipe_sm_io_doneIn_0 = x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 102:67:@36679.4]
  assign x825_outr_UnitPipe_sm_io_ctrCopyDone_0 = x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 132:80:@36721.4]
  assign RetimeWrapper_clock = clock; // @[:@36688.4]
  assign RetimeWrapper_reset = reset; // @[:@36689.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@36691.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@36690.4]
  assign RetimeWrapper_1_clock = clock; // @[:@36696.4]
  assign RetimeWrapper_1_reset = reset; // @[:@36697.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@36699.4]
  assign RetimeWrapper_1_io_in = x825_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@36698.4]
  assign x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_clock = clock; // @[:@36723.4]
  assign x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_reset = reset; // @[:@36724.4]
  assign x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_io_in_x426_TVALID = io_in_x426_TVALID; // @[sm_x825_outr_UnitPipe.scala 48:23:@36778.4]
  assign x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_io_in_x426_TDATA = io_in_x426_TDATA; // @[sm_x825_outr_UnitPipe.scala 48:23:@36776.4]
  assign x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_io_in_x426_TID = io_in_x426_TID; // @[sm_x825_outr_UnitPipe.scala 48:23:@36772.4]
  assign x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_io_in_x426_TDEST = io_in_x426_TDEST; // @[sm_x825_outr_UnitPipe.scala 48:23:@36771.4]
  assign x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_io_in_x427_TREADY = io_in_x427_TREADY; // @[sm_x825_outr_UnitPipe.scala 49:23:@36786.4]
  assign x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x825_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x825_outr_UnitPipe.scala 79:22:@36796.4]
  assign x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x825_outr_UnitPipe_sm_io_childAck_0; // @[sm_x825_outr_UnitPipe.scala 79:22:@36794.4]
  assign x825_outr_UnitPipe_kernelx825_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x825_outr_UnitPipe.scala 78:18:@36788.4]
endmodule
module AccelUnit( // @[:@36815.2]
  input          clock, // @[:@36816.4]
  input          reset, // @[:@36817.4]
  input          io_enable, // @[:@36818.4]
  output         io_done, // @[:@36818.4]
  input          io_reset, // @[:@36818.4]
  input          io_memStreams_loads_0_cmd_ready, // @[:@36818.4]
  output         io_memStreams_loads_0_cmd_valid, // @[:@36818.4]
  output [63:0]  io_memStreams_loads_0_cmd_bits_addr, // @[:@36818.4]
  output [31:0]  io_memStreams_loads_0_cmd_bits_size, // @[:@36818.4]
  output         io_memStreams_loads_0_data_ready, // @[:@36818.4]
  input          io_memStreams_loads_0_data_valid, // @[:@36818.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_0, // @[:@36818.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_1, // @[:@36818.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_2, // @[:@36818.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_3, // @[:@36818.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_4, // @[:@36818.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_5, // @[:@36818.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_6, // @[:@36818.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_7, // @[:@36818.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_8, // @[:@36818.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_9, // @[:@36818.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_10, // @[:@36818.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_11, // @[:@36818.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_12, // @[:@36818.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_13, // @[:@36818.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_14, // @[:@36818.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_15, // @[:@36818.4]
  input          io_memStreams_stores_0_cmd_ready, // @[:@36818.4]
  output         io_memStreams_stores_0_cmd_valid, // @[:@36818.4]
  output [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@36818.4]
  output [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@36818.4]
  input          io_memStreams_stores_0_data_ready, // @[:@36818.4]
  output         io_memStreams_stores_0_data_valid, // @[:@36818.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_0, // @[:@36818.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_1, // @[:@36818.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_2, // @[:@36818.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_3, // @[:@36818.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_4, // @[:@36818.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_5, // @[:@36818.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_6, // @[:@36818.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_7, // @[:@36818.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_8, // @[:@36818.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_9, // @[:@36818.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_10, // @[:@36818.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_11, // @[:@36818.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_12, // @[:@36818.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_13, // @[:@36818.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_14, // @[:@36818.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_15, // @[:@36818.4]
  output [15:0]  io_memStreams_stores_0_data_bits_wstrb, // @[:@36818.4]
  output         io_memStreams_stores_0_wresp_ready, // @[:@36818.4]
  input          io_memStreams_stores_0_wresp_valid, // @[:@36818.4]
  input          io_memStreams_stores_0_wresp_bits, // @[:@36818.4]
  input          io_memStreams_gathers_0_cmd_ready, // @[:@36818.4]
  output         io_memStreams_gathers_0_cmd_valid, // @[:@36818.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_0, // @[:@36818.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_1, // @[:@36818.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_2, // @[:@36818.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_3, // @[:@36818.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_4, // @[:@36818.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_5, // @[:@36818.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_6, // @[:@36818.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_7, // @[:@36818.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_8, // @[:@36818.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_9, // @[:@36818.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_10, // @[:@36818.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_11, // @[:@36818.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_12, // @[:@36818.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_13, // @[:@36818.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_14, // @[:@36818.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_15, // @[:@36818.4]
  output         io_memStreams_gathers_0_data_ready, // @[:@36818.4]
  input          io_memStreams_gathers_0_data_valid, // @[:@36818.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_0, // @[:@36818.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_1, // @[:@36818.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_2, // @[:@36818.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_3, // @[:@36818.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_4, // @[:@36818.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_5, // @[:@36818.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_6, // @[:@36818.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_7, // @[:@36818.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_8, // @[:@36818.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_9, // @[:@36818.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_10, // @[:@36818.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_11, // @[:@36818.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_12, // @[:@36818.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_13, // @[:@36818.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_14, // @[:@36818.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_15, // @[:@36818.4]
  input          io_memStreams_scatters_0_cmd_ready, // @[:@36818.4]
  output         io_memStreams_scatters_0_cmd_valid, // @[:@36818.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_0, // @[:@36818.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_1, // @[:@36818.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_2, // @[:@36818.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_3, // @[:@36818.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_4, // @[:@36818.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_5, // @[:@36818.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_6, // @[:@36818.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_7, // @[:@36818.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_8, // @[:@36818.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_9, // @[:@36818.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_10, // @[:@36818.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_11, // @[:@36818.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_12, // @[:@36818.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_13, // @[:@36818.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_14, // @[:@36818.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_15, // @[:@36818.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_0, // @[:@36818.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_1, // @[:@36818.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_2, // @[:@36818.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_3, // @[:@36818.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_4, // @[:@36818.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_5, // @[:@36818.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_6, // @[:@36818.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_7, // @[:@36818.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_8, // @[:@36818.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_9, // @[:@36818.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_10, // @[:@36818.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_11, // @[:@36818.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_12, // @[:@36818.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_13, // @[:@36818.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_14, // @[:@36818.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_15, // @[:@36818.4]
  output         io_memStreams_scatters_0_wresp_ready, // @[:@36818.4]
  input          io_memStreams_scatters_0_wresp_valid, // @[:@36818.4]
  input          io_memStreams_scatters_0_wresp_bits, // @[:@36818.4]
  input          io_axiStreamsIn_0_TVALID, // @[:@36818.4]
  output         io_axiStreamsIn_0_TREADY, // @[:@36818.4]
  input  [255:0] io_axiStreamsIn_0_TDATA, // @[:@36818.4]
  input  [31:0]  io_axiStreamsIn_0_TSTRB, // @[:@36818.4]
  input  [31:0]  io_axiStreamsIn_0_TKEEP, // @[:@36818.4]
  input          io_axiStreamsIn_0_TLAST, // @[:@36818.4]
  input  [7:0]   io_axiStreamsIn_0_TID, // @[:@36818.4]
  input  [7:0]   io_axiStreamsIn_0_TDEST, // @[:@36818.4]
  input  [31:0]  io_axiStreamsIn_0_TUSER, // @[:@36818.4]
  output         io_axiStreamsOut_0_TVALID, // @[:@36818.4]
  input          io_axiStreamsOut_0_TREADY, // @[:@36818.4]
  output [255:0] io_axiStreamsOut_0_TDATA, // @[:@36818.4]
  output [31:0]  io_axiStreamsOut_0_TSTRB, // @[:@36818.4]
  output [31:0]  io_axiStreamsOut_0_TKEEP, // @[:@36818.4]
  output         io_axiStreamsOut_0_TLAST, // @[:@36818.4]
  output [7:0]   io_axiStreamsOut_0_TID, // @[:@36818.4]
  output [7:0]   io_axiStreamsOut_0_TDEST, // @[:@36818.4]
  output [31:0]  io_axiStreamsOut_0_TUSER, // @[:@36818.4]
  output         io_heap_0_req_valid, // @[:@36818.4]
  output         io_heap_0_req_bits_allocDealloc, // @[:@36818.4]
  output [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@36818.4]
  input          io_heap_0_resp_valid, // @[:@36818.4]
  input          io_heap_0_resp_bits_allocDealloc, // @[:@36818.4]
  input  [63:0]  io_heap_0_resp_bits_sizeAddr, // @[:@36818.4]
  input  [63:0]  io_argIns_0, // @[:@36818.4]
  input  [63:0]  io_argIns_1, // @[:@36818.4]
  input          io_argOuts_0_port_ready, // @[:@36818.4]
  output         io_argOuts_0_port_valid, // @[:@36818.4]
  output [63:0]  io_argOuts_0_port_bits, // @[:@36818.4]
  input  [63:0]  io_argOuts_0_echo // @[:@36818.4]
);
  wire  SingleCounter_clock; // @[Main.scala 35:32:@36981.4]
  wire  SingleCounter_reset; // @[Main.scala 35:32:@36981.4]
  wire  SingleCounter_io_input_reset; // @[Main.scala 35:32:@36981.4]
  wire  SingleCounter_io_output_done; // @[Main.scala 35:32:@36981.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@36999.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@36999.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@36999.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@36999.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@36999.4]
  wire  SRFF_clock; // @[Main.scala 39:28:@37008.4]
  wire  SRFF_reset; // @[Main.scala 39:28:@37008.4]
  wire  SRFF_io_input_set; // @[Main.scala 39:28:@37008.4]
  wire  SRFF_io_input_reset; // @[Main.scala 39:28:@37008.4]
  wire  SRFF_io_input_asyn_reset; // @[Main.scala 39:28:@37008.4]
  wire  SRFF_io_output; // @[Main.scala 39:28:@37008.4]
  wire  RootController_sm_clock; // @[sm_RootController.scala 32:18:@37046.4]
  wire  RootController_sm_reset; // @[sm_RootController.scala 32:18:@37046.4]
  wire  RootController_sm_io_enable; // @[sm_RootController.scala 32:18:@37046.4]
  wire  RootController_sm_io_done; // @[sm_RootController.scala 32:18:@37046.4]
  wire  RootController_sm_io_rst; // @[sm_RootController.scala 32:18:@37046.4]
  wire  RootController_sm_io_ctrDone; // @[sm_RootController.scala 32:18:@37046.4]
  wire  RootController_sm_io_ctrInc; // @[sm_RootController.scala 32:18:@37046.4]
  wire  RootController_sm_io_doneIn_0; // @[sm_RootController.scala 32:18:@37046.4]
  wire  RootController_sm_io_enableOut_0; // @[sm_RootController.scala 32:18:@37046.4]
  wire  RootController_sm_io_childAck_0; // @[sm_RootController.scala 32:18:@37046.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@37078.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@37078.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@37078.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@37078.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@37078.4]
  wire  RootController_kernelRootController_concrete1_clock; // @[sm_RootController.scala 73:24:@37137.4]
  wire  RootController_kernelRootController_concrete1_reset; // @[sm_RootController.scala 73:24:@37137.4]
  wire  RootController_kernelRootController_concrete1_io_in_x426_TVALID; // @[sm_RootController.scala 73:24:@37137.4]
  wire  RootController_kernelRootController_concrete1_io_in_x426_TREADY; // @[sm_RootController.scala 73:24:@37137.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x426_TDATA; // @[sm_RootController.scala 73:24:@37137.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x426_TID; // @[sm_RootController.scala 73:24:@37137.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x426_TDEST; // @[sm_RootController.scala 73:24:@37137.4]
  wire  RootController_kernelRootController_concrete1_io_in_x427_TVALID; // @[sm_RootController.scala 73:24:@37137.4]
  wire  RootController_kernelRootController_concrete1_io_in_x427_TREADY; // @[sm_RootController.scala 73:24:@37137.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x427_TDATA; // @[sm_RootController.scala 73:24:@37137.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_RootController.scala 73:24:@37137.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0; // @[sm_RootController.scala 73:24:@37137.4]
  wire  RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[sm_RootController.scala 73:24:@37137.4]
  wire  RootController_kernelRootController_concrete1_io_rr; // @[sm_RootController.scala 73:24:@37137.4]
  wire  _T_599; // @[package.scala 96:25:@37004.4 package.scala 96:25:@37005.4]
  wire  _T_664; // @[Main.scala 41:50:@37074.4]
  wire  _T_665; // @[Main.scala 41:59:@37075.4]
  wire  _T_677; // @[package.scala 100:49:@37095.4]
  reg  _T_680; // @[package.scala 48:56:@37096.4]
  reg [31:0] _RAND_0;
  SingleCounter SingleCounter ( // @[Main.scala 35:32:@36981.4]
    .clock(SingleCounter_clock),
    .reset(SingleCounter_reset),
    .io_input_reset(SingleCounter_io_input_reset),
    .io_output_done(SingleCounter_io_output_done)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@36999.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  SRFF SRFF ( // @[Main.scala 39:28:@37008.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  RootController_sm RootController_sm ( // @[sm_RootController.scala 32:18:@37046.4]
    .clock(RootController_sm_clock),
    .reset(RootController_sm_reset),
    .io_enable(RootController_sm_io_enable),
    .io_done(RootController_sm_io_done),
    .io_rst(RootController_sm_io_rst),
    .io_ctrDone(RootController_sm_io_ctrDone),
    .io_ctrInc(RootController_sm_io_ctrInc),
    .io_doneIn_0(RootController_sm_io_doneIn_0),
    .io_enableOut_0(RootController_sm_io_enableOut_0),
    .io_childAck_0(RootController_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@37078.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RootController_kernelRootController_concrete1 RootController_kernelRootController_concrete1 ( // @[sm_RootController.scala 73:24:@37137.4]
    .clock(RootController_kernelRootController_concrete1_clock),
    .reset(RootController_kernelRootController_concrete1_reset),
    .io_in_x426_TVALID(RootController_kernelRootController_concrete1_io_in_x426_TVALID),
    .io_in_x426_TREADY(RootController_kernelRootController_concrete1_io_in_x426_TREADY),
    .io_in_x426_TDATA(RootController_kernelRootController_concrete1_io_in_x426_TDATA),
    .io_in_x426_TID(RootController_kernelRootController_concrete1_io_in_x426_TID),
    .io_in_x426_TDEST(RootController_kernelRootController_concrete1_io_in_x426_TDEST),
    .io_in_x427_TVALID(RootController_kernelRootController_concrete1_io_in_x427_TVALID),
    .io_in_x427_TREADY(RootController_kernelRootController_concrete1_io_in_x427_TREADY),
    .io_in_x427_TDATA(RootController_kernelRootController_concrete1_io_in_x427_TDATA),
    .io_sigsIn_smEnableOuts_0(RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(RootController_kernelRootController_concrete1_io_rr)
  );
  assign _T_599 = RetimeWrapper_io_out; // @[package.scala 96:25:@37004.4 package.scala 96:25:@37005.4]
  assign _T_664 = io_enable & _T_599; // @[Main.scala 41:50:@37074.4]
  assign _T_665 = ~ SRFF_io_output; // @[Main.scala 41:59:@37075.4]
  assign _T_677 = RootController_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@37095.4]
  assign io_done = SRFF_io_output; // @[Main.scala 48:23:@37094.4]
  assign io_memStreams_loads_0_cmd_valid = 1'h0;
  assign io_memStreams_loads_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_loads_0_cmd_bits_size = 32'h0;
  assign io_memStreams_loads_0_data_ready = 1'h0;
  assign io_memStreams_stores_0_cmd_valid = 1'h0;
  assign io_memStreams_stores_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_stores_0_cmd_bits_size = 32'h0;
  assign io_memStreams_stores_0_data_valid = 1'h0;
  assign io_memStreams_stores_0_data_bits_wdata_0 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_1 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_2 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_3 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_4 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_5 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_6 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_7 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_8 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_9 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_10 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_11 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_12 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_13 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_14 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_15 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wstrb = 16'h0;
  assign io_memStreams_stores_0_wresp_ready = 1'h0;
  assign io_memStreams_gathers_0_cmd_valid = 1'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_0 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_1 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_2 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_3 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_4 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_5 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_6 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_7 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_8 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_9 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_10 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_11 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_12 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_13 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_14 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_15 = 64'h0;
  assign io_memStreams_gathers_0_data_ready = 1'h0;
  assign io_memStreams_scatters_0_cmd_valid = 1'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_0 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_1 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_2 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_3 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_4 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_5 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_6 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_7 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_8 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_9 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_10 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_11 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_12 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_13 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_14 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_15 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_0 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_1 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_2 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_3 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_4 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_5 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_6 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_7 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_8 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_9 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_10 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_11 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_12 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_13 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_14 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_15 = 32'h0;
  assign io_memStreams_scatters_0_wresp_ready = 1'h0;
  assign io_axiStreamsIn_0_TREADY = RootController_kernelRootController_concrete1_io_in_x426_TREADY; // @[sm_RootController.scala 48:23:@37192.4]
  assign io_axiStreamsOut_0_TVALID = RootController_kernelRootController_concrete1_io_in_x427_TVALID; // @[sm_RootController.scala 49:23:@37202.4]
  assign io_axiStreamsOut_0_TDATA = RootController_kernelRootController_concrete1_io_in_x427_TDATA; // @[sm_RootController.scala 49:23:@37200.4]
  assign io_axiStreamsOut_0_TSTRB = 32'hffffffff; // @[sm_RootController.scala 49:23:@37199.4]
  assign io_axiStreamsOut_0_TKEEP = 32'hffffffff; // @[sm_RootController.scala 49:23:@37198.4]
  assign io_axiStreamsOut_0_TLAST = 1'h0; // @[sm_RootController.scala 49:23:@37197.4]
  assign io_axiStreamsOut_0_TID = 8'h0; // @[sm_RootController.scala 49:23:@37196.4]
  assign io_axiStreamsOut_0_TDEST = 8'h0; // @[sm_RootController.scala 49:23:@37195.4]
  assign io_axiStreamsOut_0_TUSER = 32'h4; // @[sm_RootController.scala 49:23:@37194.4]
  assign io_heap_0_req_valid = 1'h0;
  assign io_heap_0_req_bits_allocDealloc = 1'h0;
  assign io_heap_0_req_bits_sizeAddr = 64'h0;
  assign io_argOuts_0_port_valid = 1'h0;
  assign io_argOuts_0_port_bits = 64'h0;
  assign SingleCounter_clock = clock; // @[:@36982.4]
  assign SingleCounter_reset = reset; // @[:@36983.4]
  assign SingleCounter_io_input_reset = reset; // @[Main.scala 36:79:@36997.4]
  assign RetimeWrapper_clock = clock; // @[:@37000.4]
  assign RetimeWrapper_reset = reset; // @[:@37001.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@37003.4]
  assign RetimeWrapper_io_in = SingleCounter_io_output_done; // @[package.scala 94:16:@37002.4]
  assign SRFF_clock = clock; // @[:@37009.4]
  assign SRFF_reset = reset; // @[:@37010.4]
  assign SRFF_io_input_set = RootController_sm_io_done; // @[Main.scala 57:29:@37229.4]
  assign SRFF_io_input_reset = RetimeWrapper_1_io_out; // @[Main.scala 46:31:@37092.4]
  assign SRFF_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[Main.scala 47:36:@37093.4]
  assign RootController_sm_clock = clock; // @[:@37047.4]
  assign RootController_sm_reset = reset; // @[:@37048.4]
  assign RootController_sm_io_enable = _T_664 & _T_665; // @[Main.scala 45:33:@37091.4 SpatialBlocks.scala 112:18:@37125.4]
  assign RootController_sm_io_rst = RetimeWrapper_1_io_out; // @[SpatialBlocks.scala 106:15:@37119.4]
  assign RootController_sm_io_ctrDone = RootController_sm_io_ctrInc & _T_680; // @[Main.scala 49:34:@37099.4]
  assign RootController_sm_io_doneIn_0 = RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 102:67:@37116.4]
  assign RetimeWrapper_1_clock = clock; // @[:@37079.4]
  assign RetimeWrapper_1_reset = reset; // @[:@37080.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@37082.4]
  assign RetimeWrapper_1_io_in = reset | io_reset; // @[package.scala 94:16:@37081.4]
  assign RootController_kernelRootController_concrete1_clock = clock; // @[:@37138.4]
  assign RootController_kernelRootController_concrete1_reset = reset; // @[:@37139.4]
  assign RootController_kernelRootController_concrete1_io_in_x426_TVALID = io_axiStreamsIn_0_TVALID; // @[sm_RootController.scala 48:23:@37193.4]
  assign RootController_kernelRootController_concrete1_io_in_x426_TDATA = io_axiStreamsIn_0_TDATA; // @[sm_RootController.scala 48:23:@37191.4]
  assign RootController_kernelRootController_concrete1_io_in_x426_TID = io_axiStreamsIn_0_TID; // @[sm_RootController.scala 48:23:@37187.4]
  assign RootController_kernelRootController_concrete1_io_in_x426_TDEST = io_axiStreamsIn_0_TDEST; // @[sm_RootController.scala 48:23:@37186.4]
  assign RootController_kernelRootController_concrete1_io_in_x427_TREADY = io_axiStreamsOut_0_TREADY; // @[sm_RootController.scala 49:23:@37201.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0 = RootController_sm_io_enableOut_0; // @[sm_RootController.scala 77:22:@37211.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0 = RootController_sm_io_childAck_0; // @[sm_RootController.scala 77:22:@37209.4]
  assign RootController_kernelRootController_concrete1_io_rr = RetimeWrapper_io_out; // @[sm_RootController.scala 76:18:@37203.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_680 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_680 <= 1'h0;
    end else begin
      _T_680 <= _T_677;
    end
  end
endmodule
module SpatialIP( // @[:@37231.2]
  input         clock, // @[:@37232.4]
  input         reset, // @[:@37233.4]
  input  [31:0] io_raddr, // @[:@37234.4]
  input         io_wen, // @[:@37234.4]
  input  [31:0] io_waddr, // @[:@37234.4]
  input  [63:0] io_wdata, // @[:@37234.4]
  output [63:0] io_rdata // @[:@37234.4]
);
  wire  accel_clock; // @[Instantiator.scala 53:44:@37236.4]
  wire  accel_reset; // @[Instantiator.scala 53:44:@37236.4]
  wire  accel_io_enable; // @[Instantiator.scala 53:44:@37236.4]
  wire  accel_io_done; // @[Instantiator.scala 53:44:@37236.4]
  wire  accel_io_reset; // @[Instantiator.scala 53:44:@37236.4]
  wire  accel_io_memStreams_loads_0_cmd_ready; // @[Instantiator.scala 53:44:@37236.4]
  wire  accel_io_memStreams_loads_0_cmd_valid; // @[Instantiator.scala 53:44:@37236.4]
  wire [63:0] accel_io_memStreams_loads_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_loads_0_cmd_bits_size; // @[Instantiator.scala 53:44:@37236.4]
  wire  accel_io_memStreams_loads_0_data_ready; // @[Instantiator.scala 53:44:@37236.4]
  wire  accel_io_memStreams_loads_0_data_valid; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_0; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_1; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_2; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_3; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_4; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_5; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_6; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_7; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_8; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_9; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_10; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_11; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_12; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_13; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_14; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_15; // @[Instantiator.scala 53:44:@37236.4]
  wire  accel_io_memStreams_stores_0_cmd_ready; // @[Instantiator.scala 53:44:@37236.4]
  wire  accel_io_memStreams_stores_0_cmd_valid; // @[Instantiator.scala 53:44:@37236.4]
  wire [63:0] accel_io_memStreams_stores_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_stores_0_cmd_bits_size; // @[Instantiator.scala 53:44:@37236.4]
  wire  accel_io_memStreams_stores_0_data_ready; // @[Instantiator.scala 53:44:@37236.4]
  wire  accel_io_memStreams_stores_0_data_valid; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_1; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_2; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_3; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_4; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_5; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_6; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_7; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_8; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_9; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_10; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_11; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_12; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_13; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_14; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_15; // @[Instantiator.scala 53:44:@37236.4]
  wire [15:0] accel_io_memStreams_stores_0_data_bits_wstrb; // @[Instantiator.scala 53:44:@37236.4]
  wire  accel_io_memStreams_stores_0_wresp_ready; // @[Instantiator.scala 53:44:@37236.4]
  wire  accel_io_memStreams_stores_0_wresp_valid; // @[Instantiator.scala 53:44:@37236.4]
  wire  accel_io_memStreams_stores_0_wresp_bits; // @[Instantiator.scala 53:44:@37236.4]
  wire  accel_io_memStreams_gathers_0_cmd_ready; // @[Instantiator.scala 53:44:@37236.4]
  wire  accel_io_memStreams_gathers_0_cmd_valid; // @[Instantiator.scala 53:44:@37236.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_0; // @[Instantiator.scala 53:44:@37236.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_1; // @[Instantiator.scala 53:44:@37236.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_2; // @[Instantiator.scala 53:44:@37236.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_3; // @[Instantiator.scala 53:44:@37236.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_4; // @[Instantiator.scala 53:44:@37236.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_5; // @[Instantiator.scala 53:44:@37236.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_6; // @[Instantiator.scala 53:44:@37236.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_7; // @[Instantiator.scala 53:44:@37236.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_8; // @[Instantiator.scala 53:44:@37236.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_9; // @[Instantiator.scala 53:44:@37236.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_10; // @[Instantiator.scala 53:44:@37236.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_11; // @[Instantiator.scala 53:44:@37236.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_12; // @[Instantiator.scala 53:44:@37236.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_13; // @[Instantiator.scala 53:44:@37236.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_14; // @[Instantiator.scala 53:44:@37236.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_15; // @[Instantiator.scala 53:44:@37236.4]
  wire  accel_io_memStreams_gathers_0_data_ready; // @[Instantiator.scala 53:44:@37236.4]
  wire  accel_io_memStreams_gathers_0_data_valid; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_0; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_1; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_2; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_3; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_4; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_5; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_6; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_7; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_8; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_9; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_10; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_11; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_12; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_13; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_14; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_15; // @[Instantiator.scala 53:44:@37236.4]
  wire  accel_io_memStreams_scatters_0_cmd_ready; // @[Instantiator.scala 53:44:@37236.4]
  wire  accel_io_memStreams_scatters_0_cmd_valid; // @[Instantiator.scala 53:44:@37236.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0; // @[Instantiator.scala 53:44:@37236.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1; // @[Instantiator.scala 53:44:@37236.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2; // @[Instantiator.scala 53:44:@37236.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3; // @[Instantiator.scala 53:44:@37236.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4; // @[Instantiator.scala 53:44:@37236.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5; // @[Instantiator.scala 53:44:@37236.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6; // @[Instantiator.scala 53:44:@37236.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7; // @[Instantiator.scala 53:44:@37236.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8; // @[Instantiator.scala 53:44:@37236.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9; // @[Instantiator.scala 53:44:@37236.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10; // @[Instantiator.scala 53:44:@37236.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11; // @[Instantiator.scala 53:44:@37236.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12; // @[Instantiator.scala 53:44:@37236.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13; // @[Instantiator.scala 53:44:@37236.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14; // @[Instantiator.scala 53:44:@37236.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_0; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_1; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_2; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_3; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_4; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_5; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_6; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_7; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_8; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_9; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_10; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_11; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_12; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_13; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_14; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_15; // @[Instantiator.scala 53:44:@37236.4]
  wire  accel_io_memStreams_scatters_0_wresp_ready; // @[Instantiator.scala 53:44:@37236.4]
  wire  accel_io_memStreams_scatters_0_wresp_valid; // @[Instantiator.scala 53:44:@37236.4]
  wire  accel_io_memStreams_scatters_0_wresp_bits; // @[Instantiator.scala 53:44:@37236.4]
  wire  accel_io_axiStreamsIn_0_TVALID; // @[Instantiator.scala 53:44:@37236.4]
  wire  accel_io_axiStreamsIn_0_TREADY; // @[Instantiator.scala 53:44:@37236.4]
  wire [255:0] accel_io_axiStreamsIn_0_TDATA; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_axiStreamsIn_0_TSTRB; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_axiStreamsIn_0_TKEEP; // @[Instantiator.scala 53:44:@37236.4]
  wire  accel_io_axiStreamsIn_0_TLAST; // @[Instantiator.scala 53:44:@37236.4]
  wire [7:0] accel_io_axiStreamsIn_0_TID; // @[Instantiator.scala 53:44:@37236.4]
  wire [7:0] accel_io_axiStreamsIn_0_TDEST; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_axiStreamsIn_0_TUSER; // @[Instantiator.scala 53:44:@37236.4]
  wire  accel_io_axiStreamsOut_0_TVALID; // @[Instantiator.scala 53:44:@37236.4]
  wire  accel_io_axiStreamsOut_0_TREADY; // @[Instantiator.scala 53:44:@37236.4]
  wire [255:0] accel_io_axiStreamsOut_0_TDATA; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_axiStreamsOut_0_TSTRB; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_axiStreamsOut_0_TKEEP; // @[Instantiator.scala 53:44:@37236.4]
  wire  accel_io_axiStreamsOut_0_TLAST; // @[Instantiator.scala 53:44:@37236.4]
  wire [7:0] accel_io_axiStreamsOut_0_TID; // @[Instantiator.scala 53:44:@37236.4]
  wire [7:0] accel_io_axiStreamsOut_0_TDEST; // @[Instantiator.scala 53:44:@37236.4]
  wire [31:0] accel_io_axiStreamsOut_0_TUSER; // @[Instantiator.scala 53:44:@37236.4]
  wire  accel_io_heap_0_req_valid; // @[Instantiator.scala 53:44:@37236.4]
  wire  accel_io_heap_0_req_bits_allocDealloc; // @[Instantiator.scala 53:44:@37236.4]
  wire [63:0] accel_io_heap_0_req_bits_sizeAddr; // @[Instantiator.scala 53:44:@37236.4]
  wire  accel_io_heap_0_resp_valid; // @[Instantiator.scala 53:44:@37236.4]
  wire  accel_io_heap_0_resp_bits_allocDealloc; // @[Instantiator.scala 53:44:@37236.4]
  wire [63:0] accel_io_heap_0_resp_bits_sizeAddr; // @[Instantiator.scala 53:44:@37236.4]
  wire [63:0] accel_io_argIns_0; // @[Instantiator.scala 53:44:@37236.4]
  wire [63:0] accel_io_argIns_1; // @[Instantiator.scala 53:44:@37236.4]
  wire  accel_io_argOuts_0_port_ready; // @[Instantiator.scala 53:44:@37236.4]
  wire  accel_io_argOuts_0_port_valid; // @[Instantiator.scala 53:44:@37236.4]
  wire [63:0] accel_io_argOuts_0_port_bits; // @[Instantiator.scala 53:44:@37236.4]
  wire [63:0] accel_io_argOuts_0_echo; // @[Instantiator.scala 53:44:@37236.4]
  AccelUnit accel ( // @[Instantiator.scala 53:44:@37236.4]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_enable(accel_io_enable),
    .io_done(accel_io_done),
    .io_reset(accel_io_reset),
    .io_memStreams_loads_0_cmd_ready(accel_io_memStreams_loads_0_cmd_ready),
    .io_memStreams_loads_0_cmd_valid(accel_io_memStreams_loads_0_cmd_valid),
    .io_memStreams_loads_0_cmd_bits_addr(accel_io_memStreams_loads_0_cmd_bits_addr),
    .io_memStreams_loads_0_cmd_bits_size(accel_io_memStreams_loads_0_cmd_bits_size),
    .io_memStreams_loads_0_data_ready(accel_io_memStreams_loads_0_data_ready),
    .io_memStreams_loads_0_data_valid(accel_io_memStreams_loads_0_data_valid),
    .io_memStreams_loads_0_data_bits_rdata_0(accel_io_memStreams_loads_0_data_bits_rdata_0),
    .io_memStreams_loads_0_data_bits_rdata_1(accel_io_memStreams_loads_0_data_bits_rdata_1),
    .io_memStreams_loads_0_data_bits_rdata_2(accel_io_memStreams_loads_0_data_bits_rdata_2),
    .io_memStreams_loads_0_data_bits_rdata_3(accel_io_memStreams_loads_0_data_bits_rdata_3),
    .io_memStreams_loads_0_data_bits_rdata_4(accel_io_memStreams_loads_0_data_bits_rdata_4),
    .io_memStreams_loads_0_data_bits_rdata_5(accel_io_memStreams_loads_0_data_bits_rdata_5),
    .io_memStreams_loads_0_data_bits_rdata_6(accel_io_memStreams_loads_0_data_bits_rdata_6),
    .io_memStreams_loads_0_data_bits_rdata_7(accel_io_memStreams_loads_0_data_bits_rdata_7),
    .io_memStreams_loads_0_data_bits_rdata_8(accel_io_memStreams_loads_0_data_bits_rdata_8),
    .io_memStreams_loads_0_data_bits_rdata_9(accel_io_memStreams_loads_0_data_bits_rdata_9),
    .io_memStreams_loads_0_data_bits_rdata_10(accel_io_memStreams_loads_0_data_bits_rdata_10),
    .io_memStreams_loads_0_data_bits_rdata_11(accel_io_memStreams_loads_0_data_bits_rdata_11),
    .io_memStreams_loads_0_data_bits_rdata_12(accel_io_memStreams_loads_0_data_bits_rdata_12),
    .io_memStreams_loads_0_data_bits_rdata_13(accel_io_memStreams_loads_0_data_bits_rdata_13),
    .io_memStreams_loads_0_data_bits_rdata_14(accel_io_memStreams_loads_0_data_bits_rdata_14),
    .io_memStreams_loads_0_data_bits_rdata_15(accel_io_memStreams_loads_0_data_bits_rdata_15),
    .io_memStreams_stores_0_cmd_ready(accel_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(accel_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(accel_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(accel_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(accel_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(accel_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(accel_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wdata_1(accel_io_memStreams_stores_0_data_bits_wdata_1),
    .io_memStreams_stores_0_data_bits_wdata_2(accel_io_memStreams_stores_0_data_bits_wdata_2),
    .io_memStreams_stores_0_data_bits_wdata_3(accel_io_memStreams_stores_0_data_bits_wdata_3),
    .io_memStreams_stores_0_data_bits_wdata_4(accel_io_memStreams_stores_0_data_bits_wdata_4),
    .io_memStreams_stores_0_data_bits_wdata_5(accel_io_memStreams_stores_0_data_bits_wdata_5),
    .io_memStreams_stores_0_data_bits_wdata_6(accel_io_memStreams_stores_0_data_bits_wdata_6),
    .io_memStreams_stores_0_data_bits_wdata_7(accel_io_memStreams_stores_0_data_bits_wdata_7),
    .io_memStreams_stores_0_data_bits_wdata_8(accel_io_memStreams_stores_0_data_bits_wdata_8),
    .io_memStreams_stores_0_data_bits_wdata_9(accel_io_memStreams_stores_0_data_bits_wdata_9),
    .io_memStreams_stores_0_data_bits_wdata_10(accel_io_memStreams_stores_0_data_bits_wdata_10),
    .io_memStreams_stores_0_data_bits_wdata_11(accel_io_memStreams_stores_0_data_bits_wdata_11),
    .io_memStreams_stores_0_data_bits_wdata_12(accel_io_memStreams_stores_0_data_bits_wdata_12),
    .io_memStreams_stores_0_data_bits_wdata_13(accel_io_memStreams_stores_0_data_bits_wdata_13),
    .io_memStreams_stores_0_data_bits_wdata_14(accel_io_memStreams_stores_0_data_bits_wdata_14),
    .io_memStreams_stores_0_data_bits_wdata_15(accel_io_memStreams_stores_0_data_bits_wdata_15),
    .io_memStreams_stores_0_data_bits_wstrb(accel_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(accel_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(accel_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(accel_io_memStreams_stores_0_wresp_bits),
    .io_memStreams_gathers_0_cmd_ready(accel_io_memStreams_gathers_0_cmd_ready),
    .io_memStreams_gathers_0_cmd_valid(accel_io_memStreams_gathers_0_cmd_valid),
    .io_memStreams_gathers_0_cmd_bits_addr_0(accel_io_memStreams_gathers_0_cmd_bits_addr_0),
    .io_memStreams_gathers_0_cmd_bits_addr_1(accel_io_memStreams_gathers_0_cmd_bits_addr_1),
    .io_memStreams_gathers_0_cmd_bits_addr_2(accel_io_memStreams_gathers_0_cmd_bits_addr_2),
    .io_memStreams_gathers_0_cmd_bits_addr_3(accel_io_memStreams_gathers_0_cmd_bits_addr_3),
    .io_memStreams_gathers_0_cmd_bits_addr_4(accel_io_memStreams_gathers_0_cmd_bits_addr_4),
    .io_memStreams_gathers_0_cmd_bits_addr_5(accel_io_memStreams_gathers_0_cmd_bits_addr_5),
    .io_memStreams_gathers_0_cmd_bits_addr_6(accel_io_memStreams_gathers_0_cmd_bits_addr_6),
    .io_memStreams_gathers_0_cmd_bits_addr_7(accel_io_memStreams_gathers_0_cmd_bits_addr_7),
    .io_memStreams_gathers_0_cmd_bits_addr_8(accel_io_memStreams_gathers_0_cmd_bits_addr_8),
    .io_memStreams_gathers_0_cmd_bits_addr_9(accel_io_memStreams_gathers_0_cmd_bits_addr_9),
    .io_memStreams_gathers_0_cmd_bits_addr_10(accel_io_memStreams_gathers_0_cmd_bits_addr_10),
    .io_memStreams_gathers_0_cmd_bits_addr_11(accel_io_memStreams_gathers_0_cmd_bits_addr_11),
    .io_memStreams_gathers_0_cmd_bits_addr_12(accel_io_memStreams_gathers_0_cmd_bits_addr_12),
    .io_memStreams_gathers_0_cmd_bits_addr_13(accel_io_memStreams_gathers_0_cmd_bits_addr_13),
    .io_memStreams_gathers_0_cmd_bits_addr_14(accel_io_memStreams_gathers_0_cmd_bits_addr_14),
    .io_memStreams_gathers_0_cmd_bits_addr_15(accel_io_memStreams_gathers_0_cmd_bits_addr_15),
    .io_memStreams_gathers_0_data_ready(accel_io_memStreams_gathers_0_data_ready),
    .io_memStreams_gathers_0_data_valid(accel_io_memStreams_gathers_0_data_valid),
    .io_memStreams_gathers_0_data_bits_0(accel_io_memStreams_gathers_0_data_bits_0),
    .io_memStreams_gathers_0_data_bits_1(accel_io_memStreams_gathers_0_data_bits_1),
    .io_memStreams_gathers_0_data_bits_2(accel_io_memStreams_gathers_0_data_bits_2),
    .io_memStreams_gathers_0_data_bits_3(accel_io_memStreams_gathers_0_data_bits_3),
    .io_memStreams_gathers_0_data_bits_4(accel_io_memStreams_gathers_0_data_bits_4),
    .io_memStreams_gathers_0_data_bits_5(accel_io_memStreams_gathers_0_data_bits_5),
    .io_memStreams_gathers_0_data_bits_6(accel_io_memStreams_gathers_0_data_bits_6),
    .io_memStreams_gathers_0_data_bits_7(accel_io_memStreams_gathers_0_data_bits_7),
    .io_memStreams_gathers_0_data_bits_8(accel_io_memStreams_gathers_0_data_bits_8),
    .io_memStreams_gathers_0_data_bits_9(accel_io_memStreams_gathers_0_data_bits_9),
    .io_memStreams_gathers_0_data_bits_10(accel_io_memStreams_gathers_0_data_bits_10),
    .io_memStreams_gathers_0_data_bits_11(accel_io_memStreams_gathers_0_data_bits_11),
    .io_memStreams_gathers_0_data_bits_12(accel_io_memStreams_gathers_0_data_bits_12),
    .io_memStreams_gathers_0_data_bits_13(accel_io_memStreams_gathers_0_data_bits_13),
    .io_memStreams_gathers_0_data_bits_14(accel_io_memStreams_gathers_0_data_bits_14),
    .io_memStreams_gathers_0_data_bits_15(accel_io_memStreams_gathers_0_data_bits_15),
    .io_memStreams_scatters_0_cmd_ready(accel_io_memStreams_scatters_0_cmd_ready),
    .io_memStreams_scatters_0_cmd_valid(accel_io_memStreams_scatters_0_cmd_valid),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_0(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_1(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_2(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_3(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_4(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_5(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_6(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_7(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_8(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_9(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_10(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_11(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_12(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_13(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_14(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_15(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15),
    .io_memStreams_scatters_0_cmd_bits_wdata_0(accel_io_memStreams_scatters_0_cmd_bits_wdata_0),
    .io_memStreams_scatters_0_cmd_bits_wdata_1(accel_io_memStreams_scatters_0_cmd_bits_wdata_1),
    .io_memStreams_scatters_0_cmd_bits_wdata_2(accel_io_memStreams_scatters_0_cmd_bits_wdata_2),
    .io_memStreams_scatters_0_cmd_bits_wdata_3(accel_io_memStreams_scatters_0_cmd_bits_wdata_3),
    .io_memStreams_scatters_0_cmd_bits_wdata_4(accel_io_memStreams_scatters_0_cmd_bits_wdata_4),
    .io_memStreams_scatters_0_cmd_bits_wdata_5(accel_io_memStreams_scatters_0_cmd_bits_wdata_5),
    .io_memStreams_scatters_0_cmd_bits_wdata_6(accel_io_memStreams_scatters_0_cmd_bits_wdata_6),
    .io_memStreams_scatters_0_cmd_bits_wdata_7(accel_io_memStreams_scatters_0_cmd_bits_wdata_7),
    .io_memStreams_scatters_0_cmd_bits_wdata_8(accel_io_memStreams_scatters_0_cmd_bits_wdata_8),
    .io_memStreams_scatters_0_cmd_bits_wdata_9(accel_io_memStreams_scatters_0_cmd_bits_wdata_9),
    .io_memStreams_scatters_0_cmd_bits_wdata_10(accel_io_memStreams_scatters_0_cmd_bits_wdata_10),
    .io_memStreams_scatters_0_cmd_bits_wdata_11(accel_io_memStreams_scatters_0_cmd_bits_wdata_11),
    .io_memStreams_scatters_0_cmd_bits_wdata_12(accel_io_memStreams_scatters_0_cmd_bits_wdata_12),
    .io_memStreams_scatters_0_cmd_bits_wdata_13(accel_io_memStreams_scatters_0_cmd_bits_wdata_13),
    .io_memStreams_scatters_0_cmd_bits_wdata_14(accel_io_memStreams_scatters_0_cmd_bits_wdata_14),
    .io_memStreams_scatters_0_cmd_bits_wdata_15(accel_io_memStreams_scatters_0_cmd_bits_wdata_15),
    .io_memStreams_scatters_0_wresp_ready(accel_io_memStreams_scatters_0_wresp_ready),
    .io_memStreams_scatters_0_wresp_valid(accel_io_memStreams_scatters_0_wresp_valid),
    .io_memStreams_scatters_0_wresp_bits(accel_io_memStreams_scatters_0_wresp_bits),
    .io_axiStreamsIn_0_TVALID(accel_io_axiStreamsIn_0_TVALID),
    .io_axiStreamsIn_0_TREADY(accel_io_axiStreamsIn_0_TREADY),
    .io_axiStreamsIn_0_TDATA(accel_io_axiStreamsIn_0_TDATA),
    .io_axiStreamsIn_0_TSTRB(accel_io_axiStreamsIn_0_TSTRB),
    .io_axiStreamsIn_0_TKEEP(accel_io_axiStreamsIn_0_TKEEP),
    .io_axiStreamsIn_0_TLAST(accel_io_axiStreamsIn_0_TLAST),
    .io_axiStreamsIn_0_TID(accel_io_axiStreamsIn_0_TID),
    .io_axiStreamsIn_0_TDEST(accel_io_axiStreamsIn_0_TDEST),
    .io_axiStreamsIn_0_TUSER(accel_io_axiStreamsIn_0_TUSER),
    .io_axiStreamsOut_0_TVALID(accel_io_axiStreamsOut_0_TVALID),
    .io_axiStreamsOut_0_TREADY(accel_io_axiStreamsOut_0_TREADY),
    .io_axiStreamsOut_0_TDATA(accel_io_axiStreamsOut_0_TDATA),
    .io_axiStreamsOut_0_TSTRB(accel_io_axiStreamsOut_0_TSTRB),
    .io_axiStreamsOut_0_TKEEP(accel_io_axiStreamsOut_0_TKEEP),
    .io_axiStreamsOut_0_TLAST(accel_io_axiStreamsOut_0_TLAST),
    .io_axiStreamsOut_0_TID(accel_io_axiStreamsOut_0_TID),
    .io_axiStreamsOut_0_TDEST(accel_io_axiStreamsOut_0_TDEST),
    .io_axiStreamsOut_0_TUSER(accel_io_axiStreamsOut_0_TUSER),
    .io_heap_0_req_valid(accel_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(accel_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(accel_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(accel_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(accel_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(accel_io_heap_0_resp_bits_sizeAddr),
    .io_argIns_0(accel_io_argIns_0),
    .io_argIns_1(accel_io_argIns_1),
    .io_argOuts_0_port_ready(accel_io_argOuts_0_port_ready),
    .io_argOuts_0_port_valid(accel_io_argOuts_0_port_valid),
    .io_argOuts_0_port_bits(accel_io_argOuts_0_port_bits),
    .io_argOuts_0_echo(accel_io_argOuts_0_echo)
  );
  assign io_rdata = 64'h0;
  assign accel_clock = clock; // @[:@37237.4]
  assign accel_reset = reset; // @[:@37238.4]
  assign accel_io_enable = 1'h0;
  assign accel_io_reset = 1'h0;
  assign accel_io_memStreams_loads_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_loads_0_data_valid = 1'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_0 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_1 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_2 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_3 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_4 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_5 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_6 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_7 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_8 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_9 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_10 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_11 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_12 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_13 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_14 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_15 = 32'h0;
  assign accel_io_memStreams_stores_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_stores_0_data_ready = 1'h0;
  assign accel_io_memStreams_stores_0_wresp_valid = 1'h0;
  assign accel_io_memStreams_stores_0_wresp_bits = 1'h0;
  assign accel_io_memStreams_gathers_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_gathers_0_data_valid = 1'h0;
  assign accel_io_memStreams_gathers_0_data_bits_0 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_1 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_2 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_3 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_4 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_5 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_6 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_7 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_8 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_9 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_10 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_11 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_12 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_13 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_14 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_15 = 32'h0;
  assign accel_io_memStreams_scatters_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_scatters_0_wresp_valid = 1'h0;
  assign accel_io_memStreams_scatters_0_wresp_bits = 1'h0;
  assign accel_io_axiStreamsIn_0_TVALID = 1'h0;
  assign accel_io_axiStreamsIn_0_TDATA = 256'h0;
  assign accel_io_axiStreamsIn_0_TSTRB = 32'h0;
  assign accel_io_axiStreamsIn_0_TKEEP = 32'h0;
  assign accel_io_axiStreamsIn_0_TLAST = 1'h0;
  assign accel_io_axiStreamsIn_0_TID = 8'h0;
  assign accel_io_axiStreamsIn_0_TDEST = 8'h0;
  assign accel_io_axiStreamsIn_0_TUSER = 32'h0;
  assign accel_io_axiStreamsOut_0_TREADY = 1'h0;
  assign accel_io_heap_0_resp_valid = 1'h0;
  assign accel_io_heap_0_resp_bits_allocDealloc = 1'h0;
  assign accel_io_heap_0_resp_bits_sizeAddr = 64'h0;
  assign accel_io_argIns_0 = 64'h0;
  assign accel_io_argIns_1 = 64'h0;
  assign accel_io_argOuts_0_port_ready = 1'h0;
  assign accel_io_argOuts_0_echo = 64'h0;
endmodule
