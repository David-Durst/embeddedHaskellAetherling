// Latency = 4
module top(
  input CLK/*verilator public*/, 
  input [7:0] I/*verilator public*/, 
  output [7:0] O/*verilator public*/, 
  output valid_down/*verilator public*/, 
  input valid_up/*verilator public*/
);
  wire dontcare;
  wire [31:0] io_output_counts_1;
  wire [31:0] io_output_counts_0;

  x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1 sampler_box ( // @[m_x55_ctr_0.scala 26:17:@1721.4]
    .clock(CLK), // @[:@1296.4]
    .reset('b0), // @[:@1297.4]
    .io_in_x270_TREADY(dontcare), // @[:@1298.4]
    .io_in_x270_TDATA(I), // @[:@1298.4]
    .io_in_x270_TID(8'h0),
    .io_in_x270_TDEST(8'h0),
    .io_in_x271_TVALID(valid_down), // @[:@1298.4]
    .io_in_x271_TDATA(O), // @[:@1298.4]
    .io_in_x271_TREADY(1'b1), // @[:@1298.4]
    .io_sigsIn_datapathEn(valid_up), // @[:@1298.4]
    .io_sigsIn_backpressure(1'b0), // @[:@20563.4]
    .io_sigsIn_break(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_1(io_output_counts_1), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_0(io_output_counts_0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_0(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_1(1'b0), // @[:@20563.4]
    .io_rr('b1) // @[:@1298.4]
  );

  wire dontcare2;

  wire io_output_oobs_0;
  wire io_output_oobs_1;
  x278_ctrchain cchain ( // @[:@2879.2]
    .clock(CLK), // @[:@2880.4]
    .reset(1'b0), // @[:@2881.4]
    .io_input_reset(1'b0), // @[:@2882.4]
    .io_input_enable(valid_up), // @[:@2882.4]
    .io_output_counts_1(io_output_counts_1), // @[:@2882.4]
    .io_output_counts_0(io_output_counts_0), // @[:@2882.4]
    .io_output_oobs_0(io_output_oobs_0), // @[:@2882.4]
    .io_output_oobs_1(io_output_oobs_1), // @[:@2882.4]
    .io_output_done(dontcare2) // @[:@2882.4]
  );

endmodule

module RetimeShiftRegister
#(
    parameter WIDTH = 1,
    parameter STAGES = 1)
(
    input clock,
    input reset,
    input flow,
    input [WIDTH-1:0] init,
    input [WIDTH-1:0] in,
    output reg [WIDTH-1:0] out
);
  integer i;
  reg [WIDTH-1:0] sr[STAGES:0]; // Create 'STAGES' number of register, each 'WIDTH' bits wide

   /* synopsys dc_tcl_script_begin
    set_ungroup [current_design] true
    set_flatten true -effort high -phase true -design [current_design]
    set_dont_retime [current_design] false
    set_optimize_registers true -design [current_design]
    */
  always @(posedge clock) begin
    if (reset) begin
      for(i=0; i<STAGES; i=i+1) begin
        sr[i] <= init;
      end
    end else begin
      if (flow) begin 
        sr[0] <= in;
        for(i=1; i<STAGES; i=i+1) begin
          sr[i] <= sr[i-1];
        end
      end
    end
  end

  always @(*) begin
    out = sr[STAGES-1];
  end
endmodule
module FF( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  output [31:0] io_rPort_0_output_0, // @[:@6.4]
  input  [31:0] io_wPort_0_data_0, // @[:@6.4]
  input         io_wPort_0_reset, // @[:@6.4]
  input  [31:0] io_wPort_0_init, // @[:@6.4]
  input         io_wPort_0_en_0, // @[:@6.4]
  input         io_reset // @[:@6.4]
);
  reg [31:0] ff; // @[MemPrimitives.scala 173:19:@21.4]
  reg [31:0] _RAND_0;
  wire  anyReset; // @[MemPrimitives.scala 174:65:@22.4]
  wire [31:0] _T_68; // @[MemPrimitives.scala 177:32:@23.4]
  wire [31:0] _T_69; // @[MemPrimitives.scala 177:12:@24.4]
  assign anyReset = io_wPort_0_reset | io_reset; // @[MemPrimitives.scala 174:65:@22.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 177:32:@23.4]
  assign _T_69 = anyReset ? io_wPort_0_init : _T_68; // @[MemPrimitives.scala 177:12:@24.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 178:34:@26.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= io_wPort_0_init;
    end else begin
      if (anyReset) begin
        ff <= io_wPort_0_init;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SRFF( // @[:@28.2]
  input   clock, // @[:@29.4]
  input   reset, // @[:@30.4]
  input   io_input_set, // @[:@31.4]
  input   io_input_reset, // @[:@31.4]
  input   io_input_asyn_reset, // @[:@31.4]
  output  io_output // @[:@31.4]
);
  reg  _T_15; // @[SRFF.scala 20:21:@33.4]
  reg [31:0] _RAND_0;
  wire  _T_19; // @[SRFF.scala 21:74:@34.4]
  wire  _T_20; // @[SRFF.scala 21:48:@35.4]
  wire  _T_21; // @[SRFF.scala 21:14:@36.4]
  assign _T_19 = io_input_reset ? 1'h0 : _T_15; // @[SRFF.scala 21:74:@34.4]
  assign _T_20 = io_input_set ? 1'h1 : _T_19; // @[SRFF.scala 21:48:@35.4]
  assign _T_21 = io_input_asyn_reset ? 1'h0 : _T_20; // @[SRFF.scala 21:14:@36.4]
  assign io_output = io_input_asyn_reset ? 1'h0 : _T_15; // @[SRFF.scala 22:15:@39.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_15 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_15 <= 1'h0;
    end else begin
      if (io_input_asyn_reset) begin
        _T_15 <= 1'h0;
      end else begin
        if (io_input_set) begin
          _T_15 <= 1'h1;
        end else begin
          if (io_input_reset) begin
            _T_15 <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module SingleCounter( // @[:@41.2]
  input   clock, // @[:@42.4]
  input   reset, // @[:@43.4]
  input   io_input_reset, // @[:@44.4]
  output  io_output_done // @[:@44.4]
);
  wire  bases_0_clock; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_reset; // @[Counter.scala 253:53:@57.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 253:53:@57.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 253:53:@57.4]
  wire [31:0] bases_0_io_wPort_0_init; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_io_reset; // @[Counter.scala 253:53:@57.4]
  wire  SRFF_clock; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_set; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_output; // @[Counter.scala 255:22:@73.4]
  wire [31:0] _T_48; // @[Counter.scala 279:52:@101.4]
  wire [32:0] _T_50; // @[Counter.scala 283:33:@102.4]
  wire [31:0] _T_51; // @[Counter.scala 283:33:@103.4]
  wire [31:0] _T_52; // @[Counter.scala 283:33:@104.4]
  wire  _T_57; // @[Counter.scala 285:18:@106.4]
  wire [31:0] _T_68; // @[Counter.scala 291:115:@114.4]
  wire [31:0] _T_71; // @[Counter.scala 291:152:@117.4]
  wire [31:0] _T_72; // @[Counter.scala 291:74:@118.4]
  FF bases_0 ( // @[Counter.scala 253:53:@57.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_init(bases_0_io_wPort_0_init),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0),
    .io_reset(bases_0_io_reset)
  );
  SRFF SRFF ( // @[Counter.scala 255:22:@73.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 279:52:@101.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@102.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@103.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 283:33:@104.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'shc); // @[Counter.scala 285:18:@106.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 291:115:@114.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 291:152:@117.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 291:74:@118.4]
  assign io_output_done = $signed(_T_52) >= $signed(32'shc); // @[Counter.scala 325:20:@127.4]
  assign bases_0_clock = clock; // @[:@58.4]
  assign bases_0_reset = reset; // @[:@59.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 291:31:@120.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 273:27:@99.4]
  assign bases_0_io_wPort_0_init = 32'h0; // @[Counter.scala 272:26:@96.4]
  assign bases_0_io_wPort_0_en_0 = 1'h1; // @[Counter.scala 276:29:@100.4]
  assign bases_0_io_reset = 1'h0; // @[Counter.scala 271:18:@94.4]
  assign SRFF_clock = clock; // @[:@74.4]
  assign SRFF_reset = reset; // @[:@75.4]
  assign SRFF_io_input_set = io_input_reset == 1'h0; // @[Counter.scala 256:23:@78.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 257:25:@80.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 258:30:@81.4]
endmodule
module RetimeWrapper( // @[:@144.2]
  input   clock, // @[:@145.4]
  input   reset, // @[:@146.4]
  input   io_flow, // @[:@147.4]
  input   io_in, // @[:@147.4]
  output  io_out // @[:@147.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@149.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@149.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@162.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@161.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@160.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@159.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@158.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@156.4]
endmodule
module RootController_sm( // @[:@312.2]
  input   clock, // @[:@313.4]
  input   reset, // @[:@314.4]
  input   io_enable, // @[:@315.4]
  output  io_done, // @[:@315.4]
  input   io_rst, // @[:@315.4]
  input   io_ctrDone, // @[:@315.4]
  output  io_ctrInc, // @[:@315.4]
  input   io_doneIn_0, // @[:@315.4]
  output  io_enableOut_0, // @[:@315.4]
  output  io_childAck_0 // @[:@315.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@318.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@321.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@338.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@433.4]
  wire  finished; // @[Controllers.scala 81:26:@324.4]
  wire  synchronize; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  wire  _T_122; // @[Controllers.scala 128:33:@371.4]
  wire  _T_124; // @[Controllers.scala 128:54:@372.4]
  wire  _T_125; // @[Controllers.scala 128:52:@373.4]
  wire  _T_126; // @[Controllers.scala 128:66:@374.4]
  wire  _T_128; // @[Controllers.scala 128:98:@376.4]
  wire  _T_129; // @[Controllers.scala 128:96:@377.4]
  wire  _T_131; // @[Controllers.scala 128:123:@378.4]
  wire  _T_133; // @[Controllers.scala 129:48:@381.4]
  wire  _T_138; // @[Controllers.scala 130:52:@386.4]
  wire  _T_139; // @[Controllers.scala 130:50:@387.4]
  wire  _T_147; // @[Controllers.scala 130:129:@393.4]
  wire  _T_150; // @[Controllers.scala 131:45:@396.4]
  wire  _T_154; // @[Controllers.scala 213:68:@402.4]
  wire  _T_156; // @[Controllers.scala 213:90:@404.4]
  wire  _T_158; // @[Controllers.scala 213:132:@406.4]
  wire  _T_159; // @[Controllers.scala 213:130:@407.4]
  wire  _T_160; // @[Controllers.scala 213:156:@408.4]
  reg  _T_166; // @[package.scala 48:56:@412.4]
  reg [31:0] _RAND_0;
  reg  _T_180; // @[package.scala 48:56:@430.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@318.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@321.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@338.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@357.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@416.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@433.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  assign finished = done_0_io_output | io_done; // @[Controllers.scala 81:26:@324.4]
  assign synchronize = RetimeWrapper_io_out; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  assign _T_122 = done_0_io_output == 1'h0; // @[Controllers.scala 128:33:@371.4]
  assign _T_124 = io_ctrDone == 1'h0; // @[Controllers.scala 128:54:@372.4]
  assign _T_125 = _T_122 & _T_124; // @[Controllers.scala 128:52:@373.4]
  assign _T_126 = _T_125 & io_enable; // @[Controllers.scala 128:66:@374.4]
  assign _T_128 = ~ iterDone_0_io_output; // @[Controllers.scala 128:98:@376.4]
  assign _T_129 = _T_126 & _T_128; // @[Controllers.scala 128:96:@377.4]
  assign _T_131 = io_doneIn_0 == 1'h0; // @[Controllers.scala 128:123:@378.4]
  assign _T_133 = io_doneIn_0 | io_rst; // @[Controllers.scala 129:48:@381.4]
  assign _T_138 = synchronize == 1'h0; // @[Controllers.scala 130:52:@386.4]
  assign _T_139 = io_doneIn_0 & _T_138; // @[Controllers.scala 130:50:@387.4]
  assign _T_147 = finished == 1'h0; // @[Controllers.scala 130:129:@393.4]
  assign _T_150 = io_rst == 1'h0; // @[Controllers.scala 131:45:@396.4]
  assign _T_154 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@402.4]
  assign _T_156 = _T_154 & _T_128; // @[Controllers.scala 213:90:@404.4]
  assign _T_158 = ~ done_0_io_output; // @[Controllers.scala 213:132:@406.4]
  assign _T_159 = _T_156 & _T_158; // @[Controllers.scala 213:130:@407.4]
  assign _T_160 = ~ io_ctrDone; // @[Controllers.scala 213:156:@408.4]
  assign io_done = RetimeWrapper_2_io_out; // @[Controllers.scala 245:13:@440.4]
  assign io_ctrInc = io_doneIn_0; // @[Controllers.scala 122:17:@356.4]
  assign io_enableOut_0 = _T_159 & _T_160; // @[Controllers.scala 213:55:@410.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@401.4]
  assign active_0_clock = clock; // @[:@319.4]
  assign active_0_reset = reset; // @[:@320.4]
  assign active_0_io_input_set = _T_129 & _T_131; // @[Controllers.scala 128:30:@380.4]
  assign active_0_io_input_reset = _T_133 | done_0_io_output; // @[Controllers.scala 129:32:@385.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@326.4]
  assign done_0_clock = clock; // @[:@322.4]
  assign done_0_reset = reset; // @[:@323.4]
  assign done_0_io_input_set = io_ctrDone & _T_150; // @[Controllers.scala 131:28:@399.4]
  assign done_0_io_input_reset = io_rst | done_0_io_output; // @[Controllers.scala 86:33:@336.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@327.4]
  assign iterDone_0_clock = clock; // @[:@339.4]
  assign iterDone_0_reset = reset; // @[:@340.4]
  assign iterDone_0_io_input_set = _T_139 & _T_147; // @[Controllers.scala 130:32:@395.4]
  assign iterDone_0_io_input_reset = synchronize | io_rst; // @[Controllers.scala 92:37:@350.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@341.4]
  assign RetimeWrapper_clock = clock; // @[:@358.4]
  assign RetimeWrapper_reset = reset; // @[:@359.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@361.4]
  assign RetimeWrapper_io_in = io_doneIn_0; // @[package.scala 94:16:@360.4]
  assign RetimeWrapper_1_clock = clock; // @[:@417.4]
  assign RetimeWrapper_1_reset = reset; // @[:@418.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@420.4]
  assign RetimeWrapper_1_io_in = done_0_io_output & _T_166; // @[package.scala 94:16:@419.4]
  assign RetimeWrapper_2_clock = clock; // @[:@434.4]
  assign RetimeWrapper_2_reset = reset; // @[:@435.4]
  assign RetimeWrapper_2_io_flow = io_enable; // @[package.scala 95:18:@437.4]
  assign RetimeWrapper_2_io_in = done_0_io_output & _T_180; // @[package.scala 94:16:@436.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_166 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_180 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_166 <= 1'h0;
    end else begin
      _T_166 <= _T_122;
    end
    if (reset) begin
      _T_180 <= 1'h0;
    end else begin
      _T_180 <= _T_122;
    end
  end
endmodule
module x486_outr_UnitPipe_sm( // @[:@2389.2]
  input   clock, // @[:@2390.4]
  input   reset, // @[:@2391.4]
  input   io_enable, // @[:@2392.4]
  output  io_done, // @[:@2392.4]
  input   io_parentAck, // @[:@2392.4]
  input   io_doneIn_0, // @[:@2392.4]
  output  io_enableOut_0, // @[:@2392.4]
  output  io_childAck_0, // @[:@2392.4]
  input   io_ctrCopyDone_0 // @[:@2392.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@2395.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@2395.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@2395.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@2395.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@2395.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@2395.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@2398.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@2398.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@2398.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@2398.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@2398.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@2398.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@2415.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@2415.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@2415.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@2415.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@2415.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@2415.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@2446.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@2446.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@2446.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@2446.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@2446.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@2460.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@2460.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@2460.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@2460.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@2460.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@2478.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@2478.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@2478.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@2478.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@2478.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@2515.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@2515.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@2515.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@2515.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@2515.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@2532.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@2532.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@2532.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@2532.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@2532.4]
  wire  _T_105; // @[Controllers.scala 165:35:@2430.4]
  wire  _T_107; // @[Controllers.scala 165:60:@2431.4]
  wire  _T_108; // @[Controllers.scala 165:58:@2432.4]
  wire  _T_110; // @[Controllers.scala 165:76:@2433.4]
  wire  _T_111; // @[Controllers.scala 165:74:@2434.4]
  wire  _T_115; // @[Controllers.scala 165:109:@2437.4]
  wire  _T_118; // @[Controllers.scala 165:141:@2439.4]
  wire  _T_126; // @[package.scala 96:25:@2451.4 package.scala 96:25:@2452.4]
  wire  _T_130; // @[Controllers.scala 167:54:@2454.4]
  wire  _T_131; // @[Controllers.scala 167:52:@2455.4]
  wire  _T_138; // @[package.scala 96:25:@2465.4 package.scala 96:25:@2466.4]
  wire  _T_156; // @[package.scala 96:25:@2483.4 package.scala 96:25:@2484.4]
  wire  _T_160; // @[Controllers.scala 169:67:@2486.4]
  wire  _T_161; // @[Controllers.scala 169:86:@2487.4]
  wire  _T_174; // @[Controllers.scala 213:68:@2501.4]
  wire  _T_176; // @[Controllers.scala 213:90:@2503.4]
  wire  _T_178; // @[Controllers.scala 213:132:@2505.4]
  reg  _T_186; // @[package.scala 48:56:@2511.4]
  reg [31:0] _RAND_0;
  wire  _T_187; // @[package.scala 100:41:@2513.4]
  reg  _T_200; // @[package.scala 48:56:@2529.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@2395.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@2398.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@2415.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@2446.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@2460.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@2478.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@2515.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@2532.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_105 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@2430.4]
  assign _T_107 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@2431.4]
  assign _T_108 = _T_105 & _T_107; // @[Controllers.scala 165:58:@2432.4]
  assign _T_110 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@2433.4]
  assign _T_111 = _T_108 & _T_110; // @[Controllers.scala 165:74:@2434.4]
  assign _T_115 = _T_111 & io_enable; // @[Controllers.scala 165:109:@2437.4]
  assign _T_118 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@2439.4]
  assign _T_126 = RetimeWrapper_io_out; // @[package.scala 96:25:@2451.4 package.scala 96:25:@2452.4]
  assign _T_130 = _T_126 == 1'h0; // @[Controllers.scala 167:54:@2454.4]
  assign _T_131 = io_doneIn_0 | _T_130; // @[Controllers.scala 167:52:@2455.4]
  assign _T_138 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@2465.4 package.scala 96:25:@2466.4]
  assign _T_156 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@2483.4 package.scala 96:25:@2484.4]
  assign _T_160 = _T_156 == 1'h0; // @[Controllers.scala 169:67:@2486.4]
  assign _T_161 = _T_160 & io_enable; // @[Controllers.scala 169:86:@2487.4]
  assign _T_174 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@2501.4]
  assign _T_176 = _T_174 & _T_105; // @[Controllers.scala 213:90:@2503.4]
  assign _T_178 = ~ done_0_io_output; // @[Controllers.scala 213:132:@2505.4]
  assign _T_187 = done_0_io_output & _T_186; // @[package.scala 100:41:@2513.4]
  assign io_done = RetimeWrapper_4_io_out; // @[Controllers.scala 245:13:@2539.4]
  assign io_enableOut_0 = _T_176 & _T_178; // @[Controllers.scala 213:55:@2509.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@2500.4]
  assign active_0_clock = clock; // @[:@2396.4]
  assign active_0_reset = reset; // @[:@2397.4]
  assign active_0_io_input_set = _T_115 & _T_118; // @[Controllers.scala 165:32:@2441.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@2445.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@2403.4]
  assign done_0_clock = clock; // @[:@2399.4]
  assign done_0_reset = reset; // @[:@2400.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_161; // @[Controllers.scala 169:30:@2491.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@2413.4 Controllers.scala 170:32:@2498.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@2404.4]
  assign iterDone_0_clock = clock; // @[:@2416.4]
  assign iterDone_0_reset = reset; // @[:@2417.4]
  assign iterDone_0_io_input_set = _T_131 & io_enable; // @[Controllers.scala 167:34:@2459.4]
  assign iterDone_0_io_input_reset = _T_138 | io_parentAck; // @[Controllers.scala 92:37:@2427.4 Controllers.scala 168:36:@2475.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@2418.4]
  assign RetimeWrapper_clock = clock; // @[:@2447.4]
  assign RetimeWrapper_reset = reset; // @[:@2448.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@2450.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@2449.4]
  assign RetimeWrapper_1_clock = clock; // @[:@2461.4]
  assign RetimeWrapper_1_reset = reset; // @[:@2462.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@2464.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@2463.4]
  assign RetimeWrapper_2_clock = clock; // @[:@2479.4]
  assign RetimeWrapper_2_reset = reset; // @[:@2480.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@2482.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@2481.4]
  assign RetimeWrapper_3_clock = clock; // @[:@2516.4]
  assign RetimeWrapper_3_reset = reset; // @[:@2517.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@2519.4]
  assign RetimeWrapper_3_io_in = _T_187 | io_parentAck; // @[package.scala 94:16:@2518.4]
  assign RetimeWrapper_4_clock = clock; // @[:@2533.4]
  assign RetimeWrapper_4_reset = reset; // @[:@2534.4]
  assign RetimeWrapper_4_io_flow = io_enable; // @[package.scala 95:18:@2536.4]
  assign RetimeWrapper_4_io_in = done_0_io_output & _T_200; // @[package.scala 94:16:@2535.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_186 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_200 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_186 <= 1'h0;
    end else begin
      _T_186 <= _T_110;
    end
    if (reset) begin
      _T_200 <= 1'h0;
    end else begin
      _T_200 <= _T_110;
    end
  end
endmodule
module SingleCounter_1( // @[:@2659.2]
  input         clock, // @[:@2660.4]
  input         reset, // @[:@2661.4]
  input         io_setup_saturate, // @[:@2662.4]
  input         io_input_reset, // @[:@2662.4]
  input         io_input_enable, // @[:@2662.4]
  output [31:0] io_output_count_0, // @[:@2662.4]
  output        io_output_oobs_0, // @[:@2662.4]
  output        io_output_done, // @[:@2662.4]
  output        io_output_saturated // @[:@2662.4]
);
  wire  bases_0_clock; // @[Counter.scala 253:53:@2675.4]
  wire  bases_0_reset; // @[Counter.scala 253:53:@2675.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 253:53:@2675.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 253:53:@2675.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 253:53:@2675.4]
  wire [31:0] bases_0_io_wPort_0_init; // @[Counter.scala 253:53:@2675.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 253:53:@2675.4]
  wire  bases_0_io_reset; // @[Counter.scala 253:53:@2675.4]
  wire  SRFF_clock; // @[Counter.scala 255:22:@2691.4]
  wire  SRFF_reset; // @[Counter.scala 255:22:@2691.4]
  wire  SRFF_io_input_set; // @[Counter.scala 255:22:@2691.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 255:22:@2691.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 255:22:@2691.4]
  wire  SRFF_io_output; // @[Counter.scala 255:22:@2691.4]
  wire  _T_36; // @[Counter.scala 256:45:@2694.4]
  wire [31:0] _T_48; // @[Counter.scala 279:52:@2719.4]
  wire [32:0] _T_50; // @[Counter.scala 283:33:@2720.4]
  wire [31:0] _T_51; // @[Counter.scala 283:33:@2721.4]
  wire [31:0] _T_52; // @[Counter.scala 283:33:@2722.4]
  wire  _T_57; // @[Counter.scala 285:18:@2724.4]
  wire [31:0] _T_68; // @[Counter.scala 291:115:@2732.4]
  wire [31:0] _T_70; // @[Counter.scala 291:85:@2734.4]
  wire [31:0] _T_71; // @[Counter.scala 291:152:@2735.4]
  wire [31:0] _T_72; // @[Counter.scala 291:74:@2736.4]
  wire  _T_75; // @[Counter.scala 314:102:@2740.4]
  wire  _T_77; // @[Counter.scala 314:130:@2741.4]
  FF bases_0 ( // @[Counter.scala 253:53:@2675.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_init(bases_0_io_wPort_0_init),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0),
    .io_reset(bases_0_io_reset)
  );
  SRFF SRFF ( // @[Counter.scala 255:22:@2691.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 256:45:@2694.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 279:52:@2719.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@2720.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@2721.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 283:33:@2722.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh4); // @[Counter.scala 285:18:@2724.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 291:115:@2732.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 32'h0; // @[Counter.scala 291:85:@2734.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 291:152:@2735.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 291:74:@2736.4]
  assign _T_75 = $signed(_T_48) < $signed(32'sh0); // @[Counter.scala 314:102:@2740.4]
  assign _T_77 = $signed(_T_48) >= $signed(32'sh4); // @[Counter.scala 314:130:@2741.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 296:28:@2739.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 314:60:@2743.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 325:20:@2745.4]
  assign io_output_saturated = io_setup_saturate & _T_57; // @[Counter.scala 332:25:@2748.4]
  assign bases_0_clock = clock; // @[:@2676.4]
  assign bases_0_reset = reset; // @[:@2677.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 291:31:@2738.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 273:27:@2717.4]
  assign bases_0_io_wPort_0_init = 32'h0; // @[Counter.scala 272:26:@2714.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 276:29:@2718.4]
  assign bases_0_io_reset = 1'h0; // @[Counter.scala 271:18:@2712.4]
  assign SRFF_clock = clock; // @[:@2692.4]
  assign SRFF_reset = reset; // @[:@2693.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 256:23:@2696.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 257:25:@2698.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 258:30:@2699.4]
endmodule
module x278_ctrchain( // @[:@2879.2]
  input         clock, // @[:@2880.4]
  input         reset, // @[:@2881.4]
  input         io_input_reset, // @[:@2882.4]
  input         io_input_enable, // @[:@2882.4]
  output [31:0] io_output_counts_1, // @[:@2882.4]
  output [31:0] io_output_counts_0, // @[:@2882.4]
  output        io_output_oobs_0, // @[:@2882.4]
  output        io_output_oobs_1, // @[:@2882.4]
  output        io_output_done // @[:@2882.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_reset; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_io_setup_saturate; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 505:46:@2884.4]
  wire [31:0] ctrs_0_io_output_count_0; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_io_output_saturated; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_1_clock; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_reset; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_io_setup_saturate; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_io_input_reset; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_io_input_enable; // @[Counter.scala 505:46:@2887.4]
  wire [31:0] ctrs_1_io_output_count_0; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_io_output_oobs_0; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_io_output_done; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_io_output_saturated; // @[Counter.scala 505:46:@2887.4]
  wire  isDone; // @[Counter.scala 533:51:@2904.4]
  reg  wasDone; // @[Counter.scala 534:24:@2905.4]
  reg [31:0] _RAND_0;
  wire  _T_64; // @[Counter.scala 538:69:@2913.4]
  wire  _T_66; // @[Counter.scala 538:80:@2914.4]
  reg  doneLatch; // @[Counter.scala 542:26:@2919.4]
  reg [31:0] _RAND_1;
  wire  _T_73; // @[Counter.scala 543:48:@2920.4]
  wire  _T_74; // @[Counter.scala 543:19:@2921.4]
  SingleCounter_1 ctrs_0 ( // @[Counter.scala 505:46:@2884.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_setup_saturate(ctrs_0_io_setup_saturate),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done),
    .io_output_saturated(ctrs_0_io_output_saturated)
  );
  SingleCounter_1 ctrs_1 ( // @[Counter.scala 505:46:@2887.4]
    .clock(ctrs_1_clock),
    .reset(ctrs_1_reset),
    .io_setup_saturate(ctrs_1_io_setup_saturate),
    .io_input_reset(ctrs_1_io_input_reset),
    .io_input_enable(ctrs_1_io_input_enable),
    .io_output_count_0(ctrs_1_io_output_count_0),
    .io_output_oobs_0(ctrs_1_io_output_oobs_0),
    .io_output_done(ctrs_1_io_output_done),
    .io_output_saturated(ctrs_1_io_output_saturated)
  );
  assign isDone = ctrs_0_io_output_done & ctrs_1_io_output_done; // @[Counter.scala 533:51:@2904.4]
  assign _T_64 = io_input_enable & isDone; // @[Counter.scala 538:69:@2913.4]
  assign _T_66 = wasDone == 1'h0; // @[Counter.scala 538:80:@2914.4]
  assign _T_73 = isDone ? 1'h1 : doneLatch; // @[Counter.scala 543:48:@2920.4]
  assign _T_74 = io_input_reset ? 1'h0 : _T_73; // @[Counter.scala 543:19:@2921.4]
  assign io_output_counts_1 = ctrs_1_io_output_count_0; // @[Counter.scala 549:32:@2926.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 549:32:@2923.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 550:30:@2925.4]
  assign io_output_oobs_1 = ctrs_1_io_output_oobs_0 | doneLatch; // @[Counter.scala 550:30:@2928.4]
  assign io_output_done = _T_64 & _T_66; // @[Counter.scala 538:18:@2916.4]
  assign ctrs_0_clock = clock; // @[:@2885.4]
  assign ctrs_0_reset = reset; // @[:@2886.4]
  assign ctrs_0_io_setup_saturate = 1'h1; // @[Counter.scala 522:29:@2901.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 512:24:@2893.4]
  assign ctrs_0_io_input_enable = ctrs_1_io_output_done & io_input_enable; // @[Counter.scala 518:29:@2900.4]
  assign ctrs_1_clock = clock; // @[:@2888.4]
  assign ctrs_1_reset = reset; // @[:@2889.4]
  assign ctrs_1_io_setup_saturate = ctrs_0_io_output_saturated; // @[Counter.scala 524:31:@2903.4]
  assign ctrs_1_io_input_reset = io_input_reset; // @[Counter.scala 512:24:@2897.4]
  assign ctrs_1_io_input_enable = io_input_enable; // @[Counter.scala 516:33:@2898.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= isDone;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (isDone) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module RetimeWrapper_12( // @[:@2968.2]
  input   clock, // @[:@2969.4]
  input   reset, // @[:@2970.4]
  input   io_flow, // @[:@2971.4]
  input   io_in, // @[:@2971.4]
  output  io_out // @[:@2971.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(12)) sr ( // @[RetimeShiftRegister.scala 15:20:@2973.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@2986.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@2985.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@2984.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@2983.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@2982.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@2980.4]
endmodule
module RetimeWrapper_16( // @[:@3096.2]
  input   clock, // @[:@3097.4]
  input   reset, // @[:@3098.4]
  input   io_flow, // @[:@3099.4]
  input   io_in, // @[:@3099.4]
  output  io_out // @[:@3099.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(11)) sr ( // @[RetimeShiftRegister.scala 15:20:@3101.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3114.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3113.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3112.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3111.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3110.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3108.4]
endmodule
module x485_inr_Foreach_SAMPLER_BOX_sm( // @[:@3116.2]
  input   clock, // @[:@3117.4]
  input   reset, // @[:@3118.4]
  input   io_enable, // @[:@3119.4]
  output  io_done, // @[:@3119.4]
  output  io_doneLatch, // @[:@3119.4]
  input   io_ctrDone, // @[:@3119.4]
  output  io_datapathEn, // @[:@3119.4]
  output  io_ctrInc, // @[:@3119.4]
  output  io_ctrRst, // @[:@3119.4]
  input   io_parentAck, // @[:@3119.4]
  input   io_backpressure, // @[:@3119.4]
  input   io_break // @[:@3119.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@3121.4]
  wire  active_reset; // @[Controllers.scala 261:22:@3121.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@3121.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@3121.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@3121.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@3121.4]
  wire  done_clock; // @[Controllers.scala 262:20:@3124.4]
  wire  done_reset; // @[Controllers.scala 262:20:@3124.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@3124.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@3124.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@3124.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@3124.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3158.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3158.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3158.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@3158.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@3158.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@3180.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@3180.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@3180.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@3180.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@3180.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@3192.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@3192.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@3192.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@3192.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@3192.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@3200.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@3200.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@3200.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@3200.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@3200.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@3216.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@3216.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@3216.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@3216.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@3216.4]
  wire  _T_80; // @[Controllers.scala 264:48:@3129.4]
  wire  _T_81; // @[Controllers.scala 264:46:@3130.4]
  wire  _T_82; // @[Controllers.scala 264:62:@3131.4]
  wire  _T_83; // @[Controllers.scala 264:60:@3132.4]
  wire  _T_100; // @[package.scala 100:49:@3149.4]
  reg  _T_103; // @[package.scala 48:56:@3150.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@3163.4 package.scala 96:25:@3164.4]
  wire  _T_110; // @[package.scala 100:49:@3165.4]
  reg  _T_113; // @[package.scala 48:56:@3166.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@3168.4]
  wire  _T_118; // @[Controllers.scala 283:41:@3173.4]
  wire  _T_119; // @[Controllers.scala 283:59:@3174.4]
  wire  _T_121; // @[Controllers.scala 284:37:@3177.4]
  wire  _T_124; // @[package.scala 96:25:@3185.4 package.scala 96:25:@3186.4]
  wire  _T_126; // @[package.scala 100:49:@3187.4]
  reg  _T_129; // @[package.scala 48:56:@3188.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@3210.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@3212.4]
  reg  _T_153; // @[package.scala 48:56:@3213.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@3221.4 package.scala 96:25:@3222.4]
  wire  _T_158; // @[Controllers.scala 292:61:@3223.4]
  wire  _T_159; // @[Controllers.scala 292:24:@3224.4]
  SRFF active ( // @[Controllers.scala 261:22:@3121.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@3124.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_12 RetimeWrapper ( // @[package.scala 93:22:@3158.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_12 RetimeWrapper_1 ( // @[package.scala 93:22:@3180.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@3192.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@3200.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_16 RetimeWrapper_4 ( // @[package.scala 93:22:@3216.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@3129.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@3130.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@3131.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@3132.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@3149.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@3163.4 package.scala 96:25:@3164.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@3165.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@3168.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@3173.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@3174.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@3177.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@3185.4 package.scala 96:25:@3186.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@3187.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@3212.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@3221.4 package.scala 96:25:@3222.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@3223.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@3224.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@3191.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@3226.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@3176.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@3179.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@3171.4]
  assign active_clock = clock; // @[:@3122.4]
  assign active_reset = reset; // @[:@3123.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@3134.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@3138.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@3139.4]
  assign done_clock = clock; // @[:@3125.4]
  assign done_reset = reset; // @[:@3126.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@3154.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@3147.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@3148.4]
  assign RetimeWrapper_clock = clock; // @[:@3159.4]
  assign RetimeWrapper_reset = reset; // @[:@3160.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@3162.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@3161.4]
  assign RetimeWrapper_1_clock = clock; // @[:@3181.4]
  assign RetimeWrapper_1_reset = reset; // @[:@3182.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@3184.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@3183.4]
  assign RetimeWrapper_2_clock = clock; // @[:@3193.4]
  assign RetimeWrapper_2_reset = reset; // @[:@3194.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@3196.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@3195.4]
  assign RetimeWrapper_3_clock = clock; // @[:@3201.4]
  assign RetimeWrapper_3_reset = reset; // @[:@3202.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@3204.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@3203.4]
  assign RetimeWrapper_4_clock = clock; // @[:@3217.4]
  assign RetimeWrapper_4_reset = reset; // @[:@3218.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@3220.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@3219.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module SimBlackBoxesfix2fixBox( // @[:@3332.2]
  input  [31:0] io_a, // @[:@3335.4]
  output [31:0] io_b // @[:@3335.4]
);
  assign io_b = io_a; // @[SimBlackBoxes.scala 99:40:@3345.4]
endmodule
module _( // @[:@3347.2]
  input  [31:0] io_b, // @[:@3350.4]
  output [31:0] io_result // @[:@3350.4]
);
  wire [31:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@3355.4]
  wire [31:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@3355.4]
  SimBlackBoxesfix2fixBox SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@3355.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@3368.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@3363.4]
endmodule
module RetimeWrapper_21( // @[:@3452.2]
  input        clock, // @[:@3453.4]
  input        reset, // @[:@3454.4]
  input        io_flow, // @[:@3455.4]
  input  [7:0] io_in, // @[:@3455.4]
  output [7:0] io_out // @[:@3455.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@3457.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3470.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3469.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@3468.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3467.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3466.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3464.4]
endmodule
module Mem1D_4( // @[:@3472.2]
  input        clock, // @[:@3473.4]
  input        reset, // @[:@3474.4]
  input        io_r_ofs_0, // @[:@3475.4]
  input        io_r_backpressure, // @[:@3475.4]
  input        io_w_ofs_0, // @[:@3475.4]
  input  [7:0] io_w_data_0, // @[:@3475.4]
  input        io_w_en_0, // @[:@3475.4]
  output [7:0] io_output // @[:@3475.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3485.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3485.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3485.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@3485.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@3485.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@3494.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@3494.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@3494.4]
  wire [7:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@3494.4]
  wire [7:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@3494.4]
  reg [7:0] _T_127; // @[MemPrimitives.scala 560:26:@3479.4]
  reg [31:0] _RAND_0;
  wire  _T_130; // @[MemPrimitives.scala 561:61:@3481.4]
  wire  _T_131; // @[MemPrimitives.scala 561:44:@3482.4]
  wire [7:0] _T_132; // @[MemPrimitives.scala 561:19:@3483.4]
  wire  _T_135; // @[package.scala 96:25:@3490.4 package.scala 96:25:@3491.4]
  wire  _T_137; // @[Mux.scala 46:19:@3492.4]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@3485.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_1 ( // @[package.scala 93:22:@3494.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign _T_130 = io_w_ofs_0 == 1'h0; // @[MemPrimitives.scala 561:61:@3481.4]
  assign _T_131 = io_w_en_0 & _T_130; // @[MemPrimitives.scala 561:44:@3482.4]
  assign _T_132 = _T_131 ? io_w_data_0 : _T_127; // @[MemPrimitives.scala 561:19:@3483.4]
  assign _T_135 = RetimeWrapper_io_out; // @[package.scala 96:25:@3490.4 package.scala 96:25:@3491.4]
  assign _T_137 = 1'h0 == _T_135; // @[Mux.scala 46:19:@3492.4]
  assign io_output = RetimeWrapper_1_io_out; // @[MemPrimitives.scala 565:17:@3501.4]
  assign RetimeWrapper_clock = clock; // @[:@3486.4]
  assign RetimeWrapper_reset = reset; // @[:@3487.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@3489.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@3488.4]
  assign RetimeWrapper_1_clock = clock; // @[:@3495.4]
  assign RetimeWrapper_1_reset = reset; // @[:@3496.4]
  assign RetimeWrapper_1_io_flow = io_r_backpressure; // @[package.scala 95:18:@3498.4]
  assign RetimeWrapper_1_io_in = _T_137 ? _T_127 : 8'h0; // @[package.scala 94:16:@3497.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_127 = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_127 <= 8'h0;
    end else begin
      if (_T_131) begin
        _T_127 <= io_w_data_0;
      end
    end
  end
endmodule
module StickySelects( // @[:@4928.2]
  input   clock, // @[:@4929.4]
  input   reset, // @[:@4930.4]
  input   io_ins_0, // @[:@4931.4]
  input   io_ins_1, // @[:@4931.4]
  input   io_ins_2, // @[:@4931.4]
  input   io_ins_3, // @[:@4931.4]
  input   io_ins_4, // @[:@4931.4]
  input   io_ins_5, // @[:@4931.4]
  input   io_ins_6, // @[:@4931.4]
  input   io_ins_7, // @[:@4931.4]
  input   io_ins_8, // @[:@4931.4]
  output  io_outs_0, // @[:@4931.4]
  output  io_outs_1, // @[:@4931.4]
  output  io_outs_2, // @[:@4931.4]
  output  io_outs_3, // @[:@4931.4]
  output  io_outs_4, // @[:@4931.4]
  output  io_outs_5, // @[:@4931.4]
  output  io_outs_6, // @[:@4931.4]
  output  io_outs_7, // @[:@4931.4]
  output  io_outs_8 // @[:@4931.4]
);
  reg  _T_19; // @[StickySelects.scala 21:22:@4933.4]
  reg [31:0] _RAND_0;
  wire  _T_20; // @[StickySelects.scala 22:54:@4934.4]
  wire  _T_21; // @[StickySelects.scala 22:54:@4935.4]
  wire  _T_22; // @[StickySelects.scala 22:54:@4936.4]
  wire  _T_23; // @[StickySelects.scala 22:54:@4937.4]
  wire  _T_24; // @[StickySelects.scala 22:54:@4938.4]
  wire  _T_25; // @[StickySelects.scala 22:54:@4939.4]
  wire  _T_26; // @[StickySelects.scala 22:54:@4940.4]
  wire  _T_28; // @[StickySelects.scala 24:52:@4941.4]
  wire  _T_29; // @[StickySelects.scala 24:21:@4942.4]
  reg  _T_32; // @[StickySelects.scala 21:22:@4944.4]
  reg [31:0] _RAND_1;
  wire  _T_33; // @[StickySelects.scala 22:54:@4945.4]
  wire  _T_34; // @[StickySelects.scala 22:54:@4946.4]
  wire  _T_35; // @[StickySelects.scala 22:54:@4947.4]
  wire  _T_36; // @[StickySelects.scala 22:54:@4948.4]
  wire  _T_37; // @[StickySelects.scala 22:54:@4949.4]
  wire  _T_38; // @[StickySelects.scala 22:54:@4950.4]
  wire  _T_39; // @[StickySelects.scala 22:54:@4951.4]
  wire  _T_41; // @[StickySelects.scala 24:52:@4952.4]
  wire  _T_42; // @[StickySelects.scala 24:21:@4953.4]
  reg  _T_45; // @[StickySelects.scala 21:22:@4955.4]
  reg [31:0] _RAND_2;
  wire  _T_46; // @[StickySelects.scala 22:54:@4956.4]
  wire  _T_47; // @[StickySelects.scala 22:54:@4957.4]
  wire  _T_48; // @[StickySelects.scala 22:54:@4958.4]
  wire  _T_49; // @[StickySelects.scala 22:54:@4959.4]
  wire  _T_50; // @[StickySelects.scala 22:54:@4960.4]
  wire  _T_51; // @[StickySelects.scala 22:54:@4961.4]
  wire  _T_52; // @[StickySelects.scala 22:54:@4962.4]
  wire  _T_54; // @[StickySelects.scala 24:52:@4963.4]
  wire  _T_55; // @[StickySelects.scala 24:21:@4964.4]
  reg  _T_58; // @[StickySelects.scala 21:22:@4966.4]
  reg [31:0] _RAND_3;
  wire  _T_60; // @[StickySelects.scala 22:54:@4968.4]
  wire  _T_61; // @[StickySelects.scala 22:54:@4969.4]
  wire  _T_62; // @[StickySelects.scala 22:54:@4970.4]
  wire  _T_63; // @[StickySelects.scala 22:54:@4971.4]
  wire  _T_64; // @[StickySelects.scala 22:54:@4972.4]
  wire  _T_65; // @[StickySelects.scala 22:54:@4973.4]
  wire  _T_67; // @[StickySelects.scala 24:52:@4974.4]
  wire  _T_68; // @[StickySelects.scala 24:21:@4975.4]
  reg  _T_71; // @[StickySelects.scala 21:22:@4977.4]
  reg [31:0] _RAND_4;
  wire  _T_74; // @[StickySelects.scala 22:54:@4980.4]
  wire  _T_75; // @[StickySelects.scala 22:54:@4981.4]
  wire  _T_76; // @[StickySelects.scala 22:54:@4982.4]
  wire  _T_77; // @[StickySelects.scala 22:54:@4983.4]
  wire  _T_78; // @[StickySelects.scala 22:54:@4984.4]
  wire  _T_80; // @[StickySelects.scala 24:52:@4985.4]
  wire  _T_81; // @[StickySelects.scala 24:21:@4986.4]
  reg  _T_84; // @[StickySelects.scala 21:22:@4988.4]
  reg [31:0] _RAND_5;
  wire  _T_88; // @[StickySelects.scala 22:54:@4992.4]
  wire  _T_89; // @[StickySelects.scala 22:54:@4993.4]
  wire  _T_90; // @[StickySelects.scala 22:54:@4994.4]
  wire  _T_91; // @[StickySelects.scala 22:54:@4995.4]
  wire  _T_93; // @[StickySelects.scala 24:52:@4996.4]
  wire  _T_94; // @[StickySelects.scala 24:21:@4997.4]
  reg  _T_97; // @[StickySelects.scala 21:22:@4999.4]
  reg [31:0] _RAND_6;
  wire  _T_102; // @[StickySelects.scala 22:54:@5004.4]
  wire  _T_103; // @[StickySelects.scala 22:54:@5005.4]
  wire  _T_104; // @[StickySelects.scala 22:54:@5006.4]
  wire  _T_106; // @[StickySelects.scala 24:52:@5007.4]
  wire  _T_107; // @[StickySelects.scala 24:21:@5008.4]
  reg  _T_110; // @[StickySelects.scala 21:22:@5010.4]
  reg [31:0] _RAND_7;
  wire  _T_116; // @[StickySelects.scala 22:54:@5016.4]
  wire  _T_117; // @[StickySelects.scala 22:54:@5017.4]
  wire  _T_119; // @[StickySelects.scala 24:52:@5018.4]
  wire  _T_120; // @[StickySelects.scala 24:21:@5019.4]
  reg  _T_123; // @[StickySelects.scala 21:22:@5021.4]
  reg [31:0] _RAND_8;
  wire  _T_130; // @[StickySelects.scala 22:54:@5028.4]
  wire  _T_132; // @[StickySelects.scala 24:52:@5029.4]
  wire  _T_133; // @[StickySelects.scala 24:21:@5030.4]
  assign _T_20 = io_ins_1 | io_ins_2; // @[StickySelects.scala 22:54:@4934.4]
  assign _T_21 = _T_20 | io_ins_3; // @[StickySelects.scala 22:54:@4935.4]
  assign _T_22 = _T_21 | io_ins_4; // @[StickySelects.scala 22:54:@4936.4]
  assign _T_23 = _T_22 | io_ins_5; // @[StickySelects.scala 22:54:@4937.4]
  assign _T_24 = _T_23 | io_ins_6; // @[StickySelects.scala 22:54:@4938.4]
  assign _T_25 = _T_24 | io_ins_7; // @[StickySelects.scala 22:54:@4939.4]
  assign _T_26 = _T_25 | io_ins_8; // @[StickySelects.scala 22:54:@4940.4]
  assign _T_28 = io_ins_0 | _T_19; // @[StickySelects.scala 24:52:@4941.4]
  assign _T_29 = _T_26 ? 1'h0 : _T_28; // @[StickySelects.scala 24:21:@4942.4]
  assign _T_33 = io_ins_0 | io_ins_2; // @[StickySelects.scala 22:54:@4945.4]
  assign _T_34 = _T_33 | io_ins_3; // @[StickySelects.scala 22:54:@4946.4]
  assign _T_35 = _T_34 | io_ins_4; // @[StickySelects.scala 22:54:@4947.4]
  assign _T_36 = _T_35 | io_ins_5; // @[StickySelects.scala 22:54:@4948.4]
  assign _T_37 = _T_36 | io_ins_6; // @[StickySelects.scala 22:54:@4949.4]
  assign _T_38 = _T_37 | io_ins_7; // @[StickySelects.scala 22:54:@4950.4]
  assign _T_39 = _T_38 | io_ins_8; // @[StickySelects.scala 22:54:@4951.4]
  assign _T_41 = io_ins_1 | _T_32; // @[StickySelects.scala 24:52:@4952.4]
  assign _T_42 = _T_39 ? 1'h0 : _T_41; // @[StickySelects.scala 24:21:@4953.4]
  assign _T_46 = io_ins_0 | io_ins_1; // @[StickySelects.scala 22:54:@4956.4]
  assign _T_47 = _T_46 | io_ins_3; // @[StickySelects.scala 22:54:@4957.4]
  assign _T_48 = _T_47 | io_ins_4; // @[StickySelects.scala 22:54:@4958.4]
  assign _T_49 = _T_48 | io_ins_5; // @[StickySelects.scala 22:54:@4959.4]
  assign _T_50 = _T_49 | io_ins_6; // @[StickySelects.scala 22:54:@4960.4]
  assign _T_51 = _T_50 | io_ins_7; // @[StickySelects.scala 22:54:@4961.4]
  assign _T_52 = _T_51 | io_ins_8; // @[StickySelects.scala 22:54:@4962.4]
  assign _T_54 = io_ins_2 | _T_45; // @[StickySelects.scala 24:52:@4963.4]
  assign _T_55 = _T_52 ? 1'h0 : _T_54; // @[StickySelects.scala 24:21:@4964.4]
  assign _T_60 = _T_46 | io_ins_2; // @[StickySelects.scala 22:54:@4968.4]
  assign _T_61 = _T_60 | io_ins_4; // @[StickySelects.scala 22:54:@4969.4]
  assign _T_62 = _T_61 | io_ins_5; // @[StickySelects.scala 22:54:@4970.4]
  assign _T_63 = _T_62 | io_ins_6; // @[StickySelects.scala 22:54:@4971.4]
  assign _T_64 = _T_63 | io_ins_7; // @[StickySelects.scala 22:54:@4972.4]
  assign _T_65 = _T_64 | io_ins_8; // @[StickySelects.scala 22:54:@4973.4]
  assign _T_67 = io_ins_3 | _T_58; // @[StickySelects.scala 24:52:@4974.4]
  assign _T_68 = _T_65 ? 1'h0 : _T_67; // @[StickySelects.scala 24:21:@4975.4]
  assign _T_74 = _T_60 | io_ins_3; // @[StickySelects.scala 22:54:@4980.4]
  assign _T_75 = _T_74 | io_ins_5; // @[StickySelects.scala 22:54:@4981.4]
  assign _T_76 = _T_75 | io_ins_6; // @[StickySelects.scala 22:54:@4982.4]
  assign _T_77 = _T_76 | io_ins_7; // @[StickySelects.scala 22:54:@4983.4]
  assign _T_78 = _T_77 | io_ins_8; // @[StickySelects.scala 22:54:@4984.4]
  assign _T_80 = io_ins_4 | _T_71; // @[StickySelects.scala 24:52:@4985.4]
  assign _T_81 = _T_78 ? 1'h0 : _T_80; // @[StickySelects.scala 24:21:@4986.4]
  assign _T_88 = _T_74 | io_ins_4; // @[StickySelects.scala 22:54:@4992.4]
  assign _T_89 = _T_88 | io_ins_6; // @[StickySelects.scala 22:54:@4993.4]
  assign _T_90 = _T_89 | io_ins_7; // @[StickySelects.scala 22:54:@4994.4]
  assign _T_91 = _T_90 | io_ins_8; // @[StickySelects.scala 22:54:@4995.4]
  assign _T_93 = io_ins_5 | _T_84; // @[StickySelects.scala 24:52:@4996.4]
  assign _T_94 = _T_91 ? 1'h0 : _T_93; // @[StickySelects.scala 24:21:@4997.4]
  assign _T_102 = _T_88 | io_ins_5; // @[StickySelects.scala 22:54:@5004.4]
  assign _T_103 = _T_102 | io_ins_7; // @[StickySelects.scala 22:54:@5005.4]
  assign _T_104 = _T_103 | io_ins_8; // @[StickySelects.scala 22:54:@5006.4]
  assign _T_106 = io_ins_6 | _T_97; // @[StickySelects.scala 24:52:@5007.4]
  assign _T_107 = _T_104 ? 1'h0 : _T_106; // @[StickySelects.scala 24:21:@5008.4]
  assign _T_116 = _T_102 | io_ins_6; // @[StickySelects.scala 22:54:@5016.4]
  assign _T_117 = _T_116 | io_ins_8; // @[StickySelects.scala 22:54:@5017.4]
  assign _T_119 = io_ins_7 | _T_110; // @[StickySelects.scala 24:52:@5018.4]
  assign _T_120 = _T_117 ? 1'h0 : _T_119; // @[StickySelects.scala 24:21:@5019.4]
  assign _T_130 = _T_116 | io_ins_7; // @[StickySelects.scala 22:54:@5028.4]
  assign _T_132 = io_ins_8 | _T_123; // @[StickySelects.scala 24:52:@5029.4]
  assign _T_133 = _T_130 ? 1'h0 : _T_132; // @[StickySelects.scala 24:21:@5030.4]
  assign io_outs_0 = _T_26 ? 1'h0 : _T_28; // @[StickySelects.scala 28:52:@5032.4]
  assign io_outs_1 = _T_39 ? 1'h0 : _T_41; // @[StickySelects.scala 28:52:@5033.4]
  assign io_outs_2 = _T_52 ? 1'h0 : _T_54; // @[StickySelects.scala 28:52:@5034.4]
  assign io_outs_3 = _T_65 ? 1'h0 : _T_67; // @[StickySelects.scala 28:52:@5035.4]
  assign io_outs_4 = _T_78 ? 1'h0 : _T_80; // @[StickySelects.scala 28:52:@5036.4]
  assign io_outs_5 = _T_91 ? 1'h0 : _T_93; // @[StickySelects.scala 28:52:@5037.4]
  assign io_outs_6 = _T_104 ? 1'h0 : _T_106; // @[StickySelects.scala 28:52:@5038.4]
  assign io_outs_7 = _T_117 ? 1'h0 : _T_119; // @[StickySelects.scala 28:52:@5039.4]
  assign io_outs_8 = _T_130 ? 1'h0 : _T_132; // @[StickySelects.scala 28:52:@5040.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_32 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_45 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_58 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_71 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_84 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_97 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_110 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_123 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (_T_26) begin
        _T_19 <= 1'h0;
      end else begin
        _T_19 <= _T_28;
      end
    end
    if (reset) begin
      _T_32 <= 1'h0;
    end else begin
      if (_T_39) begin
        _T_32 <= 1'h0;
      end else begin
        _T_32 <= _T_41;
      end
    end
    if (reset) begin
      _T_45 <= 1'h0;
    end else begin
      if (_T_52) begin
        _T_45 <= 1'h0;
      end else begin
        _T_45 <= _T_54;
      end
    end
    if (reset) begin
      _T_58 <= 1'h0;
    end else begin
      if (_T_65) begin
        _T_58 <= 1'h0;
      end else begin
        _T_58 <= _T_67;
      end
    end
    if (reset) begin
      _T_71 <= 1'h0;
    end else begin
      if (_T_78) begin
        _T_71 <= 1'h0;
      end else begin
        _T_71 <= _T_80;
      end
    end
    if (reset) begin
      _T_84 <= 1'h0;
    end else begin
      if (_T_91) begin
        _T_84 <= 1'h0;
      end else begin
        _T_84 <= _T_93;
      end
    end
    if (reset) begin
      _T_97 <= 1'h0;
    end else begin
      if (_T_104) begin
        _T_97 <= 1'h0;
      end else begin
        _T_97 <= _T_106;
      end
    end
    if (reset) begin
      _T_110 <= 1'h0;
    end else begin
      if (_T_117) begin
        _T_110 <= 1'h0;
      end else begin
        _T_110 <= _T_119;
      end
    end
    if (reset) begin
      _T_123 <= 1'h0;
    end else begin
      if (_T_130) begin
        _T_123 <= 1'h0;
      end else begin
        _T_123 <= _T_132;
      end
    end
  end
endmodule
module RetimeWrapper_52( // @[:@6764.2]
  input   clock, // @[:@6765.4]
  input   reset, // @[:@6766.4]
  input   io_flow, // @[:@6767.4]
  input   io_in, // @[:@6767.4]
  output  io_out // @[:@6767.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@6769.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@6769.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@6769.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@6769.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@6769.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@6769.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@6769.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@6782.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@6781.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@6780.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@6779.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@6778.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@6776.4]
endmodule
module x283_lb_0( // @[:@11360.2]
  input        clock, // @[:@11361.4]
  input        reset, // @[:@11362.4]
  input  [2:0] io_rPort_8_banks_1, // @[:@11363.4]
  input  [2:0] io_rPort_8_banks_0, // @[:@11363.4]
  input        io_rPort_8_ofs_0, // @[:@11363.4]
  input        io_rPort_8_en_0, // @[:@11363.4]
  input        io_rPort_8_backpressure, // @[:@11363.4]
  output [7:0] io_rPort_8_output_0, // @[:@11363.4]
  input  [2:0] io_rPort_7_banks_1, // @[:@11363.4]
  input  [2:0] io_rPort_7_banks_0, // @[:@11363.4]
  input        io_rPort_7_ofs_0, // @[:@11363.4]
  input        io_rPort_7_en_0, // @[:@11363.4]
  input        io_rPort_7_backpressure, // @[:@11363.4]
  output [7:0] io_rPort_7_output_0, // @[:@11363.4]
  input  [2:0] io_rPort_6_banks_1, // @[:@11363.4]
  input  [2:0] io_rPort_6_banks_0, // @[:@11363.4]
  input        io_rPort_6_ofs_0, // @[:@11363.4]
  input        io_rPort_6_en_0, // @[:@11363.4]
  input        io_rPort_6_backpressure, // @[:@11363.4]
  output [7:0] io_rPort_6_output_0, // @[:@11363.4]
  input  [2:0] io_rPort_5_banks_1, // @[:@11363.4]
  input  [2:0] io_rPort_5_banks_0, // @[:@11363.4]
  input        io_rPort_5_ofs_0, // @[:@11363.4]
  input        io_rPort_5_en_0, // @[:@11363.4]
  input        io_rPort_5_backpressure, // @[:@11363.4]
  output [7:0] io_rPort_5_output_0, // @[:@11363.4]
  input  [2:0] io_rPort_4_banks_1, // @[:@11363.4]
  input  [2:0] io_rPort_4_banks_0, // @[:@11363.4]
  input        io_rPort_4_ofs_0, // @[:@11363.4]
  input        io_rPort_4_en_0, // @[:@11363.4]
  input        io_rPort_4_backpressure, // @[:@11363.4]
  output [7:0] io_rPort_4_output_0, // @[:@11363.4]
  input  [2:0] io_rPort_3_banks_1, // @[:@11363.4]
  input  [2:0] io_rPort_3_banks_0, // @[:@11363.4]
  input        io_rPort_3_ofs_0, // @[:@11363.4]
  input        io_rPort_3_en_0, // @[:@11363.4]
  input        io_rPort_3_backpressure, // @[:@11363.4]
  output [7:0] io_rPort_3_output_0, // @[:@11363.4]
  input  [2:0] io_rPort_2_banks_1, // @[:@11363.4]
  input  [2:0] io_rPort_2_banks_0, // @[:@11363.4]
  input        io_rPort_2_ofs_0, // @[:@11363.4]
  input        io_rPort_2_en_0, // @[:@11363.4]
  input        io_rPort_2_backpressure, // @[:@11363.4]
  output [7:0] io_rPort_2_output_0, // @[:@11363.4]
  input  [2:0] io_rPort_1_banks_1, // @[:@11363.4]
  input  [2:0] io_rPort_1_banks_0, // @[:@11363.4]
  input        io_rPort_1_ofs_0, // @[:@11363.4]
  input        io_rPort_1_en_0, // @[:@11363.4]
  input        io_rPort_1_backpressure, // @[:@11363.4]
  output [7:0] io_rPort_1_output_0, // @[:@11363.4]
  input  [2:0] io_rPort_0_banks_1, // @[:@11363.4]
  input  [2:0] io_rPort_0_banks_0, // @[:@11363.4]
  input        io_rPort_0_ofs_0, // @[:@11363.4]
  input        io_rPort_0_en_0, // @[:@11363.4]
  input        io_rPort_0_backpressure, // @[:@11363.4]
  output [7:0] io_rPort_0_output_0, // @[:@11363.4]
  input  [2:0] io_wPort_0_banks_1, // @[:@11363.4]
  input  [2:0] io_wPort_0_banks_0, // @[:@11363.4]
  input        io_wPort_0_ofs_0, // @[:@11363.4]
  input  [7:0] io_wPort_0_data_0, // @[:@11363.4]
  input        io_wPort_0_en_0 // @[:@11363.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@11428.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@11428.4]
  wire  Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@11428.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@11428.4]
  wire  Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@11428.4]
  wire [7:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@11428.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@11428.4]
  wire [7:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@11428.4]
  wire  Mem1D_1_clock; // @[MemPrimitives.scala 64:21:@11444.4]
  wire  Mem1D_1_reset; // @[MemPrimitives.scala 64:21:@11444.4]
  wire  Mem1D_1_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@11444.4]
  wire  Mem1D_1_io_r_backpressure; // @[MemPrimitives.scala 64:21:@11444.4]
  wire  Mem1D_1_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@11444.4]
  wire [7:0] Mem1D_1_io_w_data_0; // @[MemPrimitives.scala 64:21:@11444.4]
  wire  Mem1D_1_io_w_en_0; // @[MemPrimitives.scala 64:21:@11444.4]
  wire [7:0] Mem1D_1_io_output; // @[MemPrimitives.scala 64:21:@11444.4]
  wire  Mem1D_2_clock; // @[MemPrimitives.scala 64:21:@11460.4]
  wire  Mem1D_2_reset; // @[MemPrimitives.scala 64:21:@11460.4]
  wire  Mem1D_2_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@11460.4]
  wire  Mem1D_2_io_r_backpressure; // @[MemPrimitives.scala 64:21:@11460.4]
  wire  Mem1D_2_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@11460.4]
  wire [7:0] Mem1D_2_io_w_data_0; // @[MemPrimitives.scala 64:21:@11460.4]
  wire  Mem1D_2_io_w_en_0; // @[MemPrimitives.scala 64:21:@11460.4]
  wire [7:0] Mem1D_2_io_output; // @[MemPrimitives.scala 64:21:@11460.4]
  wire  Mem1D_3_clock; // @[MemPrimitives.scala 64:21:@11476.4]
  wire  Mem1D_3_reset; // @[MemPrimitives.scala 64:21:@11476.4]
  wire  Mem1D_3_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@11476.4]
  wire  Mem1D_3_io_r_backpressure; // @[MemPrimitives.scala 64:21:@11476.4]
  wire  Mem1D_3_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@11476.4]
  wire [7:0] Mem1D_3_io_w_data_0; // @[MemPrimitives.scala 64:21:@11476.4]
  wire  Mem1D_3_io_w_en_0; // @[MemPrimitives.scala 64:21:@11476.4]
  wire [7:0] Mem1D_3_io_output; // @[MemPrimitives.scala 64:21:@11476.4]
  wire  Mem1D_4_clock; // @[MemPrimitives.scala 64:21:@11492.4]
  wire  Mem1D_4_reset; // @[MemPrimitives.scala 64:21:@11492.4]
  wire  Mem1D_4_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@11492.4]
  wire  Mem1D_4_io_r_backpressure; // @[MemPrimitives.scala 64:21:@11492.4]
  wire  Mem1D_4_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@11492.4]
  wire [7:0] Mem1D_4_io_w_data_0; // @[MemPrimitives.scala 64:21:@11492.4]
  wire  Mem1D_4_io_w_en_0; // @[MemPrimitives.scala 64:21:@11492.4]
  wire [7:0] Mem1D_4_io_output; // @[MemPrimitives.scala 64:21:@11492.4]
  wire  Mem1D_5_clock; // @[MemPrimitives.scala 64:21:@11508.4]
  wire  Mem1D_5_reset; // @[MemPrimitives.scala 64:21:@11508.4]
  wire  Mem1D_5_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@11508.4]
  wire  Mem1D_5_io_r_backpressure; // @[MemPrimitives.scala 64:21:@11508.4]
  wire  Mem1D_5_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@11508.4]
  wire [7:0] Mem1D_5_io_w_data_0; // @[MemPrimitives.scala 64:21:@11508.4]
  wire  Mem1D_5_io_w_en_0; // @[MemPrimitives.scala 64:21:@11508.4]
  wire [7:0] Mem1D_5_io_output; // @[MemPrimitives.scala 64:21:@11508.4]
  wire  Mem1D_6_clock; // @[MemPrimitives.scala 64:21:@11524.4]
  wire  Mem1D_6_reset; // @[MemPrimitives.scala 64:21:@11524.4]
  wire  Mem1D_6_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@11524.4]
  wire  Mem1D_6_io_r_backpressure; // @[MemPrimitives.scala 64:21:@11524.4]
  wire  Mem1D_6_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@11524.4]
  wire [7:0] Mem1D_6_io_w_data_0; // @[MemPrimitives.scala 64:21:@11524.4]
  wire  Mem1D_6_io_w_en_0; // @[MemPrimitives.scala 64:21:@11524.4]
  wire [7:0] Mem1D_6_io_output; // @[MemPrimitives.scala 64:21:@11524.4]
  wire  Mem1D_7_clock; // @[MemPrimitives.scala 64:21:@11540.4]
  wire  Mem1D_7_reset; // @[MemPrimitives.scala 64:21:@11540.4]
  wire  Mem1D_7_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@11540.4]
  wire  Mem1D_7_io_r_backpressure; // @[MemPrimitives.scala 64:21:@11540.4]
  wire  Mem1D_7_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@11540.4]
  wire [7:0] Mem1D_7_io_w_data_0; // @[MemPrimitives.scala 64:21:@11540.4]
  wire  Mem1D_7_io_w_en_0; // @[MemPrimitives.scala 64:21:@11540.4]
  wire [7:0] Mem1D_7_io_output; // @[MemPrimitives.scala 64:21:@11540.4]
  wire  Mem1D_8_clock; // @[MemPrimitives.scala 64:21:@11556.4]
  wire  Mem1D_8_reset; // @[MemPrimitives.scala 64:21:@11556.4]
  wire  Mem1D_8_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@11556.4]
  wire  Mem1D_8_io_r_backpressure; // @[MemPrimitives.scala 64:21:@11556.4]
  wire  Mem1D_8_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@11556.4]
  wire [7:0] Mem1D_8_io_w_data_0; // @[MemPrimitives.scala 64:21:@11556.4]
  wire  Mem1D_8_io_w_en_0; // @[MemPrimitives.scala 64:21:@11556.4]
  wire [7:0] Mem1D_8_io_output; // @[MemPrimitives.scala 64:21:@11556.4]
  wire  Mem1D_9_clock; // @[MemPrimitives.scala 64:21:@11572.4]
  wire  Mem1D_9_reset; // @[MemPrimitives.scala 64:21:@11572.4]
  wire  Mem1D_9_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@11572.4]
  wire  Mem1D_9_io_r_backpressure; // @[MemPrimitives.scala 64:21:@11572.4]
  wire  Mem1D_9_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@11572.4]
  wire [7:0] Mem1D_9_io_w_data_0; // @[MemPrimitives.scala 64:21:@11572.4]
  wire  Mem1D_9_io_w_en_0; // @[MemPrimitives.scala 64:21:@11572.4]
  wire [7:0] Mem1D_9_io_output; // @[MemPrimitives.scala 64:21:@11572.4]
  wire  Mem1D_10_clock; // @[MemPrimitives.scala 64:21:@11588.4]
  wire  Mem1D_10_reset; // @[MemPrimitives.scala 64:21:@11588.4]
  wire  Mem1D_10_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@11588.4]
  wire  Mem1D_10_io_r_backpressure; // @[MemPrimitives.scala 64:21:@11588.4]
  wire  Mem1D_10_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@11588.4]
  wire [7:0] Mem1D_10_io_w_data_0; // @[MemPrimitives.scala 64:21:@11588.4]
  wire  Mem1D_10_io_w_en_0; // @[MemPrimitives.scala 64:21:@11588.4]
  wire [7:0] Mem1D_10_io_output; // @[MemPrimitives.scala 64:21:@11588.4]
  wire  Mem1D_11_clock; // @[MemPrimitives.scala 64:21:@11604.4]
  wire  Mem1D_11_reset; // @[MemPrimitives.scala 64:21:@11604.4]
  wire  Mem1D_11_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@11604.4]
  wire  Mem1D_11_io_r_backpressure; // @[MemPrimitives.scala 64:21:@11604.4]
  wire  Mem1D_11_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@11604.4]
  wire [7:0] Mem1D_11_io_w_data_0; // @[MemPrimitives.scala 64:21:@11604.4]
  wire  Mem1D_11_io_w_en_0; // @[MemPrimitives.scala 64:21:@11604.4]
  wire [7:0] Mem1D_11_io_output; // @[MemPrimitives.scala 64:21:@11604.4]
  wire  Mem1D_12_clock; // @[MemPrimitives.scala 64:21:@11620.4]
  wire  Mem1D_12_reset; // @[MemPrimitives.scala 64:21:@11620.4]
  wire  Mem1D_12_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@11620.4]
  wire  Mem1D_12_io_r_backpressure; // @[MemPrimitives.scala 64:21:@11620.4]
  wire  Mem1D_12_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@11620.4]
  wire [7:0] Mem1D_12_io_w_data_0; // @[MemPrimitives.scala 64:21:@11620.4]
  wire  Mem1D_12_io_w_en_0; // @[MemPrimitives.scala 64:21:@11620.4]
  wire [7:0] Mem1D_12_io_output; // @[MemPrimitives.scala 64:21:@11620.4]
  wire  Mem1D_13_clock; // @[MemPrimitives.scala 64:21:@11636.4]
  wire  Mem1D_13_reset; // @[MemPrimitives.scala 64:21:@11636.4]
  wire  Mem1D_13_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@11636.4]
  wire  Mem1D_13_io_r_backpressure; // @[MemPrimitives.scala 64:21:@11636.4]
  wire  Mem1D_13_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@11636.4]
  wire [7:0] Mem1D_13_io_w_data_0; // @[MemPrimitives.scala 64:21:@11636.4]
  wire  Mem1D_13_io_w_en_0; // @[MemPrimitives.scala 64:21:@11636.4]
  wire [7:0] Mem1D_13_io_output; // @[MemPrimitives.scala 64:21:@11636.4]
  wire  Mem1D_14_clock; // @[MemPrimitives.scala 64:21:@11652.4]
  wire  Mem1D_14_reset; // @[MemPrimitives.scala 64:21:@11652.4]
  wire  Mem1D_14_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@11652.4]
  wire  Mem1D_14_io_r_backpressure; // @[MemPrimitives.scala 64:21:@11652.4]
  wire  Mem1D_14_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@11652.4]
  wire [7:0] Mem1D_14_io_w_data_0; // @[MemPrimitives.scala 64:21:@11652.4]
  wire  Mem1D_14_io_w_en_0; // @[MemPrimitives.scala 64:21:@11652.4]
  wire [7:0] Mem1D_14_io_output; // @[MemPrimitives.scala 64:21:@11652.4]
  wire  Mem1D_15_clock; // @[MemPrimitives.scala 64:21:@11668.4]
  wire  Mem1D_15_reset; // @[MemPrimitives.scala 64:21:@11668.4]
  wire  Mem1D_15_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@11668.4]
  wire  Mem1D_15_io_r_backpressure; // @[MemPrimitives.scala 64:21:@11668.4]
  wire  Mem1D_15_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@11668.4]
  wire [7:0] Mem1D_15_io_w_data_0; // @[MemPrimitives.scala 64:21:@11668.4]
  wire  Mem1D_15_io_w_en_0; // @[MemPrimitives.scala 64:21:@11668.4]
  wire [7:0] Mem1D_15_io_output; // @[MemPrimitives.scala 64:21:@11668.4]
  wire  StickySelects_clock; // @[MemPrimitives.scala 121:29:@11912.4]
  wire  StickySelects_reset; // @[MemPrimitives.scala 121:29:@11912.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 121:29:@11912.4]
  wire  StickySelects_io_ins_1; // @[MemPrimitives.scala 121:29:@11912.4]
  wire  StickySelects_io_ins_2; // @[MemPrimitives.scala 121:29:@11912.4]
  wire  StickySelects_io_ins_3; // @[MemPrimitives.scala 121:29:@11912.4]
  wire  StickySelects_io_ins_4; // @[MemPrimitives.scala 121:29:@11912.4]
  wire  StickySelects_io_ins_5; // @[MemPrimitives.scala 121:29:@11912.4]
  wire  StickySelects_io_ins_6; // @[MemPrimitives.scala 121:29:@11912.4]
  wire  StickySelects_io_ins_7; // @[MemPrimitives.scala 121:29:@11912.4]
  wire  StickySelects_io_ins_8; // @[MemPrimitives.scala 121:29:@11912.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 121:29:@11912.4]
  wire  StickySelects_io_outs_1; // @[MemPrimitives.scala 121:29:@11912.4]
  wire  StickySelects_io_outs_2; // @[MemPrimitives.scala 121:29:@11912.4]
  wire  StickySelects_io_outs_3; // @[MemPrimitives.scala 121:29:@11912.4]
  wire  StickySelects_io_outs_4; // @[MemPrimitives.scala 121:29:@11912.4]
  wire  StickySelects_io_outs_5; // @[MemPrimitives.scala 121:29:@11912.4]
  wire  StickySelects_io_outs_6; // @[MemPrimitives.scala 121:29:@11912.4]
  wire  StickySelects_io_outs_7; // @[MemPrimitives.scala 121:29:@11912.4]
  wire  StickySelects_io_outs_8; // @[MemPrimitives.scala 121:29:@11912.4]
  wire  StickySelects_1_clock; // @[MemPrimitives.scala 121:29:@12001.4]
  wire  StickySelects_1_reset; // @[MemPrimitives.scala 121:29:@12001.4]
  wire  StickySelects_1_io_ins_0; // @[MemPrimitives.scala 121:29:@12001.4]
  wire  StickySelects_1_io_ins_1; // @[MemPrimitives.scala 121:29:@12001.4]
  wire  StickySelects_1_io_ins_2; // @[MemPrimitives.scala 121:29:@12001.4]
  wire  StickySelects_1_io_ins_3; // @[MemPrimitives.scala 121:29:@12001.4]
  wire  StickySelects_1_io_ins_4; // @[MemPrimitives.scala 121:29:@12001.4]
  wire  StickySelects_1_io_ins_5; // @[MemPrimitives.scala 121:29:@12001.4]
  wire  StickySelects_1_io_ins_6; // @[MemPrimitives.scala 121:29:@12001.4]
  wire  StickySelects_1_io_ins_7; // @[MemPrimitives.scala 121:29:@12001.4]
  wire  StickySelects_1_io_ins_8; // @[MemPrimitives.scala 121:29:@12001.4]
  wire  StickySelects_1_io_outs_0; // @[MemPrimitives.scala 121:29:@12001.4]
  wire  StickySelects_1_io_outs_1; // @[MemPrimitives.scala 121:29:@12001.4]
  wire  StickySelects_1_io_outs_2; // @[MemPrimitives.scala 121:29:@12001.4]
  wire  StickySelects_1_io_outs_3; // @[MemPrimitives.scala 121:29:@12001.4]
  wire  StickySelects_1_io_outs_4; // @[MemPrimitives.scala 121:29:@12001.4]
  wire  StickySelects_1_io_outs_5; // @[MemPrimitives.scala 121:29:@12001.4]
  wire  StickySelects_1_io_outs_6; // @[MemPrimitives.scala 121:29:@12001.4]
  wire  StickySelects_1_io_outs_7; // @[MemPrimitives.scala 121:29:@12001.4]
  wire  StickySelects_1_io_outs_8; // @[MemPrimitives.scala 121:29:@12001.4]
  wire  StickySelects_2_clock; // @[MemPrimitives.scala 121:29:@12090.4]
  wire  StickySelects_2_reset; // @[MemPrimitives.scala 121:29:@12090.4]
  wire  StickySelects_2_io_ins_0; // @[MemPrimitives.scala 121:29:@12090.4]
  wire  StickySelects_2_io_ins_1; // @[MemPrimitives.scala 121:29:@12090.4]
  wire  StickySelects_2_io_ins_2; // @[MemPrimitives.scala 121:29:@12090.4]
  wire  StickySelects_2_io_ins_3; // @[MemPrimitives.scala 121:29:@12090.4]
  wire  StickySelects_2_io_ins_4; // @[MemPrimitives.scala 121:29:@12090.4]
  wire  StickySelects_2_io_ins_5; // @[MemPrimitives.scala 121:29:@12090.4]
  wire  StickySelects_2_io_ins_6; // @[MemPrimitives.scala 121:29:@12090.4]
  wire  StickySelects_2_io_ins_7; // @[MemPrimitives.scala 121:29:@12090.4]
  wire  StickySelects_2_io_ins_8; // @[MemPrimitives.scala 121:29:@12090.4]
  wire  StickySelects_2_io_outs_0; // @[MemPrimitives.scala 121:29:@12090.4]
  wire  StickySelects_2_io_outs_1; // @[MemPrimitives.scala 121:29:@12090.4]
  wire  StickySelects_2_io_outs_2; // @[MemPrimitives.scala 121:29:@12090.4]
  wire  StickySelects_2_io_outs_3; // @[MemPrimitives.scala 121:29:@12090.4]
  wire  StickySelects_2_io_outs_4; // @[MemPrimitives.scala 121:29:@12090.4]
  wire  StickySelects_2_io_outs_5; // @[MemPrimitives.scala 121:29:@12090.4]
  wire  StickySelects_2_io_outs_6; // @[MemPrimitives.scala 121:29:@12090.4]
  wire  StickySelects_2_io_outs_7; // @[MemPrimitives.scala 121:29:@12090.4]
  wire  StickySelects_2_io_outs_8; // @[MemPrimitives.scala 121:29:@12090.4]
  wire  StickySelects_3_clock; // @[MemPrimitives.scala 121:29:@12179.4]
  wire  StickySelects_3_reset; // @[MemPrimitives.scala 121:29:@12179.4]
  wire  StickySelects_3_io_ins_0; // @[MemPrimitives.scala 121:29:@12179.4]
  wire  StickySelects_3_io_ins_1; // @[MemPrimitives.scala 121:29:@12179.4]
  wire  StickySelects_3_io_ins_2; // @[MemPrimitives.scala 121:29:@12179.4]
  wire  StickySelects_3_io_ins_3; // @[MemPrimitives.scala 121:29:@12179.4]
  wire  StickySelects_3_io_ins_4; // @[MemPrimitives.scala 121:29:@12179.4]
  wire  StickySelects_3_io_ins_5; // @[MemPrimitives.scala 121:29:@12179.4]
  wire  StickySelects_3_io_ins_6; // @[MemPrimitives.scala 121:29:@12179.4]
  wire  StickySelects_3_io_ins_7; // @[MemPrimitives.scala 121:29:@12179.4]
  wire  StickySelects_3_io_ins_8; // @[MemPrimitives.scala 121:29:@12179.4]
  wire  StickySelects_3_io_outs_0; // @[MemPrimitives.scala 121:29:@12179.4]
  wire  StickySelects_3_io_outs_1; // @[MemPrimitives.scala 121:29:@12179.4]
  wire  StickySelects_3_io_outs_2; // @[MemPrimitives.scala 121:29:@12179.4]
  wire  StickySelects_3_io_outs_3; // @[MemPrimitives.scala 121:29:@12179.4]
  wire  StickySelects_3_io_outs_4; // @[MemPrimitives.scala 121:29:@12179.4]
  wire  StickySelects_3_io_outs_5; // @[MemPrimitives.scala 121:29:@12179.4]
  wire  StickySelects_3_io_outs_6; // @[MemPrimitives.scala 121:29:@12179.4]
  wire  StickySelects_3_io_outs_7; // @[MemPrimitives.scala 121:29:@12179.4]
  wire  StickySelects_3_io_outs_8; // @[MemPrimitives.scala 121:29:@12179.4]
  wire  StickySelects_4_clock; // @[MemPrimitives.scala 121:29:@12268.4]
  wire  StickySelects_4_reset; // @[MemPrimitives.scala 121:29:@12268.4]
  wire  StickySelects_4_io_ins_0; // @[MemPrimitives.scala 121:29:@12268.4]
  wire  StickySelects_4_io_ins_1; // @[MemPrimitives.scala 121:29:@12268.4]
  wire  StickySelects_4_io_ins_2; // @[MemPrimitives.scala 121:29:@12268.4]
  wire  StickySelects_4_io_ins_3; // @[MemPrimitives.scala 121:29:@12268.4]
  wire  StickySelects_4_io_ins_4; // @[MemPrimitives.scala 121:29:@12268.4]
  wire  StickySelects_4_io_ins_5; // @[MemPrimitives.scala 121:29:@12268.4]
  wire  StickySelects_4_io_ins_6; // @[MemPrimitives.scala 121:29:@12268.4]
  wire  StickySelects_4_io_ins_7; // @[MemPrimitives.scala 121:29:@12268.4]
  wire  StickySelects_4_io_ins_8; // @[MemPrimitives.scala 121:29:@12268.4]
  wire  StickySelects_4_io_outs_0; // @[MemPrimitives.scala 121:29:@12268.4]
  wire  StickySelects_4_io_outs_1; // @[MemPrimitives.scala 121:29:@12268.4]
  wire  StickySelects_4_io_outs_2; // @[MemPrimitives.scala 121:29:@12268.4]
  wire  StickySelects_4_io_outs_3; // @[MemPrimitives.scala 121:29:@12268.4]
  wire  StickySelects_4_io_outs_4; // @[MemPrimitives.scala 121:29:@12268.4]
  wire  StickySelects_4_io_outs_5; // @[MemPrimitives.scala 121:29:@12268.4]
  wire  StickySelects_4_io_outs_6; // @[MemPrimitives.scala 121:29:@12268.4]
  wire  StickySelects_4_io_outs_7; // @[MemPrimitives.scala 121:29:@12268.4]
  wire  StickySelects_4_io_outs_8; // @[MemPrimitives.scala 121:29:@12268.4]
  wire  StickySelects_5_clock; // @[MemPrimitives.scala 121:29:@12357.4]
  wire  StickySelects_5_reset; // @[MemPrimitives.scala 121:29:@12357.4]
  wire  StickySelects_5_io_ins_0; // @[MemPrimitives.scala 121:29:@12357.4]
  wire  StickySelects_5_io_ins_1; // @[MemPrimitives.scala 121:29:@12357.4]
  wire  StickySelects_5_io_ins_2; // @[MemPrimitives.scala 121:29:@12357.4]
  wire  StickySelects_5_io_ins_3; // @[MemPrimitives.scala 121:29:@12357.4]
  wire  StickySelects_5_io_ins_4; // @[MemPrimitives.scala 121:29:@12357.4]
  wire  StickySelects_5_io_ins_5; // @[MemPrimitives.scala 121:29:@12357.4]
  wire  StickySelects_5_io_ins_6; // @[MemPrimitives.scala 121:29:@12357.4]
  wire  StickySelects_5_io_ins_7; // @[MemPrimitives.scala 121:29:@12357.4]
  wire  StickySelects_5_io_ins_8; // @[MemPrimitives.scala 121:29:@12357.4]
  wire  StickySelects_5_io_outs_0; // @[MemPrimitives.scala 121:29:@12357.4]
  wire  StickySelects_5_io_outs_1; // @[MemPrimitives.scala 121:29:@12357.4]
  wire  StickySelects_5_io_outs_2; // @[MemPrimitives.scala 121:29:@12357.4]
  wire  StickySelects_5_io_outs_3; // @[MemPrimitives.scala 121:29:@12357.4]
  wire  StickySelects_5_io_outs_4; // @[MemPrimitives.scala 121:29:@12357.4]
  wire  StickySelects_5_io_outs_5; // @[MemPrimitives.scala 121:29:@12357.4]
  wire  StickySelects_5_io_outs_6; // @[MemPrimitives.scala 121:29:@12357.4]
  wire  StickySelects_5_io_outs_7; // @[MemPrimitives.scala 121:29:@12357.4]
  wire  StickySelects_5_io_outs_8; // @[MemPrimitives.scala 121:29:@12357.4]
  wire  StickySelects_6_clock; // @[MemPrimitives.scala 121:29:@12446.4]
  wire  StickySelects_6_reset; // @[MemPrimitives.scala 121:29:@12446.4]
  wire  StickySelects_6_io_ins_0; // @[MemPrimitives.scala 121:29:@12446.4]
  wire  StickySelects_6_io_ins_1; // @[MemPrimitives.scala 121:29:@12446.4]
  wire  StickySelects_6_io_ins_2; // @[MemPrimitives.scala 121:29:@12446.4]
  wire  StickySelects_6_io_ins_3; // @[MemPrimitives.scala 121:29:@12446.4]
  wire  StickySelects_6_io_ins_4; // @[MemPrimitives.scala 121:29:@12446.4]
  wire  StickySelects_6_io_ins_5; // @[MemPrimitives.scala 121:29:@12446.4]
  wire  StickySelects_6_io_ins_6; // @[MemPrimitives.scala 121:29:@12446.4]
  wire  StickySelects_6_io_ins_7; // @[MemPrimitives.scala 121:29:@12446.4]
  wire  StickySelects_6_io_ins_8; // @[MemPrimitives.scala 121:29:@12446.4]
  wire  StickySelects_6_io_outs_0; // @[MemPrimitives.scala 121:29:@12446.4]
  wire  StickySelects_6_io_outs_1; // @[MemPrimitives.scala 121:29:@12446.4]
  wire  StickySelects_6_io_outs_2; // @[MemPrimitives.scala 121:29:@12446.4]
  wire  StickySelects_6_io_outs_3; // @[MemPrimitives.scala 121:29:@12446.4]
  wire  StickySelects_6_io_outs_4; // @[MemPrimitives.scala 121:29:@12446.4]
  wire  StickySelects_6_io_outs_5; // @[MemPrimitives.scala 121:29:@12446.4]
  wire  StickySelects_6_io_outs_6; // @[MemPrimitives.scala 121:29:@12446.4]
  wire  StickySelects_6_io_outs_7; // @[MemPrimitives.scala 121:29:@12446.4]
  wire  StickySelects_6_io_outs_8; // @[MemPrimitives.scala 121:29:@12446.4]
  wire  StickySelects_7_clock; // @[MemPrimitives.scala 121:29:@12535.4]
  wire  StickySelects_7_reset; // @[MemPrimitives.scala 121:29:@12535.4]
  wire  StickySelects_7_io_ins_0; // @[MemPrimitives.scala 121:29:@12535.4]
  wire  StickySelects_7_io_ins_1; // @[MemPrimitives.scala 121:29:@12535.4]
  wire  StickySelects_7_io_ins_2; // @[MemPrimitives.scala 121:29:@12535.4]
  wire  StickySelects_7_io_ins_3; // @[MemPrimitives.scala 121:29:@12535.4]
  wire  StickySelects_7_io_ins_4; // @[MemPrimitives.scala 121:29:@12535.4]
  wire  StickySelects_7_io_ins_5; // @[MemPrimitives.scala 121:29:@12535.4]
  wire  StickySelects_7_io_ins_6; // @[MemPrimitives.scala 121:29:@12535.4]
  wire  StickySelects_7_io_ins_7; // @[MemPrimitives.scala 121:29:@12535.4]
  wire  StickySelects_7_io_ins_8; // @[MemPrimitives.scala 121:29:@12535.4]
  wire  StickySelects_7_io_outs_0; // @[MemPrimitives.scala 121:29:@12535.4]
  wire  StickySelects_7_io_outs_1; // @[MemPrimitives.scala 121:29:@12535.4]
  wire  StickySelects_7_io_outs_2; // @[MemPrimitives.scala 121:29:@12535.4]
  wire  StickySelects_7_io_outs_3; // @[MemPrimitives.scala 121:29:@12535.4]
  wire  StickySelects_7_io_outs_4; // @[MemPrimitives.scala 121:29:@12535.4]
  wire  StickySelects_7_io_outs_5; // @[MemPrimitives.scala 121:29:@12535.4]
  wire  StickySelects_7_io_outs_6; // @[MemPrimitives.scala 121:29:@12535.4]
  wire  StickySelects_7_io_outs_7; // @[MemPrimitives.scala 121:29:@12535.4]
  wire  StickySelects_7_io_outs_8; // @[MemPrimitives.scala 121:29:@12535.4]
  wire  StickySelects_8_clock; // @[MemPrimitives.scala 121:29:@12624.4]
  wire  StickySelects_8_reset; // @[MemPrimitives.scala 121:29:@12624.4]
  wire  StickySelects_8_io_ins_0; // @[MemPrimitives.scala 121:29:@12624.4]
  wire  StickySelects_8_io_ins_1; // @[MemPrimitives.scala 121:29:@12624.4]
  wire  StickySelects_8_io_ins_2; // @[MemPrimitives.scala 121:29:@12624.4]
  wire  StickySelects_8_io_ins_3; // @[MemPrimitives.scala 121:29:@12624.4]
  wire  StickySelects_8_io_ins_4; // @[MemPrimitives.scala 121:29:@12624.4]
  wire  StickySelects_8_io_ins_5; // @[MemPrimitives.scala 121:29:@12624.4]
  wire  StickySelects_8_io_ins_6; // @[MemPrimitives.scala 121:29:@12624.4]
  wire  StickySelects_8_io_ins_7; // @[MemPrimitives.scala 121:29:@12624.4]
  wire  StickySelects_8_io_ins_8; // @[MemPrimitives.scala 121:29:@12624.4]
  wire  StickySelects_8_io_outs_0; // @[MemPrimitives.scala 121:29:@12624.4]
  wire  StickySelects_8_io_outs_1; // @[MemPrimitives.scala 121:29:@12624.4]
  wire  StickySelects_8_io_outs_2; // @[MemPrimitives.scala 121:29:@12624.4]
  wire  StickySelects_8_io_outs_3; // @[MemPrimitives.scala 121:29:@12624.4]
  wire  StickySelects_8_io_outs_4; // @[MemPrimitives.scala 121:29:@12624.4]
  wire  StickySelects_8_io_outs_5; // @[MemPrimitives.scala 121:29:@12624.4]
  wire  StickySelects_8_io_outs_6; // @[MemPrimitives.scala 121:29:@12624.4]
  wire  StickySelects_8_io_outs_7; // @[MemPrimitives.scala 121:29:@12624.4]
  wire  StickySelects_8_io_outs_8; // @[MemPrimitives.scala 121:29:@12624.4]
  wire  StickySelects_9_clock; // @[MemPrimitives.scala 121:29:@12713.4]
  wire  StickySelects_9_reset; // @[MemPrimitives.scala 121:29:@12713.4]
  wire  StickySelects_9_io_ins_0; // @[MemPrimitives.scala 121:29:@12713.4]
  wire  StickySelects_9_io_ins_1; // @[MemPrimitives.scala 121:29:@12713.4]
  wire  StickySelects_9_io_ins_2; // @[MemPrimitives.scala 121:29:@12713.4]
  wire  StickySelects_9_io_ins_3; // @[MemPrimitives.scala 121:29:@12713.4]
  wire  StickySelects_9_io_ins_4; // @[MemPrimitives.scala 121:29:@12713.4]
  wire  StickySelects_9_io_ins_5; // @[MemPrimitives.scala 121:29:@12713.4]
  wire  StickySelects_9_io_ins_6; // @[MemPrimitives.scala 121:29:@12713.4]
  wire  StickySelects_9_io_ins_7; // @[MemPrimitives.scala 121:29:@12713.4]
  wire  StickySelects_9_io_ins_8; // @[MemPrimitives.scala 121:29:@12713.4]
  wire  StickySelects_9_io_outs_0; // @[MemPrimitives.scala 121:29:@12713.4]
  wire  StickySelects_9_io_outs_1; // @[MemPrimitives.scala 121:29:@12713.4]
  wire  StickySelects_9_io_outs_2; // @[MemPrimitives.scala 121:29:@12713.4]
  wire  StickySelects_9_io_outs_3; // @[MemPrimitives.scala 121:29:@12713.4]
  wire  StickySelects_9_io_outs_4; // @[MemPrimitives.scala 121:29:@12713.4]
  wire  StickySelects_9_io_outs_5; // @[MemPrimitives.scala 121:29:@12713.4]
  wire  StickySelects_9_io_outs_6; // @[MemPrimitives.scala 121:29:@12713.4]
  wire  StickySelects_9_io_outs_7; // @[MemPrimitives.scala 121:29:@12713.4]
  wire  StickySelects_9_io_outs_8; // @[MemPrimitives.scala 121:29:@12713.4]
  wire  StickySelects_10_clock; // @[MemPrimitives.scala 121:29:@12802.4]
  wire  StickySelects_10_reset; // @[MemPrimitives.scala 121:29:@12802.4]
  wire  StickySelects_10_io_ins_0; // @[MemPrimitives.scala 121:29:@12802.4]
  wire  StickySelects_10_io_ins_1; // @[MemPrimitives.scala 121:29:@12802.4]
  wire  StickySelects_10_io_ins_2; // @[MemPrimitives.scala 121:29:@12802.4]
  wire  StickySelects_10_io_ins_3; // @[MemPrimitives.scala 121:29:@12802.4]
  wire  StickySelects_10_io_ins_4; // @[MemPrimitives.scala 121:29:@12802.4]
  wire  StickySelects_10_io_ins_5; // @[MemPrimitives.scala 121:29:@12802.4]
  wire  StickySelects_10_io_ins_6; // @[MemPrimitives.scala 121:29:@12802.4]
  wire  StickySelects_10_io_ins_7; // @[MemPrimitives.scala 121:29:@12802.4]
  wire  StickySelects_10_io_ins_8; // @[MemPrimitives.scala 121:29:@12802.4]
  wire  StickySelects_10_io_outs_0; // @[MemPrimitives.scala 121:29:@12802.4]
  wire  StickySelects_10_io_outs_1; // @[MemPrimitives.scala 121:29:@12802.4]
  wire  StickySelects_10_io_outs_2; // @[MemPrimitives.scala 121:29:@12802.4]
  wire  StickySelects_10_io_outs_3; // @[MemPrimitives.scala 121:29:@12802.4]
  wire  StickySelects_10_io_outs_4; // @[MemPrimitives.scala 121:29:@12802.4]
  wire  StickySelects_10_io_outs_5; // @[MemPrimitives.scala 121:29:@12802.4]
  wire  StickySelects_10_io_outs_6; // @[MemPrimitives.scala 121:29:@12802.4]
  wire  StickySelects_10_io_outs_7; // @[MemPrimitives.scala 121:29:@12802.4]
  wire  StickySelects_10_io_outs_8; // @[MemPrimitives.scala 121:29:@12802.4]
  wire  StickySelects_11_clock; // @[MemPrimitives.scala 121:29:@12891.4]
  wire  StickySelects_11_reset; // @[MemPrimitives.scala 121:29:@12891.4]
  wire  StickySelects_11_io_ins_0; // @[MemPrimitives.scala 121:29:@12891.4]
  wire  StickySelects_11_io_ins_1; // @[MemPrimitives.scala 121:29:@12891.4]
  wire  StickySelects_11_io_ins_2; // @[MemPrimitives.scala 121:29:@12891.4]
  wire  StickySelects_11_io_ins_3; // @[MemPrimitives.scala 121:29:@12891.4]
  wire  StickySelects_11_io_ins_4; // @[MemPrimitives.scala 121:29:@12891.4]
  wire  StickySelects_11_io_ins_5; // @[MemPrimitives.scala 121:29:@12891.4]
  wire  StickySelects_11_io_ins_6; // @[MemPrimitives.scala 121:29:@12891.4]
  wire  StickySelects_11_io_ins_7; // @[MemPrimitives.scala 121:29:@12891.4]
  wire  StickySelects_11_io_ins_8; // @[MemPrimitives.scala 121:29:@12891.4]
  wire  StickySelects_11_io_outs_0; // @[MemPrimitives.scala 121:29:@12891.4]
  wire  StickySelects_11_io_outs_1; // @[MemPrimitives.scala 121:29:@12891.4]
  wire  StickySelects_11_io_outs_2; // @[MemPrimitives.scala 121:29:@12891.4]
  wire  StickySelects_11_io_outs_3; // @[MemPrimitives.scala 121:29:@12891.4]
  wire  StickySelects_11_io_outs_4; // @[MemPrimitives.scala 121:29:@12891.4]
  wire  StickySelects_11_io_outs_5; // @[MemPrimitives.scala 121:29:@12891.4]
  wire  StickySelects_11_io_outs_6; // @[MemPrimitives.scala 121:29:@12891.4]
  wire  StickySelects_11_io_outs_7; // @[MemPrimitives.scala 121:29:@12891.4]
  wire  StickySelects_11_io_outs_8; // @[MemPrimitives.scala 121:29:@12891.4]
  wire  StickySelects_12_clock; // @[MemPrimitives.scala 121:29:@12980.4]
  wire  StickySelects_12_reset; // @[MemPrimitives.scala 121:29:@12980.4]
  wire  StickySelects_12_io_ins_0; // @[MemPrimitives.scala 121:29:@12980.4]
  wire  StickySelects_12_io_ins_1; // @[MemPrimitives.scala 121:29:@12980.4]
  wire  StickySelects_12_io_ins_2; // @[MemPrimitives.scala 121:29:@12980.4]
  wire  StickySelects_12_io_ins_3; // @[MemPrimitives.scala 121:29:@12980.4]
  wire  StickySelects_12_io_ins_4; // @[MemPrimitives.scala 121:29:@12980.4]
  wire  StickySelects_12_io_ins_5; // @[MemPrimitives.scala 121:29:@12980.4]
  wire  StickySelects_12_io_ins_6; // @[MemPrimitives.scala 121:29:@12980.4]
  wire  StickySelects_12_io_ins_7; // @[MemPrimitives.scala 121:29:@12980.4]
  wire  StickySelects_12_io_ins_8; // @[MemPrimitives.scala 121:29:@12980.4]
  wire  StickySelects_12_io_outs_0; // @[MemPrimitives.scala 121:29:@12980.4]
  wire  StickySelects_12_io_outs_1; // @[MemPrimitives.scala 121:29:@12980.4]
  wire  StickySelects_12_io_outs_2; // @[MemPrimitives.scala 121:29:@12980.4]
  wire  StickySelects_12_io_outs_3; // @[MemPrimitives.scala 121:29:@12980.4]
  wire  StickySelects_12_io_outs_4; // @[MemPrimitives.scala 121:29:@12980.4]
  wire  StickySelects_12_io_outs_5; // @[MemPrimitives.scala 121:29:@12980.4]
  wire  StickySelects_12_io_outs_6; // @[MemPrimitives.scala 121:29:@12980.4]
  wire  StickySelects_12_io_outs_7; // @[MemPrimitives.scala 121:29:@12980.4]
  wire  StickySelects_12_io_outs_8; // @[MemPrimitives.scala 121:29:@12980.4]
  wire  StickySelects_13_clock; // @[MemPrimitives.scala 121:29:@13069.4]
  wire  StickySelects_13_reset; // @[MemPrimitives.scala 121:29:@13069.4]
  wire  StickySelects_13_io_ins_0; // @[MemPrimitives.scala 121:29:@13069.4]
  wire  StickySelects_13_io_ins_1; // @[MemPrimitives.scala 121:29:@13069.4]
  wire  StickySelects_13_io_ins_2; // @[MemPrimitives.scala 121:29:@13069.4]
  wire  StickySelects_13_io_ins_3; // @[MemPrimitives.scala 121:29:@13069.4]
  wire  StickySelects_13_io_ins_4; // @[MemPrimitives.scala 121:29:@13069.4]
  wire  StickySelects_13_io_ins_5; // @[MemPrimitives.scala 121:29:@13069.4]
  wire  StickySelects_13_io_ins_6; // @[MemPrimitives.scala 121:29:@13069.4]
  wire  StickySelects_13_io_ins_7; // @[MemPrimitives.scala 121:29:@13069.4]
  wire  StickySelects_13_io_ins_8; // @[MemPrimitives.scala 121:29:@13069.4]
  wire  StickySelects_13_io_outs_0; // @[MemPrimitives.scala 121:29:@13069.4]
  wire  StickySelects_13_io_outs_1; // @[MemPrimitives.scala 121:29:@13069.4]
  wire  StickySelects_13_io_outs_2; // @[MemPrimitives.scala 121:29:@13069.4]
  wire  StickySelects_13_io_outs_3; // @[MemPrimitives.scala 121:29:@13069.4]
  wire  StickySelects_13_io_outs_4; // @[MemPrimitives.scala 121:29:@13069.4]
  wire  StickySelects_13_io_outs_5; // @[MemPrimitives.scala 121:29:@13069.4]
  wire  StickySelects_13_io_outs_6; // @[MemPrimitives.scala 121:29:@13069.4]
  wire  StickySelects_13_io_outs_7; // @[MemPrimitives.scala 121:29:@13069.4]
  wire  StickySelects_13_io_outs_8; // @[MemPrimitives.scala 121:29:@13069.4]
  wire  StickySelects_14_clock; // @[MemPrimitives.scala 121:29:@13158.4]
  wire  StickySelects_14_reset; // @[MemPrimitives.scala 121:29:@13158.4]
  wire  StickySelects_14_io_ins_0; // @[MemPrimitives.scala 121:29:@13158.4]
  wire  StickySelects_14_io_ins_1; // @[MemPrimitives.scala 121:29:@13158.4]
  wire  StickySelects_14_io_ins_2; // @[MemPrimitives.scala 121:29:@13158.4]
  wire  StickySelects_14_io_ins_3; // @[MemPrimitives.scala 121:29:@13158.4]
  wire  StickySelects_14_io_ins_4; // @[MemPrimitives.scala 121:29:@13158.4]
  wire  StickySelects_14_io_ins_5; // @[MemPrimitives.scala 121:29:@13158.4]
  wire  StickySelects_14_io_ins_6; // @[MemPrimitives.scala 121:29:@13158.4]
  wire  StickySelects_14_io_ins_7; // @[MemPrimitives.scala 121:29:@13158.4]
  wire  StickySelects_14_io_ins_8; // @[MemPrimitives.scala 121:29:@13158.4]
  wire  StickySelects_14_io_outs_0; // @[MemPrimitives.scala 121:29:@13158.4]
  wire  StickySelects_14_io_outs_1; // @[MemPrimitives.scala 121:29:@13158.4]
  wire  StickySelects_14_io_outs_2; // @[MemPrimitives.scala 121:29:@13158.4]
  wire  StickySelects_14_io_outs_3; // @[MemPrimitives.scala 121:29:@13158.4]
  wire  StickySelects_14_io_outs_4; // @[MemPrimitives.scala 121:29:@13158.4]
  wire  StickySelects_14_io_outs_5; // @[MemPrimitives.scala 121:29:@13158.4]
  wire  StickySelects_14_io_outs_6; // @[MemPrimitives.scala 121:29:@13158.4]
  wire  StickySelects_14_io_outs_7; // @[MemPrimitives.scala 121:29:@13158.4]
  wire  StickySelects_14_io_outs_8; // @[MemPrimitives.scala 121:29:@13158.4]
  wire  StickySelects_15_clock; // @[MemPrimitives.scala 121:29:@13247.4]
  wire  StickySelects_15_reset; // @[MemPrimitives.scala 121:29:@13247.4]
  wire  StickySelects_15_io_ins_0; // @[MemPrimitives.scala 121:29:@13247.4]
  wire  StickySelects_15_io_ins_1; // @[MemPrimitives.scala 121:29:@13247.4]
  wire  StickySelects_15_io_ins_2; // @[MemPrimitives.scala 121:29:@13247.4]
  wire  StickySelects_15_io_ins_3; // @[MemPrimitives.scala 121:29:@13247.4]
  wire  StickySelects_15_io_ins_4; // @[MemPrimitives.scala 121:29:@13247.4]
  wire  StickySelects_15_io_ins_5; // @[MemPrimitives.scala 121:29:@13247.4]
  wire  StickySelects_15_io_ins_6; // @[MemPrimitives.scala 121:29:@13247.4]
  wire  StickySelects_15_io_ins_7; // @[MemPrimitives.scala 121:29:@13247.4]
  wire  StickySelects_15_io_ins_8; // @[MemPrimitives.scala 121:29:@13247.4]
  wire  StickySelects_15_io_outs_0; // @[MemPrimitives.scala 121:29:@13247.4]
  wire  StickySelects_15_io_outs_1; // @[MemPrimitives.scala 121:29:@13247.4]
  wire  StickySelects_15_io_outs_2; // @[MemPrimitives.scala 121:29:@13247.4]
  wire  StickySelects_15_io_outs_3; // @[MemPrimitives.scala 121:29:@13247.4]
  wire  StickySelects_15_io_outs_4; // @[MemPrimitives.scala 121:29:@13247.4]
  wire  StickySelects_15_io_outs_5; // @[MemPrimitives.scala 121:29:@13247.4]
  wire  StickySelects_15_io_outs_6; // @[MemPrimitives.scala 121:29:@13247.4]
  wire  StickySelects_15_io_outs_7; // @[MemPrimitives.scala 121:29:@13247.4]
  wire  StickySelects_15_io_outs_8; // @[MemPrimitives.scala 121:29:@13247.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@13349.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@13349.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@13349.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@13349.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@13349.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@13357.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@13357.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@13357.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@13357.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@13357.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@13365.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@13365.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@13365.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@13365.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@13365.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@13373.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@13373.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@13373.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@13373.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@13373.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@13381.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@13381.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@13381.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@13381.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@13381.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@13389.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@13389.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@13389.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@13389.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@13389.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@13397.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@13397.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@13397.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@13397.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@13397.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@13405.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@13405.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@13405.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@13405.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@13405.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@13413.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@13413.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@13413.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@13413.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@13413.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@13421.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@13421.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@13421.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@13421.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@13421.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@13429.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@13429.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@13429.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@13429.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@13429.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@13437.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@13437.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@13437.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@13437.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@13437.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@13445.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@13445.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@13445.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@13445.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@13445.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@13453.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@13453.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@13453.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@13453.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@13453.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@13461.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@13461.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@13461.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@13461.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@13461.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@13469.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@13469.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@13469.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@13469.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@13469.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@13541.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@13541.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@13541.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@13541.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@13541.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@13549.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@13549.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@13549.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@13549.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@13549.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@13557.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@13557.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@13557.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@13557.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@13557.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@13565.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@13565.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@13565.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@13565.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@13565.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@13573.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@13573.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@13573.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@13573.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@13573.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@13581.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@13581.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@13581.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@13581.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@13581.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@13589.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@13589.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@13589.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@13589.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@13589.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@13597.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@13597.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@13597.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@13597.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@13597.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@13605.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@13605.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@13605.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@13605.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@13605.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@13613.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@13613.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@13613.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@13613.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@13613.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@13621.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@13621.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@13621.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@13621.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@13621.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@13629.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@13629.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@13629.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@13629.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@13629.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@13637.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@13637.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@13637.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@13637.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@13637.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@13645.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@13645.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@13645.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@13645.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@13645.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@13653.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@13653.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@13653.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@13653.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@13653.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@13661.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@13661.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@13661.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@13661.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@13661.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@13733.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@13733.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@13733.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@13733.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@13733.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@13741.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@13741.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@13741.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@13741.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@13741.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@13749.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@13749.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@13749.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@13749.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@13749.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@13757.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@13757.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@13757.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@13757.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@13757.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@13765.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@13765.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@13765.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@13765.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@13765.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@13773.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@13773.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@13773.4]
  wire  RetimeWrapper_37_io_in; // @[package.scala 93:22:@13773.4]
  wire  RetimeWrapper_37_io_out; // @[package.scala 93:22:@13773.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@13781.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@13781.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@13781.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@13781.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@13781.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@13789.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@13789.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@13789.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@13789.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@13789.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@13797.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@13797.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@13797.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@13797.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@13797.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@13805.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@13805.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@13805.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@13805.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@13805.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@13813.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@13813.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@13813.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@13813.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@13813.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@13821.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@13821.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@13821.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@13821.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@13821.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@13829.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@13829.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@13829.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@13829.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@13829.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@13837.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@13837.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@13837.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@13837.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@13837.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@13845.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@13845.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@13845.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@13845.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@13845.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@13853.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@13853.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@13853.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@13853.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@13853.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@13925.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@13925.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@13925.4]
  wire  RetimeWrapper_48_io_in; // @[package.scala 93:22:@13925.4]
  wire  RetimeWrapper_48_io_out; // @[package.scala 93:22:@13925.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@13933.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@13933.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@13933.4]
  wire  RetimeWrapper_49_io_in; // @[package.scala 93:22:@13933.4]
  wire  RetimeWrapper_49_io_out; // @[package.scala 93:22:@13933.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@13941.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@13941.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@13941.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@13941.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@13941.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@13949.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@13949.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@13949.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@13949.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@13949.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@13957.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@13957.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@13957.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@13957.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@13957.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@13965.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@13965.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@13965.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@13965.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@13965.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@13973.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@13973.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@13973.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@13973.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@13973.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@13981.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@13981.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@13981.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@13981.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@13981.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@13989.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@13989.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@13989.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@13989.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@13989.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@13997.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@13997.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@13997.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@13997.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@13997.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@14005.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@14005.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@14005.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@14005.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@14005.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@14013.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@14013.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@14013.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@14013.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@14013.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@14021.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@14021.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@14021.4]
  wire  RetimeWrapper_60_io_in; // @[package.scala 93:22:@14021.4]
  wire  RetimeWrapper_60_io_out; // @[package.scala 93:22:@14021.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@14029.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@14029.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@14029.4]
  wire  RetimeWrapper_61_io_in; // @[package.scala 93:22:@14029.4]
  wire  RetimeWrapper_61_io_out; // @[package.scala 93:22:@14029.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@14037.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@14037.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@14037.4]
  wire  RetimeWrapper_62_io_in; // @[package.scala 93:22:@14037.4]
  wire  RetimeWrapper_62_io_out; // @[package.scala 93:22:@14037.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@14045.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@14045.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@14045.4]
  wire  RetimeWrapper_63_io_in; // @[package.scala 93:22:@14045.4]
  wire  RetimeWrapper_63_io_out; // @[package.scala 93:22:@14045.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@14117.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@14117.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@14117.4]
  wire  RetimeWrapper_64_io_in; // @[package.scala 93:22:@14117.4]
  wire  RetimeWrapper_64_io_out; // @[package.scala 93:22:@14117.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@14125.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@14125.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@14125.4]
  wire  RetimeWrapper_65_io_in; // @[package.scala 93:22:@14125.4]
  wire  RetimeWrapper_65_io_out; // @[package.scala 93:22:@14125.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@14133.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@14133.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@14133.4]
  wire  RetimeWrapper_66_io_in; // @[package.scala 93:22:@14133.4]
  wire  RetimeWrapper_66_io_out; // @[package.scala 93:22:@14133.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@14141.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@14141.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@14141.4]
  wire  RetimeWrapper_67_io_in; // @[package.scala 93:22:@14141.4]
  wire  RetimeWrapper_67_io_out; // @[package.scala 93:22:@14141.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@14149.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@14149.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@14149.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@14149.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@14149.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@14157.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@14157.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@14157.4]
  wire  RetimeWrapper_69_io_in; // @[package.scala 93:22:@14157.4]
  wire  RetimeWrapper_69_io_out; // @[package.scala 93:22:@14157.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@14165.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@14165.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@14165.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@14165.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@14165.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@14173.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@14173.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@14173.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@14173.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@14173.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@14181.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@14181.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@14181.4]
  wire  RetimeWrapper_72_io_in; // @[package.scala 93:22:@14181.4]
  wire  RetimeWrapper_72_io_out; // @[package.scala 93:22:@14181.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@14189.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@14189.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@14189.4]
  wire  RetimeWrapper_73_io_in; // @[package.scala 93:22:@14189.4]
  wire  RetimeWrapper_73_io_out; // @[package.scala 93:22:@14189.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@14197.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@14197.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@14197.4]
  wire  RetimeWrapper_74_io_in; // @[package.scala 93:22:@14197.4]
  wire  RetimeWrapper_74_io_out; // @[package.scala 93:22:@14197.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@14205.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@14205.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@14205.4]
  wire  RetimeWrapper_75_io_in; // @[package.scala 93:22:@14205.4]
  wire  RetimeWrapper_75_io_out; // @[package.scala 93:22:@14205.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@14213.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@14213.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@14213.4]
  wire  RetimeWrapper_76_io_in; // @[package.scala 93:22:@14213.4]
  wire  RetimeWrapper_76_io_out; // @[package.scala 93:22:@14213.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@14221.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@14221.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@14221.4]
  wire  RetimeWrapper_77_io_in; // @[package.scala 93:22:@14221.4]
  wire  RetimeWrapper_77_io_out; // @[package.scala 93:22:@14221.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@14229.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@14229.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@14229.4]
  wire  RetimeWrapper_78_io_in; // @[package.scala 93:22:@14229.4]
  wire  RetimeWrapper_78_io_out; // @[package.scala 93:22:@14229.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@14237.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@14237.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@14237.4]
  wire  RetimeWrapper_79_io_in; // @[package.scala 93:22:@14237.4]
  wire  RetimeWrapper_79_io_out; // @[package.scala 93:22:@14237.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@14309.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@14309.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@14309.4]
  wire  RetimeWrapper_80_io_in; // @[package.scala 93:22:@14309.4]
  wire  RetimeWrapper_80_io_out; // @[package.scala 93:22:@14309.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@14317.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@14317.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@14317.4]
  wire  RetimeWrapper_81_io_in; // @[package.scala 93:22:@14317.4]
  wire  RetimeWrapper_81_io_out; // @[package.scala 93:22:@14317.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@14325.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@14325.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@14325.4]
  wire  RetimeWrapper_82_io_in; // @[package.scala 93:22:@14325.4]
  wire  RetimeWrapper_82_io_out; // @[package.scala 93:22:@14325.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@14333.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@14333.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@14333.4]
  wire  RetimeWrapper_83_io_in; // @[package.scala 93:22:@14333.4]
  wire  RetimeWrapper_83_io_out; // @[package.scala 93:22:@14333.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@14341.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@14341.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@14341.4]
  wire  RetimeWrapper_84_io_in; // @[package.scala 93:22:@14341.4]
  wire  RetimeWrapper_84_io_out; // @[package.scala 93:22:@14341.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@14349.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@14349.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@14349.4]
  wire  RetimeWrapper_85_io_in; // @[package.scala 93:22:@14349.4]
  wire  RetimeWrapper_85_io_out; // @[package.scala 93:22:@14349.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@14357.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@14357.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@14357.4]
  wire  RetimeWrapper_86_io_in; // @[package.scala 93:22:@14357.4]
  wire  RetimeWrapper_86_io_out; // @[package.scala 93:22:@14357.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@14365.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@14365.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@14365.4]
  wire  RetimeWrapper_87_io_in; // @[package.scala 93:22:@14365.4]
  wire  RetimeWrapper_87_io_out; // @[package.scala 93:22:@14365.4]
  wire  RetimeWrapper_88_clock; // @[package.scala 93:22:@14373.4]
  wire  RetimeWrapper_88_reset; // @[package.scala 93:22:@14373.4]
  wire  RetimeWrapper_88_io_flow; // @[package.scala 93:22:@14373.4]
  wire  RetimeWrapper_88_io_in; // @[package.scala 93:22:@14373.4]
  wire  RetimeWrapper_88_io_out; // @[package.scala 93:22:@14373.4]
  wire  RetimeWrapper_89_clock; // @[package.scala 93:22:@14381.4]
  wire  RetimeWrapper_89_reset; // @[package.scala 93:22:@14381.4]
  wire  RetimeWrapper_89_io_flow; // @[package.scala 93:22:@14381.4]
  wire  RetimeWrapper_89_io_in; // @[package.scala 93:22:@14381.4]
  wire  RetimeWrapper_89_io_out; // @[package.scala 93:22:@14381.4]
  wire  RetimeWrapper_90_clock; // @[package.scala 93:22:@14389.4]
  wire  RetimeWrapper_90_reset; // @[package.scala 93:22:@14389.4]
  wire  RetimeWrapper_90_io_flow; // @[package.scala 93:22:@14389.4]
  wire  RetimeWrapper_90_io_in; // @[package.scala 93:22:@14389.4]
  wire  RetimeWrapper_90_io_out; // @[package.scala 93:22:@14389.4]
  wire  RetimeWrapper_91_clock; // @[package.scala 93:22:@14397.4]
  wire  RetimeWrapper_91_reset; // @[package.scala 93:22:@14397.4]
  wire  RetimeWrapper_91_io_flow; // @[package.scala 93:22:@14397.4]
  wire  RetimeWrapper_91_io_in; // @[package.scala 93:22:@14397.4]
  wire  RetimeWrapper_91_io_out; // @[package.scala 93:22:@14397.4]
  wire  RetimeWrapper_92_clock; // @[package.scala 93:22:@14405.4]
  wire  RetimeWrapper_92_reset; // @[package.scala 93:22:@14405.4]
  wire  RetimeWrapper_92_io_flow; // @[package.scala 93:22:@14405.4]
  wire  RetimeWrapper_92_io_in; // @[package.scala 93:22:@14405.4]
  wire  RetimeWrapper_92_io_out; // @[package.scala 93:22:@14405.4]
  wire  RetimeWrapper_93_clock; // @[package.scala 93:22:@14413.4]
  wire  RetimeWrapper_93_reset; // @[package.scala 93:22:@14413.4]
  wire  RetimeWrapper_93_io_flow; // @[package.scala 93:22:@14413.4]
  wire  RetimeWrapper_93_io_in; // @[package.scala 93:22:@14413.4]
  wire  RetimeWrapper_93_io_out; // @[package.scala 93:22:@14413.4]
  wire  RetimeWrapper_94_clock; // @[package.scala 93:22:@14421.4]
  wire  RetimeWrapper_94_reset; // @[package.scala 93:22:@14421.4]
  wire  RetimeWrapper_94_io_flow; // @[package.scala 93:22:@14421.4]
  wire  RetimeWrapper_94_io_in; // @[package.scala 93:22:@14421.4]
  wire  RetimeWrapper_94_io_out; // @[package.scala 93:22:@14421.4]
  wire  RetimeWrapper_95_clock; // @[package.scala 93:22:@14429.4]
  wire  RetimeWrapper_95_reset; // @[package.scala 93:22:@14429.4]
  wire  RetimeWrapper_95_io_flow; // @[package.scala 93:22:@14429.4]
  wire  RetimeWrapper_95_io_in; // @[package.scala 93:22:@14429.4]
  wire  RetimeWrapper_95_io_out; // @[package.scala 93:22:@14429.4]
  wire  RetimeWrapper_96_clock; // @[package.scala 93:22:@14501.4]
  wire  RetimeWrapper_96_reset; // @[package.scala 93:22:@14501.4]
  wire  RetimeWrapper_96_io_flow; // @[package.scala 93:22:@14501.4]
  wire  RetimeWrapper_96_io_in; // @[package.scala 93:22:@14501.4]
  wire  RetimeWrapper_96_io_out; // @[package.scala 93:22:@14501.4]
  wire  RetimeWrapper_97_clock; // @[package.scala 93:22:@14509.4]
  wire  RetimeWrapper_97_reset; // @[package.scala 93:22:@14509.4]
  wire  RetimeWrapper_97_io_flow; // @[package.scala 93:22:@14509.4]
  wire  RetimeWrapper_97_io_in; // @[package.scala 93:22:@14509.4]
  wire  RetimeWrapper_97_io_out; // @[package.scala 93:22:@14509.4]
  wire  RetimeWrapper_98_clock; // @[package.scala 93:22:@14517.4]
  wire  RetimeWrapper_98_reset; // @[package.scala 93:22:@14517.4]
  wire  RetimeWrapper_98_io_flow; // @[package.scala 93:22:@14517.4]
  wire  RetimeWrapper_98_io_in; // @[package.scala 93:22:@14517.4]
  wire  RetimeWrapper_98_io_out; // @[package.scala 93:22:@14517.4]
  wire  RetimeWrapper_99_clock; // @[package.scala 93:22:@14525.4]
  wire  RetimeWrapper_99_reset; // @[package.scala 93:22:@14525.4]
  wire  RetimeWrapper_99_io_flow; // @[package.scala 93:22:@14525.4]
  wire  RetimeWrapper_99_io_in; // @[package.scala 93:22:@14525.4]
  wire  RetimeWrapper_99_io_out; // @[package.scala 93:22:@14525.4]
  wire  RetimeWrapper_100_clock; // @[package.scala 93:22:@14533.4]
  wire  RetimeWrapper_100_reset; // @[package.scala 93:22:@14533.4]
  wire  RetimeWrapper_100_io_flow; // @[package.scala 93:22:@14533.4]
  wire  RetimeWrapper_100_io_in; // @[package.scala 93:22:@14533.4]
  wire  RetimeWrapper_100_io_out; // @[package.scala 93:22:@14533.4]
  wire  RetimeWrapper_101_clock; // @[package.scala 93:22:@14541.4]
  wire  RetimeWrapper_101_reset; // @[package.scala 93:22:@14541.4]
  wire  RetimeWrapper_101_io_flow; // @[package.scala 93:22:@14541.4]
  wire  RetimeWrapper_101_io_in; // @[package.scala 93:22:@14541.4]
  wire  RetimeWrapper_101_io_out; // @[package.scala 93:22:@14541.4]
  wire  RetimeWrapper_102_clock; // @[package.scala 93:22:@14549.4]
  wire  RetimeWrapper_102_reset; // @[package.scala 93:22:@14549.4]
  wire  RetimeWrapper_102_io_flow; // @[package.scala 93:22:@14549.4]
  wire  RetimeWrapper_102_io_in; // @[package.scala 93:22:@14549.4]
  wire  RetimeWrapper_102_io_out; // @[package.scala 93:22:@14549.4]
  wire  RetimeWrapper_103_clock; // @[package.scala 93:22:@14557.4]
  wire  RetimeWrapper_103_reset; // @[package.scala 93:22:@14557.4]
  wire  RetimeWrapper_103_io_flow; // @[package.scala 93:22:@14557.4]
  wire  RetimeWrapper_103_io_in; // @[package.scala 93:22:@14557.4]
  wire  RetimeWrapper_103_io_out; // @[package.scala 93:22:@14557.4]
  wire  RetimeWrapper_104_clock; // @[package.scala 93:22:@14565.4]
  wire  RetimeWrapper_104_reset; // @[package.scala 93:22:@14565.4]
  wire  RetimeWrapper_104_io_flow; // @[package.scala 93:22:@14565.4]
  wire  RetimeWrapper_104_io_in; // @[package.scala 93:22:@14565.4]
  wire  RetimeWrapper_104_io_out; // @[package.scala 93:22:@14565.4]
  wire  RetimeWrapper_105_clock; // @[package.scala 93:22:@14573.4]
  wire  RetimeWrapper_105_reset; // @[package.scala 93:22:@14573.4]
  wire  RetimeWrapper_105_io_flow; // @[package.scala 93:22:@14573.4]
  wire  RetimeWrapper_105_io_in; // @[package.scala 93:22:@14573.4]
  wire  RetimeWrapper_105_io_out; // @[package.scala 93:22:@14573.4]
  wire  RetimeWrapper_106_clock; // @[package.scala 93:22:@14581.4]
  wire  RetimeWrapper_106_reset; // @[package.scala 93:22:@14581.4]
  wire  RetimeWrapper_106_io_flow; // @[package.scala 93:22:@14581.4]
  wire  RetimeWrapper_106_io_in; // @[package.scala 93:22:@14581.4]
  wire  RetimeWrapper_106_io_out; // @[package.scala 93:22:@14581.4]
  wire  RetimeWrapper_107_clock; // @[package.scala 93:22:@14589.4]
  wire  RetimeWrapper_107_reset; // @[package.scala 93:22:@14589.4]
  wire  RetimeWrapper_107_io_flow; // @[package.scala 93:22:@14589.4]
  wire  RetimeWrapper_107_io_in; // @[package.scala 93:22:@14589.4]
  wire  RetimeWrapper_107_io_out; // @[package.scala 93:22:@14589.4]
  wire  RetimeWrapper_108_clock; // @[package.scala 93:22:@14597.4]
  wire  RetimeWrapper_108_reset; // @[package.scala 93:22:@14597.4]
  wire  RetimeWrapper_108_io_flow; // @[package.scala 93:22:@14597.4]
  wire  RetimeWrapper_108_io_in; // @[package.scala 93:22:@14597.4]
  wire  RetimeWrapper_108_io_out; // @[package.scala 93:22:@14597.4]
  wire  RetimeWrapper_109_clock; // @[package.scala 93:22:@14605.4]
  wire  RetimeWrapper_109_reset; // @[package.scala 93:22:@14605.4]
  wire  RetimeWrapper_109_io_flow; // @[package.scala 93:22:@14605.4]
  wire  RetimeWrapper_109_io_in; // @[package.scala 93:22:@14605.4]
  wire  RetimeWrapper_109_io_out; // @[package.scala 93:22:@14605.4]
  wire  RetimeWrapper_110_clock; // @[package.scala 93:22:@14613.4]
  wire  RetimeWrapper_110_reset; // @[package.scala 93:22:@14613.4]
  wire  RetimeWrapper_110_io_flow; // @[package.scala 93:22:@14613.4]
  wire  RetimeWrapper_110_io_in; // @[package.scala 93:22:@14613.4]
  wire  RetimeWrapper_110_io_out; // @[package.scala 93:22:@14613.4]
  wire  RetimeWrapper_111_clock; // @[package.scala 93:22:@14621.4]
  wire  RetimeWrapper_111_reset; // @[package.scala 93:22:@14621.4]
  wire  RetimeWrapper_111_io_flow; // @[package.scala 93:22:@14621.4]
  wire  RetimeWrapper_111_io_in; // @[package.scala 93:22:@14621.4]
  wire  RetimeWrapper_111_io_out; // @[package.scala 93:22:@14621.4]
  wire  RetimeWrapper_112_clock; // @[package.scala 93:22:@14693.4]
  wire  RetimeWrapper_112_reset; // @[package.scala 93:22:@14693.4]
  wire  RetimeWrapper_112_io_flow; // @[package.scala 93:22:@14693.4]
  wire  RetimeWrapper_112_io_in; // @[package.scala 93:22:@14693.4]
  wire  RetimeWrapper_112_io_out; // @[package.scala 93:22:@14693.4]
  wire  RetimeWrapper_113_clock; // @[package.scala 93:22:@14701.4]
  wire  RetimeWrapper_113_reset; // @[package.scala 93:22:@14701.4]
  wire  RetimeWrapper_113_io_flow; // @[package.scala 93:22:@14701.4]
  wire  RetimeWrapper_113_io_in; // @[package.scala 93:22:@14701.4]
  wire  RetimeWrapper_113_io_out; // @[package.scala 93:22:@14701.4]
  wire  RetimeWrapper_114_clock; // @[package.scala 93:22:@14709.4]
  wire  RetimeWrapper_114_reset; // @[package.scala 93:22:@14709.4]
  wire  RetimeWrapper_114_io_flow; // @[package.scala 93:22:@14709.4]
  wire  RetimeWrapper_114_io_in; // @[package.scala 93:22:@14709.4]
  wire  RetimeWrapper_114_io_out; // @[package.scala 93:22:@14709.4]
  wire  RetimeWrapper_115_clock; // @[package.scala 93:22:@14717.4]
  wire  RetimeWrapper_115_reset; // @[package.scala 93:22:@14717.4]
  wire  RetimeWrapper_115_io_flow; // @[package.scala 93:22:@14717.4]
  wire  RetimeWrapper_115_io_in; // @[package.scala 93:22:@14717.4]
  wire  RetimeWrapper_115_io_out; // @[package.scala 93:22:@14717.4]
  wire  RetimeWrapper_116_clock; // @[package.scala 93:22:@14725.4]
  wire  RetimeWrapper_116_reset; // @[package.scala 93:22:@14725.4]
  wire  RetimeWrapper_116_io_flow; // @[package.scala 93:22:@14725.4]
  wire  RetimeWrapper_116_io_in; // @[package.scala 93:22:@14725.4]
  wire  RetimeWrapper_116_io_out; // @[package.scala 93:22:@14725.4]
  wire  RetimeWrapper_117_clock; // @[package.scala 93:22:@14733.4]
  wire  RetimeWrapper_117_reset; // @[package.scala 93:22:@14733.4]
  wire  RetimeWrapper_117_io_flow; // @[package.scala 93:22:@14733.4]
  wire  RetimeWrapper_117_io_in; // @[package.scala 93:22:@14733.4]
  wire  RetimeWrapper_117_io_out; // @[package.scala 93:22:@14733.4]
  wire  RetimeWrapper_118_clock; // @[package.scala 93:22:@14741.4]
  wire  RetimeWrapper_118_reset; // @[package.scala 93:22:@14741.4]
  wire  RetimeWrapper_118_io_flow; // @[package.scala 93:22:@14741.4]
  wire  RetimeWrapper_118_io_in; // @[package.scala 93:22:@14741.4]
  wire  RetimeWrapper_118_io_out; // @[package.scala 93:22:@14741.4]
  wire  RetimeWrapper_119_clock; // @[package.scala 93:22:@14749.4]
  wire  RetimeWrapper_119_reset; // @[package.scala 93:22:@14749.4]
  wire  RetimeWrapper_119_io_flow; // @[package.scala 93:22:@14749.4]
  wire  RetimeWrapper_119_io_in; // @[package.scala 93:22:@14749.4]
  wire  RetimeWrapper_119_io_out; // @[package.scala 93:22:@14749.4]
  wire  RetimeWrapper_120_clock; // @[package.scala 93:22:@14757.4]
  wire  RetimeWrapper_120_reset; // @[package.scala 93:22:@14757.4]
  wire  RetimeWrapper_120_io_flow; // @[package.scala 93:22:@14757.4]
  wire  RetimeWrapper_120_io_in; // @[package.scala 93:22:@14757.4]
  wire  RetimeWrapper_120_io_out; // @[package.scala 93:22:@14757.4]
  wire  RetimeWrapper_121_clock; // @[package.scala 93:22:@14765.4]
  wire  RetimeWrapper_121_reset; // @[package.scala 93:22:@14765.4]
  wire  RetimeWrapper_121_io_flow; // @[package.scala 93:22:@14765.4]
  wire  RetimeWrapper_121_io_in; // @[package.scala 93:22:@14765.4]
  wire  RetimeWrapper_121_io_out; // @[package.scala 93:22:@14765.4]
  wire  RetimeWrapper_122_clock; // @[package.scala 93:22:@14773.4]
  wire  RetimeWrapper_122_reset; // @[package.scala 93:22:@14773.4]
  wire  RetimeWrapper_122_io_flow; // @[package.scala 93:22:@14773.4]
  wire  RetimeWrapper_122_io_in; // @[package.scala 93:22:@14773.4]
  wire  RetimeWrapper_122_io_out; // @[package.scala 93:22:@14773.4]
  wire  RetimeWrapper_123_clock; // @[package.scala 93:22:@14781.4]
  wire  RetimeWrapper_123_reset; // @[package.scala 93:22:@14781.4]
  wire  RetimeWrapper_123_io_flow; // @[package.scala 93:22:@14781.4]
  wire  RetimeWrapper_123_io_in; // @[package.scala 93:22:@14781.4]
  wire  RetimeWrapper_123_io_out; // @[package.scala 93:22:@14781.4]
  wire  RetimeWrapper_124_clock; // @[package.scala 93:22:@14789.4]
  wire  RetimeWrapper_124_reset; // @[package.scala 93:22:@14789.4]
  wire  RetimeWrapper_124_io_flow; // @[package.scala 93:22:@14789.4]
  wire  RetimeWrapper_124_io_in; // @[package.scala 93:22:@14789.4]
  wire  RetimeWrapper_124_io_out; // @[package.scala 93:22:@14789.4]
  wire  RetimeWrapper_125_clock; // @[package.scala 93:22:@14797.4]
  wire  RetimeWrapper_125_reset; // @[package.scala 93:22:@14797.4]
  wire  RetimeWrapper_125_io_flow; // @[package.scala 93:22:@14797.4]
  wire  RetimeWrapper_125_io_in; // @[package.scala 93:22:@14797.4]
  wire  RetimeWrapper_125_io_out; // @[package.scala 93:22:@14797.4]
  wire  RetimeWrapper_126_clock; // @[package.scala 93:22:@14805.4]
  wire  RetimeWrapper_126_reset; // @[package.scala 93:22:@14805.4]
  wire  RetimeWrapper_126_io_flow; // @[package.scala 93:22:@14805.4]
  wire  RetimeWrapper_126_io_in; // @[package.scala 93:22:@14805.4]
  wire  RetimeWrapper_126_io_out; // @[package.scala 93:22:@14805.4]
  wire  RetimeWrapper_127_clock; // @[package.scala 93:22:@14813.4]
  wire  RetimeWrapper_127_reset; // @[package.scala 93:22:@14813.4]
  wire  RetimeWrapper_127_io_flow; // @[package.scala 93:22:@14813.4]
  wire  RetimeWrapper_127_io_in; // @[package.scala 93:22:@14813.4]
  wire  RetimeWrapper_127_io_out; // @[package.scala 93:22:@14813.4]
  wire  RetimeWrapper_128_clock; // @[package.scala 93:22:@14885.4]
  wire  RetimeWrapper_128_reset; // @[package.scala 93:22:@14885.4]
  wire  RetimeWrapper_128_io_flow; // @[package.scala 93:22:@14885.4]
  wire  RetimeWrapper_128_io_in; // @[package.scala 93:22:@14885.4]
  wire  RetimeWrapper_128_io_out; // @[package.scala 93:22:@14885.4]
  wire  RetimeWrapper_129_clock; // @[package.scala 93:22:@14893.4]
  wire  RetimeWrapper_129_reset; // @[package.scala 93:22:@14893.4]
  wire  RetimeWrapper_129_io_flow; // @[package.scala 93:22:@14893.4]
  wire  RetimeWrapper_129_io_in; // @[package.scala 93:22:@14893.4]
  wire  RetimeWrapper_129_io_out; // @[package.scala 93:22:@14893.4]
  wire  RetimeWrapper_130_clock; // @[package.scala 93:22:@14901.4]
  wire  RetimeWrapper_130_reset; // @[package.scala 93:22:@14901.4]
  wire  RetimeWrapper_130_io_flow; // @[package.scala 93:22:@14901.4]
  wire  RetimeWrapper_130_io_in; // @[package.scala 93:22:@14901.4]
  wire  RetimeWrapper_130_io_out; // @[package.scala 93:22:@14901.4]
  wire  RetimeWrapper_131_clock; // @[package.scala 93:22:@14909.4]
  wire  RetimeWrapper_131_reset; // @[package.scala 93:22:@14909.4]
  wire  RetimeWrapper_131_io_flow; // @[package.scala 93:22:@14909.4]
  wire  RetimeWrapper_131_io_in; // @[package.scala 93:22:@14909.4]
  wire  RetimeWrapper_131_io_out; // @[package.scala 93:22:@14909.4]
  wire  RetimeWrapper_132_clock; // @[package.scala 93:22:@14917.4]
  wire  RetimeWrapper_132_reset; // @[package.scala 93:22:@14917.4]
  wire  RetimeWrapper_132_io_flow; // @[package.scala 93:22:@14917.4]
  wire  RetimeWrapper_132_io_in; // @[package.scala 93:22:@14917.4]
  wire  RetimeWrapper_132_io_out; // @[package.scala 93:22:@14917.4]
  wire  RetimeWrapper_133_clock; // @[package.scala 93:22:@14925.4]
  wire  RetimeWrapper_133_reset; // @[package.scala 93:22:@14925.4]
  wire  RetimeWrapper_133_io_flow; // @[package.scala 93:22:@14925.4]
  wire  RetimeWrapper_133_io_in; // @[package.scala 93:22:@14925.4]
  wire  RetimeWrapper_133_io_out; // @[package.scala 93:22:@14925.4]
  wire  RetimeWrapper_134_clock; // @[package.scala 93:22:@14933.4]
  wire  RetimeWrapper_134_reset; // @[package.scala 93:22:@14933.4]
  wire  RetimeWrapper_134_io_flow; // @[package.scala 93:22:@14933.4]
  wire  RetimeWrapper_134_io_in; // @[package.scala 93:22:@14933.4]
  wire  RetimeWrapper_134_io_out; // @[package.scala 93:22:@14933.4]
  wire  RetimeWrapper_135_clock; // @[package.scala 93:22:@14941.4]
  wire  RetimeWrapper_135_reset; // @[package.scala 93:22:@14941.4]
  wire  RetimeWrapper_135_io_flow; // @[package.scala 93:22:@14941.4]
  wire  RetimeWrapper_135_io_in; // @[package.scala 93:22:@14941.4]
  wire  RetimeWrapper_135_io_out; // @[package.scala 93:22:@14941.4]
  wire  RetimeWrapper_136_clock; // @[package.scala 93:22:@14949.4]
  wire  RetimeWrapper_136_reset; // @[package.scala 93:22:@14949.4]
  wire  RetimeWrapper_136_io_flow; // @[package.scala 93:22:@14949.4]
  wire  RetimeWrapper_136_io_in; // @[package.scala 93:22:@14949.4]
  wire  RetimeWrapper_136_io_out; // @[package.scala 93:22:@14949.4]
  wire  RetimeWrapper_137_clock; // @[package.scala 93:22:@14957.4]
  wire  RetimeWrapper_137_reset; // @[package.scala 93:22:@14957.4]
  wire  RetimeWrapper_137_io_flow; // @[package.scala 93:22:@14957.4]
  wire  RetimeWrapper_137_io_in; // @[package.scala 93:22:@14957.4]
  wire  RetimeWrapper_137_io_out; // @[package.scala 93:22:@14957.4]
  wire  RetimeWrapper_138_clock; // @[package.scala 93:22:@14965.4]
  wire  RetimeWrapper_138_reset; // @[package.scala 93:22:@14965.4]
  wire  RetimeWrapper_138_io_flow; // @[package.scala 93:22:@14965.4]
  wire  RetimeWrapper_138_io_in; // @[package.scala 93:22:@14965.4]
  wire  RetimeWrapper_138_io_out; // @[package.scala 93:22:@14965.4]
  wire  RetimeWrapper_139_clock; // @[package.scala 93:22:@14973.4]
  wire  RetimeWrapper_139_reset; // @[package.scala 93:22:@14973.4]
  wire  RetimeWrapper_139_io_flow; // @[package.scala 93:22:@14973.4]
  wire  RetimeWrapper_139_io_in; // @[package.scala 93:22:@14973.4]
  wire  RetimeWrapper_139_io_out; // @[package.scala 93:22:@14973.4]
  wire  RetimeWrapper_140_clock; // @[package.scala 93:22:@14981.4]
  wire  RetimeWrapper_140_reset; // @[package.scala 93:22:@14981.4]
  wire  RetimeWrapper_140_io_flow; // @[package.scala 93:22:@14981.4]
  wire  RetimeWrapper_140_io_in; // @[package.scala 93:22:@14981.4]
  wire  RetimeWrapper_140_io_out; // @[package.scala 93:22:@14981.4]
  wire  RetimeWrapper_141_clock; // @[package.scala 93:22:@14989.4]
  wire  RetimeWrapper_141_reset; // @[package.scala 93:22:@14989.4]
  wire  RetimeWrapper_141_io_flow; // @[package.scala 93:22:@14989.4]
  wire  RetimeWrapper_141_io_in; // @[package.scala 93:22:@14989.4]
  wire  RetimeWrapper_141_io_out; // @[package.scala 93:22:@14989.4]
  wire  RetimeWrapper_142_clock; // @[package.scala 93:22:@14997.4]
  wire  RetimeWrapper_142_reset; // @[package.scala 93:22:@14997.4]
  wire  RetimeWrapper_142_io_flow; // @[package.scala 93:22:@14997.4]
  wire  RetimeWrapper_142_io_in; // @[package.scala 93:22:@14997.4]
  wire  RetimeWrapper_142_io_out; // @[package.scala 93:22:@14997.4]
  wire  RetimeWrapper_143_clock; // @[package.scala 93:22:@15005.4]
  wire  RetimeWrapper_143_reset; // @[package.scala 93:22:@15005.4]
  wire  RetimeWrapper_143_io_flow; // @[package.scala 93:22:@15005.4]
  wire  RetimeWrapper_143_io_in; // @[package.scala 93:22:@15005.4]
  wire  RetimeWrapper_143_io_out; // @[package.scala 93:22:@15005.4]
  wire  _T_316; // @[MemPrimitives.scala 82:210:@11684.4]
  wire  _T_318; // @[MemPrimitives.scala 82:210:@11685.4]
  wire  _T_319; // @[MemPrimitives.scala 82:228:@11686.4]
  wire  _T_320; // @[MemPrimitives.scala 83:102:@11687.4]
  wire [9:0] _T_322; // @[Cat.scala 30:58:@11689.4]
  wire  _T_329; // @[MemPrimitives.scala 82:210:@11697.4]
  wire  _T_330; // @[MemPrimitives.scala 82:228:@11698.4]
  wire  _T_331; // @[MemPrimitives.scala 83:102:@11699.4]
  wire [9:0] _T_333; // @[Cat.scala 30:58:@11701.4]
  wire  _T_340; // @[MemPrimitives.scala 82:210:@11709.4]
  wire  _T_341; // @[MemPrimitives.scala 82:228:@11710.4]
  wire  _T_342; // @[MemPrimitives.scala 83:102:@11711.4]
  wire [9:0] _T_344; // @[Cat.scala 30:58:@11713.4]
  wire  _T_351; // @[MemPrimitives.scala 82:210:@11721.4]
  wire  _T_352; // @[MemPrimitives.scala 82:228:@11722.4]
  wire  _T_353; // @[MemPrimitives.scala 83:102:@11723.4]
  wire [9:0] _T_355; // @[Cat.scala 30:58:@11725.4]
  wire  _T_360; // @[MemPrimitives.scala 82:210:@11732.4]
  wire  _T_363; // @[MemPrimitives.scala 82:228:@11734.4]
  wire  _T_364; // @[MemPrimitives.scala 83:102:@11735.4]
  wire [9:0] _T_366; // @[Cat.scala 30:58:@11737.4]
  wire  _T_374; // @[MemPrimitives.scala 82:228:@11746.4]
  wire  _T_375; // @[MemPrimitives.scala 83:102:@11747.4]
  wire [9:0] _T_377; // @[Cat.scala 30:58:@11749.4]
  wire  _T_385; // @[MemPrimitives.scala 82:228:@11758.4]
  wire  _T_386; // @[MemPrimitives.scala 83:102:@11759.4]
  wire [9:0] _T_388; // @[Cat.scala 30:58:@11761.4]
  wire  _T_396; // @[MemPrimitives.scala 82:228:@11770.4]
  wire  _T_397; // @[MemPrimitives.scala 83:102:@11771.4]
  wire [9:0] _T_399; // @[Cat.scala 30:58:@11773.4]
  wire  _T_404; // @[MemPrimitives.scala 82:210:@11780.4]
  wire  _T_407; // @[MemPrimitives.scala 82:228:@11782.4]
  wire  _T_408; // @[MemPrimitives.scala 83:102:@11783.4]
  wire [9:0] _T_410; // @[Cat.scala 30:58:@11785.4]
  wire  _T_418; // @[MemPrimitives.scala 82:228:@11794.4]
  wire  _T_419; // @[MemPrimitives.scala 83:102:@11795.4]
  wire [9:0] _T_421; // @[Cat.scala 30:58:@11797.4]
  wire  _T_429; // @[MemPrimitives.scala 82:228:@11806.4]
  wire  _T_430; // @[MemPrimitives.scala 83:102:@11807.4]
  wire [9:0] _T_432; // @[Cat.scala 30:58:@11809.4]
  wire  _T_440; // @[MemPrimitives.scala 82:228:@11818.4]
  wire  _T_441; // @[MemPrimitives.scala 83:102:@11819.4]
  wire [9:0] _T_443; // @[Cat.scala 30:58:@11821.4]
  wire  _T_448; // @[MemPrimitives.scala 82:210:@11828.4]
  wire  _T_451; // @[MemPrimitives.scala 82:228:@11830.4]
  wire  _T_452; // @[MemPrimitives.scala 83:102:@11831.4]
  wire [9:0] _T_454; // @[Cat.scala 30:58:@11833.4]
  wire  _T_462; // @[MemPrimitives.scala 82:228:@11842.4]
  wire  _T_463; // @[MemPrimitives.scala 83:102:@11843.4]
  wire [9:0] _T_465; // @[Cat.scala 30:58:@11845.4]
  wire  _T_473; // @[MemPrimitives.scala 82:228:@11854.4]
  wire  _T_474; // @[MemPrimitives.scala 83:102:@11855.4]
  wire [9:0] _T_476; // @[Cat.scala 30:58:@11857.4]
  wire  _T_484; // @[MemPrimitives.scala 82:228:@11866.4]
  wire  _T_485; // @[MemPrimitives.scala 83:102:@11867.4]
  wire [9:0] _T_487; // @[Cat.scala 30:58:@11869.4]
  wire  _T_492; // @[MemPrimitives.scala 110:210:@11876.4]
  wire  _T_494; // @[MemPrimitives.scala 110:210:@11877.4]
  wire  _T_495; // @[MemPrimitives.scala 110:228:@11878.4]
  wire  _T_498; // @[MemPrimitives.scala 110:210:@11880.4]
  wire  _T_500; // @[MemPrimitives.scala 110:210:@11881.4]
  wire  _T_501; // @[MemPrimitives.scala 110:228:@11882.4]
  wire  _T_504; // @[MemPrimitives.scala 110:210:@11884.4]
  wire  _T_506; // @[MemPrimitives.scala 110:210:@11885.4]
  wire  _T_507; // @[MemPrimitives.scala 110:228:@11886.4]
  wire  _T_510; // @[MemPrimitives.scala 110:210:@11888.4]
  wire  _T_512; // @[MemPrimitives.scala 110:210:@11889.4]
  wire  _T_513; // @[MemPrimitives.scala 110:228:@11890.4]
  wire  _T_516; // @[MemPrimitives.scala 110:210:@11892.4]
  wire  _T_518; // @[MemPrimitives.scala 110:210:@11893.4]
  wire  _T_519; // @[MemPrimitives.scala 110:228:@11894.4]
  wire  _T_522; // @[MemPrimitives.scala 110:210:@11896.4]
  wire  _T_524; // @[MemPrimitives.scala 110:210:@11897.4]
  wire  _T_525; // @[MemPrimitives.scala 110:228:@11898.4]
  wire  _T_528; // @[MemPrimitives.scala 110:210:@11900.4]
  wire  _T_530; // @[MemPrimitives.scala 110:210:@11901.4]
  wire  _T_531; // @[MemPrimitives.scala 110:228:@11902.4]
  wire  _T_534; // @[MemPrimitives.scala 110:210:@11904.4]
  wire  _T_536; // @[MemPrimitives.scala 110:210:@11905.4]
  wire  _T_537; // @[MemPrimitives.scala 110:228:@11906.4]
  wire  _T_540; // @[MemPrimitives.scala 110:210:@11908.4]
  wire  _T_542; // @[MemPrimitives.scala 110:210:@11909.4]
  wire  _T_543; // @[MemPrimitives.scala 110:228:@11910.4]
  wire  _T_545; // @[MemPrimitives.scala 123:41:@11924.4]
  wire  _T_546; // @[MemPrimitives.scala 123:41:@11925.4]
  wire  _T_547; // @[MemPrimitives.scala 123:41:@11926.4]
  wire  _T_548; // @[MemPrimitives.scala 123:41:@11927.4]
  wire  _T_549; // @[MemPrimitives.scala 123:41:@11928.4]
  wire  _T_550; // @[MemPrimitives.scala 123:41:@11929.4]
  wire  _T_551; // @[MemPrimitives.scala 123:41:@11930.4]
  wire  _T_552; // @[MemPrimitives.scala 123:41:@11931.4]
  wire  _T_553; // @[MemPrimitives.scala 123:41:@11932.4]
  wire [2:0] _T_555; // @[Cat.scala 30:58:@11934.4]
  wire [2:0] _T_557; // @[Cat.scala 30:58:@11936.4]
  wire [2:0] _T_559; // @[Cat.scala 30:58:@11938.4]
  wire [2:0] _T_561; // @[Cat.scala 30:58:@11940.4]
  wire [2:0] _T_563; // @[Cat.scala 30:58:@11942.4]
  wire [2:0] _T_565; // @[Cat.scala 30:58:@11944.4]
  wire [2:0] _T_567; // @[Cat.scala 30:58:@11946.4]
  wire [2:0] _T_569; // @[Cat.scala 30:58:@11948.4]
  wire [2:0] _T_571; // @[Cat.scala 30:58:@11950.4]
  wire [2:0] _T_572; // @[Mux.scala 31:69:@11951.4]
  wire [2:0] _T_573; // @[Mux.scala 31:69:@11952.4]
  wire [2:0] _T_574; // @[Mux.scala 31:69:@11953.4]
  wire [2:0] _T_575; // @[Mux.scala 31:69:@11954.4]
  wire [2:0] _T_576; // @[Mux.scala 31:69:@11955.4]
  wire [2:0] _T_577; // @[Mux.scala 31:69:@11956.4]
  wire [2:0] _T_578; // @[Mux.scala 31:69:@11957.4]
  wire [2:0] _T_579; // @[Mux.scala 31:69:@11958.4]
  wire  _T_586; // @[MemPrimitives.scala 110:210:@11966.4]
  wire  _T_587; // @[MemPrimitives.scala 110:228:@11967.4]
  wire  _T_592; // @[MemPrimitives.scala 110:210:@11970.4]
  wire  _T_593; // @[MemPrimitives.scala 110:228:@11971.4]
  wire  _T_598; // @[MemPrimitives.scala 110:210:@11974.4]
  wire  _T_599; // @[MemPrimitives.scala 110:228:@11975.4]
  wire  _T_604; // @[MemPrimitives.scala 110:210:@11978.4]
  wire  _T_605; // @[MemPrimitives.scala 110:228:@11979.4]
  wire  _T_610; // @[MemPrimitives.scala 110:210:@11982.4]
  wire  _T_611; // @[MemPrimitives.scala 110:228:@11983.4]
  wire  _T_616; // @[MemPrimitives.scala 110:210:@11986.4]
  wire  _T_617; // @[MemPrimitives.scala 110:228:@11987.4]
  wire  _T_622; // @[MemPrimitives.scala 110:210:@11990.4]
  wire  _T_623; // @[MemPrimitives.scala 110:228:@11991.4]
  wire  _T_628; // @[MemPrimitives.scala 110:210:@11994.4]
  wire  _T_629; // @[MemPrimitives.scala 110:228:@11995.4]
  wire  _T_634; // @[MemPrimitives.scala 110:210:@11998.4]
  wire  _T_635; // @[MemPrimitives.scala 110:228:@11999.4]
  wire  _T_637; // @[MemPrimitives.scala 123:41:@12013.4]
  wire  _T_638; // @[MemPrimitives.scala 123:41:@12014.4]
  wire  _T_639; // @[MemPrimitives.scala 123:41:@12015.4]
  wire  _T_640; // @[MemPrimitives.scala 123:41:@12016.4]
  wire  _T_641; // @[MemPrimitives.scala 123:41:@12017.4]
  wire  _T_642; // @[MemPrimitives.scala 123:41:@12018.4]
  wire  _T_643; // @[MemPrimitives.scala 123:41:@12019.4]
  wire  _T_644; // @[MemPrimitives.scala 123:41:@12020.4]
  wire  _T_645; // @[MemPrimitives.scala 123:41:@12021.4]
  wire [2:0] _T_647; // @[Cat.scala 30:58:@12023.4]
  wire [2:0] _T_649; // @[Cat.scala 30:58:@12025.4]
  wire [2:0] _T_651; // @[Cat.scala 30:58:@12027.4]
  wire [2:0] _T_653; // @[Cat.scala 30:58:@12029.4]
  wire [2:0] _T_655; // @[Cat.scala 30:58:@12031.4]
  wire [2:0] _T_657; // @[Cat.scala 30:58:@12033.4]
  wire [2:0] _T_659; // @[Cat.scala 30:58:@12035.4]
  wire [2:0] _T_661; // @[Cat.scala 30:58:@12037.4]
  wire [2:0] _T_663; // @[Cat.scala 30:58:@12039.4]
  wire [2:0] _T_664; // @[Mux.scala 31:69:@12040.4]
  wire [2:0] _T_665; // @[Mux.scala 31:69:@12041.4]
  wire [2:0] _T_666; // @[Mux.scala 31:69:@12042.4]
  wire [2:0] _T_667; // @[Mux.scala 31:69:@12043.4]
  wire [2:0] _T_668; // @[Mux.scala 31:69:@12044.4]
  wire [2:0] _T_669; // @[Mux.scala 31:69:@12045.4]
  wire [2:0] _T_670; // @[Mux.scala 31:69:@12046.4]
  wire [2:0] _T_671; // @[Mux.scala 31:69:@12047.4]
  wire  _T_678; // @[MemPrimitives.scala 110:210:@12055.4]
  wire  _T_679; // @[MemPrimitives.scala 110:228:@12056.4]
  wire  _T_684; // @[MemPrimitives.scala 110:210:@12059.4]
  wire  _T_685; // @[MemPrimitives.scala 110:228:@12060.4]
  wire  _T_690; // @[MemPrimitives.scala 110:210:@12063.4]
  wire  _T_691; // @[MemPrimitives.scala 110:228:@12064.4]
  wire  _T_696; // @[MemPrimitives.scala 110:210:@12067.4]
  wire  _T_697; // @[MemPrimitives.scala 110:228:@12068.4]
  wire  _T_702; // @[MemPrimitives.scala 110:210:@12071.4]
  wire  _T_703; // @[MemPrimitives.scala 110:228:@12072.4]
  wire  _T_708; // @[MemPrimitives.scala 110:210:@12075.4]
  wire  _T_709; // @[MemPrimitives.scala 110:228:@12076.4]
  wire  _T_714; // @[MemPrimitives.scala 110:210:@12079.4]
  wire  _T_715; // @[MemPrimitives.scala 110:228:@12080.4]
  wire  _T_720; // @[MemPrimitives.scala 110:210:@12083.4]
  wire  _T_721; // @[MemPrimitives.scala 110:228:@12084.4]
  wire  _T_726; // @[MemPrimitives.scala 110:210:@12087.4]
  wire  _T_727; // @[MemPrimitives.scala 110:228:@12088.4]
  wire  _T_729; // @[MemPrimitives.scala 123:41:@12102.4]
  wire  _T_730; // @[MemPrimitives.scala 123:41:@12103.4]
  wire  _T_731; // @[MemPrimitives.scala 123:41:@12104.4]
  wire  _T_732; // @[MemPrimitives.scala 123:41:@12105.4]
  wire  _T_733; // @[MemPrimitives.scala 123:41:@12106.4]
  wire  _T_734; // @[MemPrimitives.scala 123:41:@12107.4]
  wire  _T_735; // @[MemPrimitives.scala 123:41:@12108.4]
  wire  _T_736; // @[MemPrimitives.scala 123:41:@12109.4]
  wire  _T_737; // @[MemPrimitives.scala 123:41:@12110.4]
  wire [2:0] _T_739; // @[Cat.scala 30:58:@12112.4]
  wire [2:0] _T_741; // @[Cat.scala 30:58:@12114.4]
  wire [2:0] _T_743; // @[Cat.scala 30:58:@12116.4]
  wire [2:0] _T_745; // @[Cat.scala 30:58:@12118.4]
  wire [2:0] _T_747; // @[Cat.scala 30:58:@12120.4]
  wire [2:0] _T_749; // @[Cat.scala 30:58:@12122.4]
  wire [2:0] _T_751; // @[Cat.scala 30:58:@12124.4]
  wire [2:0] _T_753; // @[Cat.scala 30:58:@12126.4]
  wire [2:0] _T_755; // @[Cat.scala 30:58:@12128.4]
  wire [2:0] _T_756; // @[Mux.scala 31:69:@12129.4]
  wire [2:0] _T_757; // @[Mux.scala 31:69:@12130.4]
  wire [2:0] _T_758; // @[Mux.scala 31:69:@12131.4]
  wire [2:0] _T_759; // @[Mux.scala 31:69:@12132.4]
  wire [2:0] _T_760; // @[Mux.scala 31:69:@12133.4]
  wire [2:0] _T_761; // @[Mux.scala 31:69:@12134.4]
  wire [2:0] _T_762; // @[Mux.scala 31:69:@12135.4]
  wire [2:0] _T_763; // @[Mux.scala 31:69:@12136.4]
  wire  _T_770; // @[MemPrimitives.scala 110:210:@12144.4]
  wire  _T_771; // @[MemPrimitives.scala 110:228:@12145.4]
  wire  _T_776; // @[MemPrimitives.scala 110:210:@12148.4]
  wire  _T_777; // @[MemPrimitives.scala 110:228:@12149.4]
  wire  _T_782; // @[MemPrimitives.scala 110:210:@12152.4]
  wire  _T_783; // @[MemPrimitives.scala 110:228:@12153.4]
  wire  _T_788; // @[MemPrimitives.scala 110:210:@12156.4]
  wire  _T_789; // @[MemPrimitives.scala 110:228:@12157.4]
  wire  _T_794; // @[MemPrimitives.scala 110:210:@12160.4]
  wire  _T_795; // @[MemPrimitives.scala 110:228:@12161.4]
  wire  _T_800; // @[MemPrimitives.scala 110:210:@12164.4]
  wire  _T_801; // @[MemPrimitives.scala 110:228:@12165.4]
  wire  _T_806; // @[MemPrimitives.scala 110:210:@12168.4]
  wire  _T_807; // @[MemPrimitives.scala 110:228:@12169.4]
  wire  _T_812; // @[MemPrimitives.scala 110:210:@12172.4]
  wire  _T_813; // @[MemPrimitives.scala 110:228:@12173.4]
  wire  _T_818; // @[MemPrimitives.scala 110:210:@12176.4]
  wire  _T_819; // @[MemPrimitives.scala 110:228:@12177.4]
  wire  _T_821; // @[MemPrimitives.scala 123:41:@12191.4]
  wire  _T_822; // @[MemPrimitives.scala 123:41:@12192.4]
  wire  _T_823; // @[MemPrimitives.scala 123:41:@12193.4]
  wire  _T_824; // @[MemPrimitives.scala 123:41:@12194.4]
  wire  _T_825; // @[MemPrimitives.scala 123:41:@12195.4]
  wire  _T_826; // @[MemPrimitives.scala 123:41:@12196.4]
  wire  _T_827; // @[MemPrimitives.scala 123:41:@12197.4]
  wire  _T_828; // @[MemPrimitives.scala 123:41:@12198.4]
  wire  _T_829; // @[MemPrimitives.scala 123:41:@12199.4]
  wire [2:0] _T_831; // @[Cat.scala 30:58:@12201.4]
  wire [2:0] _T_833; // @[Cat.scala 30:58:@12203.4]
  wire [2:0] _T_835; // @[Cat.scala 30:58:@12205.4]
  wire [2:0] _T_837; // @[Cat.scala 30:58:@12207.4]
  wire [2:0] _T_839; // @[Cat.scala 30:58:@12209.4]
  wire [2:0] _T_841; // @[Cat.scala 30:58:@12211.4]
  wire [2:0] _T_843; // @[Cat.scala 30:58:@12213.4]
  wire [2:0] _T_845; // @[Cat.scala 30:58:@12215.4]
  wire [2:0] _T_847; // @[Cat.scala 30:58:@12217.4]
  wire [2:0] _T_848; // @[Mux.scala 31:69:@12218.4]
  wire [2:0] _T_849; // @[Mux.scala 31:69:@12219.4]
  wire [2:0] _T_850; // @[Mux.scala 31:69:@12220.4]
  wire [2:0] _T_851; // @[Mux.scala 31:69:@12221.4]
  wire [2:0] _T_852; // @[Mux.scala 31:69:@12222.4]
  wire [2:0] _T_853; // @[Mux.scala 31:69:@12223.4]
  wire [2:0] _T_854; // @[Mux.scala 31:69:@12224.4]
  wire [2:0] _T_855; // @[Mux.scala 31:69:@12225.4]
  wire  _T_860; // @[MemPrimitives.scala 110:210:@12232.4]
  wire  _T_863; // @[MemPrimitives.scala 110:228:@12234.4]
  wire  _T_866; // @[MemPrimitives.scala 110:210:@12236.4]
  wire  _T_869; // @[MemPrimitives.scala 110:228:@12238.4]
  wire  _T_872; // @[MemPrimitives.scala 110:210:@12240.4]
  wire  _T_875; // @[MemPrimitives.scala 110:228:@12242.4]
  wire  _T_878; // @[MemPrimitives.scala 110:210:@12244.4]
  wire  _T_881; // @[MemPrimitives.scala 110:228:@12246.4]
  wire  _T_884; // @[MemPrimitives.scala 110:210:@12248.4]
  wire  _T_887; // @[MemPrimitives.scala 110:228:@12250.4]
  wire  _T_890; // @[MemPrimitives.scala 110:210:@12252.4]
  wire  _T_893; // @[MemPrimitives.scala 110:228:@12254.4]
  wire  _T_896; // @[MemPrimitives.scala 110:210:@12256.4]
  wire  _T_899; // @[MemPrimitives.scala 110:228:@12258.4]
  wire  _T_902; // @[MemPrimitives.scala 110:210:@12260.4]
  wire  _T_905; // @[MemPrimitives.scala 110:228:@12262.4]
  wire  _T_908; // @[MemPrimitives.scala 110:210:@12264.4]
  wire  _T_911; // @[MemPrimitives.scala 110:228:@12266.4]
  wire  _T_913; // @[MemPrimitives.scala 123:41:@12280.4]
  wire  _T_914; // @[MemPrimitives.scala 123:41:@12281.4]
  wire  _T_915; // @[MemPrimitives.scala 123:41:@12282.4]
  wire  _T_916; // @[MemPrimitives.scala 123:41:@12283.4]
  wire  _T_917; // @[MemPrimitives.scala 123:41:@12284.4]
  wire  _T_918; // @[MemPrimitives.scala 123:41:@12285.4]
  wire  _T_919; // @[MemPrimitives.scala 123:41:@12286.4]
  wire  _T_920; // @[MemPrimitives.scala 123:41:@12287.4]
  wire  _T_921; // @[MemPrimitives.scala 123:41:@12288.4]
  wire [2:0] _T_923; // @[Cat.scala 30:58:@12290.4]
  wire [2:0] _T_925; // @[Cat.scala 30:58:@12292.4]
  wire [2:0] _T_927; // @[Cat.scala 30:58:@12294.4]
  wire [2:0] _T_929; // @[Cat.scala 30:58:@12296.4]
  wire [2:0] _T_931; // @[Cat.scala 30:58:@12298.4]
  wire [2:0] _T_933; // @[Cat.scala 30:58:@12300.4]
  wire [2:0] _T_935; // @[Cat.scala 30:58:@12302.4]
  wire [2:0] _T_937; // @[Cat.scala 30:58:@12304.4]
  wire [2:0] _T_939; // @[Cat.scala 30:58:@12306.4]
  wire [2:0] _T_940; // @[Mux.scala 31:69:@12307.4]
  wire [2:0] _T_941; // @[Mux.scala 31:69:@12308.4]
  wire [2:0] _T_942; // @[Mux.scala 31:69:@12309.4]
  wire [2:0] _T_943; // @[Mux.scala 31:69:@12310.4]
  wire [2:0] _T_944; // @[Mux.scala 31:69:@12311.4]
  wire [2:0] _T_945; // @[Mux.scala 31:69:@12312.4]
  wire [2:0] _T_946; // @[Mux.scala 31:69:@12313.4]
  wire [2:0] _T_947; // @[Mux.scala 31:69:@12314.4]
  wire  _T_955; // @[MemPrimitives.scala 110:228:@12323.4]
  wire  _T_961; // @[MemPrimitives.scala 110:228:@12327.4]
  wire  _T_967; // @[MemPrimitives.scala 110:228:@12331.4]
  wire  _T_973; // @[MemPrimitives.scala 110:228:@12335.4]
  wire  _T_979; // @[MemPrimitives.scala 110:228:@12339.4]
  wire  _T_985; // @[MemPrimitives.scala 110:228:@12343.4]
  wire  _T_991; // @[MemPrimitives.scala 110:228:@12347.4]
  wire  _T_997; // @[MemPrimitives.scala 110:228:@12351.4]
  wire  _T_1003; // @[MemPrimitives.scala 110:228:@12355.4]
  wire  _T_1005; // @[MemPrimitives.scala 123:41:@12369.4]
  wire  _T_1006; // @[MemPrimitives.scala 123:41:@12370.4]
  wire  _T_1007; // @[MemPrimitives.scala 123:41:@12371.4]
  wire  _T_1008; // @[MemPrimitives.scala 123:41:@12372.4]
  wire  _T_1009; // @[MemPrimitives.scala 123:41:@12373.4]
  wire  _T_1010; // @[MemPrimitives.scala 123:41:@12374.4]
  wire  _T_1011; // @[MemPrimitives.scala 123:41:@12375.4]
  wire  _T_1012; // @[MemPrimitives.scala 123:41:@12376.4]
  wire  _T_1013; // @[MemPrimitives.scala 123:41:@12377.4]
  wire [2:0] _T_1015; // @[Cat.scala 30:58:@12379.4]
  wire [2:0] _T_1017; // @[Cat.scala 30:58:@12381.4]
  wire [2:0] _T_1019; // @[Cat.scala 30:58:@12383.4]
  wire [2:0] _T_1021; // @[Cat.scala 30:58:@12385.4]
  wire [2:0] _T_1023; // @[Cat.scala 30:58:@12387.4]
  wire [2:0] _T_1025; // @[Cat.scala 30:58:@12389.4]
  wire [2:0] _T_1027; // @[Cat.scala 30:58:@12391.4]
  wire [2:0] _T_1029; // @[Cat.scala 30:58:@12393.4]
  wire [2:0] _T_1031; // @[Cat.scala 30:58:@12395.4]
  wire [2:0] _T_1032; // @[Mux.scala 31:69:@12396.4]
  wire [2:0] _T_1033; // @[Mux.scala 31:69:@12397.4]
  wire [2:0] _T_1034; // @[Mux.scala 31:69:@12398.4]
  wire [2:0] _T_1035; // @[Mux.scala 31:69:@12399.4]
  wire [2:0] _T_1036; // @[Mux.scala 31:69:@12400.4]
  wire [2:0] _T_1037; // @[Mux.scala 31:69:@12401.4]
  wire [2:0] _T_1038; // @[Mux.scala 31:69:@12402.4]
  wire [2:0] _T_1039; // @[Mux.scala 31:69:@12403.4]
  wire  _T_1047; // @[MemPrimitives.scala 110:228:@12412.4]
  wire  _T_1053; // @[MemPrimitives.scala 110:228:@12416.4]
  wire  _T_1059; // @[MemPrimitives.scala 110:228:@12420.4]
  wire  _T_1065; // @[MemPrimitives.scala 110:228:@12424.4]
  wire  _T_1071; // @[MemPrimitives.scala 110:228:@12428.4]
  wire  _T_1077; // @[MemPrimitives.scala 110:228:@12432.4]
  wire  _T_1083; // @[MemPrimitives.scala 110:228:@12436.4]
  wire  _T_1089; // @[MemPrimitives.scala 110:228:@12440.4]
  wire  _T_1095; // @[MemPrimitives.scala 110:228:@12444.4]
  wire  _T_1097; // @[MemPrimitives.scala 123:41:@12458.4]
  wire  _T_1098; // @[MemPrimitives.scala 123:41:@12459.4]
  wire  _T_1099; // @[MemPrimitives.scala 123:41:@12460.4]
  wire  _T_1100; // @[MemPrimitives.scala 123:41:@12461.4]
  wire  _T_1101; // @[MemPrimitives.scala 123:41:@12462.4]
  wire  _T_1102; // @[MemPrimitives.scala 123:41:@12463.4]
  wire  _T_1103; // @[MemPrimitives.scala 123:41:@12464.4]
  wire  _T_1104; // @[MemPrimitives.scala 123:41:@12465.4]
  wire  _T_1105; // @[MemPrimitives.scala 123:41:@12466.4]
  wire [2:0] _T_1107; // @[Cat.scala 30:58:@12468.4]
  wire [2:0] _T_1109; // @[Cat.scala 30:58:@12470.4]
  wire [2:0] _T_1111; // @[Cat.scala 30:58:@12472.4]
  wire [2:0] _T_1113; // @[Cat.scala 30:58:@12474.4]
  wire [2:0] _T_1115; // @[Cat.scala 30:58:@12476.4]
  wire [2:0] _T_1117; // @[Cat.scala 30:58:@12478.4]
  wire [2:0] _T_1119; // @[Cat.scala 30:58:@12480.4]
  wire [2:0] _T_1121; // @[Cat.scala 30:58:@12482.4]
  wire [2:0] _T_1123; // @[Cat.scala 30:58:@12484.4]
  wire [2:0] _T_1124; // @[Mux.scala 31:69:@12485.4]
  wire [2:0] _T_1125; // @[Mux.scala 31:69:@12486.4]
  wire [2:0] _T_1126; // @[Mux.scala 31:69:@12487.4]
  wire [2:0] _T_1127; // @[Mux.scala 31:69:@12488.4]
  wire [2:0] _T_1128; // @[Mux.scala 31:69:@12489.4]
  wire [2:0] _T_1129; // @[Mux.scala 31:69:@12490.4]
  wire [2:0] _T_1130; // @[Mux.scala 31:69:@12491.4]
  wire [2:0] _T_1131; // @[Mux.scala 31:69:@12492.4]
  wire  _T_1139; // @[MemPrimitives.scala 110:228:@12501.4]
  wire  _T_1145; // @[MemPrimitives.scala 110:228:@12505.4]
  wire  _T_1151; // @[MemPrimitives.scala 110:228:@12509.4]
  wire  _T_1157; // @[MemPrimitives.scala 110:228:@12513.4]
  wire  _T_1163; // @[MemPrimitives.scala 110:228:@12517.4]
  wire  _T_1169; // @[MemPrimitives.scala 110:228:@12521.4]
  wire  _T_1175; // @[MemPrimitives.scala 110:228:@12525.4]
  wire  _T_1181; // @[MemPrimitives.scala 110:228:@12529.4]
  wire  _T_1187; // @[MemPrimitives.scala 110:228:@12533.4]
  wire  _T_1189; // @[MemPrimitives.scala 123:41:@12547.4]
  wire  _T_1190; // @[MemPrimitives.scala 123:41:@12548.4]
  wire  _T_1191; // @[MemPrimitives.scala 123:41:@12549.4]
  wire  _T_1192; // @[MemPrimitives.scala 123:41:@12550.4]
  wire  _T_1193; // @[MemPrimitives.scala 123:41:@12551.4]
  wire  _T_1194; // @[MemPrimitives.scala 123:41:@12552.4]
  wire  _T_1195; // @[MemPrimitives.scala 123:41:@12553.4]
  wire  _T_1196; // @[MemPrimitives.scala 123:41:@12554.4]
  wire  _T_1197; // @[MemPrimitives.scala 123:41:@12555.4]
  wire [2:0] _T_1199; // @[Cat.scala 30:58:@12557.4]
  wire [2:0] _T_1201; // @[Cat.scala 30:58:@12559.4]
  wire [2:0] _T_1203; // @[Cat.scala 30:58:@12561.4]
  wire [2:0] _T_1205; // @[Cat.scala 30:58:@12563.4]
  wire [2:0] _T_1207; // @[Cat.scala 30:58:@12565.4]
  wire [2:0] _T_1209; // @[Cat.scala 30:58:@12567.4]
  wire [2:0] _T_1211; // @[Cat.scala 30:58:@12569.4]
  wire [2:0] _T_1213; // @[Cat.scala 30:58:@12571.4]
  wire [2:0] _T_1215; // @[Cat.scala 30:58:@12573.4]
  wire [2:0] _T_1216; // @[Mux.scala 31:69:@12574.4]
  wire [2:0] _T_1217; // @[Mux.scala 31:69:@12575.4]
  wire [2:0] _T_1218; // @[Mux.scala 31:69:@12576.4]
  wire [2:0] _T_1219; // @[Mux.scala 31:69:@12577.4]
  wire [2:0] _T_1220; // @[Mux.scala 31:69:@12578.4]
  wire [2:0] _T_1221; // @[Mux.scala 31:69:@12579.4]
  wire [2:0] _T_1222; // @[Mux.scala 31:69:@12580.4]
  wire [2:0] _T_1223; // @[Mux.scala 31:69:@12581.4]
  wire  _T_1228; // @[MemPrimitives.scala 110:210:@12588.4]
  wire  _T_1231; // @[MemPrimitives.scala 110:228:@12590.4]
  wire  _T_1234; // @[MemPrimitives.scala 110:210:@12592.4]
  wire  _T_1237; // @[MemPrimitives.scala 110:228:@12594.4]
  wire  _T_1240; // @[MemPrimitives.scala 110:210:@12596.4]
  wire  _T_1243; // @[MemPrimitives.scala 110:228:@12598.4]
  wire  _T_1246; // @[MemPrimitives.scala 110:210:@12600.4]
  wire  _T_1249; // @[MemPrimitives.scala 110:228:@12602.4]
  wire  _T_1252; // @[MemPrimitives.scala 110:210:@12604.4]
  wire  _T_1255; // @[MemPrimitives.scala 110:228:@12606.4]
  wire  _T_1258; // @[MemPrimitives.scala 110:210:@12608.4]
  wire  _T_1261; // @[MemPrimitives.scala 110:228:@12610.4]
  wire  _T_1264; // @[MemPrimitives.scala 110:210:@12612.4]
  wire  _T_1267; // @[MemPrimitives.scala 110:228:@12614.4]
  wire  _T_1270; // @[MemPrimitives.scala 110:210:@12616.4]
  wire  _T_1273; // @[MemPrimitives.scala 110:228:@12618.4]
  wire  _T_1276; // @[MemPrimitives.scala 110:210:@12620.4]
  wire  _T_1279; // @[MemPrimitives.scala 110:228:@12622.4]
  wire  _T_1281; // @[MemPrimitives.scala 123:41:@12636.4]
  wire  _T_1282; // @[MemPrimitives.scala 123:41:@12637.4]
  wire  _T_1283; // @[MemPrimitives.scala 123:41:@12638.4]
  wire  _T_1284; // @[MemPrimitives.scala 123:41:@12639.4]
  wire  _T_1285; // @[MemPrimitives.scala 123:41:@12640.4]
  wire  _T_1286; // @[MemPrimitives.scala 123:41:@12641.4]
  wire  _T_1287; // @[MemPrimitives.scala 123:41:@12642.4]
  wire  _T_1288; // @[MemPrimitives.scala 123:41:@12643.4]
  wire  _T_1289; // @[MemPrimitives.scala 123:41:@12644.4]
  wire [2:0] _T_1291; // @[Cat.scala 30:58:@12646.4]
  wire [2:0] _T_1293; // @[Cat.scala 30:58:@12648.4]
  wire [2:0] _T_1295; // @[Cat.scala 30:58:@12650.4]
  wire [2:0] _T_1297; // @[Cat.scala 30:58:@12652.4]
  wire [2:0] _T_1299; // @[Cat.scala 30:58:@12654.4]
  wire [2:0] _T_1301; // @[Cat.scala 30:58:@12656.4]
  wire [2:0] _T_1303; // @[Cat.scala 30:58:@12658.4]
  wire [2:0] _T_1305; // @[Cat.scala 30:58:@12660.4]
  wire [2:0] _T_1307; // @[Cat.scala 30:58:@12662.4]
  wire [2:0] _T_1308; // @[Mux.scala 31:69:@12663.4]
  wire [2:0] _T_1309; // @[Mux.scala 31:69:@12664.4]
  wire [2:0] _T_1310; // @[Mux.scala 31:69:@12665.4]
  wire [2:0] _T_1311; // @[Mux.scala 31:69:@12666.4]
  wire [2:0] _T_1312; // @[Mux.scala 31:69:@12667.4]
  wire [2:0] _T_1313; // @[Mux.scala 31:69:@12668.4]
  wire [2:0] _T_1314; // @[Mux.scala 31:69:@12669.4]
  wire [2:0] _T_1315; // @[Mux.scala 31:69:@12670.4]
  wire  _T_1323; // @[MemPrimitives.scala 110:228:@12679.4]
  wire  _T_1329; // @[MemPrimitives.scala 110:228:@12683.4]
  wire  _T_1335; // @[MemPrimitives.scala 110:228:@12687.4]
  wire  _T_1341; // @[MemPrimitives.scala 110:228:@12691.4]
  wire  _T_1347; // @[MemPrimitives.scala 110:228:@12695.4]
  wire  _T_1353; // @[MemPrimitives.scala 110:228:@12699.4]
  wire  _T_1359; // @[MemPrimitives.scala 110:228:@12703.4]
  wire  _T_1365; // @[MemPrimitives.scala 110:228:@12707.4]
  wire  _T_1371; // @[MemPrimitives.scala 110:228:@12711.4]
  wire  _T_1373; // @[MemPrimitives.scala 123:41:@12725.4]
  wire  _T_1374; // @[MemPrimitives.scala 123:41:@12726.4]
  wire  _T_1375; // @[MemPrimitives.scala 123:41:@12727.4]
  wire  _T_1376; // @[MemPrimitives.scala 123:41:@12728.4]
  wire  _T_1377; // @[MemPrimitives.scala 123:41:@12729.4]
  wire  _T_1378; // @[MemPrimitives.scala 123:41:@12730.4]
  wire  _T_1379; // @[MemPrimitives.scala 123:41:@12731.4]
  wire  _T_1380; // @[MemPrimitives.scala 123:41:@12732.4]
  wire  _T_1381; // @[MemPrimitives.scala 123:41:@12733.4]
  wire [2:0] _T_1383; // @[Cat.scala 30:58:@12735.4]
  wire [2:0] _T_1385; // @[Cat.scala 30:58:@12737.4]
  wire [2:0] _T_1387; // @[Cat.scala 30:58:@12739.4]
  wire [2:0] _T_1389; // @[Cat.scala 30:58:@12741.4]
  wire [2:0] _T_1391; // @[Cat.scala 30:58:@12743.4]
  wire [2:0] _T_1393; // @[Cat.scala 30:58:@12745.4]
  wire [2:0] _T_1395; // @[Cat.scala 30:58:@12747.4]
  wire [2:0] _T_1397; // @[Cat.scala 30:58:@12749.4]
  wire [2:0] _T_1399; // @[Cat.scala 30:58:@12751.4]
  wire [2:0] _T_1400; // @[Mux.scala 31:69:@12752.4]
  wire [2:0] _T_1401; // @[Mux.scala 31:69:@12753.4]
  wire [2:0] _T_1402; // @[Mux.scala 31:69:@12754.4]
  wire [2:0] _T_1403; // @[Mux.scala 31:69:@12755.4]
  wire [2:0] _T_1404; // @[Mux.scala 31:69:@12756.4]
  wire [2:0] _T_1405; // @[Mux.scala 31:69:@12757.4]
  wire [2:0] _T_1406; // @[Mux.scala 31:69:@12758.4]
  wire [2:0] _T_1407; // @[Mux.scala 31:69:@12759.4]
  wire  _T_1415; // @[MemPrimitives.scala 110:228:@12768.4]
  wire  _T_1421; // @[MemPrimitives.scala 110:228:@12772.4]
  wire  _T_1427; // @[MemPrimitives.scala 110:228:@12776.4]
  wire  _T_1433; // @[MemPrimitives.scala 110:228:@12780.4]
  wire  _T_1439; // @[MemPrimitives.scala 110:228:@12784.4]
  wire  _T_1445; // @[MemPrimitives.scala 110:228:@12788.4]
  wire  _T_1451; // @[MemPrimitives.scala 110:228:@12792.4]
  wire  _T_1457; // @[MemPrimitives.scala 110:228:@12796.4]
  wire  _T_1463; // @[MemPrimitives.scala 110:228:@12800.4]
  wire  _T_1465; // @[MemPrimitives.scala 123:41:@12814.4]
  wire  _T_1466; // @[MemPrimitives.scala 123:41:@12815.4]
  wire  _T_1467; // @[MemPrimitives.scala 123:41:@12816.4]
  wire  _T_1468; // @[MemPrimitives.scala 123:41:@12817.4]
  wire  _T_1469; // @[MemPrimitives.scala 123:41:@12818.4]
  wire  _T_1470; // @[MemPrimitives.scala 123:41:@12819.4]
  wire  _T_1471; // @[MemPrimitives.scala 123:41:@12820.4]
  wire  _T_1472; // @[MemPrimitives.scala 123:41:@12821.4]
  wire  _T_1473; // @[MemPrimitives.scala 123:41:@12822.4]
  wire [2:0] _T_1475; // @[Cat.scala 30:58:@12824.4]
  wire [2:0] _T_1477; // @[Cat.scala 30:58:@12826.4]
  wire [2:0] _T_1479; // @[Cat.scala 30:58:@12828.4]
  wire [2:0] _T_1481; // @[Cat.scala 30:58:@12830.4]
  wire [2:0] _T_1483; // @[Cat.scala 30:58:@12832.4]
  wire [2:0] _T_1485; // @[Cat.scala 30:58:@12834.4]
  wire [2:0] _T_1487; // @[Cat.scala 30:58:@12836.4]
  wire [2:0] _T_1489; // @[Cat.scala 30:58:@12838.4]
  wire [2:0] _T_1491; // @[Cat.scala 30:58:@12840.4]
  wire [2:0] _T_1492; // @[Mux.scala 31:69:@12841.4]
  wire [2:0] _T_1493; // @[Mux.scala 31:69:@12842.4]
  wire [2:0] _T_1494; // @[Mux.scala 31:69:@12843.4]
  wire [2:0] _T_1495; // @[Mux.scala 31:69:@12844.4]
  wire [2:0] _T_1496; // @[Mux.scala 31:69:@12845.4]
  wire [2:0] _T_1497; // @[Mux.scala 31:69:@12846.4]
  wire [2:0] _T_1498; // @[Mux.scala 31:69:@12847.4]
  wire [2:0] _T_1499; // @[Mux.scala 31:69:@12848.4]
  wire  _T_1507; // @[MemPrimitives.scala 110:228:@12857.4]
  wire  _T_1513; // @[MemPrimitives.scala 110:228:@12861.4]
  wire  _T_1519; // @[MemPrimitives.scala 110:228:@12865.4]
  wire  _T_1525; // @[MemPrimitives.scala 110:228:@12869.4]
  wire  _T_1531; // @[MemPrimitives.scala 110:228:@12873.4]
  wire  _T_1537; // @[MemPrimitives.scala 110:228:@12877.4]
  wire  _T_1543; // @[MemPrimitives.scala 110:228:@12881.4]
  wire  _T_1549; // @[MemPrimitives.scala 110:228:@12885.4]
  wire  _T_1555; // @[MemPrimitives.scala 110:228:@12889.4]
  wire  _T_1557; // @[MemPrimitives.scala 123:41:@12903.4]
  wire  _T_1558; // @[MemPrimitives.scala 123:41:@12904.4]
  wire  _T_1559; // @[MemPrimitives.scala 123:41:@12905.4]
  wire  _T_1560; // @[MemPrimitives.scala 123:41:@12906.4]
  wire  _T_1561; // @[MemPrimitives.scala 123:41:@12907.4]
  wire  _T_1562; // @[MemPrimitives.scala 123:41:@12908.4]
  wire  _T_1563; // @[MemPrimitives.scala 123:41:@12909.4]
  wire  _T_1564; // @[MemPrimitives.scala 123:41:@12910.4]
  wire  _T_1565; // @[MemPrimitives.scala 123:41:@12911.4]
  wire [2:0] _T_1567; // @[Cat.scala 30:58:@12913.4]
  wire [2:0] _T_1569; // @[Cat.scala 30:58:@12915.4]
  wire [2:0] _T_1571; // @[Cat.scala 30:58:@12917.4]
  wire [2:0] _T_1573; // @[Cat.scala 30:58:@12919.4]
  wire [2:0] _T_1575; // @[Cat.scala 30:58:@12921.4]
  wire [2:0] _T_1577; // @[Cat.scala 30:58:@12923.4]
  wire [2:0] _T_1579; // @[Cat.scala 30:58:@12925.4]
  wire [2:0] _T_1581; // @[Cat.scala 30:58:@12927.4]
  wire [2:0] _T_1583; // @[Cat.scala 30:58:@12929.4]
  wire [2:0] _T_1584; // @[Mux.scala 31:69:@12930.4]
  wire [2:0] _T_1585; // @[Mux.scala 31:69:@12931.4]
  wire [2:0] _T_1586; // @[Mux.scala 31:69:@12932.4]
  wire [2:0] _T_1587; // @[Mux.scala 31:69:@12933.4]
  wire [2:0] _T_1588; // @[Mux.scala 31:69:@12934.4]
  wire [2:0] _T_1589; // @[Mux.scala 31:69:@12935.4]
  wire [2:0] _T_1590; // @[Mux.scala 31:69:@12936.4]
  wire [2:0] _T_1591; // @[Mux.scala 31:69:@12937.4]
  wire  _T_1596; // @[MemPrimitives.scala 110:210:@12944.4]
  wire  _T_1599; // @[MemPrimitives.scala 110:228:@12946.4]
  wire  _T_1602; // @[MemPrimitives.scala 110:210:@12948.4]
  wire  _T_1605; // @[MemPrimitives.scala 110:228:@12950.4]
  wire  _T_1608; // @[MemPrimitives.scala 110:210:@12952.4]
  wire  _T_1611; // @[MemPrimitives.scala 110:228:@12954.4]
  wire  _T_1614; // @[MemPrimitives.scala 110:210:@12956.4]
  wire  _T_1617; // @[MemPrimitives.scala 110:228:@12958.4]
  wire  _T_1620; // @[MemPrimitives.scala 110:210:@12960.4]
  wire  _T_1623; // @[MemPrimitives.scala 110:228:@12962.4]
  wire  _T_1626; // @[MemPrimitives.scala 110:210:@12964.4]
  wire  _T_1629; // @[MemPrimitives.scala 110:228:@12966.4]
  wire  _T_1632; // @[MemPrimitives.scala 110:210:@12968.4]
  wire  _T_1635; // @[MemPrimitives.scala 110:228:@12970.4]
  wire  _T_1638; // @[MemPrimitives.scala 110:210:@12972.4]
  wire  _T_1641; // @[MemPrimitives.scala 110:228:@12974.4]
  wire  _T_1644; // @[MemPrimitives.scala 110:210:@12976.4]
  wire  _T_1647; // @[MemPrimitives.scala 110:228:@12978.4]
  wire  _T_1649; // @[MemPrimitives.scala 123:41:@12992.4]
  wire  _T_1650; // @[MemPrimitives.scala 123:41:@12993.4]
  wire  _T_1651; // @[MemPrimitives.scala 123:41:@12994.4]
  wire  _T_1652; // @[MemPrimitives.scala 123:41:@12995.4]
  wire  _T_1653; // @[MemPrimitives.scala 123:41:@12996.4]
  wire  _T_1654; // @[MemPrimitives.scala 123:41:@12997.4]
  wire  _T_1655; // @[MemPrimitives.scala 123:41:@12998.4]
  wire  _T_1656; // @[MemPrimitives.scala 123:41:@12999.4]
  wire  _T_1657; // @[MemPrimitives.scala 123:41:@13000.4]
  wire [2:0] _T_1659; // @[Cat.scala 30:58:@13002.4]
  wire [2:0] _T_1661; // @[Cat.scala 30:58:@13004.4]
  wire [2:0] _T_1663; // @[Cat.scala 30:58:@13006.4]
  wire [2:0] _T_1665; // @[Cat.scala 30:58:@13008.4]
  wire [2:0] _T_1667; // @[Cat.scala 30:58:@13010.4]
  wire [2:0] _T_1669; // @[Cat.scala 30:58:@13012.4]
  wire [2:0] _T_1671; // @[Cat.scala 30:58:@13014.4]
  wire [2:0] _T_1673; // @[Cat.scala 30:58:@13016.4]
  wire [2:0] _T_1675; // @[Cat.scala 30:58:@13018.4]
  wire [2:0] _T_1676; // @[Mux.scala 31:69:@13019.4]
  wire [2:0] _T_1677; // @[Mux.scala 31:69:@13020.4]
  wire [2:0] _T_1678; // @[Mux.scala 31:69:@13021.4]
  wire [2:0] _T_1679; // @[Mux.scala 31:69:@13022.4]
  wire [2:0] _T_1680; // @[Mux.scala 31:69:@13023.4]
  wire [2:0] _T_1681; // @[Mux.scala 31:69:@13024.4]
  wire [2:0] _T_1682; // @[Mux.scala 31:69:@13025.4]
  wire [2:0] _T_1683; // @[Mux.scala 31:69:@13026.4]
  wire  _T_1691; // @[MemPrimitives.scala 110:228:@13035.4]
  wire  _T_1697; // @[MemPrimitives.scala 110:228:@13039.4]
  wire  _T_1703; // @[MemPrimitives.scala 110:228:@13043.4]
  wire  _T_1709; // @[MemPrimitives.scala 110:228:@13047.4]
  wire  _T_1715; // @[MemPrimitives.scala 110:228:@13051.4]
  wire  _T_1721; // @[MemPrimitives.scala 110:228:@13055.4]
  wire  _T_1727; // @[MemPrimitives.scala 110:228:@13059.4]
  wire  _T_1733; // @[MemPrimitives.scala 110:228:@13063.4]
  wire  _T_1739; // @[MemPrimitives.scala 110:228:@13067.4]
  wire  _T_1741; // @[MemPrimitives.scala 123:41:@13081.4]
  wire  _T_1742; // @[MemPrimitives.scala 123:41:@13082.4]
  wire  _T_1743; // @[MemPrimitives.scala 123:41:@13083.4]
  wire  _T_1744; // @[MemPrimitives.scala 123:41:@13084.4]
  wire  _T_1745; // @[MemPrimitives.scala 123:41:@13085.4]
  wire  _T_1746; // @[MemPrimitives.scala 123:41:@13086.4]
  wire  _T_1747; // @[MemPrimitives.scala 123:41:@13087.4]
  wire  _T_1748; // @[MemPrimitives.scala 123:41:@13088.4]
  wire  _T_1749; // @[MemPrimitives.scala 123:41:@13089.4]
  wire [2:0] _T_1751; // @[Cat.scala 30:58:@13091.4]
  wire [2:0] _T_1753; // @[Cat.scala 30:58:@13093.4]
  wire [2:0] _T_1755; // @[Cat.scala 30:58:@13095.4]
  wire [2:0] _T_1757; // @[Cat.scala 30:58:@13097.4]
  wire [2:0] _T_1759; // @[Cat.scala 30:58:@13099.4]
  wire [2:0] _T_1761; // @[Cat.scala 30:58:@13101.4]
  wire [2:0] _T_1763; // @[Cat.scala 30:58:@13103.4]
  wire [2:0] _T_1765; // @[Cat.scala 30:58:@13105.4]
  wire [2:0] _T_1767; // @[Cat.scala 30:58:@13107.4]
  wire [2:0] _T_1768; // @[Mux.scala 31:69:@13108.4]
  wire [2:0] _T_1769; // @[Mux.scala 31:69:@13109.4]
  wire [2:0] _T_1770; // @[Mux.scala 31:69:@13110.4]
  wire [2:0] _T_1771; // @[Mux.scala 31:69:@13111.4]
  wire [2:0] _T_1772; // @[Mux.scala 31:69:@13112.4]
  wire [2:0] _T_1773; // @[Mux.scala 31:69:@13113.4]
  wire [2:0] _T_1774; // @[Mux.scala 31:69:@13114.4]
  wire [2:0] _T_1775; // @[Mux.scala 31:69:@13115.4]
  wire  _T_1783; // @[MemPrimitives.scala 110:228:@13124.4]
  wire  _T_1789; // @[MemPrimitives.scala 110:228:@13128.4]
  wire  _T_1795; // @[MemPrimitives.scala 110:228:@13132.4]
  wire  _T_1801; // @[MemPrimitives.scala 110:228:@13136.4]
  wire  _T_1807; // @[MemPrimitives.scala 110:228:@13140.4]
  wire  _T_1813; // @[MemPrimitives.scala 110:228:@13144.4]
  wire  _T_1819; // @[MemPrimitives.scala 110:228:@13148.4]
  wire  _T_1825; // @[MemPrimitives.scala 110:228:@13152.4]
  wire  _T_1831; // @[MemPrimitives.scala 110:228:@13156.4]
  wire  _T_1833; // @[MemPrimitives.scala 123:41:@13170.4]
  wire  _T_1834; // @[MemPrimitives.scala 123:41:@13171.4]
  wire  _T_1835; // @[MemPrimitives.scala 123:41:@13172.4]
  wire  _T_1836; // @[MemPrimitives.scala 123:41:@13173.4]
  wire  _T_1837; // @[MemPrimitives.scala 123:41:@13174.4]
  wire  _T_1838; // @[MemPrimitives.scala 123:41:@13175.4]
  wire  _T_1839; // @[MemPrimitives.scala 123:41:@13176.4]
  wire  _T_1840; // @[MemPrimitives.scala 123:41:@13177.4]
  wire  _T_1841; // @[MemPrimitives.scala 123:41:@13178.4]
  wire [2:0] _T_1843; // @[Cat.scala 30:58:@13180.4]
  wire [2:0] _T_1845; // @[Cat.scala 30:58:@13182.4]
  wire [2:0] _T_1847; // @[Cat.scala 30:58:@13184.4]
  wire [2:0] _T_1849; // @[Cat.scala 30:58:@13186.4]
  wire [2:0] _T_1851; // @[Cat.scala 30:58:@13188.4]
  wire [2:0] _T_1853; // @[Cat.scala 30:58:@13190.4]
  wire [2:0] _T_1855; // @[Cat.scala 30:58:@13192.4]
  wire [2:0] _T_1857; // @[Cat.scala 30:58:@13194.4]
  wire [2:0] _T_1859; // @[Cat.scala 30:58:@13196.4]
  wire [2:0] _T_1860; // @[Mux.scala 31:69:@13197.4]
  wire [2:0] _T_1861; // @[Mux.scala 31:69:@13198.4]
  wire [2:0] _T_1862; // @[Mux.scala 31:69:@13199.4]
  wire [2:0] _T_1863; // @[Mux.scala 31:69:@13200.4]
  wire [2:0] _T_1864; // @[Mux.scala 31:69:@13201.4]
  wire [2:0] _T_1865; // @[Mux.scala 31:69:@13202.4]
  wire [2:0] _T_1866; // @[Mux.scala 31:69:@13203.4]
  wire [2:0] _T_1867; // @[Mux.scala 31:69:@13204.4]
  wire  _T_1875; // @[MemPrimitives.scala 110:228:@13213.4]
  wire  _T_1881; // @[MemPrimitives.scala 110:228:@13217.4]
  wire  _T_1887; // @[MemPrimitives.scala 110:228:@13221.4]
  wire  _T_1893; // @[MemPrimitives.scala 110:228:@13225.4]
  wire  _T_1899; // @[MemPrimitives.scala 110:228:@13229.4]
  wire  _T_1905; // @[MemPrimitives.scala 110:228:@13233.4]
  wire  _T_1911; // @[MemPrimitives.scala 110:228:@13237.4]
  wire  _T_1917; // @[MemPrimitives.scala 110:228:@13241.4]
  wire  _T_1923; // @[MemPrimitives.scala 110:228:@13245.4]
  wire  _T_1925; // @[MemPrimitives.scala 123:41:@13259.4]
  wire  _T_1926; // @[MemPrimitives.scala 123:41:@13260.4]
  wire  _T_1927; // @[MemPrimitives.scala 123:41:@13261.4]
  wire  _T_1928; // @[MemPrimitives.scala 123:41:@13262.4]
  wire  _T_1929; // @[MemPrimitives.scala 123:41:@13263.4]
  wire  _T_1930; // @[MemPrimitives.scala 123:41:@13264.4]
  wire  _T_1931; // @[MemPrimitives.scala 123:41:@13265.4]
  wire  _T_1932; // @[MemPrimitives.scala 123:41:@13266.4]
  wire  _T_1933; // @[MemPrimitives.scala 123:41:@13267.4]
  wire [2:0] _T_1935; // @[Cat.scala 30:58:@13269.4]
  wire [2:0] _T_1937; // @[Cat.scala 30:58:@13271.4]
  wire [2:0] _T_1939; // @[Cat.scala 30:58:@13273.4]
  wire [2:0] _T_1941; // @[Cat.scala 30:58:@13275.4]
  wire [2:0] _T_1943; // @[Cat.scala 30:58:@13277.4]
  wire [2:0] _T_1945; // @[Cat.scala 30:58:@13279.4]
  wire [2:0] _T_1947; // @[Cat.scala 30:58:@13281.4]
  wire [2:0] _T_1949; // @[Cat.scala 30:58:@13283.4]
  wire [2:0] _T_1951; // @[Cat.scala 30:58:@13285.4]
  wire [2:0] _T_1952; // @[Mux.scala 31:69:@13286.4]
  wire [2:0] _T_1953; // @[Mux.scala 31:69:@13287.4]
  wire [2:0] _T_1954; // @[Mux.scala 31:69:@13288.4]
  wire [2:0] _T_1955; // @[Mux.scala 31:69:@13289.4]
  wire [2:0] _T_1956; // @[Mux.scala 31:69:@13290.4]
  wire [2:0] _T_1957; // @[Mux.scala 31:69:@13291.4]
  wire [2:0] _T_1958; // @[Mux.scala 31:69:@13292.4]
  wire [2:0] _T_1959; // @[Mux.scala 31:69:@13293.4]
  wire  _T_2087; // @[package.scala 96:25:@13466.4 package.scala 96:25:@13467.4]
  wire [7:0] _T_2091; // @[Mux.scala 31:69:@13476.4]
  wire  _T_2084; // @[package.scala 96:25:@13458.4 package.scala 96:25:@13459.4]
  wire [7:0] _T_2092; // @[Mux.scala 31:69:@13477.4]
  wire  _T_2081; // @[package.scala 96:25:@13450.4 package.scala 96:25:@13451.4]
  wire [7:0] _T_2093; // @[Mux.scala 31:69:@13478.4]
  wire  _T_2078; // @[package.scala 96:25:@13442.4 package.scala 96:25:@13443.4]
  wire [7:0] _T_2094; // @[Mux.scala 31:69:@13479.4]
  wire  _T_2075; // @[package.scala 96:25:@13434.4 package.scala 96:25:@13435.4]
  wire [7:0] _T_2095; // @[Mux.scala 31:69:@13480.4]
  wire  _T_2072; // @[package.scala 96:25:@13426.4 package.scala 96:25:@13427.4]
  wire [7:0] _T_2096; // @[Mux.scala 31:69:@13481.4]
  wire  _T_2069; // @[package.scala 96:25:@13418.4 package.scala 96:25:@13419.4]
  wire [7:0] _T_2097; // @[Mux.scala 31:69:@13482.4]
  wire  _T_2066; // @[package.scala 96:25:@13410.4 package.scala 96:25:@13411.4]
  wire [7:0] _T_2098; // @[Mux.scala 31:69:@13483.4]
  wire  _T_2063; // @[package.scala 96:25:@13402.4 package.scala 96:25:@13403.4]
  wire [7:0] _T_2099; // @[Mux.scala 31:69:@13484.4]
  wire  _T_2060; // @[package.scala 96:25:@13394.4 package.scala 96:25:@13395.4]
  wire [7:0] _T_2100; // @[Mux.scala 31:69:@13485.4]
  wire  _T_2057; // @[package.scala 96:25:@13386.4 package.scala 96:25:@13387.4]
  wire [7:0] _T_2101; // @[Mux.scala 31:69:@13486.4]
  wire  _T_2054; // @[package.scala 96:25:@13378.4 package.scala 96:25:@13379.4]
  wire [7:0] _T_2102; // @[Mux.scala 31:69:@13487.4]
  wire  _T_2051; // @[package.scala 96:25:@13370.4 package.scala 96:25:@13371.4]
  wire [7:0] _T_2103; // @[Mux.scala 31:69:@13488.4]
  wire  _T_2048; // @[package.scala 96:25:@13362.4 package.scala 96:25:@13363.4]
  wire [7:0] _T_2104; // @[Mux.scala 31:69:@13489.4]
  wire  _T_2045; // @[package.scala 96:25:@13354.4 package.scala 96:25:@13355.4]
  wire  _T_2230; // @[package.scala 96:25:@13658.4 package.scala 96:25:@13659.4]
  wire [7:0] _T_2234; // @[Mux.scala 31:69:@13668.4]
  wire  _T_2227; // @[package.scala 96:25:@13650.4 package.scala 96:25:@13651.4]
  wire [7:0] _T_2235; // @[Mux.scala 31:69:@13669.4]
  wire  _T_2224; // @[package.scala 96:25:@13642.4 package.scala 96:25:@13643.4]
  wire [7:0] _T_2236; // @[Mux.scala 31:69:@13670.4]
  wire  _T_2221; // @[package.scala 96:25:@13634.4 package.scala 96:25:@13635.4]
  wire [7:0] _T_2237; // @[Mux.scala 31:69:@13671.4]
  wire  _T_2218; // @[package.scala 96:25:@13626.4 package.scala 96:25:@13627.4]
  wire [7:0] _T_2238; // @[Mux.scala 31:69:@13672.4]
  wire  _T_2215; // @[package.scala 96:25:@13618.4 package.scala 96:25:@13619.4]
  wire [7:0] _T_2239; // @[Mux.scala 31:69:@13673.4]
  wire  _T_2212; // @[package.scala 96:25:@13610.4 package.scala 96:25:@13611.4]
  wire [7:0] _T_2240; // @[Mux.scala 31:69:@13674.4]
  wire  _T_2209; // @[package.scala 96:25:@13602.4 package.scala 96:25:@13603.4]
  wire [7:0] _T_2241; // @[Mux.scala 31:69:@13675.4]
  wire  _T_2206; // @[package.scala 96:25:@13594.4 package.scala 96:25:@13595.4]
  wire [7:0] _T_2242; // @[Mux.scala 31:69:@13676.4]
  wire  _T_2203; // @[package.scala 96:25:@13586.4 package.scala 96:25:@13587.4]
  wire [7:0] _T_2243; // @[Mux.scala 31:69:@13677.4]
  wire  _T_2200; // @[package.scala 96:25:@13578.4 package.scala 96:25:@13579.4]
  wire [7:0] _T_2244; // @[Mux.scala 31:69:@13678.4]
  wire  _T_2197; // @[package.scala 96:25:@13570.4 package.scala 96:25:@13571.4]
  wire [7:0] _T_2245; // @[Mux.scala 31:69:@13679.4]
  wire  _T_2194; // @[package.scala 96:25:@13562.4 package.scala 96:25:@13563.4]
  wire [7:0] _T_2246; // @[Mux.scala 31:69:@13680.4]
  wire  _T_2191; // @[package.scala 96:25:@13554.4 package.scala 96:25:@13555.4]
  wire [7:0] _T_2247; // @[Mux.scala 31:69:@13681.4]
  wire  _T_2188; // @[package.scala 96:25:@13546.4 package.scala 96:25:@13547.4]
  wire  _T_2373; // @[package.scala 96:25:@13850.4 package.scala 96:25:@13851.4]
  wire [7:0] _T_2377; // @[Mux.scala 31:69:@13860.4]
  wire  _T_2370; // @[package.scala 96:25:@13842.4 package.scala 96:25:@13843.4]
  wire [7:0] _T_2378; // @[Mux.scala 31:69:@13861.4]
  wire  _T_2367; // @[package.scala 96:25:@13834.4 package.scala 96:25:@13835.4]
  wire [7:0] _T_2379; // @[Mux.scala 31:69:@13862.4]
  wire  _T_2364; // @[package.scala 96:25:@13826.4 package.scala 96:25:@13827.4]
  wire [7:0] _T_2380; // @[Mux.scala 31:69:@13863.4]
  wire  _T_2361; // @[package.scala 96:25:@13818.4 package.scala 96:25:@13819.4]
  wire [7:0] _T_2381; // @[Mux.scala 31:69:@13864.4]
  wire  _T_2358; // @[package.scala 96:25:@13810.4 package.scala 96:25:@13811.4]
  wire [7:0] _T_2382; // @[Mux.scala 31:69:@13865.4]
  wire  _T_2355; // @[package.scala 96:25:@13802.4 package.scala 96:25:@13803.4]
  wire [7:0] _T_2383; // @[Mux.scala 31:69:@13866.4]
  wire  _T_2352; // @[package.scala 96:25:@13794.4 package.scala 96:25:@13795.4]
  wire [7:0] _T_2384; // @[Mux.scala 31:69:@13867.4]
  wire  _T_2349; // @[package.scala 96:25:@13786.4 package.scala 96:25:@13787.4]
  wire [7:0] _T_2385; // @[Mux.scala 31:69:@13868.4]
  wire  _T_2346; // @[package.scala 96:25:@13778.4 package.scala 96:25:@13779.4]
  wire [7:0] _T_2386; // @[Mux.scala 31:69:@13869.4]
  wire  _T_2343; // @[package.scala 96:25:@13770.4 package.scala 96:25:@13771.4]
  wire [7:0] _T_2387; // @[Mux.scala 31:69:@13870.4]
  wire  _T_2340; // @[package.scala 96:25:@13762.4 package.scala 96:25:@13763.4]
  wire [7:0] _T_2388; // @[Mux.scala 31:69:@13871.4]
  wire  _T_2337; // @[package.scala 96:25:@13754.4 package.scala 96:25:@13755.4]
  wire [7:0] _T_2389; // @[Mux.scala 31:69:@13872.4]
  wire  _T_2334; // @[package.scala 96:25:@13746.4 package.scala 96:25:@13747.4]
  wire [7:0] _T_2390; // @[Mux.scala 31:69:@13873.4]
  wire  _T_2331; // @[package.scala 96:25:@13738.4 package.scala 96:25:@13739.4]
  wire  _T_2516; // @[package.scala 96:25:@14042.4 package.scala 96:25:@14043.4]
  wire [7:0] _T_2520; // @[Mux.scala 31:69:@14052.4]
  wire  _T_2513; // @[package.scala 96:25:@14034.4 package.scala 96:25:@14035.4]
  wire [7:0] _T_2521; // @[Mux.scala 31:69:@14053.4]
  wire  _T_2510; // @[package.scala 96:25:@14026.4 package.scala 96:25:@14027.4]
  wire [7:0] _T_2522; // @[Mux.scala 31:69:@14054.4]
  wire  _T_2507; // @[package.scala 96:25:@14018.4 package.scala 96:25:@14019.4]
  wire [7:0] _T_2523; // @[Mux.scala 31:69:@14055.4]
  wire  _T_2504; // @[package.scala 96:25:@14010.4 package.scala 96:25:@14011.4]
  wire [7:0] _T_2524; // @[Mux.scala 31:69:@14056.4]
  wire  _T_2501; // @[package.scala 96:25:@14002.4 package.scala 96:25:@14003.4]
  wire [7:0] _T_2525; // @[Mux.scala 31:69:@14057.4]
  wire  _T_2498; // @[package.scala 96:25:@13994.4 package.scala 96:25:@13995.4]
  wire [7:0] _T_2526; // @[Mux.scala 31:69:@14058.4]
  wire  _T_2495; // @[package.scala 96:25:@13986.4 package.scala 96:25:@13987.4]
  wire [7:0] _T_2527; // @[Mux.scala 31:69:@14059.4]
  wire  _T_2492; // @[package.scala 96:25:@13978.4 package.scala 96:25:@13979.4]
  wire [7:0] _T_2528; // @[Mux.scala 31:69:@14060.4]
  wire  _T_2489; // @[package.scala 96:25:@13970.4 package.scala 96:25:@13971.4]
  wire [7:0] _T_2529; // @[Mux.scala 31:69:@14061.4]
  wire  _T_2486; // @[package.scala 96:25:@13962.4 package.scala 96:25:@13963.4]
  wire [7:0] _T_2530; // @[Mux.scala 31:69:@14062.4]
  wire  _T_2483; // @[package.scala 96:25:@13954.4 package.scala 96:25:@13955.4]
  wire [7:0] _T_2531; // @[Mux.scala 31:69:@14063.4]
  wire  _T_2480; // @[package.scala 96:25:@13946.4 package.scala 96:25:@13947.4]
  wire [7:0] _T_2532; // @[Mux.scala 31:69:@14064.4]
  wire  _T_2477; // @[package.scala 96:25:@13938.4 package.scala 96:25:@13939.4]
  wire [7:0] _T_2533; // @[Mux.scala 31:69:@14065.4]
  wire  _T_2474; // @[package.scala 96:25:@13930.4 package.scala 96:25:@13931.4]
  wire  _T_2659; // @[package.scala 96:25:@14234.4 package.scala 96:25:@14235.4]
  wire [7:0] _T_2663; // @[Mux.scala 31:69:@14244.4]
  wire  _T_2656; // @[package.scala 96:25:@14226.4 package.scala 96:25:@14227.4]
  wire [7:0] _T_2664; // @[Mux.scala 31:69:@14245.4]
  wire  _T_2653; // @[package.scala 96:25:@14218.4 package.scala 96:25:@14219.4]
  wire [7:0] _T_2665; // @[Mux.scala 31:69:@14246.4]
  wire  _T_2650; // @[package.scala 96:25:@14210.4 package.scala 96:25:@14211.4]
  wire [7:0] _T_2666; // @[Mux.scala 31:69:@14247.4]
  wire  _T_2647; // @[package.scala 96:25:@14202.4 package.scala 96:25:@14203.4]
  wire [7:0] _T_2667; // @[Mux.scala 31:69:@14248.4]
  wire  _T_2644; // @[package.scala 96:25:@14194.4 package.scala 96:25:@14195.4]
  wire [7:0] _T_2668; // @[Mux.scala 31:69:@14249.4]
  wire  _T_2641; // @[package.scala 96:25:@14186.4 package.scala 96:25:@14187.4]
  wire [7:0] _T_2669; // @[Mux.scala 31:69:@14250.4]
  wire  _T_2638; // @[package.scala 96:25:@14178.4 package.scala 96:25:@14179.4]
  wire [7:0] _T_2670; // @[Mux.scala 31:69:@14251.4]
  wire  _T_2635; // @[package.scala 96:25:@14170.4 package.scala 96:25:@14171.4]
  wire [7:0] _T_2671; // @[Mux.scala 31:69:@14252.4]
  wire  _T_2632; // @[package.scala 96:25:@14162.4 package.scala 96:25:@14163.4]
  wire [7:0] _T_2672; // @[Mux.scala 31:69:@14253.4]
  wire  _T_2629; // @[package.scala 96:25:@14154.4 package.scala 96:25:@14155.4]
  wire [7:0] _T_2673; // @[Mux.scala 31:69:@14254.4]
  wire  _T_2626; // @[package.scala 96:25:@14146.4 package.scala 96:25:@14147.4]
  wire [7:0] _T_2674; // @[Mux.scala 31:69:@14255.4]
  wire  _T_2623; // @[package.scala 96:25:@14138.4 package.scala 96:25:@14139.4]
  wire [7:0] _T_2675; // @[Mux.scala 31:69:@14256.4]
  wire  _T_2620; // @[package.scala 96:25:@14130.4 package.scala 96:25:@14131.4]
  wire [7:0] _T_2676; // @[Mux.scala 31:69:@14257.4]
  wire  _T_2617; // @[package.scala 96:25:@14122.4 package.scala 96:25:@14123.4]
  wire  _T_2802; // @[package.scala 96:25:@14426.4 package.scala 96:25:@14427.4]
  wire [7:0] _T_2806; // @[Mux.scala 31:69:@14436.4]
  wire  _T_2799; // @[package.scala 96:25:@14418.4 package.scala 96:25:@14419.4]
  wire [7:0] _T_2807; // @[Mux.scala 31:69:@14437.4]
  wire  _T_2796; // @[package.scala 96:25:@14410.4 package.scala 96:25:@14411.4]
  wire [7:0] _T_2808; // @[Mux.scala 31:69:@14438.4]
  wire  _T_2793; // @[package.scala 96:25:@14402.4 package.scala 96:25:@14403.4]
  wire [7:0] _T_2809; // @[Mux.scala 31:69:@14439.4]
  wire  _T_2790; // @[package.scala 96:25:@14394.4 package.scala 96:25:@14395.4]
  wire [7:0] _T_2810; // @[Mux.scala 31:69:@14440.4]
  wire  _T_2787; // @[package.scala 96:25:@14386.4 package.scala 96:25:@14387.4]
  wire [7:0] _T_2811; // @[Mux.scala 31:69:@14441.4]
  wire  _T_2784; // @[package.scala 96:25:@14378.4 package.scala 96:25:@14379.4]
  wire [7:0] _T_2812; // @[Mux.scala 31:69:@14442.4]
  wire  _T_2781; // @[package.scala 96:25:@14370.4 package.scala 96:25:@14371.4]
  wire [7:0] _T_2813; // @[Mux.scala 31:69:@14443.4]
  wire  _T_2778; // @[package.scala 96:25:@14362.4 package.scala 96:25:@14363.4]
  wire [7:0] _T_2814; // @[Mux.scala 31:69:@14444.4]
  wire  _T_2775; // @[package.scala 96:25:@14354.4 package.scala 96:25:@14355.4]
  wire [7:0] _T_2815; // @[Mux.scala 31:69:@14445.4]
  wire  _T_2772; // @[package.scala 96:25:@14346.4 package.scala 96:25:@14347.4]
  wire [7:0] _T_2816; // @[Mux.scala 31:69:@14446.4]
  wire  _T_2769; // @[package.scala 96:25:@14338.4 package.scala 96:25:@14339.4]
  wire [7:0] _T_2817; // @[Mux.scala 31:69:@14447.4]
  wire  _T_2766; // @[package.scala 96:25:@14330.4 package.scala 96:25:@14331.4]
  wire [7:0] _T_2818; // @[Mux.scala 31:69:@14448.4]
  wire  _T_2763; // @[package.scala 96:25:@14322.4 package.scala 96:25:@14323.4]
  wire [7:0] _T_2819; // @[Mux.scala 31:69:@14449.4]
  wire  _T_2760; // @[package.scala 96:25:@14314.4 package.scala 96:25:@14315.4]
  wire  _T_2945; // @[package.scala 96:25:@14618.4 package.scala 96:25:@14619.4]
  wire [7:0] _T_2949; // @[Mux.scala 31:69:@14628.4]
  wire  _T_2942; // @[package.scala 96:25:@14610.4 package.scala 96:25:@14611.4]
  wire [7:0] _T_2950; // @[Mux.scala 31:69:@14629.4]
  wire  _T_2939; // @[package.scala 96:25:@14602.4 package.scala 96:25:@14603.4]
  wire [7:0] _T_2951; // @[Mux.scala 31:69:@14630.4]
  wire  _T_2936; // @[package.scala 96:25:@14594.4 package.scala 96:25:@14595.4]
  wire [7:0] _T_2952; // @[Mux.scala 31:69:@14631.4]
  wire  _T_2933; // @[package.scala 96:25:@14586.4 package.scala 96:25:@14587.4]
  wire [7:0] _T_2953; // @[Mux.scala 31:69:@14632.4]
  wire  _T_2930; // @[package.scala 96:25:@14578.4 package.scala 96:25:@14579.4]
  wire [7:0] _T_2954; // @[Mux.scala 31:69:@14633.4]
  wire  _T_2927; // @[package.scala 96:25:@14570.4 package.scala 96:25:@14571.4]
  wire [7:0] _T_2955; // @[Mux.scala 31:69:@14634.4]
  wire  _T_2924; // @[package.scala 96:25:@14562.4 package.scala 96:25:@14563.4]
  wire [7:0] _T_2956; // @[Mux.scala 31:69:@14635.4]
  wire  _T_2921; // @[package.scala 96:25:@14554.4 package.scala 96:25:@14555.4]
  wire [7:0] _T_2957; // @[Mux.scala 31:69:@14636.4]
  wire  _T_2918; // @[package.scala 96:25:@14546.4 package.scala 96:25:@14547.4]
  wire [7:0] _T_2958; // @[Mux.scala 31:69:@14637.4]
  wire  _T_2915; // @[package.scala 96:25:@14538.4 package.scala 96:25:@14539.4]
  wire [7:0] _T_2959; // @[Mux.scala 31:69:@14638.4]
  wire  _T_2912; // @[package.scala 96:25:@14530.4 package.scala 96:25:@14531.4]
  wire [7:0] _T_2960; // @[Mux.scala 31:69:@14639.4]
  wire  _T_2909; // @[package.scala 96:25:@14522.4 package.scala 96:25:@14523.4]
  wire [7:0] _T_2961; // @[Mux.scala 31:69:@14640.4]
  wire  _T_2906; // @[package.scala 96:25:@14514.4 package.scala 96:25:@14515.4]
  wire [7:0] _T_2962; // @[Mux.scala 31:69:@14641.4]
  wire  _T_2903; // @[package.scala 96:25:@14506.4 package.scala 96:25:@14507.4]
  wire  _T_3088; // @[package.scala 96:25:@14810.4 package.scala 96:25:@14811.4]
  wire [7:0] _T_3092; // @[Mux.scala 31:69:@14820.4]
  wire  _T_3085; // @[package.scala 96:25:@14802.4 package.scala 96:25:@14803.4]
  wire [7:0] _T_3093; // @[Mux.scala 31:69:@14821.4]
  wire  _T_3082; // @[package.scala 96:25:@14794.4 package.scala 96:25:@14795.4]
  wire [7:0] _T_3094; // @[Mux.scala 31:69:@14822.4]
  wire  _T_3079; // @[package.scala 96:25:@14786.4 package.scala 96:25:@14787.4]
  wire [7:0] _T_3095; // @[Mux.scala 31:69:@14823.4]
  wire  _T_3076; // @[package.scala 96:25:@14778.4 package.scala 96:25:@14779.4]
  wire [7:0] _T_3096; // @[Mux.scala 31:69:@14824.4]
  wire  _T_3073; // @[package.scala 96:25:@14770.4 package.scala 96:25:@14771.4]
  wire [7:0] _T_3097; // @[Mux.scala 31:69:@14825.4]
  wire  _T_3070; // @[package.scala 96:25:@14762.4 package.scala 96:25:@14763.4]
  wire [7:0] _T_3098; // @[Mux.scala 31:69:@14826.4]
  wire  _T_3067; // @[package.scala 96:25:@14754.4 package.scala 96:25:@14755.4]
  wire [7:0] _T_3099; // @[Mux.scala 31:69:@14827.4]
  wire  _T_3064; // @[package.scala 96:25:@14746.4 package.scala 96:25:@14747.4]
  wire [7:0] _T_3100; // @[Mux.scala 31:69:@14828.4]
  wire  _T_3061; // @[package.scala 96:25:@14738.4 package.scala 96:25:@14739.4]
  wire [7:0] _T_3101; // @[Mux.scala 31:69:@14829.4]
  wire  _T_3058; // @[package.scala 96:25:@14730.4 package.scala 96:25:@14731.4]
  wire [7:0] _T_3102; // @[Mux.scala 31:69:@14830.4]
  wire  _T_3055; // @[package.scala 96:25:@14722.4 package.scala 96:25:@14723.4]
  wire [7:0] _T_3103; // @[Mux.scala 31:69:@14831.4]
  wire  _T_3052; // @[package.scala 96:25:@14714.4 package.scala 96:25:@14715.4]
  wire [7:0] _T_3104; // @[Mux.scala 31:69:@14832.4]
  wire  _T_3049; // @[package.scala 96:25:@14706.4 package.scala 96:25:@14707.4]
  wire [7:0] _T_3105; // @[Mux.scala 31:69:@14833.4]
  wire  _T_3046; // @[package.scala 96:25:@14698.4 package.scala 96:25:@14699.4]
  wire  _T_3231; // @[package.scala 96:25:@15002.4 package.scala 96:25:@15003.4]
  wire [7:0] _T_3235; // @[Mux.scala 31:69:@15012.4]
  wire  _T_3228; // @[package.scala 96:25:@14994.4 package.scala 96:25:@14995.4]
  wire [7:0] _T_3236; // @[Mux.scala 31:69:@15013.4]
  wire  _T_3225; // @[package.scala 96:25:@14986.4 package.scala 96:25:@14987.4]
  wire [7:0] _T_3237; // @[Mux.scala 31:69:@15014.4]
  wire  _T_3222; // @[package.scala 96:25:@14978.4 package.scala 96:25:@14979.4]
  wire [7:0] _T_3238; // @[Mux.scala 31:69:@15015.4]
  wire  _T_3219; // @[package.scala 96:25:@14970.4 package.scala 96:25:@14971.4]
  wire [7:0] _T_3239; // @[Mux.scala 31:69:@15016.4]
  wire  _T_3216; // @[package.scala 96:25:@14962.4 package.scala 96:25:@14963.4]
  wire [7:0] _T_3240; // @[Mux.scala 31:69:@15017.4]
  wire  _T_3213; // @[package.scala 96:25:@14954.4 package.scala 96:25:@14955.4]
  wire [7:0] _T_3241; // @[Mux.scala 31:69:@15018.4]
  wire  _T_3210; // @[package.scala 96:25:@14946.4 package.scala 96:25:@14947.4]
  wire [7:0] _T_3242; // @[Mux.scala 31:69:@15019.4]
  wire  _T_3207; // @[package.scala 96:25:@14938.4 package.scala 96:25:@14939.4]
  wire [7:0] _T_3243; // @[Mux.scala 31:69:@15020.4]
  wire  _T_3204; // @[package.scala 96:25:@14930.4 package.scala 96:25:@14931.4]
  wire [7:0] _T_3244; // @[Mux.scala 31:69:@15021.4]
  wire  _T_3201; // @[package.scala 96:25:@14922.4 package.scala 96:25:@14923.4]
  wire [7:0] _T_3245; // @[Mux.scala 31:69:@15022.4]
  wire  _T_3198; // @[package.scala 96:25:@14914.4 package.scala 96:25:@14915.4]
  wire [7:0] _T_3246; // @[Mux.scala 31:69:@15023.4]
  wire  _T_3195; // @[package.scala 96:25:@14906.4 package.scala 96:25:@14907.4]
  wire [7:0] _T_3247; // @[Mux.scala 31:69:@15024.4]
  wire  _T_3192; // @[package.scala 96:25:@14898.4 package.scala 96:25:@14899.4]
  wire [7:0] _T_3248; // @[Mux.scala 31:69:@15025.4]
  wire  _T_3189; // @[package.scala 96:25:@14890.4 package.scala 96:25:@14891.4]
  Mem1D_4 Mem1D ( // @[MemPrimitives.scala 64:21:@11428.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  Mem1D_4 Mem1D_1 ( // @[MemPrimitives.scala 64:21:@11444.4]
    .clock(Mem1D_1_clock),
    .reset(Mem1D_1_reset),
    .io_r_ofs_0(Mem1D_1_io_r_ofs_0),
    .io_r_backpressure(Mem1D_1_io_r_backpressure),
    .io_w_ofs_0(Mem1D_1_io_w_ofs_0),
    .io_w_data_0(Mem1D_1_io_w_data_0),
    .io_w_en_0(Mem1D_1_io_w_en_0),
    .io_output(Mem1D_1_io_output)
  );
  Mem1D_4 Mem1D_2 ( // @[MemPrimitives.scala 64:21:@11460.4]
    .clock(Mem1D_2_clock),
    .reset(Mem1D_2_reset),
    .io_r_ofs_0(Mem1D_2_io_r_ofs_0),
    .io_r_backpressure(Mem1D_2_io_r_backpressure),
    .io_w_ofs_0(Mem1D_2_io_w_ofs_0),
    .io_w_data_0(Mem1D_2_io_w_data_0),
    .io_w_en_0(Mem1D_2_io_w_en_0),
    .io_output(Mem1D_2_io_output)
  );
  Mem1D_4 Mem1D_3 ( // @[MemPrimitives.scala 64:21:@11476.4]
    .clock(Mem1D_3_clock),
    .reset(Mem1D_3_reset),
    .io_r_ofs_0(Mem1D_3_io_r_ofs_0),
    .io_r_backpressure(Mem1D_3_io_r_backpressure),
    .io_w_ofs_0(Mem1D_3_io_w_ofs_0),
    .io_w_data_0(Mem1D_3_io_w_data_0),
    .io_w_en_0(Mem1D_3_io_w_en_0),
    .io_output(Mem1D_3_io_output)
  );
  Mem1D_4 Mem1D_4 ( // @[MemPrimitives.scala 64:21:@11492.4]
    .clock(Mem1D_4_clock),
    .reset(Mem1D_4_reset),
    .io_r_ofs_0(Mem1D_4_io_r_ofs_0),
    .io_r_backpressure(Mem1D_4_io_r_backpressure),
    .io_w_ofs_0(Mem1D_4_io_w_ofs_0),
    .io_w_data_0(Mem1D_4_io_w_data_0),
    .io_w_en_0(Mem1D_4_io_w_en_0),
    .io_output(Mem1D_4_io_output)
  );
  Mem1D_4 Mem1D_5 ( // @[MemPrimitives.scala 64:21:@11508.4]
    .clock(Mem1D_5_clock),
    .reset(Mem1D_5_reset),
    .io_r_ofs_0(Mem1D_5_io_r_ofs_0),
    .io_r_backpressure(Mem1D_5_io_r_backpressure),
    .io_w_ofs_0(Mem1D_5_io_w_ofs_0),
    .io_w_data_0(Mem1D_5_io_w_data_0),
    .io_w_en_0(Mem1D_5_io_w_en_0),
    .io_output(Mem1D_5_io_output)
  );
  Mem1D_4 Mem1D_6 ( // @[MemPrimitives.scala 64:21:@11524.4]
    .clock(Mem1D_6_clock),
    .reset(Mem1D_6_reset),
    .io_r_ofs_0(Mem1D_6_io_r_ofs_0),
    .io_r_backpressure(Mem1D_6_io_r_backpressure),
    .io_w_ofs_0(Mem1D_6_io_w_ofs_0),
    .io_w_data_0(Mem1D_6_io_w_data_0),
    .io_w_en_0(Mem1D_6_io_w_en_0),
    .io_output(Mem1D_6_io_output)
  );
  Mem1D_4 Mem1D_7 ( // @[MemPrimitives.scala 64:21:@11540.4]
    .clock(Mem1D_7_clock),
    .reset(Mem1D_7_reset),
    .io_r_ofs_0(Mem1D_7_io_r_ofs_0),
    .io_r_backpressure(Mem1D_7_io_r_backpressure),
    .io_w_ofs_0(Mem1D_7_io_w_ofs_0),
    .io_w_data_0(Mem1D_7_io_w_data_0),
    .io_w_en_0(Mem1D_7_io_w_en_0),
    .io_output(Mem1D_7_io_output)
  );
  Mem1D_4 Mem1D_8 ( // @[MemPrimitives.scala 64:21:@11556.4]
    .clock(Mem1D_8_clock),
    .reset(Mem1D_8_reset),
    .io_r_ofs_0(Mem1D_8_io_r_ofs_0),
    .io_r_backpressure(Mem1D_8_io_r_backpressure),
    .io_w_ofs_0(Mem1D_8_io_w_ofs_0),
    .io_w_data_0(Mem1D_8_io_w_data_0),
    .io_w_en_0(Mem1D_8_io_w_en_0),
    .io_output(Mem1D_8_io_output)
  );
  Mem1D_4 Mem1D_9 ( // @[MemPrimitives.scala 64:21:@11572.4]
    .clock(Mem1D_9_clock),
    .reset(Mem1D_9_reset),
    .io_r_ofs_0(Mem1D_9_io_r_ofs_0),
    .io_r_backpressure(Mem1D_9_io_r_backpressure),
    .io_w_ofs_0(Mem1D_9_io_w_ofs_0),
    .io_w_data_0(Mem1D_9_io_w_data_0),
    .io_w_en_0(Mem1D_9_io_w_en_0),
    .io_output(Mem1D_9_io_output)
  );
  Mem1D_4 Mem1D_10 ( // @[MemPrimitives.scala 64:21:@11588.4]
    .clock(Mem1D_10_clock),
    .reset(Mem1D_10_reset),
    .io_r_ofs_0(Mem1D_10_io_r_ofs_0),
    .io_r_backpressure(Mem1D_10_io_r_backpressure),
    .io_w_ofs_0(Mem1D_10_io_w_ofs_0),
    .io_w_data_0(Mem1D_10_io_w_data_0),
    .io_w_en_0(Mem1D_10_io_w_en_0),
    .io_output(Mem1D_10_io_output)
  );
  Mem1D_4 Mem1D_11 ( // @[MemPrimitives.scala 64:21:@11604.4]
    .clock(Mem1D_11_clock),
    .reset(Mem1D_11_reset),
    .io_r_ofs_0(Mem1D_11_io_r_ofs_0),
    .io_r_backpressure(Mem1D_11_io_r_backpressure),
    .io_w_ofs_0(Mem1D_11_io_w_ofs_0),
    .io_w_data_0(Mem1D_11_io_w_data_0),
    .io_w_en_0(Mem1D_11_io_w_en_0),
    .io_output(Mem1D_11_io_output)
  );
  Mem1D_4 Mem1D_12 ( // @[MemPrimitives.scala 64:21:@11620.4]
    .clock(Mem1D_12_clock),
    .reset(Mem1D_12_reset),
    .io_r_ofs_0(Mem1D_12_io_r_ofs_0),
    .io_r_backpressure(Mem1D_12_io_r_backpressure),
    .io_w_ofs_0(Mem1D_12_io_w_ofs_0),
    .io_w_data_0(Mem1D_12_io_w_data_0),
    .io_w_en_0(Mem1D_12_io_w_en_0),
    .io_output(Mem1D_12_io_output)
  );
  Mem1D_4 Mem1D_13 ( // @[MemPrimitives.scala 64:21:@11636.4]
    .clock(Mem1D_13_clock),
    .reset(Mem1D_13_reset),
    .io_r_ofs_0(Mem1D_13_io_r_ofs_0),
    .io_r_backpressure(Mem1D_13_io_r_backpressure),
    .io_w_ofs_0(Mem1D_13_io_w_ofs_0),
    .io_w_data_0(Mem1D_13_io_w_data_0),
    .io_w_en_0(Mem1D_13_io_w_en_0),
    .io_output(Mem1D_13_io_output)
  );
  Mem1D_4 Mem1D_14 ( // @[MemPrimitives.scala 64:21:@11652.4]
    .clock(Mem1D_14_clock),
    .reset(Mem1D_14_reset),
    .io_r_ofs_0(Mem1D_14_io_r_ofs_0),
    .io_r_backpressure(Mem1D_14_io_r_backpressure),
    .io_w_ofs_0(Mem1D_14_io_w_ofs_0),
    .io_w_data_0(Mem1D_14_io_w_data_0),
    .io_w_en_0(Mem1D_14_io_w_en_0),
    .io_output(Mem1D_14_io_output)
  );
  Mem1D_4 Mem1D_15 ( // @[MemPrimitives.scala 64:21:@11668.4]
    .clock(Mem1D_15_clock),
    .reset(Mem1D_15_reset),
    .io_r_ofs_0(Mem1D_15_io_r_ofs_0),
    .io_r_backpressure(Mem1D_15_io_r_backpressure),
    .io_w_ofs_0(Mem1D_15_io_w_ofs_0),
    .io_w_data_0(Mem1D_15_io_w_data_0),
    .io_w_en_0(Mem1D_15_io_w_en_0),
    .io_output(Mem1D_15_io_output)
  );
  StickySelects StickySelects ( // @[MemPrimitives.scala 121:29:@11912.4]
    .clock(StickySelects_clock),
    .reset(StickySelects_reset),
    .io_ins_0(StickySelects_io_ins_0),
    .io_ins_1(StickySelects_io_ins_1),
    .io_ins_2(StickySelects_io_ins_2),
    .io_ins_3(StickySelects_io_ins_3),
    .io_ins_4(StickySelects_io_ins_4),
    .io_ins_5(StickySelects_io_ins_5),
    .io_ins_6(StickySelects_io_ins_6),
    .io_ins_7(StickySelects_io_ins_7),
    .io_ins_8(StickySelects_io_ins_8),
    .io_outs_0(StickySelects_io_outs_0),
    .io_outs_1(StickySelects_io_outs_1),
    .io_outs_2(StickySelects_io_outs_2),
    .io_outs_3(StickySelects_io_outs_3),
    .io_outs_4(StickySelects_io_outs_4),
    .io_outs_5(StickySelects_io_outs_5),
    .io_outs_6(StickySelects_io_outs_6),
    .io_outs_7(StickySelects_io_outs_7),
    .io_outs_8(StickySelects_io_outs_8)
  );
  StickySelects StickySelects_1 ( // @[MemPrimitives.scala 121:29:@12001.4]
    .clock(StickySelects_1_clock),
    .reset(StickySelects_1_reset),
    .io_ins_0(StickySelects_1_io_ins_0),
    .io_ins_1(StickySelects_1_io_ins_1),
    .io_ins_2(StickySelects_1_io_ins_2),
    .io_ins_3(StickySelects_1_io_ins_3),
    .io_ins_4(StickySelects_1_io_ins_4),
    .io_ins_5(StickySelects_1_io_ins_5),
    .io_ins_6(StickySelects_1_io_ins_6),
    .io_ins_7(StickySelects_1_io_ins_7),
    .io_ins_8(StickySelects_1_io_ins_8),
    .io_outs_0(StickySelects_1_io_outs_0),
    .io_outs_1(StickySelects_1_io_outs_1),
    .io_outs_2(StickySelects_1_io_outs_2),
    .io_outs_3(StickySelects_1_io_outs_3),
    .io_outs_4(StickySelects_1_io_outs_4),
    .io_outs_5(StickySelects_1_io_outs_5),
    .io_outs_6(StickySelects_1_io_outs_6),
    .io_outs_7(StickySelects_1_io_outs_7),
    .io_outs_8(StickySelects_1_io_outs_8)
  );
  StickySelects StickySelects_2 ( // @[MemPrimitives.scala 121:29:@12090.4]
    .clock(StickySelects_2_clock),
    .reset(StickySelects_2_reset),
    .io_ins_0(StickySelects_2_io_ins_0),
    .io_ins_1(StickySelects_2_io_ins_1),
    .io_ins_2(StickySelects_2_io_ins_2),
    .io_ins_3(StickySelects_2_io_ins_3),
    .io_ins_4(StickySelects_2_io_ins_4),
    .io_ins_5(StickySelects_2_io_ins_5),
    .io_ins_6(StickySelects_2_io_ins_6),
    .io_ins_7(StickySelects_2_io_ins_7),
    .io_ins_8(StickySelects_2_io_ins_8),
    .io_outs_0(StickySelects_2_io_outs_0),
    .io_outs_1(StickySelects_2_io_outs_1),
    .io_outs_2(StickySelects_2_io_outs_2),
    .io_outs_3(StickySelects_2_io_outs_3),
    .io_outs_4(StickySelects_2_io_outs_4),
    .io_outs_5(StickySelects_2_io_outs_5),
    .io_outs_6(StickySelects_2_io_outs_6),
    .io_outs_7(StickySelects_2_io_outs_7),
    .io_outs_8(StickySelects_2_io_outs_8)
  );
  StickySelects StickySelects_3 ( // @[MemPrimitives.scala 121:29:@12179.4]
    .clock(StickySelects_3_clock),
    .reset(StickySelects_3_reset),
    .io_ins_0(StickySelects_3_io_ins_0),
    .io_ins_1(StickySelects_3_io_ins_1),
    .io_ins_2(StickySelects_3_io_ins_2),
    .io_ins_3(StickySelects_3_io_ins_3),
    .io_ins_4(StickySelects_3_io_ins_4),
    .io_ins_5(StickySelects_3_io_ins_5),
    .io_ins_6(StickySelects_3_io_ins_6),
    .io_ins_7(StickySelects_3_io_ins_7),
    .io_ins_8(StickySelects_3_io_ins_8),
    .io_outs_0(StickySelects_3_io_outs_0),
    .io_outs_1(StickySelects_3_io_outs_1),
    .io_outs_2(StickySelects_3_io_outs_2),
    .io_outs_3(StickySelects_3_io_outs_3),
    .io_outs_4(StickySelects_3_io_outs_4),
    .io_outs_5(StickySelects_3_io_outs_5),
    .io_outs_6(StickySelects_3_io_outs_6),
    .io_outs_7(StickySelects_3_io_outs_7),
    .io_outs_8(StickySelects_3_io_outs_8)
  );
  StickySelects StickySelects_4 ( // @[MemPrimitives.scala 121:29:@12268.4]
    .clock(StickySelects_4_clock),
    .reset(StickySelects_4_reset),
    .io_ins_0(StickySelects_4_io_ins_0),
    .io_ins_1(StickySelects_4_io_ins_1),
    .io_ins_2(StickySelects_4_io_ins_2),
    .io_ins_3(StickySelects_4_io_ins_3),
    .io_ins_4(StickySelects_4_io_ins_4),
    .io_ins_5(StickySelects_4_io_ins_5),
    .io_ins_6(StickySelects_4_io_ins_6),
    .io_ins_7(StickySelects_4_io_ins_7),
    .io_ins_8(StickySelects_4_io_ins_8),
    .io_outs_0(StickySelects_4_io_outs_0),
    .io_outs_1(StickySelects_4_io_outs_1),
    .io_outs_2(StickySelects_4_io_outs_2),
    .io_outs_3(StickySelects_4_io_outs_3),
    .io_outs_4(StickySelects_4_io_outs_4),
    .io_outs_5(StickySelects_4_io_outs_5),
    .io_outs_6(StickySelects_4_io_outs_6),
    .io_outs_7(StickySelects_4_io_outs_7),
    .io_outs_8(StickySelects_4_io_outs_8)
  );
  StickySelects StickySelects_5 ( // @[MemPrimitives.scala 121:29:@12357.4]
    .clock(StickySelects_5_clock),
    .reset(StickySelects_5_reset),
    .io_ins_0(StickySelects_5_io_ins_0),
    .io_ins_1(StickySelects_5_io_ins_1),
    .io_ins_2(StickySelects_5_io_ins_2),
    .io_ins_3(StickySelects_5_io_ins_3),
    .io_ins_4(StickySelects_5_io_ins_4),
    .io_ins_5(StickySelects_5_io_ins_5),
    .io_ins_6(StickySelects_5_io_ins_6),
    .io_ins_7(StickySelects_5_io_ins_7),
    .io_ins_8(StickySelects_5_io_ins_8),
    .io_outs_0(StickySelects_5_io_outs_0),
    .io_outs_1(StickySelects_5_io_outs_1),
    .io_outs_2(StickySelects_5_io_outs_2),
    .io_outs_3(StickySelects_5_io_outs_3),
    .io_outs_4(StickySelects_5_io_outs_4),
    .io_outs_5(StickySelects_5_io_outs_5),
    .io_outs_6(StickySelects_5_io_outs_6),
    .io_outs_7(StickySelects_5_io_outs_7),
    .io_outs_8(StickySelects_5_io_outs_8)
  );
  StickySelects StickySelects_6 ( // @[MemPrimitives.scala 121:29:@12446.4]
    .clock(StickySelects_6_clock),
    .reset(StickySelects_6_reset),
    .io_ins_0(StickySelects_6_io_ins_0),
    .io_ins_1(StickySelects_6_io_ins_1),
    .io_ins_2(StickySelects_6_io_ins_2),
    .io_ins_3(StickySelects_6_io_ins_3),
    .io_ins_4(StickySelects_6_io_ins_4),
    .io_ins_5(StickySelects_6_io_ins_5),
    .io_ins_6(StickySelects_6_io_ins_6),
    .io_ins_7(StickySelects_6_io_ins_7),
    .io_ins_8(StickySelects_6_io_ins_8),
    .io_outs_0(StickySelects_6_io_outs_0),
    .io_outs_1(StickySelects_6_io_outs_1),
    .io_outs_2(StickySelects_6_io_outs_2),
    .io_outs_3(StickySelects_6_io_outs_3),
    .io_outs_4(StickySelects_6_io_outs_4),
    .io_outs_5(StickySelects_6_io_outs_5),
    .io_outs_6(StickySelects_6_io_outs_6),
    .io_outs_7(StickySelects_6_io_outs_7),
    .io_outs_8(StickySelects_6_io_outs_8)
  );
  StickySelects StickySelects_7 ( // @[MemPrimitives.scala 121:29:@12535.4]
    .clock(StickySelects_7_clock),
    .reset(StickySelects_7_reset),
    .io_ins_0(StickySelects_7_io_ins_0),
    .io_ins_1(StickySelects_7_io_ins_1),
    .io_ins_2(StickySelects_7_io_ins_2),
    .io_ins_3(StickySelects_7_io_ins_3),
    .io_ins_4(StickySelects_7_io_ins_4),
    .io_ins_5(StickySelects_7_io_ins_5),
    .io_ins_6(StickySelects_7_io_ins_6),
    .io_ins_7(StickySelects_7_io_ins_7),
    .io_ins_8(StickySelects_7_io_ins_8),
    .io_outs_0(StickySelects_7_io_outs_0),
    .io_outs_1(StickySelects_7_io_outs_1),
    .io_outs_2(StickySelects_7_io_outs_2),
    .io_outs_3(StickySelects_7_io_outs_3),
    .io_outs_4(StickySelects_7_io_outs_4),
    .io_outs_5(StickySelects_7_io_outs_5),
    .io_outs_6(StickySelects_7_io_outs_6),
    .io_outs_7(StickySelects_7_io_outs_7),
    .io_outs_8(StickySelects_7_io_outs_8)
  );
  StickySelects StickySelects_8 ( // @[MemPrimitives.scala 121:29:@12624.4]
    .clock(StickySelects_8_clock),
    .reset(StickySelects_8_reset),
    .io_ins_0(StickySelects_8_io_ins_0),
    .io_ins_1(StickySelects_8_io_ins_1),
    .io_ins_2(StickySelects_8_io_ins_2),
    .io_ins_3(StickySelects_8_io_ins_3),
    .io_ins_4(StickySelects_8_io_ins_4),
    .io_ins_5(StickySelects_8_io_ins_5),
    .io_ins_6(StickySelects_8_io_ins_6),
    .io_ins_7(StickySelects_8_io_ins_7),
    .io_ins_8(StickySelects_8_io_ins_8),
    .io_outs_0(StickySelects_8_io_outs_0),
    .io_outs_1(StickySelects_8_io_outs_1),
    .io_outs_2(StickySelects_8_io_outs_2),
    .io_outs_3(StickySelects_8_io_outs_3),
    .io_outs_4(StickySelects_8_io_outs_4),
    .io_outs_5(StickySelects_8_io_outs_5),
    .io_outs_6(StickySelects_8_io_outs_6),
    .io_outs_7(StickySelects_8_io_outs_7),
    .io_outs_8(StickySelects_8_io_outs_8)
  );
  StickySelects StickySelects_9 ( // @[MemPrimitives.scala 121:29:@12713.4]
    .clock(StickySelects_9_clock),
    .reset(StickySelects_9_reset),
    .io_ins_0(StickySelects_9_io_ins_0),
    .io_ins_1(StickySelects_9_io_ins_1),
    .io_ins_2(StickySelects_9_io_ins_2),
    .io_ins_3(StickySelects_9_io_ins_3),
    .io_ins_4(StickySelects_9_io_ins_4),
    .io_ins_5(StickySelects_9_io_ins_5),
    .io_ins_6(StickySelects_9_io_ins_6),
    .io_ins_7(StickySelects_9_io_ins_7),
    .io_ins_8(StickySelects_9_io_ins_8),
    .io_outs_0(StickySelects_9_io_outs_0),
    .io_outs_1(StickySelects_9_io_outs_1),
    .io_outs_2(StickySelects_9_io_outs_2),
    .io_outs_3(StickySelects_9_io_outs_3),
    .io_outs_4(StickySelects_9_io_outs_4),
    .io_outs_5(StickySelects_9_io_outs_5),
    .io_outs_6(StickySelects_9_io_outs_6),
    .io_outs_7(StickySelects_9_io_outs_7),
    .io_outs_8(StickySelects_9_io_outs_8)
  );
  StickySelects StickySelects_10 ( // @[MemPrimitives.scala 121:29:@12802.4]
    .clock(StickySelects_10_clock),
    .reset(StickySelects_10_reset),
    .io_ins_0(StickySelects_10_io_ins_0),
    .io_ins_1(StickySelects_10_io_ins_1),
    .io_ins_2(StickySelects_10_io_ins_2),
    .io_ins_3(StickySelects_10_io_ins_3),
    .io_ins_4(StickySelects_10_io_ins_4),
    .io_ins_5(StickySelects_10_io_ins_5),
    .io_ins_6(StickySelects_10_io_ins_6),
    .io_ins_7(StickySelects_10_io_ins_7),
    .io_ins_8(StickySelects_10_io_ins_8),
    .io_outs_0(StickySelects_10_io_outs_0),
    .io_outs_1(StickySelects_10_io_outs_1),
    .io_outs_2(StickySelects_10_io_outs_2),
    .io_outs_3(StickySelects_10_io_outs_3),
    .io_outs_4(StickySelects_10_io_outs_4),
    .io_outs_5(StickySelects_10_io_outs_5),
    .io_outs_6(StickySelects_10_io_outs_6),
    .io_outs_7(StickySelects_10_io_outs_7),
    .io_outs_8(StickySelects_10_io_outs_8)
  );
  StickySelects StickySelects_11 ( // @[MemPrimitives.scala 121:29:@12891.4]
    .clock(StickySelects_11_clock),
    .reset(StickySelects_11_reset),
    .io_ins_0(StickySelects_11_io_ins_0),
    .io_ins_1(StickySelects_11_io_ins_1),
    .io_ins_2(StickySelects_11_io_ins_2),
    .io_ins_3(StickySelects_11_io_ins_3),
    .io_ins_4(StickySelects_11_io_ins_4),
    .io_ins_5(StickySelects_11_io_ins_5),
    .io_ins_6(StickySelects_11_io_ins_6),
    .io_ins_7(StickySelects_11_io_ins_7),
    .io_ins_8(StickySelects_11_io_ins_8),
    .io_outs_0(StickySelects_11_io_outs_0),
    .io_outs_1(StickySelects_11_io_outs_1),
    .io_outs_2(StickySelects_11_io_outs_2),
    .io_outs_3(StickySelects_11_io_outs_3),
    .io_outs_4(StickySelects_11_io_outs_4),
    .io_outs_5(StickySelects_11_io_outs_5),
    .io_outs_6(StickySelects_11_io_outs_6),
    .io_outs_7(StickySelects_11_io_outs_7),
    .io_outs_8(StickySelects_11_io_outs_8)
  );
  StickySelects StickySelects_12 ( // @[MemPrimitives.scala 121:29:@12980.4]
    .clock(StickySelects_12_clock),
    .reset(StickySelects_12_reset),
    .io_ins_0(StickySelects_12_io_ins_0),
    .io_ins_1(StickySelects_12_io_ins_1),
    .io_ins_2(StickySelects_12_io_ins_2),
    .io_ins_3(StickySelects_12_io_ins_3),
    .io_ins_4(StickySelects_12_io_ins_4),
    .io_ins_5(StickySelects_12_io_ins_5),
    .io_ins_6(StickySelects_12_io_ins_6),
    .io_ins_7(StickySelects_12_io_ins_7),
    .io_ins_8(StickySelects_12_io_ins_8),
    .io_outs_0(StickySelects_12_io_outs_0),
    .io_outs_1(StickySelects_12_io_outs_1),
    .io_outs_2(StickySelects_12_io_outs_2),
    .io_outs_3(StickySelects_12_io_outs_3),
    .io_outs_4(StickySelects_12_io_outs_4),
    .io_outs_5(StickySelects_12_io_outs_5),
    .io_outs_6(StickySelects_12_io_outs_6),
    .io_outs_7(StickySelects_12_io_outs_7),
    .io_outs_8(StickySelects_12_io_outs_8)
  );
  StickySelects StickySelects_13 ( // @[MemPrimitives.scala 121:29:@13069.4]
    .clock(StickySelects_13_clock),
    .reset(StickySelects_13_reset),
    .io_ins_0(StickySelects_13_io_ins_0),
    .io_ins_1(StickySelects_13_io_ins_1),
    .io_ins_2(StickySelects_13_io_ins_2),
    .io_ins_3(StickySelects_13_io_ins_3),
    .io_ins_4(StickySelects_13_io_ins_4),
    .io_ins_5(StickySelects_13_io_ins_5),
    .io_ins_6(StickySelects_13_io_ins_6),
    .io_ins_7(StickySelects_13_io_ins_7),
    .io_ins_8(StickySelects_13_io_ins_8),
    .io_outs_0(StickySelects_13_io_outs_0),
    .io_outs_1(StickySelects_13_io_outs_1),
    .io_outs_2(StickySelects_13_io_outs_2),
    .io_outs_3(StickySelects_13_io_outs_3),
    .io_outs_4(StickySelects_13_io_outs_4),
    .io_outs_5(StickySelects_13_io_outs_5),
    .io_outs_6(StickySelects_13_io_outs_6),
    .io_outs_7(StickySelects_13_io_outs_7),
    .io_outs_8(StickySelects_13_io_outs_8)
  );
  StickySelects StickySelects_14 ( // @[MemPrimitives.scala 121:29:@13158.4]
    .clock(StickySelects_14_clock),
    .reset(StickySelects_14_reset),
    .io_ins_0(StickySelects_14_io_ins_0),
    .io_ins_1(StickySelects_14_io_ins_1),
    .io_ins_2(StickySelects_14_io_ins_2),
    .io_ins_3(StickySelects_14_io_ins_3),
    .io_ins_4(StickySelects_14_io_ins_4),
    .io_ins_5(StickySelects_14_io_ins_5),
    .io_ins_6(StickySelects_14_io_ins_6),
    .io_ins_7(StickySelects_14_io_ins_7),
    .io_ins_8(StickySelects_14_io_ins_8),
    .io_outs_0(StickySelects_14_io_outs_0),
    .io_outs_1(StickySelects_14_io_outs_1),
    .io_outs_2(StickySelects_14_io_outs_2),
    .io_outs_3(StickySelects_14_io_outs_3),
    .io_outs_4(StickySelects_14_io_outs_4),
    .io_outs_5(StickySelects_14_io_outs_5),
    .io_outs_6(StickySelects_14_io_outs_6),
    .io_outs_7(StickySelects_14_io_outs_7),
    .io_outs_8(StickySelects_14_io_outs_8)
  );
  StickySelects StickySelects_15 ( // @[MemPrimitives.scala 121:29:@13247.4]
    .clock(StickySelects_15_clock),
    .reset(StickySelects_15_reset),
    .io_ins_0(StickySelects_15_io_ins_0),
    .io_ins_1(StickySelects_15_io_ins_1),
    .io_ins_2(StickySelects_15_io_ins_2),
    .io_ins_3(StickySelects_15_io_ins_3),
    .io_ins_4(StickySelects_15_io_ins_4),
    .io_ins_5(StickySelects_15_io_ins_5),
    .io_ins_6(StickySelects_15_io_ins_6),
    .io_ins_7(StickySelects_15_io_ins_7),
    .io_ins_8(StickySelects_15_io_ins_8),
    .io_outs_0(StickySelects_15_io_outs_0),
    .io_outs_1(StickySelects_15_io_outs_1),
    .io_outs_2(StickySelects_15_io_outs_2),
    .io_outs_3(StickySelects_15_io_outs_3),
    .io_outs_4(StickySelects_15_io_outs_4),
    .io_outs_5(StickySelects_15_io_outs_5),
    .io_outs_6(StickySelects_15_io_outs_6),
    .io_outs_7(StickySelects_15_io_outs_7),
    .io_outs_8(StickySelects_15_io_outs_8)
  );
  RetimeWrapper_52 RetimeWrapper ( // @[package.scala 93:22:@13349.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_1 ( // @[package.scala 93:22:@13357.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_2 ( // @[package.scala 93:22:@13365.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_3 ( // @[package.scala 93:22:@13373.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_4 ( // @[package.scala 93:22:@13381.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_5 ( // @[package.scala 93:22:@13389.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_6 ( // @[package.scala 93:22:@13397.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_7 ( // @[package.scala 93:22:@13405.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_8 ( // @[package.scala 93:22:@13413.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_9 ( // @[package.scala 93:22:@13421.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_10 ( // @[package.scala 93:22:@13429.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_11 ( // @[package.scala 93:22:@13437.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_12 ( // @[package.scala 93:22:@13445.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_13 ( // @[package.scala 93:22:@13453.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_14 ( // @[package.scala 93:22:@13461.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_15 ( // @[package.scala 93:22:@13469.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_16 ( // @[package.scala 93:22:@13541.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_17 ( // @[package.scala 93:22:@13549.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_18 ( // @[package.scala 93:22:@13557.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_19 ( // @[package.scala 93:22:@13565.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_20 ( // @[package.scala 93:22:@13573.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_21 ( // @[package.scala 93:22:@13581.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_22 ( // @[package.scala 93:22:@13589.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_23 ( // @[package.scala 93:22:@13597.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_24 ( // @[package.scala 93:22:@13605.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_25 ( // @[package.scala 93:22:@13613.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_26 ( // @[package.scala 93:22:@13621.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_27 ( // @[package.scala 93:22:@13629.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_28 ( // @[package.scala 93:22:@13637.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_29 ( // @[package.scala 93:22:@13645.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_30 ( // @[package.scala 93:22:@13653.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_31 ( // @[package.scala 93:22:@13661.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_32 ( // @[package.scala 93:22:@13733.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_33 ( // @[package.scala 93:22:@13741.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_34 ( // @[package.scala 93:22:@13749.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_35 ( // @[package.scala 93:22:@13757.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_36 ( // @[package.scala 93:22:@13765.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_37 ( // @[package.scala 93:22:@13773.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_38 ( // @[package.scala 93:22:@13781.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_39 ( // @[package.scala 93:22:@13789.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_40 ( // @[package.scala 93:22:@13797.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_41 ( // @[package.scala 93:22:@13805.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_42 ( // @[package.scala 93:22:@13813.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_43 ( // @[package.scala 93:22:@13821.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_44 ( // @[package.scala 93:22:@13829.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_45 ( // @[package.scala 93:22:@13837.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_46 ( // @[package.scala 93:22:@13845.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_47 ( // @[package.scala 93:22:@13853.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_48 ( // @[package.scala 93:22:@13925.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_49 ( // @[package.scala 93:22:@13933.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_50 ( // @[package.scala 93:22:@13941.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_51 ( // @[package.scala 93:22:@13949.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_52 ( // @[package.scala 93:22:@13957.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_53 ( // @[package.scala 93:22:@13965.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_54 ( // @[package.scala 93:22:@13973.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_55 ( // @[package.scala 93:22:@13981.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_56 ( // @[package.scala 93:22:@13989.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_57 ( // @[package.scala 93:22:@13997.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_58 ( // @[package.scala 93:22:@14005.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_59 ( // @[package.scala 93:22:@14013.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_60 ( // @[package.scala 93:22:@14021.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_61 ( // @[package.scala 93:22:@14029.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_62 ( // @[package.scala 93:22:@14037.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_63 ( // @[package.scala 93:22:@14045.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_64 ( // @[package.scala 93:22:@14117.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_65 ( // @[package.scala 93:22:@14125.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_66 ( // @[package.scala 93:22:@14133.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_67 ( // @[package.scala 93:22:@14141.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_68 ( // @[package.scala 93:22:@14149.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_69 ( // @[package.scala 93:22:@14157.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_70 ( // @[package.scala 93:22:@14165.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_71 ( // @[package.scala 93:22:@14173.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_72 ( // @[package.scala 93:22:@14181.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_73 ( // @[package.scala 93:22:@14189.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_74 ( // @[package.scala 93:22:@14197.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_75 ( // @[package.scala 93:22:@14205.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_76 ( // @[package.scala 93:22:@14213.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_77 ( // @[package.scala 93:22:@14221.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_78 ( // @[package.scala 93:22:@14229.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_79 ( // @[package.scala 93:22:@14237.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_80 ( // @[package.scala 93:22:@14309.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_81 ( // @[package.scala 93:22:@14317.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_82 ( // @[package.scala 93:22:@14325.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_83 ( // @[package.scala 93:22:@14333.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_84 ( // @[package.scala 93:22:@14341.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_85 ( // @[package.scala 93:22:@14349.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_86 ( // @[package.scala 93:22:@14357.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_87 ( // @[package.scala 93:22:@14365.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_88 ( // @[package.scala 93:22:@14373.4]
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_89 ( // @[package.scala 93:22:@14381.4]
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_90 ( // @[package.scala 93:22:@14389.4]
    .clock(RetimeWrapper_90_clock),
    .reset(RetimeWrapper_90_reset),
    .io_flow(RetimeWrapper_90_io_flow),
    .io_in(RetimeWrapper_90_io_in),
    .io_out(RetimeWrapper_90_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_91 ( // @[package.scala 93:22:@14397.4]
    .clock(RetimeWrapper_91_clock),
    .reset(RetimeWrapper_91_reset),
    .io_flow(RetimeWrapper_91_io_flow),
    .io_in(RetimeWrapper_91_io_in),
    .io_out(RetimeWrapper_91_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_92 ( // @[package.scala 93:22:@14405.4]
    .clock(RetimeWrapper_92_clock),
    .reset(RetimeWrapper_92_reset),
    .io_flow(RetimeWrapper_92_io_flow),
    .io_in(RetimeWrapper_92_io_in),
    .io_out(RetimeWrapper_92_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_93 ( // @[package.scala 93:22:@14413.4]
    .clock(RetimeWrapper_93_clock),
    .reset(RetimeWrapper_93_reset),
    .io_flow(RetimeWrapper_93_io_flow),
    .io_in(RetimeWrapper_93_io_in),
    .io_out(RetimeWrapper_93_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_94 ( // @[package.scala 93:22:@14421.4]
    .clock(RetimeWrapper_94_clock),
    .reset(RetimeWrapper_94_reset),
    .io_flow(RetimeWrapper_94_io_flow),
    .io_in(RetimeWrapper_94_io_in),
    .io_out(RetimeWrapper_94_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_95 ( // @[package.scala 93:22:@14429.4]
    .clock(RetimeWrapper_95_clock),
    .reset(RetimeWrapper_95_reset),
    .io_flow(RetimeWrapper_95_io_flow),
    .io_in(RetimeWrapper_95_io_in),
    .io_out(RetimeWrapper_95_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_96 ( // @[package.scala 93:22:@14501.4]
    .clock(RetimeWrapper_96_clock),
    .reset(RetimeWrapper_96_reset),
    .io_flow(RetimeWrapper_96_io_flow),
    .io_in(RetimeWrapper_96_io_in),
    .io_out(RetimeWrapper_96_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_97 ( // @[package.scala 93:22:@14509.4]
    .clock(RetimeWrapper_97_clock),
    .reset(RetimeWrapper_97_reset),
    .io_flow(RetimeWrapper_97_io_flow),
    .io_in(RetimeWrapper_97_io_in),
    .io_out(RetimeWrapper_97_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_98 ( // @[package.scala 93:22:@14517.4]
    .clock(RetimeWrapper_98_clock),
    .reset(RetimeWrapper_98_reset),
    .io_flow(RetimeWrapper_98_io_flow),
    .io_in(RetimeWrapper_98_io_in),
    .io_out(RetimeWrapper_98_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_99 ( // @[package.scala 93:22:@14525.4]
    .clock(RetimeWrapper_99_clock),
    .reset(RetimeWrapper_99_reset),
    .io_flow(RetimeWrapper_99_io_flow),
    .io_in(RetimeWrapper_99_io_in),
    .io_out(RetimeWrapper_99_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_100 ( // @[package.scala 93:22:@14533.4]
    .clock(RetimeWrapper_100_clock),
    .reset(RetimeWrapper_100_reset),
    .io_flow(RetimeWrapper_100_io_flow),
    .io_in(RetimeWrapper_100_io_in),
    .io_out(RetimeWrapper_100_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_101 ( // @[package.scala 93:22:@14541.4]
    .clock(RetimeWrapper_101_clock),
    .reset(RetimeWrapper_101_reset),
    .io_flow(RetimeWrapper_101_io_flow),
    .io_in(RetimeWrapper_101_io_in),
    .io_out(RetimeWrapper_101_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_102 ( // @[package.scala 93:22:@14549.4]
    .clock(RetimeWrapper_102_clock),
    .reset(RetimeWrapper_102_reset),
    .io_flow(RetimeWrapper_102_io_flow),
    .io_in(RetimeWrapper_102_io_in),
    .io_out(RetimeWrapper_102_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_103 ( // @[package.scala 93:22:@14557.4]
    .clock(RetimeWrapper_103_clock),
    .reset(RetimeWrapper_103_reset),
    .io_flow(RetimeWrapper_103_io_flow),
    .io_in(RetimeWrapper_103_io_in),
    .io_out(RetimeWrapper_103_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_104 ( // @[package.scala 93:22:@14565.4]
    .clock(RetimeWrapper_104_clock),
    .reset(RetimeWrapper_104_reset),
    .io_flow(RetimeWrapper_104_io_flow),
    .io_in(RetimeWrapper_104_io_in),
    .io_out(RetimeWrapper_104_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_105 ( // @[package.scala 93:22:@14573.4]
    .clock(RetimeWrapper_105_clock),
    .reset(RetimeWrapper_105_reset),
    .io_flow(RetimeWrapper_105_io_flow),
    .io_in(RetimeWrapper_105_io_in),
    .io_out(RetimeWrapper_105_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_106 ( // @[package.scala 93:22:@14581.4]
    .clock(RetimeWrapper_106_clock),
    .reset(RetimeWrapper_106_reset),
    .io_flow(RetimeWrapper_106_io_flow),
    .io_in(RetimeWrapper_106_io_in),
    .io_out(RetimeWrapper_106_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_107 ( // @[package.scala 93:22:@14589.4]
    .clock(RetimeWrapper_107_clock),
    .reset(RetimeWrapper_107_reset),
    .io_flow(RetimeWrapper_107_io_flow),
    .io_in(RetimeWrapper_107_io_in),
    .io_out(RetimeWrapper_107_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_108 ( // @[package.scala 93:22:@14597.4]
    .clock(RetimeWrapper_108_clock),
    .reset(RetimeWrapper_108_reset),
    .io_flow(RetimeWrapper_108_io_flow),
    .io_in(RetimeWrapper_108_io_in),
    .io_out(RetimeWrapper_108_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_109 ( // @[package.scala 93:22:@14605.4]
    .clock(RetimeWrapper_109_clock),
    .reset(RetimeWrapper_109_reset),
    .io_flow(RetimeWrapper_109_io_flow),
    .io_in(RetimeWrapper_109_io_in),
    .io_out(RetimeWrapper_109_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_110 ( // @[package.scala 93:22:@14613.4]
    .clock(RetimeWrapper_110_clock),
    .reset(RetimeWrapper_110_reset),
    .io_flow(RetimeWrapper_110_io_flow),
    .io_in(RetimeWrapper_110_io_in),
    .io_out(RetimeWrapper_110_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_111 ( // @[package.scala 93:22:@14621.4]
    .clock(RetimeWrapper_111_clock),
    .reset(RetimeWrapper_111_reset),
    .io_flow(RetimeWrapper_111_io_flow),
    .io_in(RetimeWrapper_111_io_in),
    .io_out(RetimeWrapper_111_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_112 ( // @[package.scala 93:22:@14693.4]
    .clock(RetimeWrapper_112_clock),
    .reset(RetimeWrapper_112_reset),
    .io_flow(RetimeWrapper_112_io_flow),
    .io_in(RetimeWrapper_112_io_in),
    .io_out(RetimeWrapper_112_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_113 ( // @[package.scala 93:22:@14701.4]
    .clock(RetimeWrapper_113_clock),
    .reset(RetimeWrapper_113_reset),
    .io_flow(RetimeWrapper_113_io_flow),
    .io_in(RetimeWrapper_113_io_in),
    .io_out(RetimeWrapper_113_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_114 ( // @[package.scala 93:22:@14709.4]
    .clock(RetimeWrapper_114_clock),
    .reset(RetimeWrapper_114_reset),
    .io_flow(RetimeWrapper_114_io_flow),
    .io_in(RetimeWrapper_114_io_in),
    .io_out(RetimeWrapper_114_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_115 ( // @[package.scala 93:22:@14717.4]
    .clock(RetimeWrapper_115_clock),
    .reset(RetimeWrapper_115_reset),
    .io_flow(RetimeWrapper_115_io_flow),
    .io_in(RetimeWrapper_115_io_in),
    .io_out(RetimeWrapper_115_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_116 ( // @[package.scala 93:22:@14725.4]
    .clock(RetimeWrapper_116_clock),
    .reset(RetimeWrapper_116_reset),
    .io_flow(RetimeWrapper_116_io_flow),
    .io_in(RetimeWrapper_116_io_in),
    .io_out(RetimeWrapper_116_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_117 ( // @[package.scala 93:22:@14733.4]
    .clock(RetimeWrapper_117_clock),
    .reset(RetimeWrapper_117_reset),
    .io_flow(RetimeWrapper_117_io_flow),
    .io_in(RetimeWrapper_117_io_in),
    .io_out(RetimeWrapper_117_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_118 ( // @[package.scala 93:22:@14741.4]
    .clock(RetimeWrapper_118_clock),
    .reset(RetimeWrapper_118_reset),
    .io_flow(RetimeWrapper_118_io_flow),
    .io_in(RetimeWrapper_118_io_in),
    .io_out(RetimeWrapper_118_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_119 ( // @[package.scala 93:22:@14749.4]
    .clock(RetimeWrapper_119_clock),
    .reset(RetimeWrapper_119_reset),
    .io_flow(RetimeWrapper_119_io_flow),
    .io_in(RetimeWrapper_119_io_in),
    .io_out(RetimeWrapper_119_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_120 ( // @[package.scala 93:22:@14757.4]
    .clock(RetimeWrapper_120_clock),
    .reset(RetimeWrapper_120_reset),
    .io_flow(RetimeWrapper_120_io_flow),
    .io_in(RetimeWrapper_120_io_in),
    .io_out(RetimeWrapper_120_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_121 ( // @[package.scala 93:22:@14765.4]
    .clock(RetimeWrapper_121_clock),
    .reset(RetimeWrapper_121_reset),
    .io_flow(RetimeWrapper_121_io_flow),
    .io_in(RetimeWrapper_121_io_in),
    .io_out(RetimeWrapper_121_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_122 ( // @[package.scala 93:22:@14773.4]
    .clock(RetimeWrapper_122_clock),
    .reset(RetimeWrapper_122_reset),
    .io_flow(RetimeWrapper_122_io_flow),
    .io_in(RetimeWrapper_122_io_in),
    .io_out(RetimeWrapper_122_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_123 ( // @[package.scala 93:22:@14781.4]
    .clock(RetimeWrapper_123_clock),
    .reset(RetimeWrapper_123_reset),
    .io_flow(RetimeWrapper_123_io_flow),
    .io_in(RetimeWrapper_123_io_in),
    .io_out(RetimeWrapper_123_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_124 ( // @[package.scala 93:22:@14789.4]
    .clock(RetimeWrapper_124_clock),
    .reset(RetimeWrapper_124_reset),
    .io_flow(RetimeWrapper_124_io_flow),
    .io_in(RetimeWrapper_124_io_in),
    .io_out(RetimeWrapper_124_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_125 ( // @[package.scala 93:22:@14797.4]
    .clock(RetimeWrapper_125_clock),
    .reset(RetimeWrapper_125_reset),
    .io_flow(RetimeWrapper_125_io_flow),
    .io_in(RetimeWrapper_125_io_in),
    .io_out(RetimeWrapper_125_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_126 ( // @[package.scala 93:22:@14805.4]
    .clock(RetimeWrapper_126_clock),
    .reset(RetimeWrapper_126_reset),
    .io_flow(RetimeWrapper_126_io_flow),
    .io_in(RetimeWrapper_126_io_in),
    .io_out(RetimeWrapper_126_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_127 ( // @[package.scala 93:22:@14813.4]
    .clock(RetimeWrapper_127_clock),
    .reset(RetimeWrapper_127_reset),
    .io_flow(RetimeWrapper_127_io_flow),
    .io_in(RetimeWrapper_127_io_in),
    .io_out(RetimeWrapper_127_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_128 ( // @[package.scala 93:22:@14885.4]
    .clock(RetimeWrapper_128_clock),
    .reset(RetimeWrapper_128_reset),
    .io_flow(RetimeWrapper_128_io_flow),
    .io_in(RetimeWrapper_128_io_in),
    .io_out(RetimeWrapper_128_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_129 ( // @[package.scala 93:22:@14893.4]
    .clock(RetimeWrapper_129_clock),
    .reset(RetimeWrapper_129_reset),
    .io_flow(RetimeWrapper_129_io_flow),
    .io_in(RetimeWrapper_129_io_in),
    .io_out(RetimeWrapper_129_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_130 ( // @[package.scala 93:22:@14901.4]
    .clock(RetimeWrapper_130_clock),
    .reset(RetimeWrapper_130_reset),
    .io_flow(RetimeWrapper_130_io_flow),
    .io_in(RetimeWrapper_130_io_in),
    .io_out(RetimeWrapper_130_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_131 ( // @[package.scala 93:22:@14909.4]
    .clock(RetimeWrapper_131_clock),
    .reset(RetimeWrapper_131_reset),
    .io_flow(RetimeWrapper_131_io_flow),
    .io_in(RetimeWrapper_131_io_in),
    .io_out(RetimeWrapper_131_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_132 ( // @[package.scala 93:22:@14917.4]
    .clock(RetimeWrapper_132_clock),
    .reset(RetimeWrapper_132_reset),
    .io_flow(RetimeWrapper_132_io_flow),
    .io_in(RetimeWrapper_132_io_in),
    .io_out(RetimeWrapper_132_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_133 ( // @[package.scala 93:22:@14925.4]
    .clock(RetimeWrapper_133_clock),
    .reset(RetimeWrapper_133_reset),
    .io_flow(RetimeWrapper_133_io_flow),
    .io_in(RetimeWrapper_133_io_in),
    .io_out(RetimeWrapper_133_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_134 ( // @[package.scala 93:22:@14933.4]
    .clock(RetimeWrapper_134_clock),
    .reset(RetimeWrapper_134_reset),
    .io_flow(RetimeWrapper_134_io_flow),
    .io_in(RetimeWrapper_134_io_in),
    .io_out(RetimeWrapper_134_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_135 ( // @[package.scala 93:22:@14941.4]
    .clock(RetimeWrapper_135_clock),
    .reset(RetimeWrapper_135_reset),
    .io_flow(RetimeWrapper_135_io_flow),
    .io_in(RetimeWrapper_135_io_in),
    .io_out(RetimeWrapper_135_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_136 ( // @[package.scala 93:22:@14949.4]
    .clock(RetimeWrapper_136_clock),
    .reset(RetimeWrapper_136_reset),
    .io_flow(RetimeWrapper_136_io_flow),
    .io_in(RetimeWrapper_136_io_in),
    .io_out(RetimeWrapper_136_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_137 ( // @[package.scala 93:22:@14957.4]
    .clock(RetimeWrapper_137_clock),
    .reset(RetimeWrapper_137_reset),
    .io_flow(RetimeWrapper_137_io_flow),
    .io_in(RetimeWrapper_137_io_in),
    .io_out(RetimeWrapper_137_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_138 ( // @[package.scala 93:22:@14965.4]
    .clock(RetimeWrapper_138_clock),
    .reset(RetimeWrapper_138_reset),
    .io_flow(RetimeWrapper_138_io_flow),
    .io_in(RetimeWrapper_138_io_in),
    .io_out(RetimeWrapper_138_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_139 ( // @[package.scala 93:22:@14973.4]
    .clock(RetimeWrapper_139_clock),
    .reset(RetimeWrapper_139_reset),
    .io_flow(RetimeWrapper_139_io_flow),
    .io_in(RetimeWrapper_139_io_in),
    .io_out(RetimeWrapper_139_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_140 ( // @[package.scala 93:22:@14981.4]
    .clock(RetimeWrapper_140_clock),
    .reset(RetimeWrapper_140_reset),
    .io_flow(RetimeWrapper_140_io_flow),
    .io_in(RetimeWrapper_140_io_in),
    .io_out(RetimeWrapper_140_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_141 ( // @[package.scala 93:22:@14989.4]
    .clock(RetimeWrapper_141_clock),
    .reset(RetimeWrapper_141_reset),
    .io_flow(RetimeWrapper_141_io_flow),
    .io_in(RetimeWrapper_141_io_in),
    .io_out(RetimeWrapper_141_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_142 ( // @[package.scala 93:22:@14997.4]
    .clock(RetimeWrapper_142_clock),
    .reset(RetimeWrapper_142_reset),
    .io_flow(RetimeWrapper_142_io_flow),
    .io_in(RetimeWrapper_142_io_in),
    .io_out(RetimeWrapper_142_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_143 ( // @[package.scala 93:22:@15005.4]
    .clock(RetimeWrapper_143_clock),
    .reset(RetimeWrapper_143_reset),
    .io_flow(RetimeWrapper_143_io_flow),
    .io_in(RetimeWrapper_143_io_in),
    .io_out(RetimeWrapper_143_io_out)
  );
  assign _T_316 = io_wPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@11684.4]
  assign _T_318 = io_wPort_0_banks_1 == 3'h0; // @[MemPrimitives.scala 82:210:@11685.4]
  assign _T_319 = _T_316 & _T_318; // @[MemPrimitives.scala 82:228:@11686.4]
  assign _T_320 = io_wPort_0_en_0 & _T_319; // @[MemPrimitives.scala 83:102:@11687.4]
  assign _T_322 = {_T_320,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@11689.4]
  assign _T_329 = io_wPort_0_banks_1 == 3'h1; // @[MemPrimitives.scala 82:210:@11697.4]
  assign _T_330 = _T_316 & _T_329; // @[MemPrimitives.scala 82:228:@11698.4]
  assign _T_331 = io_wPort_0_en_0 & _T_330; // @[MemPrimitives.scala 83:102:@11699.4]
  assign _T_333 = {_T_331,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@11701.4]
  assign _T_340 = io_wPort_0_banks_1 == 3'h2; // @[MemPrimitives.scala 82:210:@11709.4]
  assign _T_341 = _T_316 & _T_340; // @[MemPrimitives.scala 82:228:@11710.4]
  assign _T_342 = io_wPort_0_en_0 & _T_341; // @[MemPrimitives.scala 83:102:@11711.4]
  assign _T_344 = {_T_342,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@11713.4]
  assign _T_351 = io_wPort_0_banks_1 == 3'h3; // @[MemPrimitives.scala 82:210:@11721.4]
  assign _T_352 = _T_316 & _T_351; // @[MemPrimitives.scala 82:228:@11722.4]
  assign _T_353 = io_wPort_0_en_0 & _T_352; // @[MemPrimitives.scala 83:102:@11723.4]
  assign _T_355 = {_T_353,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@11725.4]
  assign _T_360 = io_wPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@11732.4]
  assign _T_363 = _T_360 & _T_318; // @[MemPrimitives.scala 82:228:@11734.4]
  assign _T_364 = io_wPort_0_en_0 & _T_363; // @[MemPrimitives.scala 83:102:@11735.4]
  assign _T_366 = {_T_364,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@11737.4]
  assign _T_374 = _T_360 & _T_329; // @[MemPrimitives.scala 82:228:@11746.4]
  assign _T_375 = io_wPort_0_en_0 & _T_374; // @[MemPrimitives.scala 83:102:@11747.4]
  assign _T_377 = {_T_375,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@11749.4]
  assign _T_385 = _T_360 & _T_340; // @[MemPrimitives.scala 82:228:@11758.4]
  assign _T_386 = io_wPort_0_en_0 & _T_385; // @[MemPrimitives.scala 83:102:@11759.4]
  assign _T_388 = {_T_386,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@11761.4]
  assign _T_396 = _T_360 & _T_351; // @[MemPrimitives.scala 82:228:@11770.4]
  assign _T_397 = io_wPort_0_en_0 & _T_396; // @[MemPrimitives.scala 83:102:@11771.4]
  assign _T_399 = {_T_397,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@11773.4]
  assign _T_404 = io_wPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@11780.4]
  assign _T_407 = _T_404 & _T_318; // @[MemPrimitives.scala 82:228:@11782.4]
  assign _T_408 = io_wPort_0_en_0 & _T_407; // @[MemPrimitives.scala 83:102:@11783.4]
  assign _T_410 = {_T_408,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@11785.4]
  assign _T_418 = _T_404 & _T_329; // @[MemPrimitives.scala 82:228:@11794.4]
  assign _T_419 = io_wPort_0_en_0 & _T_418; // @[MemPrimitives.scala 83:102:@11795.4]
  assign _T_421 = {_T_419,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@11797.4]
  assign _T_429 = _T_404 & _T_340; // @[MemPrimitives.scala 82:228:@11806.4]
  assign _T_430 = io_wPort_0_en_0 & _T_429; // @[MemPrimitives.scala 83:102:@11807.4]
  assign _T_432 = {_T_430,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@11809.4]
  assign _T_440 = _T_404 & _T_351; // @[MemPrimitives.scala 82:228:@11818.4]
  assign _T_441 = io_wPort_0_en_0 & _T_440; // @[MemPrimitives.scala 83:102:@11819.4]
  assign _T_443 = {_T_441,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@11821.4]
  assign _T_448 = io_wPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@11828.4]
  assign _T_451 = _T_448 & _T_318; // @[MemPrimitives.scala 82:228:@11830.4]
  assign _T_452 = io_wPort_0_en_0 & _T_451; // @[MemPrimitives.scala 83:102:@11831.4]
  assign _T_454 = {_T_452,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@11833.4]
  assign _T_462 = _T_448 & _T_329; // @[MemPrimitives.scala 82:228:@11842.4]
  assign _T_463 = io_wPort_0_en_0 & _T_462; // @[MemPrimitives.scala 83:102:@11843.4]
  assign _T_465 = {_T_463,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@11845.4]
  assign _T_473 = _T_448 & _T_340; // @[MemPrimitives.scala 82:228:@11854.4]
  assign _T_474 = io_wPort_0_en_0 & _T_473; // @[MemPrimitives.scala 83:102:@11855.4]
  assign _T_476 = {_T_474,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@11857.4]
  assign _T_484 = _T_448 & _T_351; // @[MemPrimitives.scala 82:228:@11866.4]
  assign _T_485 = io_wPort_0_en_0 & _T_484; // @[MemPrimitives.scala 83:102:@11867.4]
  assign _T_487 = {_T_485,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@11869.4]
  assign _T_492 = io_rPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@11876.4]
  assign _T_494 = io_rPort_0_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@11877.4]
  assign _T_495 = _T_492 & _T_494; // @[MemPrimitives.scala 110:228:@11878.4]
  assign _T_498 = io_rPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@11880.4]
  assign _T_500 = io_rPort_1_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@11881.4]
  assign _T_501 = _T_498 & _T_500; // @[MemPrimitives.scala 110:228:@11882.4]
  assign _T_504 = io_rPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@11884.4]
  assign _T_506 = io_rPort_2_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@11885.4]
  assign _T_507 = _T_504 & _T_506; // @[MemPrimitives.scala 110:228:@11886.4]
  assign _T_510 = io_rPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@11888.4]
  assign _T_512 = io_rPort_3_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@11889.4]
  assign _T_513 = _T_510 & _T_512; // @[MemPrimitives.scala 110:228:@11890.4]
  assign _T_516 = io_rPort_4_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@11892.4]
  assign _T_518 = io_rPort_4_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@11893.4]
  assign _T_519 = _T_516 & _T_518; // @[MemPrimitives.scala 110:228:@11894.4]
  assign _T_522 = io_rPort_5_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@11896.4]
  assign _T_524 = io_rPort_5_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@11897.4]
  assign _T_525 = _T_522 & _T_524; // @[MemPrimitives.scala 110:228:@11898.4]
  assign _T_528 = io_rPort_6_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@11900.4]
  assign _T_530 = io_rPort_6_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@11901.4]
  assign _T_531 = _T_528 & _T_530; // @[MemPrimitives.scala 110:228:@11902.4]
  assign _T_534 = io_rPort_7_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@11904.4]
  assign _T_536 = io_rPort_7_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@11905.4]
  assign _T_537 = _T_534 & _T_536; // @[MemPrimitives.scala 110:228:@11906.4]
  assign _T_540 = io_rPort_8_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@11908.4]
  assign _T_542 = io_rPort_8_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@11909.4]
  assign _T_543 = _T_540 & _T_542; // @[MemPrimitives.scala 110:228:@11910.4]
  assign _T_545 = StickySelects_io_outs_0; // @[MemPrimitives.scala 123:41:@11924.4]
  assign _T_546 = StickySelects_io_outs_1; // @[MemPrimitives.scala 123:41:@11925.4]
  assign _T_547 = StickySelects_io_outs_2; // @[MemPrimitives.scala 123:41:@11926.4]
  assign _T_548 = StickySelects_io_outs_3; // @[MemPrimitives.scala 123:41:@11927.4]
  assign _T_549 = StickySelects_io_outs_4; // @[MemPrimitives.scala 123:41:@11928.4]
  assign _T_550 = StickySelects_io_outs_5; // @[MemPrimitives.scala 123:41:@11929.4]
  assign _T_551 = StickySelects_io_outs_6; // @[MemPrimitives.scala 123:41:@11930.4]
  assign _T_552 = StickySelects_io_outs_7; // @[MemPrimitives.scala 123:41:@11931.4]
  assign _T_553 = StickySelects_io_outs_8; // @[MemPrimitives.scala 123:41:@11932.4]
  assign _T_555 = {_T_545,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@11934.4]
  assign _T_557 = {_T_546,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@11936.4]
  assign _T_559 = {_T_547,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@11938.4]
  assign _T_561 = {_T_548,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@11940.4]
  assign _T_563 = {_T_549,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@11942.4]
  assign _T_565 = {_T_550,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@11944.4]
  assign _T_567 = {_T_551,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@11946.4]
  assign _T_569 = {_T_552,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@11948.4]
  assign _T_571 = {_T_553,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@11950.4]
  assign _T_572 = _T_552 ? _T_569 : _T_571; // @[Mux.scala 31:69:@11951.4]
  assign _T_573 = _T_551 ? _T_567 : _T_572; // @[Mux.scala 31:69:@11952.4]
  assign _T_574 = _T_550 ? _T_565 : _T_573; // @[Mux.scala 31:69:@11953.4]
  assign _T_575 = _T_549 ? _T_563 : _T_574; // @[Mux.scala 31:69:@11954.4]
  assign _T_576 = _T_548 ? _T_561 : _T_575; // @[Mux.scala 31:69:@11955.4]
  assign _T_577 = _T_547 ? _T_559 : _T_576; // @[Mux.scala 31:69:@11956.4]
  assign _T_578 = _T_546 ? _T_557 : _T_577; // @[Mux.scala 31:69:@11957.4]
  assign _T_579 = _T_545 ? _T_555 : _T_578; // @[Mux.scala 31:69:@11958.4]
  assign _T_586 = io_rPort_0_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@11966.4]
  assign _T_587 = _T_492 & _T_586; // @[MemPrimitives.scala 110:228:@11967.4]
  assign _T_592 = io_rPort_1_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@11970.4]
  assign _T_593 = _T_498 & _T_592; // @[MemPrimitives.scala 110:228:@11971.4]
  assign _T_598 = io_rPort_2_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@11974.4]
  assign _T_599 = _T_504 & _T_598; // @[MemPrimitives.scala 110:228:@11975.4]
  assign _T_604 = io_rPort_3_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@11978.4]
  assign _T_605 = _T_510 & _T_604; // @[MemPrimitives.scala 110:228:@11979.4]
  assign _T_610 = io_rPort_4_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@11982.4]
  assign _T_611 = _T_516 & _T_610; // @[MemPrimitives.scala 110:228:@11983.4]
  assign _T_616 = io_rPort_5_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@11986.4]
  assign _T_617 = _T_522 & _T_616; // @[MemPrimitives.scala 110:228:@11987.4]
  assign _T_622 = io_rPort_6_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@11990.4]
  assign _T_623 = _T_528 & _T_622; // @[MemPrimitives.scala 110:228:@11991.4]
  assign _T_628 = io_rPort_7_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@11994.4]
  assign _T_629 = _T_534 & _T_628; // @[MemPrimitives.scala 110:228:@11995.4]
  assign _T_634 = io_rPort_8_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@11998.4]
  assign _T_635 = _T_540 & _T_634; // @[MemPrimitives.scala 110:228:@11999.4]
  assign _T_637 = StickySelects_1_io_outs_0; // @[MemPrimitives.scala 123:41:@12013.4]
  assign _T_638 = StickySelects_1_io_outs_1; // @[MemPrimitives.scala 123:41:@12014.4]
  assign _T_639 = StickySelects_1_io_outs_2; // @[MemPrimitives.scala 123:41:@12015.4]
  assign _T_640 = StickySelects_1_io_outs_3; // @[MemPrimitives.scala 123:41:@12016.4]
  assign _T_641 = StickySelects_1_io_outs_4; // @[MemPrimitives.scala 123:41:@12017.4]
  assign _T_642 = StickySelects_1_io_outs_5; // @[MemPrimitives.scala 123:41:@12018.4]
  assign _T_643 = StickySelects_1_io_outs_6; // @[MemPrimitives.scala 123:41:@12019.4]
  assign _T_644 = StickySelects_1_io_outs_7; // @[MemPrimitives.scala 123:41:@12020.4]
  assign _T_645 = StickySelects_1_io_outs_8; // @[MemPrimitives.scala 123:41:@12021.4]
  assign _T_647 = {_T_637,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@12023.4]
  assign _T_649 = {_T_638,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@12025.4]
  assign _T_651 = {_T_639,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@12027.4]
  assign _T_653 = {_T_640,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@12029.4]
  assign _T_655 = {_T_641,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@12031.4]
  assign _T_657 = {_T_642,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@12033.4]
  assign _T_659 = {_T_643,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@12035.4]
  assign _T_661 = {_T_644,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@12037.4]
  assign _T_663 = {_T_645,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@12039.4]
  assign _T_664 = _T_644 ? _T_661 : _T_663; // @[Mux.scala 31:69:@12040.4]
  assign _T_665 = _T_643 ? _T_659 : _T_664; // @[Mux.scala 31:69:@12041.4]
  assign _T_666 = _T_642 ? _T_657 : _T_665; // @[Mux.scala 31:69:@12042.4]
  assign _T_667 = _T_641 ? _T_655 : _T_666; // @[Mux.scala 31:69:@12043.4]
  assign _T_668 = _T_640 ? _T_653 : _T_667; // @[Mux.scala 31:69:@12044.4]
  assign _T_669 = _T_639 ? _T_651 : _T_668; // @[Mux.scala 31:69:@12045.4]
  assign _T_670 = _T_638 ? _T_649 : _T_669; // @[Mux.scala 31:69:@12046.4]
  assign _T_671 = _T_637 ? _T_647 : _T_670; // @[Mux.scala 31:69:@12047.4]
  assign _T_678 = io_rPort_0_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@12055.4]
  assign _T_679 = _T_492 & _T_678; // @[MemPrimitives.scala 110:228:@12056.4]
  assign _T_684 = io_rPort_1_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@12059.4]
  assign _T_685 = _T_498 & _T_684; // @[MemPrimitives.scala 110:228:@12060.4]
  assign _T_690 = io_rPort_2_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@12063.4]
  assign _T_691 = _T_504 & _T_690; // @[MemPrimitives.scala 110:228:@12064.4]
  assign _T_696 = io_rPort_3_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@12067.4]
  assign _T_697 = _T_510 & _T_696; // @[MemPrimitives.scala 110:228:@12068.4]
  assign _T_702 = io_rPort_4_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@12071.4]
  assign _T_703 = _T_516 & _T_702; // @[MemPrimitives.scala 110:228:@12072.4]
  assign _T_708 = io_rPort_5_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@12075.4]
  assign _T_709 = _T_522 & _T_708; // @[MemPrimitives.scala 110:228:@12076.4]
  assign _T_714 = io_rPort_6_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@12079.4]
  assign _T_715 = _T_528 & _T_714; // @[MemPrimitives.scala 110:228:@12080.4]
  assign _T_720 = io_rPort_7_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@12083.4]
  assign _T_721 = _T_534 & _T_720; // @[MemPrimitives.scala 110:228:@12084.4]
  assign _T_726 = io_rPort_8_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@12087.4]
  assign _T_727 = _T_540 & _T_726; // @[MemPrimitives.scala 110:228:@12088.4]
  assign _T_729 = StickySelects_2_io_outs_0; // @[MemPrimitives.scala 123:41:@12102.4]
  assign _T_730 = StickySelects_2_io_outs_1; // @[MemPrimitives.scala 123:41:@12103.4]
  assign _T_731 = StickySelects_2_io_outs_2; // @[MemPrimitives.scala 123:41:@12104.4]
  assign _T_732 = StickySelects_2_io_outs_3; // @[MemPrimitives.scala 123:41:@12105.4]
  assign _T_733 = StickySelects_2_io_outs_4; // @[MemPrimitives.scala 123:41:@12106.4]
  assign _T_734 = StickySelects_2_io_outs_5; // @[MemPrimitives.scala 123:41:@12107.4]
  assign _T_735 = StickySelects_2_io_outs_6; // @[MemPrimitives.scala 123:41:@12108.4]
  assign _T_736 = StickySelects_2_io_outs_7; // @[MemPrimitives.scala 123:41:@12109.4]
  assign _T_737 = StickySelects_2_io_outs_8; // @[MemPrimitives.scala 123:41:@12110.4]
  assign _T_739 = {_T_729,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@12112.4]
  assign _T_741 = {_T_730,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@12114.4]
  assign _T_743 = {_T_731,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@12116.4]
  assign _T_745 = {_T_732,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@12118.4]
  assign _T_747 = {_T_733,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@12120.4]
  assign _T_749 = {_T_734,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@12122.4]
  assign _T_751 = {_T_735,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@12124.4]
  assign _T_753 = {_T_736,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@12126.4]
  assign _T_755 = {_T_737,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@12128.4]
  assign _T_756 = _T_736 ? _T_753 : _T_755; // @[Mux.scala 31:69:@12129.4]
  assign _T_757 = _T_735 ? _T_751 : _T_756; // @[Mux.scala 31:69:@12130.4]
  assign _T_758 = _T_734 ? _T_749 : _T_757; // @[Mux.scala 31:69:@12131.4]
  assign _T_759 = _T_733 ? _T_747 : _T_758; // @[Mux.scala 31:69:@12132.4]
  assign _T_760 = _T_732 ? _T_745 : _T_759; // @[Mux.scala 31:69:@12133.4]
  assign _T_761 = _T_731 ? _T_743 : _T_760; // @[Mux.scala 31:69:@12134.4]
  assign _T_762 = _T_730 ? _T_741 : _T_761; // @[Mux.scala 31:69:@12135.4]
  assign _T_763 = _T_729 ? _T_739 : _T_762; // @[Mux.scala 31:69:@12136.4]
  assign _T_770 = io_rPort_0_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@12144.4]
  assign _T_771 = _T_492 & _T_770; // @[MemPrimitives.scala 110:228:@12145.4]
  assign _T_776 = io_rPort_1_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@12148.4]
  assign _T_777 = _T_498 & _T_776; // @[MemPrimitives.scala 110:228:@12149.4]
  assign _T_782 = io_rPort_2_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@12152.4]
  assign _T_783 = _T_504 & _T_782; // @[MemPrimitives.scala 110:228:@12153.4]
  assign _T_788 = io_rPort_3_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@12156.4]
  assign _T_789 = _T_510 & _T_788; // @[MemPrimitives.scala 110:228:@12157.4]
  assign _T_794 = io_rPort_4_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@12160.4]
  assign _T_795 = _T_516 & _T_794; // @[MemPrimitives.scala 110:228:@12161.4]
  assign _T_800 = io_rPort_5_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@12164.4]
  assign _T_801 = _T_522 & _T_800; // @[MemPrimitives.scala 110:228:@12165.4]
  assign _T_806 = io_rPort_6_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@12168.4]
  assign _T_807 = _T_528 & _T_806; // @[MemPrimitives.scala 110:228:@12169.4]
  assign _T_812 = io_rPort_7_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@12172.4]
  assign _T_813 = _T_534 & _T_812; // @[MemPrimitives.scala 110:228:@12173.4]
  assign _T_818 = io_rPort_8_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@12176.4]
  assign _T_819 = _T_540 & _T_818; // @[MemPrimitives.scala 110:228:@12177.4]
  assign _T_821 = StickySelects_3_io_outs_0; // @[MemPrimitives.scala 123:41:@12191.4]
  assign _T_822 = StickySelects_3_io_outs_1; // @[MemPrimitives.scala 123:41:@12192.4]
  assign _T_823 = StickySelects_3_io_outs_2; // @[MemPrimitives.scala 123:41:@12193.4]
  assign _T_824 = StickySelects_3_io_outs_3; // @[MemPrimitives.scala 123:41:@12194.4]
  assign _T_825 = StickySelects_3_io_outs_4; // @[MemPrimitives.scala 123:41:@12195.4]
  assign _T_826 = StickySelects_3_io_outs_5; // @[MemPrimitives.scala 123:41:@12196.4]
  assign _T_827 = StickySelects_3_io_outs_6; // @[MemPrimitives.scala 123:41:@12197.4]
  assign _T_828 = StickySelects_3_io_outs_7; // @[MemPrimitives.scala 123:41:@12198.4]
  assign _T_829 = StickySelects_3_io_outs_8; // @[MemPrimitives.scala 123:41:@12199.4]
  assign _T_831 = {_T_821,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@12201.4]
  assign _T_833 = {_T_822,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@12203.4]
  assign _T_835 = {_T_823,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@12205.4]
  assign _T_837 = {_T_824,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@12207.4]
  assign _T_839 = {_T_825,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@12209.4]
  assign _T_841 = {_T_826,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@12211.4]
  assign _T_843 = {_T_827,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@12213.4]
  assign _T_845 = {_T_828,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@12215.4]
  assign _T_847 = {_T_829,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@12217.4]
  assign _T_848 = _T_828 ? _T_845 : _T_847; // @[Mux.scala 31:69:@12218.4]
  assign _T_849 = _T_827 ? _T_843 : _T_848; // @[Mux.scala 31:69:@12219.4]
  assign _T_850 = _T_826 ? _T_841 : _T_849; // @[Mux.scala 31:69:@12220.4]
  assign _T_851 = _T_825 ? _T_839 : _T_850; // @[Mux.scala 31:69:@12221.4]
  assign _T_852 = _T_824 ? _T_837 : _T_851; // @[Mux.scala 31:69:@12222.4]
  assign _T_853 = _T_823 ? _T_835 : _T_852; // @[Mux.scala 31:69:@12223.4]
  assign _T_854 = _T_822 ? _T_833 : _T_853; // @[Mux.scala 31:69:@12224.4]
  assign _T_855 = _T_821 ? _T_831 : _T_854; // @[Mux.scala 31:69:@12225.4]
  assign _T_860 = io_rPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@12232.4]
  assign _T_863 = _T_860 & _T_494; // @[MemPrimitives.scala 110:228:@12234.4]
  assign _T_866 = io_rPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@12236.4]
  assign _T_869 = _T_866 & _T_500; // @[MemPrimitives.scala 110:228:@12238.4]
  assign _T_872 = io_rPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@12240.4]
  assign _T_875 = _T_872 & _T_506; // @[MemPrimitives.scala 110:228:@12242.4]
  assign _T_878 = io_rPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@12244.4]
  assign _T_881 = _T_878 & _T_512; // @[MemPrimitives.scala 110:228:@12246.4]
  assign _T_884 = io_rPort_4_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@12248.4]
  assign _T_887 = _T_884 & _T_518; // @[MemPrimitives.scala 110:228:@12250.4]
  assign _T_890 = io_rPort_5_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@12252.4]
  assign _T_893 = _T_890 & _T_524; // @[MemPrimitives.scala 110:228:@12254.4]
  assign _T_896 = io_rPort_6_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@12256.4]
  assign _T_899 = _T_896 & _T_530; // @[MemPrimitives.scala 110:228:@12258.4]
  assign _T_902 = io_rPort_7_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@12260.4]
  assign _T_905 = _T_902 & _T_536; // @[MemPrimitives.scala 110:228:@12262.4]
  assign _T_908 = io_rPort_8_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@12264.4]
  assign _T_911 = _T_908 & _T_542; // @[MemPrimitives.scala 110:228:@12266.4]
  assign _T_913 = StickySelects_4_io_outs_0; // @[MemPrimitives.scala 123:41:@12280.4]
  assign _T_914 = StickySelects_4_io_outs_1; // @[MemPrimitives.scala 123:41:@12281.4]
  assign _T_915 = StickySelects_4_io_outs_2; // @[MemPrimitives.scala 123:41:@12282.4]
  assign _T_916 = StickySelects_4_io_outs_3; // @[MemPrimitives.scala 123:41:@12283.4]
  assign _T_917 = StickySelects_4_io_outs_4; // @[MemPrimitives.scala 123:41:@12284.4]
  assign _T_918 = StickySelects_4_io_outs_5; // @[MemPrimitives.scala 123:41:@12285.4]
  assign _T_919 = StickySelects_4_io_outs_6; // @[MemPrimitives.scala 123:41:@12286.4]
  assign _T_920 = StickySelects_4_io_outs_7; // @[MemPrimitives.scala 123:41:@12287.4]
  assign _T_921 = StickySelects_4_io_outs_8; // @[MemPrimitives.scala 123:41:@12288.4]
  assign _T_923 = {_T_913,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@12290.4]
  assign _T_925 = {_T_914,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@12292.4]
  assign _T_927 = {_T_915,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@12294.4]
  assign _T_929 = {_T_916,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@12296.4]
  assign _T_931 = {_T_917,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@12298.4]
  assign _T_933 = {_T_918,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@12300.4]
  assign _T_935 = {_T_919,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@12302.4]
  assign _T_937 = {_T_920,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@12304.4]
  assign _T_939 = {_T_921,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@12306.4]
  assign _T_940 = _T_920 ? _T_937 : _T_939; // @[Mux.scala 31:69:@12307.4]
  assign _T_941 = _T_919 ? _T_935 : _T_940; // @[Mux.scala 31:69:@12308.4]
  assign _T_942 = _T_918 ? _T_933 : _T_941; // @[Mux.scala 31:69:@12309.4]
  assign _T_943 = _T_917 ? _T_931 : _T_942; // @[Mux.scala 31:69:@12310.4]
  assign _T_944 = _T_916 ? _T_929 : _T_943; // @[Mux.scala 31:69:@12311.4]
  assign _T_945 = _T_915 ? _T_927 : _T_944; // @[Mux.scala 31:69:@12312.4]
  assign _T_946 = _T_914 ? _T_925 : _T_945; // @[Mux.scala 31:69:@12313.4]
  assign _T_947 = _T_913 ? _T_923 : _T_946; // @[Mux.scala 31:69:@12314.4]
  assign _T_955 = _T_860 & _T_586; // @[MemPrimitives.scala 110:228:@12323.4]
  assign _T_961 = _T_866 & _T_592; // @[MemPrimitives.scala 110:228:@12327.4]
  assign _T_967 = _T_872 & _T_598; // @[MemPrimitives.scala 110:228:@12331.4]
  assign _T_973 = _T_878 & _T_604; // @[MemPrimitives.scala 110:228:@12335.4]
  assign _T_979 = _T_884 & _T_610; // @[MemPrimitives.scala 110:228:@12339.4]
  assign _T_985 = _T_890 & _T_616; // @[MemPrimitives.scala 110:228:@12343.4]
  assign _T_991 = _T_896 & _T_622; // @[MemPrimitives.scala 110:228:@12347.4]
  assign _T_997 = _T_902 & _T_628; // @[MemPrimitives.scala 110:228:@12351.4]
  assign _T_1003 = _T_908 & _T_634; // @[MemPrimitives.scala 110:228:@12355.4]
  assign _T_1005 = StickySelects_5_io_outs_0; // @[MemPrimitives.scala 123:41:@12369.4]
  assign _T_1006 = StickySelects_5_io_outs_1; // @[MemPrimitives.scala 123:41:@12370.4]
  assign _T_1007 = StickySelects_5_io_outs_2; // @[MemPrimitives.scala 123:41:@12371.4]
  assign _T_1008 = StickySelects_5_io_outs_3; // @[MemPrimitives.scala 123:41:@12372.4]
  assign _T_1009 = StickySelects_5_io_outs_4; // @[MemPrimitives.scala 123:41:@12373.4]
  assign _T_1010 = StickySelects_5_io_outs_5; // @[MemPrimitives.scala 123:41:@12374.4]
  assign _T_1011 = StickySelects_5_io_outs_6; // @[MemPrimitives.scala 123:41:@12375.4]
  assign _T_1012 = StickySelects_5_io_outs_7; // @[MemPrimitives.scala 123:41:@12376.4]
  assign _T_1013 = StickySelects_5_io_outs_8; // @[MemPrimitives.scala 123:41:@12377.4]
  assign _T_1015 = {_T_1005,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@12379.4]
  assign _T_1017 = {_T_1006,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@12381.4]
  assign _T_1019 = {_T_1007,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@12383.4]
  assign _T_1021 = {_T_1008,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@12385.4]
  assign _T_1023 = {_T_1009,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@12387.4]
  assign _T_1025 = {_T_1010,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@12389.4]
  assign _T_1027 = {_T_1011,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@12391.4]
  assign _T_1029 = {_T_1012,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@12393.4]
  assign _T_1031 = {_T_1013,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@12395.4]
  assign _T_1032 = _T_1012 ? _T_1029 : _T_1031; // @[Mux.scala 31:69:@12396.4]
  assign _T_1033 = _T_1011 ? _T_1027 : _T_1032; // @[Mux.scala 31:69:@12397.4]
  assign _T_1034 = _T_1010 ? _T_1025 : _T_1033; // @[Mux.scala 31:69:@12398.4]
  assign _T_1035 = _T_1009 ? _T_1023 : _T_1034; // @[Mux.scala 31:69:@12399.4]
  assign _T_1036 = _T_1008 ? _T_1021 : _T_1035; // @[Mux.scala 31:69:@12400.4]
  assign _T_1037 = _T_1007 ? _T_1019 : _T_1036; // @[Mux.scala 31:69:@12401.4]
  assign _T_1038 = _T_1006 ? _T_1017 : _T_1037; // @[Mux.scala 31:69:@12402.4]
  assign _T_1039 = _T_1005 ? _T_1015 : _T_1038; // @[Mux.scala 31:69:@12403.4]
  assign _T_1047 = _T_860 & _T_678; // @[MemPrimitives.scala 110:228:@12412.4]
  assign _T_1053 = _T_866 & _T_684; // @[MemPrimitives.scala 110:228:@12416.4]
  assign _T_1059 = _T_872 & _T_690; // @[MemPrimitives.scala 110:228:@12420.4]
  assign _T_1065 = _T_878 & _T_696; // @[MemPrimitives.scala 110:228:@12424.4]
  assign _T_1071 = _T_884 & _T_702; // @[MemPrimitives.scala 110:228:@12428.4]
  assign _T_1077 = _T_890 & _T_708; // @[MemPrimitives.scala 110:228:@12432.4]
  assign _T_1083 = _T_896 & _T_714; // @[MemPrimitives.scala 110:228:@12436.4]
  assign _T_1089 = _T_902 & _T_720; // @[MemPrimitives.scala 110:228:@12440.4]
  assign _T_1095 = _T_908 & _T_726; // @[MemPrimitives.scala 110:228:@12444.4]
  assign _T_1097 = StickySelects_6_io_outs_0; // @[MemPrimitives.scala 123:41:@12458.4]
  assign _T_1098 = StickySelects_6_io_outs_1; // @[MemPrimitives.scala 123:41:@12459.4]
  assign _T_1099 = StickySelects_6_io_outs_2; // @[MemPrimitives.scala 123:41:@12460.4]
  assign _T_1100 = StickySelects_6_io_outs_3; // @[MemPrimitives.scala 123:41:@12461.4]
  assign _T_1101 = StickySelects_6_io_outs_4; // @[MemPrimitives.scala 123:41:@12462.4]
  assign _T_1102 = StickySelects_6_io_outs_5; // @[MemPrimitives.scala 123:41:@12463.4]
  assign _T_1103 = StickySelects_6_io_outs_6; // @[MemPrimitives.scala 123:41:@12464.4]
  assign _T_1104 = StickySelects_6_io_outs_7; // @[MemPrimitives.scala 123:41:@12465.4]
  assign _T_1105 = StickySelects_6_io_outs_8; // @[MemPrimitives.scala 123:41:@12466.4]
  assign _T_1107 = {_T_1097,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@12468.4]
  assign _T_1109 = {_T_1098,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@12470.4]
  assign _T_1111 = {_T_1099,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@12472.4]
  assign _T_1113 = {_T_1100,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@12474.4]
  assign _T_1115 = {_T_1101,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@12476.4]
  assign _T_1117 = {_T_1102,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@12478.4]
  assign _T_1119 = {_T_1103,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@12480.4]
  assign _T_1121 = {_T_1104,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@12482.4]
  assign _T_1123 = {_T_1105,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@12484.4]
  assign _T_1124 = _T_1104 ? _T_1121 : _T_1123; // @[Mux.scala 31:69:@12485.4]
  assign _T_1125 = _T_1103 ? _T_1119 : _T_1124; // @[Mux.scala 31:69:@12486.4]
  assign _T_1126 = _T_1102 ? _T_1117 : _T_1125; // @[Mux.scala 31:69:@12487.4]
  assign _T_1127 = _T_1101 ? _T_1115 : _T_1126; // @[Mux.scala 31:69:@12488.4]
  assign _T_1128 = _T_1100 ? _T_1113 : _T_1127; // @[Mux.scala 31:69:@12489.4]
  assign _T_1129 = _T_1099 ? _T_1111 : _T_1128; // @[Mux.scala 31:69:@12490.4]
  assign _T_1130 = _T_1098 ? _T_1109 : _T_1129; // @[Mux.scala 31:69:@12491.4]
  assign _T_1131 = _T_1097 ? _T_1107 : _T_1130; // @[Mux.scala 31:69:@12492.4]
  assign _T_1139 = _T_860 & _T_770; // @[MemPrimitives.scala 110:228:@12501.4]
  assign _T_1145 = _T_866 & _T_776; // @[MemPrimitives.scala 110:228:@12505.4]
  assign _T_1151 = _T_872 & _T_782; // @[MemPrimitives.scala 110:228:@12509.4]
  assign _T_1157 = _T_878 & _T_788; // @[MemPrimitives.scala 110:228:@12513.4]
  assign _T_1163 = _T_884 & _T_794; // @[MemPrimitives.scala 110:228:@12517.4]
  assign _T_1169 = _T_890 & _T_800; // @[MemPrimitives.scala 110:228:@12521.4]
  assign _T_1175 = _T_896 & _T_806; // @[MemPrimitives.scala 110:228:@12525.4]
  assign _T_1181 = _T_902 & _T_812; // @[MemPrimitives.scala 110:228:@12529.4]
  assign _T_1187 = _T_908 & _T_818; // @[MemPrimitives.scala 110:228:@12533.4]
  assign _T_1189 = StickySelects_7_io_outs_0; // @[MemPrimitives.scala 123:41:@12547.4]
  assign _T_1190 = StickySelects_7_io_outs_1; // @[MemPrimitives.scala 123:41:@12548.4]
  assign _T_1191 = StickySelects_7_io_outs_2; // @[MemPrimitives.scala 123:41:@12549.4]
  assign _T_1192 = StickySelects_7_io_outs_3; // @[MemPrimitives.scala 123:41:@12550.4]
  assign _T_1193 = StickySelects_7_io_outs_4; // @[MemPrimitives.scala 123:41:@12551.4]
  assign _T_1194 = StickySelects_7_io_outs_5; // @[MemPrimitives.scala 123:41:@12552.4]
  assign _T_1195 = StickySelects_7_io_outs_6; // @[MemPrimitives.scala 123:41:@12553.4]
  assign _T_1196 = StickySelects_7_io_outs_7; // @[MemPrimitives.scala 123:41:@12554.4]
  assign _T_1197 = StickySelects_7_io_outs_8; // @[MemPrimitives.scala 123:41:@12555.4]
  assign _T_1199 = {_T_1189,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@12557.4]
  assign _T_1201 = {_T_1190,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@12559.4]
  assign _T_1203 = {_T_1191,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@12561.4]
  assign _T_1205 = {_T_1192,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@12563.4]
  assign _T_1207 = {_T_1193,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@12565.4]
  assign _T_1209 = {_T_1194,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@12567.4]
  assign _T_1211 = {_T_1195,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@12569.4]
  assign _T_1213 = {_T_1196,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@12571.4]
  assign _T_1215 = {_T_1197,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@12573.4]
  assign _T_1216 = _T_1196 ? _T_1213 : _T_1215; // @[Mux.scala 31:69:@12574.4]
  assign _T_1217 = _T_1195 ? _T_1211 : _T_1216; // @[Mux.scala 31:69:@12575.4]
  assign _T_1218 = _T_1194 ? _T_1209 : _T_1217; // @[Mux.scala 31:69:@12576.4]
  assign _T_1219 = _T_1193 ? _T_1207 : _T_1218; // @[Mux.scala 31:69:@12577.4]
  assign _T_1220 = _T_1192 ? _T_1205 : _T_1219; // @[Mux.scala 31:69:@12578.4]
  assign _T_1221 = _T_1191 ? _T_1203 : _T_1220; // @[Mux.scala 31:69:@12579.4]
  assign _T_1222 = _T_1190 ? _T_1201 : _T_1221; // @[Mux.scala 31:69:@12580.4]
  assign _T_1223 = _T_1189 ? _T_1199 : _T_1222; // @[Mux.scala 31:69:@12581.4]
  assign _T_1228 = io_rPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@12588.4]
  assign _T_1231 = _T_1228 & _T_494; // @[MemPrimitives.scala 110:228:@12590.4]
  assign _T_1234 = io_rPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@12592.4]
  assign _T_1237 = _T_1234 & _T_500; // @[MemPrimitives.scala 110:228:@12594.4]
  assign _T_1240 = io_rPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@12596.4]
  assign _T_1243 = _T_1240 & _T_506; // @[MemPrimitives.scala 110:228:@12598.4]
  assign _T_1246 = io_rPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@12600.4]
  assign _T_1249 = _T_1246 & _T_512; // @[MemPrimitives.scala 110:228:@12602.4]
  assign _T_1252 = io_rPort_4_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@12604.4]
  assign _T_1255 = _T_1252 & _T_518; // @[MemPrimitives.scala 110:228:@12606.4]
  assign _T_1258 = io_rPort_5_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@12608.4]
  assign _T_1261 = _T_1258 & _T_524; // @[MemPrimitives.scala 110:228:@12610.4]
  assign _T_1264 = io_rPort_6_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@12612.4]
  assign _T_1267 = _T_1264 & _T_530; // @[MemPrimitives.scala 110:228:@12614.4]
  assign _T_1270 = io_rPort_7_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@12616.4]
  assign _T_1273 = _T_1270 & _T_536; // @[MemPrimitives.scala 110:228:@12618.4]
  assign _T_1276 = io_rPort_8_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@12620.4]
  assign _T_1279 = _T_1276 & _T_542; // @[MemPrimitives.scala 110:228:@12622.4]
  assign _T_1281 = StickySelects_8_io_outs_0; // @[MemPrimitives.scala 123:41:@12636.4]
  assign _T_1282 = StickySelects_8_io_outs_1; // @[MemPrimitives.scala 123:41:@12637.4]
  assign _T_1283 = StickySelects_8_io_outs_2; // @[MemPrimitives.scala 123:41:@12638.4]
  assign _T_1284 = StickySelects_8_io_outs_3; // @[MemPrimitives.scala 123:41:@12639.4]
  assign _T_1285 = StickySelects_8_io_outs_4; // @[MemPrimitives.scala 123:41:@12640.4]
  assign _T_1286 = StickySelects_8_io_outs_5; // @[MemPrimitives.scala 123:41:@12641.4]
  assign _T_1287 = StickySelects_8_io_outs_6; // @[MemPrimitives.scala 123:41:@12642.4]
  assign _T_1288 = StickySelects_8_io_outs_7; // @[MemPrimitives.scala 123:41:@12643.4]
  assign _T_1289 = StickySelects_8_io_outs_8; // @[MemPrimitives.scala 123:41:@12644.4]
  assign _T_1291 = {_T_1281,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@12646.4]
  assign _T_1293 = {_T_1282,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@12648.4]
  assign _T_1295 = {_T_1283,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@12650.4]
  assign _T_1297 = {_T_1284,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@12652.4]
  assign _T_1299 = {_T_1285,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@12654.4]
  assign _T_1301 = {_T_1286,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@12656.4]
  assign _T_1303 = {_T_1287,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@12658.4]
  assign _T_1305 = {_T_1288,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@12660.4]
  assign _T_1307 = {_T_1289,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@12662.4]
  assign _T_1308 = _T_1288 ? _T_1305 : _T_1307; // @[Mux.scala 31:69:@12663.4]
  assign _T_1309 = _T_1287 ? _T_1303 : _T_1308; // @[Mux.scala 31:69:@12664.4]
  assign _T_1310 = _T_1286 ? _T_1301 : _T_1309; // @[Mux.scala 31:69:@12665.4]
  assign _T_1311 = _T_1285 ? _T_1299 : _T_1310; // @[Mux.scala 31:69:@12666.4]
  assign _T_1312 = _T_1284 ? _T_1297 : _T_1311; // @[Mux.scala 31:69:@12667.4]
  assign _T_1313 = _T_1283 ? _T_1295 : _T_1312; // @[Mux.scala 31:69:@12668.4]
  assign _T_1314 = _T_1282 ? _T_1293 : _T_1313; // @[Mux.scala 31:69:@12669.4]
  assign _T_1315 = _T_1281 ? _T_1291 : _T_1314; // @[Mux.scala 31:69:@12670.4]
  assign _T_1323 = _T_1228 & _T_586; // @[MemPrimitives.scala 110:228:@12679.4]
  assign _T_1329 = _T_1234 & _T_592; // @[MemPrimitives.scala 110:228:@12683.4]
  assign _T_1335 = _T_1240 & _T_598; // @[MemPrimitives.scala 110:228:@12687.4]
  assign _T_1341 = _T_1246 & _T_604; // @[MemPrimitives.scala 110:228:@12691.4]
  assign _T_1347 = _T_1252 & _T_610; // @[MemPrimitives.scala 110:228:@12695.4]
  assign _T_1353 = _T_1258 & _T_616; // @[MemPrimitives.scala 110:228:@12699.4]
  assign _T_1359 = _T_1264 & _T_622; // @[MemPrimitives.scala 110:228:@12703.4]
  assign _T_1365 = _T_1270 & _T_628; // @[MemPrimitives.scala 110:228:@12707.4]
  assign _T_1371 = _T_1276 & _T_634; // @[MemPrimitives.scala 110:228:@12711.4]
  assign _T_1373 = StickySelects_9_io_outs_0; // @[MemPrimitives.scala 123:41:@12725.4]
  assign _T_1374 = StickySelects_9_io_outs_1; // @[MemPrimitives.scala 123:41:@12726.4]
  assign _T_1375 = StickySelects_9_io_outs_2; // @[MemPrimitives.scala 123:41:@12727.4]
  assign _T_1376 = StickySelects_9_io_outs_3; // @[MemPrimitives.scala 123:41:@12728.4]
  assign _T_1377 = StickySelects_9_io_outs_4; // @[MemPrimitives.scala 123:41:@12729.4]
  assign _T_1378 = StickySelects_9_io_outs_5; // @[MemPrimitives.scala 123:41:@12730.4]
  assign _T_1379 = StickySelects_9_io_outs_6; // @[MemPrimitives.scala 123:41:@12731.4]
  assign _T_1380 = StickySelects_9_io_outs_7; // @[MemPrimitives.scala 123:41:@12732.4]
  assign _T_1381 = StickySelects_9_io_outs_8; // @[MemPrimitives.scala 123:41:@12733.4]
  assign _T_1383 = {_T_1373,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@12735.4]
  assign _T_1385 = {_T_1374,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@12737.4]
  assign _T_1387 = {_T_1375,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@12739.4]
  assign _T_1389 = {_T_1376,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@12741.4]
  assign _T_1391 = {_T_1377,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@12743.4]
  assign _T_1393 = {_T_1378,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@12745.4]
  assign _T_1395 = {_T_1379,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@12747.4]
  assign _T_1397 = {_T_1380,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@12749.4]
  assign _T_1399 = {_T_1381,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@12751.4]
  assign _T_1400 = _T_1380 ? _T_1397 : _T_1399; // @[Mux.scala 31:69:@12752.4]
  assign _T_1401 = _T_1379 ? _T_1395 : _T_1400; // @[Mux.scala 31:69:@12753.4]
  assign _T_1402 = _T_1378 ? _T_1393 : _T_1401; // @[Mux.scala 31:69:@12754.4]
  assign _T_1403 = _T_1377 ? _T_1391 : _T_1402; // @[Mux.scala 31:69:@12755.4]
  assign _T_1404 = _T_1376 ? _T_1389 : _T_1403; // @[Mux.scala 31:69:@12756.4]
  assign _T_1405 = _T_1375 ? _T_1387 : _T_1404; // @[Mux.scala 31:69:@12757.4]
  assign _T_1406 = _T_1374 ? _T_1385 : _T_1405; // @[Mux.scala 31:69:@12758.4]
  assign _T_1407 = _T_1373 ? _T_1383 : _T_1406; // @[Mux.scala 31:69:@12759.4]
  assign _T_1415 = _T_1228 & _T_678; // @[MemPrimitives.scala 110:228:@12768.4]
  assign _T_1421 = _T_1234 & _T_684; // @[MemPrimitives.scala 110:228:@12772.4]
  assign _T_1427 = _T_1240 & _T_690; // @[MemPrimitives.scala 110:228:@12776.4]
  assign _T_1433 = _T_1246 & _T_696; // @[MemPrimitives.scala 110:228:@12780.4]
  assign _T_1439 = _T_1252 & _T_702; // @[MemPrimitives.scala 110:228:@12784.4]
  assign _T_1445 = _T_1258 & _T_708; // @[MemPrimitives.scala 110:228:@12788.4]
  assign _T_1451 = _T_1264 & _T_714; // @[MemPrimitives.scala 110:228:@12792.4]
  assign _T_1457 = _T_1270 & _T_720; // @[MemPrimitives.scala 110:228:@12796.4]
  assign _T_1463 = _T_1276 & _T_726; // @[MemPrimitives.scala 110:228:@12800.4]
  assign _T_1465 = StickySelects_10_io_outs_0; // @[MemPrimitives.scala 123:41:@12814.4]
  assign _T_1466 = StickySelects_10_io_outs_1; // @[MemPrimitives.scala 123:41:@12815.4]
  assign _T_1467 = StickySelects_10_io_outs_2; // @[MemPrimitives.scala 123:41:@12816.4]
  assign _T_1468 = StickySelects_10_io_outs_3; // @[MemPrimitives.scala 123:41:@12817.4]
  assign _T_1469 = StickySelects_10_io_outs_4; // @[MemPrimitives.scala 123:41:@12818.4]
  assign _T_1470 = StickySelects_10_io_outs_5; // @[MemPrimitives.scala 123:41:@12819.4]
  assign _T_1471 = StickySelects_10_io_outs_6; // @[MemPrimitives.scala 123:41:@12820.4]
  assign _T_1472 = StickySelects_10_io_outs_7; // @[MemPrimitives.scala 123:41:@12821.4]
  assign _T_1473 = StickySelects_10_io_outs_8; // @[MemPrimitives.scala 123:41:@12822.4]
  assign _T_1475 = {_T_1465,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@12824.4]
  assign _T_1477 = {_T_1466,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@12826.4]
  assign _T_1479 = {_T_1467,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@12828.4]
  assign _T_1481 = {_T_1468,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@12830.4]
  assign _T_1483 = {_T_1469,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@12832.4]
  assign _T_1485 = {_T_1470,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@12834.4]
  assign _T_1487 = {_T_1471,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@12836.4]
  assign _T_1489 = {_T_1472,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@12838.4]
  assign _T_1491 = {_T_1473,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@12840.4]
  assign _T_1492 = _T_1472 ? _T_1489 : _T_1491; // @[Mux.scala 31:69:@12841.4]
  assign _T_1493 = _T_1471 ? _T_1487 : _T_1492; // @[Mux.scala 31:69:@12842.4]
  assign _T_1494 = _T_1470 ? _T_1485 : _T_1493; // @[Mux.scala 31:69:@12843.4]
  assign _T_1495 = _T_1469 ? _T_1483 : _T_1494; // @[Mux.scala 31:69:@12844.4]
  assign _T_1496 = _T_1468 ? _T_1481 : _T_1495; // @[Mux.scala 31:69:@12845.4]
  assign _T_1497 = _T_1467 ? _T_1479 : _T_1496; // @[Mux.scala 31:69:@12846.4]
  assign _T_1498 = _T_1466 ? _T_1477 : _T_1497; // @[Mux.scala 31:69:@12847.4]
  assign _T_1499 = _T_1465 ? _T_1475 : _T_1498; // @[Mux.scala 31:69:@12848.4]
  assign _T_1507 = _T_1228 & _T_770; // @[MemPrimitives.scala 110:228:@12857.4]
  assign _T_1513 = _T_1234 & _T_776; // @[MemPrimitives.scala 110:228:@12861.4]
  assign _T_1519 = _T_1240 & _T_782; // @[MemPrimitives.scala 110:228:@12865.4]
  assign _T_1525 = _T_1246 & _T_788; // @[MemPrimitives.scala 110:228:@12869.4]
  assign _T_1531 = _T_1252 & _T_794; // @[MemPrimitives.scala 110:228:@12873.4]
  assign _T_1537 = _T_1258 & _T_800; // @[MemPrimitives.scala 110:228:@12877.4]
  assign _T_1543 = _T_1264 & _T_806; // @[MemPrimitives.scala 110:228:@12881.4]
  assign _T_1549 = _T_1270 & _T_812; // @[MemPrimitives.scala 110:228:@12885.4]
  assign _T_1555 = _T_1276 & _T_818; // @[MemPrimitives.scala 110:228:@12889.4]
  assign _T_1557 = StickySelects_11_io_outs_0; // @[MemPrimitives.scala 123:41:@12903.4]
  assign _T_1558 = StickySelects_11_io_outs_1; // @[MemPrimitives.scala 123:41:@12904.4]
  assign _T_1559 = StickySelects_11_io_outs_2; // @[MemPrimitives.scala 123:41:@12905.4]
  assign _T_1560 = StickySelects_11_io_outs_3; // @[MemPrimitives.scala 123:41:@12906.4]
  assign _T_1561 = StickySelects_11_io_outs_4; // @[MemPrimitives.scala 123:41:@12907.4]
  assign _T_1562 = StickySelects_11_io_outs_5; // @[MemPrimitives.scala 123:41:@12908.4]
  assign _T_1563 = StickySelects_11_io_outs_6; // @[MemPrimitives.scala 123:41:@12909.4]
  assign _T_1564 = StickySelects_11_io_outs_7; // @[MemPrimitives.scala 123:41:@12910.4]
  assign _T_1565 = StickySelects_11_io_outs_8; // @[MemPrimitives.scala 123:41:@12911.4]
  assign _T_1567 = {_T_1557,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@12913.4]
  assign _T_1569 = {_T_1558,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@12915.4]
  assign _T_1571 = {_T_1559,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@12917.4]
  assign _T_1573 = {_T_1560,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@12919.4]
  assign _T_1575 = {_T_1561,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@12921.4]
  assign _T_1577 = {_T_1562,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@12923.4]
  assign _T_1579 = {_T_1563,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@12925.4]
  assign _T_1581 = {_T_1564,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@12927.4]
  assign _T_1583 = {_T_1565,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@12929.4]
  assign _T_1584 = _T_1564 ? _T_1581 : _T_1583; // @[Mux.scala 31:69:@12930.4]
  assign _T_1585 = _T_1563 ? _T_1579 : _T_1584; // @[Mux.scala 31:69:@12931.4]
  assign _T_1586 = _T_1562 ? _T_1577 : _T_1585; // @[Mux.scala 31:69:@12932.4]
  assign _T_1587 = _T_1561 ? _T_1575 : _T_1586; // @[Mux.scala 31:69:@12933.4]
  assign _T_1588 = _T_1560 ? _T_1573 : _T_1587; // @[Mux.scala 31:69:@12934.4]
  assign _T_1589 = _T_1559 ? _T_1571 : _T_1588; // @[Mux.scala 31:69:@12935.4]
  assign _T_1590 = _T_1558 ? _T_1569 : _T_1589; // @[Mux.scala 31:69:@12936.4]
  assign _T_1591 = _T_1557 ? _T_1567 : _T_1590; // @[Mux.scala 31:69:@12937.4]
  assign _T_1596 = io_rPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@12944.4]
  assign _T_1599 = _T_1596 & _T_494; // @[MemPrimitives.scala 110:228:@12946.4]
  assign _T_1602 = io_rPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@12948.4]
  assign _T_1605 = _T_1602 & _T_500; // @[MemPrimitives.scala 110:228:@12950.4]
  assign _T_1608 = io_rPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@12952.4]
  assign _T_1611 = _T_1608 & _T_506; // @[MemPrimitives.scala 110:228:@12954.4]
  assign _T_1614 = io_rPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@12956.4]
  assign _T_1617 = _T_1614 & _T_512; // @[MemPrimitives.scala 110:228:@12958.4]
  assign _T_1620 = io_rPort_4_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@12960.4]
  assign _T_1623 = _T_1620 & _T_518; // @[MemPrimitives.scala 110:228:@12962.4]
  assign _T_1626 = io_rPort_5_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@12964.4]
  assign _T_1629 = _T_1626 & _T_524; // @[MemPrimitives.scala 110:228:@12966.4]
  assign _T_1632 = io_rPort_6_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@12968.4]
  assign _T_1635 = _T_1632 & _T_530; // @[MemPrimitives.scala 110:228:@12970.4]
  assign _T_1638 = io_rPort_7_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@12972.4]
  assign _T_1641 = _T_1638 & _T_536; // @[MemPrimitives.scala 110:228:@12974.4]
  assign _T_1644 = io_rPort_8_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@12976.4]
  assign _T_1647 = _T_1644 & _T_542; // @[MemPrimitives.scala 110:228:@12978.4]
  assign _T_1649 = StickySelects_12_io_outs_0; // @[MemPrimitives.scala 123:41:@12992.4]
  assign _T_1650 = StickySelects_12_io_outs_1; // @[MemPrimitives.scala 123:41:@12993.4]
  assign _T_1651 = StickySelects_12_io_outs_2; // @[MemPrimitives.scala 123:41:@12994.4]
  assign _T_1652 = StickySelects_12_io_outs_3; // @[MemPrimitives.scala 123:41:@12995.4]
  assign _T_1653 = StickySelects_12_io_outs_4; // @[MemPrimitives.scala 123:41:@12996.4]
  assign _T_1654 = StickySelects_12_io_outs_5; // @[MemPrimitives.scala 123:41:@12997.4]
  assign _T_1655 = StickySelects_12_io_outs_6; // @[MemPrimitives.scala 123:41:@12998.4]
  assign _T_1656 = StickySelects_12_io_outs_7; // @[MemPrimitives.scala 123:41:@12999.4]
  assign _T_1657 = StickySelects_12_io_outs_8; // @[MemPrimitives.scala 123:41:@13000.4]
  assign _T_1659 = {_T_1649,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13002.4]
  assign _T_1661 = {_T_1650,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13004.4]
  assign _T_1663 = {_T_1651,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13006.4]
  assign _T_1665 = {_T_1652,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13008.4]
  assign _T_1667 = {_T_1653,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13010.4]
  assign _T_1669 = {_T_1654,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13012.4]
  assign _T_1671 = {_T_1655,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13014.4]
  assign _T_1673 = {_T_1656,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13016.4]
  assign _T_1675 = {_T_1657,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13018.4]
  assign _T_1676 = _T_1656 ? _T_1673 : _T_1675; // @[Mux.scala 31:69:@13019.4]
  assign _T_1677 = _T_1655 ? _T_1671 : _T_1676; // @[Mux.scala 31:69:@13020.4]
  assign _T_1678 = _T_1654 ? _T_1669 : _T_1677; // @[Mux.scala 31:69:@13021.4]
  assign _T_1679 = _T_1653 ? _T_1667 : _T_1678; // @[Mux.scala 31:69:@13022.4]
  assign _T_1680 = _T_1652 ? _T_1665 : _T_1679; // @[Mux.scala 31:69:@13023.4]
  assign _T_1681 = _T_1651 ? _T_1663 : _T_1680; // @[Mux.scala 31:69:@13024.4]
  assign _T_1682 = _T_1650 ? _T_1661 : _T_1681; // @[Mux.scala 31:69:@13025.4]
  assign _T_1683 = _T_1649 ? _T_1659 : _T_1682; // @[Mux.scala 31:69:@13026.4]
  assign _T_1691 = _T_1596 & _T_586; // @[MemPrimitives.scala 110:228:@13035.4]
  assign _T_1697 = _T_1602 & _T_592; // @[MemPrimitives.scala 110:228:@13039.4]
  assign _T_1703 = _T_1608 & _T_598; // @[MemPrimitives.scala 110:228:@13043.4]
  assign _T_1709 = _T_1614 & _T_604; // @[MemPrimitives.scala 110:228:@13047.4]
  assign _T_1715 = _T_1620 & _T_610; // @[MemPrimitives.scala 110:228:@13051.4]
  assign _T_1721 = _T_1626 & _T_616; // @[MemPrimitives.scala 110:228:@13055.4]
  assign _T_1727 = _T_1632 & _T_622; // @[MemPrimitives.scala 110:228:@13059.4]
  assign _T_1733 = _T_1638 & _T_628; // @[MemPrimitives.scala 110:228:@13063.4]
  assign _T_1739 = _T_1644 & _T_634; // @[MemPrimitives.scala 110:228:@13067.4]
  assign _T_1741 = StickySelects_13_io_outs_0; // @[MemPrimitives.scala 123:41:@13081.4]
  assign _T_1742 = StickySelects_13_io_outs_1; // @[MemPrimitives.scala 123:41:@13082.4]
  assign _T_1743 = StickySelects_13_io_outs_2; // @[MemPrimitives.scala 123:41:@13083.4]
  assign _T_1744 = StickySelects_13_io_outs_3; // @[MemPrimitives.scala 123:41:@13084.4]
  assign _T_1745 = StickySelects_13_io_outs_4; // @[MemPrimitives.scala 123:41:@13085.4]
  assign _T_1746 = StickySelects_13_io_outs_5; // @[MemPrimitives.scala 123:41:@13086.4]
  assign _T_1747 = StickySelects_13_io_outs_6; // @[MemPrimitives.scala 123:41:@13087.4]
  assign _T_1748 = StickySelects_13_io_outs_7; // @[MemPrimitives.scala 123:41:@13088.4]
  assign _T_1749 = StickySelects_13_io_outs_8; // @[MemPrimitives.scala 123:41:@13089.4]
  assign _T_1751 = {_T_1741,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13091.4]
  assign _T_1753 = {_T_1742,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13093.4]
  assign _T_1755 = {_T_1743,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13095.4]
  assign _T_1757 = {_T_1744,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13097.4]
  assign _T_1759 = {_T_1745,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13099.4]
  assign _T_1761 = {_T_1746,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13101.4]
  assign _T_1763 = {_T_1747,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13103.4]
  assign _T_1765 = {_T_1748,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13105.4]
  assign _T_1767 = {_T_1749,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13107.4]
  assign _T_1768 = _T_1748 ? _T_1765 : _T_1767; // @[Mux.scala 31:69:@13108.4]
  assign _T_1769 = _T_1747 ? _T_1763 : _T_1768; // @[Mux.scala 31:69:@13109.4]
  assign _T_1770 = _T_1746 ? _T_1761 : _T_1769; // @[Mux.scala 31:69:@13110.4]
  assign _T_1771 = _T_1745 ? _T_1759 : _T_1770; // @[Mux.scala 31:69:@13111.4]
  assign _T_1772 = _T_1744 ? _T_1757 : _T_1771; // @[Mux.scala 31:69:@13112.4]
  assign _T_1773 = _T_1743 ? _T_1755 : _T_1772; // @[Mux.scala 31:69:@13113.4]
  assign _T_1774 = _T_1742 ? _T_1753 : _T_1773; // @[Mux.scala 31:69:@13114.4]
  assign _T_1775 = _T_1741 ? _T_1751 : _T_1774; // @[Mux.scala 31:69:@13115.4]
  assign _T_1783 = _T_1596 & _T_678; // @[MemPrimitives.scala 110:228:@13124.4]
  assign _T_1789 = _T_1602 & _T_684; // @[MemPrimitives.scala 110:228:@13128.4]
  assign _T_1795 = _T_1608 & _T_690; // @[MemPrimitives.scala 110:228:@13132.4]
  assign _T_1801 = _T_1614 & _T_696; // @[MemPrimitives.scala 110:228:@13136.4]
  assign _T_1807 = _T_1620 & _T_702; // @[MemPrimitives.scala 110:228:@13140.4]
  assign _T_1813 = _T_1626 & _T_708; // @[MemPrimitives.scala 110:228:@13144.4]
  assign _T_1819 = _T_1632 & _T_714; // @[MemPrimitives.scala 110:228:@13148.4]
  assign _T_1825 = _T_1638 & _T_720; // @[MemPrimitives.scala 110:228:@13152.4]
  assign _T_1831 = _T_1644 & _T_726; // @[MemPrimitives.scala 110:228:@13156.4]
  assign _T_1833 = StickySelects_14_io_outs_0; // @[MemPrimitives.scala 123:41:@13170.4]
  assign _T_1834 = StickySelects_14_io_outs_1; // @[MemPrimitives.scala 123:41:@13171.4]
  assign _T_1835 = StickySelects_14_io_outs_2; // @[MemPrimitives.scala 123:41:@13172.4]
  assign _T_1836 = StickySelects_14_io_outs_3; // @[MemPrimitives.scala 123:41:@13173.4]
  assign _T_1837 = StickySelects_14_io_outs_4; // @[MemPrimitives.scala 123:41:@13174.4]
  assign _T_1838 = StickySelects_14_io_outs_5; // @[MemPrimitives.scala 123:41:@13175.4]
  assign _T_1839 = StickySelects_14_io_outs_6; // @[MemPrimitives.scala 123:41:@13176.4]
  assign _T_1840 = StickySelects_14_io_outs_7; // @[MemPrimitives.scala 123:41:@13177.4]
  assign _T_1841 = StickySelects_14_io_outs_8; // @[MemPrimitives.scala 123:41:@13178.4]
  assign _T_1843 = {_T_1833,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13180.4]
  assign _T_1845 = {_T_1834,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13182.4]
  assign _T_1847 = {_T_1835,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13184.4]
  assign _T_1849 = {_T_1836,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13186.4]
  assign _T_1851 = {_T_1837,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13188.4]
  assign _T_1853 = {_T_1838,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13190.4]
  assign _T_1855 = {_T_1839,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13192.4]
  assign _T_1857 = {_T_1840,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13194.4]
  assign _T_1859 = {_T_1841,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13196.4]
  assign _T_1860 = _T_1840 ? _T_1857 : _T_1859; // @[Mux.scala 31:69:@13197.4]
  assign _T_1861 = _T_1839 ? _T_1855 : _T_1860; // @[Mux.scala 31:69:@13198.4]
  assign _T_1862 = _T_1838 ? _T_1853 : _T_1861; // @[Mux.scala 31:69:@13199.4]
  assign _T_1863 = _T_1837 ? _T_1851 : _T_1862; // @[Mux.scala 31:69:@13200.4]
  assign _T_1864 = _T_1836 ? _T_1849 : _T_1863; // @[Mux.scala 31:69:@13201.4]
  assign _T_1865 = _T_1835 ? _T_1847 : _T_1864; // @[Mux.scala 31:69:@13202.4]
  assign _T_1866 = _T_1834 ? _T_1845 : _T_1865; // @[Mux.scala 31:69:@13203.4]
  assign _T_1867 = _T_1833 ? _T_1843 : _T_1866; // @[Mux.scala 31:69:@13204.4]
  assign _T_1875 = _T_1596 & _T_770; // @[MemPrimitives.scala 110:228:@13213.4]
  assign _T_1881 = _T_1602 & _T_776; // @[MemPrimitives.scala 110:228:@13217.4]
  assign _T_1887 = _T_1608 & _T_782; // @[MemPrimitives.scala 110:228:@13221.4]
  assign _T_1893 = _T_1614 & _T_788; // @[MemPrimitives.scala 110:228:@13225.4]
  assign _T_1899 = _T_1620 & _T_794; // @[MemPrimitives.scala 110:228:@13229.4]
  assign _T_1905 = _T_1626 & _T_800; // @[MemPrimitives.scala 110:228:@13233.4]
  assign _T_1911 = _T_1632 & _T_806; // @[MemPrimitives.scala 110:228:@13237.4]
  assign _T_1917 = _T_1638 & _T_812; // @[MemPrimitives.scala 110:228:@13241.4]
  assign _T_1923 = _T_1644 & _T_818; // @[MemPrimitives.scala 110:228:@13245.4]
  assign _T_1925 = StickySelects_15_io_outs_0; // @[MemPrimitives.scala 123:41:@13259.4]
  assign _T_1926 = StickySelects_15_io_outs_1; // @[MemPrimitives.scala 123:41:@13260.4]
  assign _T_1927 = StickySelects_15_io_outs_2; // @[MemPrimitives.scala 123:41:@13261.4]
  assign _T_1928 = StickySelects_15_io_outs_3; // @[MemPrimitives.scala 123:41:@13262.4]
  assign _T_1929 = StickySelects_15_io_outs_4; // @[MemPrimitives.scala 123:41:@13263.4]
  assign _T_1930 = StickySelects_15_io_outs_5; // @[MemPrimitives.scala 123:41:@13264.4]
  assign _T_1931 = StickySelects_15_io_outs_6; // @[MemPrimitives.scala 123:41:@13265.4]
  assign _T_1932 = StickySelects_15_io_outs_7; // @[MemPrimitives.scala 123:41:@13266.4]
  assign _T_1933 = StickySelects_15_io_outs_8; // @[MemPrimitives.scala 123:41:@13267.4]
  assign _T_1935 = {_T_1925,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13269.4]
  assign _T_1937 = {_T_1926,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13271.4]
  assign _T_1939 = {_T_1927,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13273.4]
  assign _T_1941 = {_T_1928,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13275.4]
  assign _T_1943 = {_T_1929,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13277.4]
  assign _T_1945 = {_T_1930,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13279.4]
  assign _T_1947 = {_T_1931,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13281.4]
  assign _T_1949 = {_T_1932,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13283.4]
  assign _T_1951 = {_T_1933,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13285.4]
  assign _T_1952 = _T_1932 ? _T_1949 : _T_1951; // @[Mux.scala 31:69:@13286.4]
  assign _T_1953 = _T_1931 ? _T_1947 : _T_1952; // @[Mux.scala 31:69:@13287.4]
  assign _T_1954 = _T_1930 ? _T_1945 : _T_1953; // @[Mux.scala 31:69:@13288.4]
  assign _T_1955 = _T_1929 ? _T_1943 : _T_1954; // @[Mux.scala 31:69:@13289.4]
  assign _T_1956 = _T_1928 ? _T_1941 : _T_1955; // @[Mux.scala 31:69:@13290.4]
  assign _T_1957 = _T_1927 ? _T_1939 : _T_1956; // @[Mux.scala 31:69:@13291.4]
  assign _T_1958 = _T_1926 ? _T_1937 : _T_1957; // @[Mux.scala 31:69:@13292.4]
  assign _T_1959 = _T_1925 ? _T_1935 : _T_1958; // @[Mux.scala 31:69:@13293.4]
  assign _T_2087 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@13466.4 package.scala 96:25:@13467.4]
  assign _T_2091 = _T_2087 ? Mem1D_14_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@13476.4]
  assign _T_2084 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@13458.4 package.scala 96:25:@13459.4]
  assign _T_2092 = _T_2084 ? Mem1D_13_io_output : _T_2091; // @[Mux.scala 31:69:@13477.4]
  assign _T_2081 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@13450.4 package.scala 96:25:@13451.4]
  assign _T_2093 = _T_2081 ? Mem1D_12_io_output : _T_2092; // @[Mux.scala 31:69:@13478.4]
  assign _T_2078 = RetimeWrapper_11_io_out; // @[package.scala 96:25:@13442.4 package.scala 96:25:@13443.4]
  assign _T_2094 = _T_2078 ? Mem1D_11_io_output : _T_2093; // @[Mux.scala 31:69:@13479.4]
  assign _T_2075 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@13434.4 package.scala 96:25:@13435.4]
  assign _T_2095 = _T_2075 ? Mem1D_10_io_output : _T_2094; // @[Mux.scala 31:69:@13480.4]
  assign _T_2072 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@13426.4 package.scala 96:25:@13427.4]
  assign _T_2096 = _T_2072 ? Mem1D_9_io_output : _T_2095; // @[Mux.scala 31:69:@13481.4]
  assign _T_2069 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@13418.4 package.scala 96:25:@13419.4]
  assign _T_2097 = _T_2069 ? Mem1D_8_io_output : _T_2096; // @[Mux.scala 31:69:@13482.4]
  assign _T_2066 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@13410.4 package.scala 96:25:@13411.4]
  assign _T_2098 = _T_2066 ? Mem1D_7_io_output : _T_2097; // @[Mux.scala 31:69:@13483.4]
  assign _T_2063 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@13402.4 package.scala 96:25:@13403.4]
  assign _T_2099 = _T_2063 ? Mem1D_6_io_output : _T_2098; // @[Mux.scala 31:69:@13484.4]
  assign _T_2060 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@13394.4 package.scala 96:25:@13395.4]
  assign _T_2100 = _T_2060 ? Mem1D_5_io_output : _T_2099; // @[Mux.scala 31:69:@13485.4]
  assign _T_2057 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@13386.4 package.scala 96:25:@13387.4]
  assign _T_2101 = _T_2057 ? Mem1D_4_io_output : _T_2100; // @[Mux.scala 31:69:@13486.4]
  assign _T_2054 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@13378.4 package.scala 96:25:@13379.4]
  assign _T_2102 = _T_2054 ? Mem1D_3_io_output : _T_2101; // @[Mux.scala 31:69:@13487.4]
  assign _T_2051 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@13370.4 package.scala 96:25:@13371.4]
  assign _T_2103 = _T_2051 ? Mem1D_2_io_output : _T_2102; // @[Mux.scala 31:69:@13488.4]
  assign _T_2048 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@13362.4 package.scala 96:25:@13363.4]
  assign _T_2104 = _T_2048 ? Mem1D_1_io_output : _T_2103; // @[Mux.scala 31:69:@13489.4]
  assign _T_2045 = RetimeWrapper_io_out; // @[package.scala 96:25:@13354.4 package.scala 96:25:@13355.4]
  assign _T_2230 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@13658.4 package.scala 96:25:@13659.4]
  assign _T_2234 = _T_2230 ? Mem1D_14_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@13668.4]
  assign _T_2227 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@13650.4 package.scala 96:25:@13651.4]
  assign _T_2235 = _T_2227 ? Mem1D_13_io_output : _T_2234; // @[Mux.scala 31:69:@13669.4]
  assign _T_2224 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@13642.4 package.scala 96:25:@13643.4]
  assign _T_2236 = _T_2224 ? Mem1D_12_io_output : _T_2235; // @[Mux.scala 31:69:@13670.4]
  assign _T_2221 = RetimeWrapper_27_io_out; // @[package.scala 96:25:@13634.4 package.scala 96:25:@13635.4]
  assign _T_2237 = _T_2221 ? Mem1D_11_io_output : _T_2236; // @[Mux.scala 31:69:@13671.4]
  assign _T_2218 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@13626.4 package.scala 96:25:@13627.4]
  assign _T_2238 = _T_2218 ? Mem1D_10_io_output : _T_2237; // @[Mux.scala 31:69:@13672.4]
  assign _T_2215 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@13618.4 package.scala 96:25:@13619.4]
  assign _T_2239 = _T_2215 ? Mem1D_9_io_output : _T_2238; // @[Mux.scala 31:69:@13673.4]
  assign _T_2212 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@13610.4 package.scala 96:25:@13611.4]
  assign _T_2240 = _T_2212 ? Mem1D_8_io_output : _T_2239; // @[Mux.scala 31:69:@13674.4]
  assign _T_2209 = RetimeWrapper_23_io_out; // @[package.scala 96:25:@13602.4 package.scala 96:25:@13603.4]
  assign _T_2241 = _T_2209 ? Mem1D_7_io_output : _T_2240; // @[Mux.scala 31:69:@13675.4]
  assign _T_2206 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@13594.4 package.scala 96:25:@13595.4]
  assign _T_2242 = _T_2206 ? Mem1D_6_io_output : _T_2241; // @[Mux.scala 31:69:@13676.4]
  assign _T_2203 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@13586.4 package.scala 96:25:@13587.4]
  assign _T_2243 = _T_2203 ? Mem1D_5_io_output : _T_2242; // @[Mux.scala 31:69:@13677.4]
  assign _T_2200 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@13578.4 package.scala 96:25:@13579.4]
  assign _T_2244 = _T_2200 ? Mem1D_4_io_output : _T_2243; // @[Mux.scala 31:69:@13678.4]
  assign _T_2197 = RetimeWrapper_19_io_out; // @[package.scala 96:25:@13570.4 package.scala 96:25:@13571.4]
  assign _T_2245 = _T_2197 ? Mem1D_3_io_output : _T_2244; // @[Mux.scala 31:69:@13679.4]
  assign _T_2194 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@13562.4 package.scala 96:25:@13563.4]
  assign _T_2246 = _T_2194 ? Mem1D_2_io_output : _T_2245; // @[Mux.scala 31:69:@13680.4]
  assign _T_2191 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@13554.4 package.scala 96:25:@13555.4]
  assign _T_2247 = _T_2191 ? Mem1D_1_io_output : _T_2246; // @[Mux.scala 31:69:@13681.4]
  assign _T_2188 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@13546.4 package.scala 96:25:@13547.4]
  assign _T_2373 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@13850.4 package.scala 96:25:@13851.4]
  assign _T_2377 = _T_2373 ? Mem1D_14_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@13860.4]
  assign _T_2370 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@13842.4 package.scala 96:25:@13843.4]
  assign _T_2378 = _T_2370 ? Mem1D_13_io_output : _T_2377; // @[Mux.scala 31:69:@13861.4]
  assign _T_2367 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@13834.4 package.scala 96:25:@13835.4]
  assign _T_2379 = _T_2367 ? Mem1D_12_io_output : _T_2378; // @[Mux.scala 31:69:@13862.4]
  assign _T_2364 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@13826.4 package.scala 96:25:@13827.4]
  assign _T_2380 = _T_2364 ? Mem1D_11_io_output : _T_2379; // @[Mux.scala 31:69:@13863.4]
  assign _T_2361 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@13818.4 package.scala 96:25:@13819.4]
  assign _T_2381 = _T_2361 ? Mem1D_10_io_output : _T_2380; // @[Mux.scala 31:69:@13864.4]
  assign _T_2358 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@13810.4 package.scala 96:25:@13811.4]
  assign _T_2382 = _T_2358 ? Mem1D_9_io_output : _T_2381; // @[Mux.scala 31:69:@13865.4]
  assign _T_2355 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@13802.4 package.scala 96:25:@13803.4]
  assign _T_2383 = _T_2355 ? Mem1D_8_io_output : _T_2382; // @[Mux.scala 31:69:@13866.4]
  assign _T_2352 = RetimeWrapper_39_io_out; // @[package.scala 96:25:@13794.4 package.scala 96:25:@13795.4]
  assign _T_2384 = _T_2352 ? Mem1D_7_io_output : _T_2383; // @[Mux.scala 31:69:@13867.4]
  assign _T_2349 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@13786.4 package.scala 96:25:@13787.4]
  assign _T_2385 = _T_2349 ? Mem1D_6_io_output : _T_2384; // @[Mux.scala 31:69:@13868.4]
  assign _T_2346 = RetimeWrapper_37_io_out; // @[package.scala 96:25:@13778.4 package.scala 96:25:@13779.4]
  assign _T_2386 = _T_2346 ? Mem1D_5_io_output : _T_2385; // @[Mux.scala 31:69:@13869.4]
  assign _T_2343 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@13770.4 package.scala 96:25:@13771.4]
  assign _T_2387 = _T_2343 ? Mem1D_4_io_output : _T_2386; // @[Mux.scala 31:69:@13870.4]
  assign _T_2340 = RetimeWrapper_35_io_out; // @[package.scala 96:25:@13762.4 package.scala 96:25:@13763.4]
  assign _T_2388 = _T_2340 ? Mem1D_3_io_output : _T_2387; // @[Mux.scala 31:69:@13871.4]
  assign _T_2337 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@13754.4 package.scala 96:25:@13755.4]
  assign _T_2389 = _T_2337 ? Mem1D_2_io_output : _T_2388; // @[Mux.scala 31:69:@13872.4]
  assign _T_2334 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@13746.4 package.scala 96:25:@13747.4]
  assign _T_2390 = _T_2334 ? Mem1D_1_io_output : _T_2389; // @[Mux.scala 31:69:@13873.4]
  assign _T_2331 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@13738.4 package.scala 96:25:@13739.4]
  assign _T_2516 = RetimeWrapper_62_io_out; // @[package.scala 96:25:@14042.4 package.scala 96:25:@14043.4]
  assign _T_2520 = _T_2516 ? Mem1D_14_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@14052.4]
  assign _T_2513 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@14034.4 package.scala 96:25:@14035.4]
  assign _T_2521 = _T_2513 ? Mem1D_13_io_output : _T_2520; // @[Mux.scala 31:69:@14053.4]
  assign _T_2510 = RetimeWrapper_60_io_out; // @[package.scala 96:25:@14026.4 package.scala 96:25:@14027.4]
  assign _T_2522 = _T_2510 ? Mem1D_12_io_output : _T_2521; // @[Mux.scala 31:69:@14054.4]
  assign _T_2507 = RetimeWrapper_59_io_out; // @[package.scala 96:25:@14018.4 package.scala 96:25:@14019.4]
  assign _T_2523 = _T_2507 ? Mem1D_11_io_output : _T_2522; // @[Mux.scala 31:69:@14055.4]
  assign _T_2504 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@14010.4 package.scala 96:25:@14011.4]
  assign _T_2524 = _T_2504 ? Mem1D_10_io_output : _T_2523; // @[Mux.scala 31:69:@14056.4]
  assign _T_2501 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@14002.4 package.scala 96:25:@14003.4]
  assign _T_2525 = _T_2501 ? Mem1D_9_io_output : _T_2524; // @[Mux.scala 31:69:@14057.4]
  assign _T_2498 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@13994.4 package.scala 96:25:@13995.4]
  assign _T_2526 = _T_2498 ? Mem1D_8_io_output : _T_2525; // @[Mux.scala 31:69:@14058.4]
  assign _T_2495 = RetimeWrapper_55_io_out; // @[package.scala 96:25:@13986.4 package.scala 96:25:@13987.4]
  assign _T_2527 = _T_2495 ? Mem1D_7_io_output : _T_2526; // @[Mux.scala 31:69:@14059.4]
  assign _T_2492 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@13978.4 package.scala 96:25:@13979.4]
  assign _T_2528 = _T_2492 ? Mem1D_6_io_output : _T_2527; // @[Mux.scala 31:69:@14060.4]
  assign _T_2489 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@13970.4 package.scala 96:25:@13971.4]
  assign _T_2529 = _T_2489 ? Mem1D_5_io_output : _T_2528; // @[Mux.scala 31:69:@14061.4]
  assign _T_2486 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@13962.4 package.scala 96:25:@13963.4]
  assign _T_2530 = _T_2486 ? Mem1D_4_io_output : _T_2529; // @[Mux.scala 31:69:@14062.4]
  assign _T_2483 = RetimeWrapper_51_io_out; // @[package.scala 96:25:@13954.4 package.scala 96:25:@13955.4]
  assign _T_2531 = _T_2483 ? Mem1D_3_io_output : _T_2530; // @[Mux.scala 31:69:@14063.4]
  assign _T_2480 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@13946.4 package.scala 96:25:@13947.4]
  assign _T_2532 = _T_2480 ? Mem1D_2_io_output : _T_2531; // @[Mux.scala 31:69:@14064.4]
  assign _T_2477 = RetimeWrapper_49_io_out; // @[package.scala 96:25:@13938.4 package.scala 96:25:@13939.4]
  assign _T_2533 = _T_2477 ? Mem1D_1_io_output : _T_2532; // @[Mux.scala 31:69:@14065.4]
  assign _T_2474 = RetimeWrapper_48_io_out; // @[package.scala 96:25:@13930.4 package.scala 96:25:@13931.4]
  assign _T_2659 = RetimeWrapper_78_io_out; // @[package.scala 96:25:@14234.4 package.scala 96:25:@14235.4]
  assign _T_2663 = _T_2659 ? Mem1D_14_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@14244.4]
  assign _T_2656 = RetimeWrapper_77_io_out; // @[package.scala 96:25:@14226.4 package.scala 96:25:@14227.4]
  assign _T_2664 = _T_2656 ? Mem1D_13_io_output : _T_2663; // @[Mux.scala 31:69:@14245.4]
  assign _T_2653 = RetimeWrapper_76_io_out; // @[package.scala 96:25:@14218.4 package.scala 96:25:@14219.4]
  assign _T_2665 = _T_2653 ? Mem1D_12_io_output : _T_2664; // @[Mux.scala 31:69:@14246.4]
  assign _T_2650 = RetimeWrapper_75_io_out; // @[package.scala 96:25:@14210.4 package.scala 96:25:@14211.4]
  assign _T_2666 = _T_2650 ? Mem1D_11_io_output : _T_2665; // @[Mux.scala 31:69:@14247.4]
  assign _T_2647 = RetimeWrapper_74_io_out; // @[package.scala 96:25:@14202.4 package.scala 96:25:@14203.4]
  assign _T_2667 = _T_2647 ? Mem1D_10_io_output : _T_2666; // @[Mux.scala 31:69:@14248.4]
  assign _T_2644 = RetimeWrapper_73_io_out; // @[package.scala 96:25:@14194.4 package.scala 96:25:@14195.4]
  assign _T_2668 = _T_2644 ? Mem1D_9_io_output : _T_2667; // @[Mux.scala 31:69:@14249.4]
  assign _T_2641 = RetimeWrapper_72_io_out; // @[package.scala 96:25:@14186.4 package.scala 96:25:@14187.4]
  assign _T_2669 = _T_2641 ? Mem1D_8_io_output : _T_2668; // @[Mux.scala 31:69:@14250.4]
  assign _T_2638 = RetimeWrapper_71_io_out; // @[package.scala 96:25:@14178.4 package.scala 96:25:@14179.4]
  assign _T_2670 = _T_2638 ? Mem1D_7_io_output : _T_2669; // @[Mux.scala 31:69:@14251.4]
  assign _T_2635 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@14170.4 package.scala 96:25:@14171.4]
  assign _T_2671 = _T_2635 ? Mem1D_6_io_output : _T_2670; // @[Mux.scala 31:69:@14252.4]
  assign _T_2632 = RetimeWrapper_69_io_out; // @[package.scala 96:25:@14162.4 package.scala 96:25:@14163.4]
  assign _T_2672 = _T_2632 ? Mem1D_5_io_output : _T_2671; // @[Mux.scala 31:69:@14253.4]
  assign _T_2629 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@14154.4 package.scala 96:25:@14155.4]
  assign _T_2673 = _T_2629 ? Mem1D_4_io_output : _T_2672; // @[Mux.scala 31:69:@14254.4]
  assign _T_2626 = RetimeWrapper_67_io_out; // @[package.scala 96:25:@14146.4 package.scala 96:25:@14147.4]
  assign _T_2674 = _T_2626 ? Mem1D_3_io_output : _T_2673; // @[Mux.scala 31:69:@14255.4]
  assign _T_2623 = RetimeWrapper_66_io_out; // @[package.scala 96:25:@14138.4 package.scala 96:25:@14139.4]
  assign _T_2675 = _T_2623 ? Mem1D_2_io_output : _T_2674; // @[Mux.scala 31:69:@14256.4]
  assign _T_2620 = RetimeWrapper_65_io_out; // @[package.scala 96:25:@14130.4 package.scala 96:25:@14131.4]
  assign _T_2676 = _T_2620 ? Mem1D_1_io_output : _T_2675; // @[Mux.scala 31:69:@14257.4]
  assign _T_2617 = RetimeWrapper_64_io_out; // @[package.scala 96:25:@14122.4 package.scala 96:25:@14123.4]
  assign _T_2802 = RetimeWrapper_94_io_out; // @[package.scala 96:25:@14426.4 package.scala 96:25:@14427.4]
  assign _T_2806 = _T_2802 ? Mem1D_14_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@14436.4]
  assign _T_2799 = RetimeWrapper_93_io_out; // @[package.scala 96:25:@14418.4 package.scala 96:25:@14419.4]
  assign _T_2807 = _T_2799 ? Mem1D_13_io_output : _T_2806; // @[Mux.scala 31:69:@14437.4]
  assign _T_2796 = RetimeWrapper_92_io_out; // @[package.scala 96:25:@14410.4 package.scala 96:25:@14411.4]
  assign _T_2808 = _T_2796 ? Mem1D_12_io_output : _T_2807; // @[Mux.scala 31:69:@14438.4]
  assign _T_2793 = RetimeWrapper_91_io_out; // @[package.scala 96:25:@14402.4 package.scala 96:25:@14403.4]
  assign _T_2809 = _T_2793 ? Mem1D_11_io_output : _T_2808; // @[Mux.scala 31:69:@14439.4]
  assign _T_2790 = RetimeWrapper_90_io_out; // @[package.scala 96:25:@14394.4 package.scala 96:25:@14395.4]
  assign _T_2810 = _T_2790 ? Mem1D_10_io_output : _T_2809; // @[Mux.scala 31:69:@14440.4]
  assign _T_2787 = RetimeWrapper_89_io_out; // @[package.scala 96:25:@14386.4 package.scala 96:25:@14387.4]
  assign _T_2811 = _T_2787 ? Mem1D_9_io_output : _T_2810; // @[Mux.scala 31:69:@14441.4]
  assign _T_2784 = RetimeWrapper_88_io_out; // @[package.scala 96:25:@14378.4 package.scala 96:25:@14379.4]
  assign _T_2812 = _T_2784 ? Mem1D_8_io_output : _T_2811; // @[Mux.scala 31:69:@14442.4]
  assign _T_2781 = RetimeWrapper_87_io_out; // @[package.scala 96:25:@14370.4 package.scala 96:25:@14371.4]
  assign _T_2813 = _T_2781 ? Mem1D_7_io_output : _T_2812; // @[Mux.scala 31:69:@14443.4]
  assign _T_2778 = RetimeWrapper_86_io_out; // @[package.scala 96:25:@14362.4 package.scala 96:25:@14363.4]
  assign _T_2814 = _T_2778 ? Mem1D_6_io_output : _T_2813; // @[Mux.scala 31:69:@14444.4]
  assign _T_2775 = RetimeWrapper_85_io_out; // @[package.scala 96:25:@14354.4 package.scala 96:25:@14355.4]
  assign _T_2815 = _T_2775 ? Mem1D_5_io_output : _T_2814; // @[Mux.scala 31:69:@14445.4]
  assign _T_2772 = RetimeWrapper_84_io_out; // @[package.scala 96:25:@14346.4 package.scala 96:25:@14347.4]
  assign _T_2816 = _T_2772 ? Mem1D_4_io_output : _T_2815; // @[Mux.scala 31:69:@14446.4]
  assign _T_2769 = RetimeWrapper_83_io_out; // @[package.scala 96:25:@14338.4 package.scala 96:25:@14339.4]
  assign _T_2817 = _T_2769 ? Mem1D_3_io_output : _T_2816; // @[Mux.scala 31:69:@14447.4]
  assign _T_2766 = RetimeWrapper_82_io_out; // @[package.scala 96:25:@14330.4 package.scala 96:25:@14331.4]
  assign _T_2818 = _T_2766 ? Mem1D_2_io_output : _T_2817; // @[Mux.scala 31:69:@14448.4]
  assign _T_2763 = RetimeWrapper_81_io_out; // @[package.scala 96:25:@14322.4 package.scala 96:25:@14323.4]
  assign _T_2819 = _T_2763 ? Mem1D_1_io_output : _T_2818; // @[Mux.scala 31:69:@14449.4]
  assign _T_2760 = RetimeWrapper_80_io_out; // @[package.scala 96:25:@14314.4 package.scala 96:25:@14315.4]
  assign _T_2945 = RetimeWrapper_110_io_out; // @[package.scala 96:25:@14618.4 package.scala 96:25:@14619.4]
  assign _T_2949 = _T_2945 ? Mem1D_14_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@14628.4]
  assign _T_2942 = RetimeWrapper_109_io_out; // @[package.scala 96:25:@14610.4 package.scala 96:25:@14611.4]
  assign _T_2950 = _T_2942 ? Mem1D_13_io_output : _T_2949; // @[Mux.scala 31:69:@14629.4]
  assign _T_2939 = RetimeWrapper_108_io_out; // @[package.scala 96:25:@14602.4 package.scala 96:25:@14603.4]
  assign _T_2951 = _T_2939 ? Mem1D_12_io_output : _T_2950; // @[Mux.scala 31:69:@14630.4]
  assign _T_2936 = RetimeWrapper_107_io_out; // @[package.scala 96:25:@14594.4 package.scala 96:25:@14595.4]
  assign _T_2952 = _T_2936 ? Mem1D_11_io_output : _T_2951; // @[Mux.scala 31:69:@14631.4]
  assign _T_2933 = RetimeWrapper_106_io_out; // @[package.scala 96:25:@14586.4 package.scala 96:25:@14587.4]
  assign _T_2953 = _T_2933 ? Mem1D_10_io_output : _T_2952; // @[Mux.scala 31:69:@14632.4]
  assign _T_2930 = RetimeWrapper_105_io_out; // @[package.scala 96:25:@14578.4 package.scala 96:25:@14579.4]
  assign _T_2954 = _T_2930 ? Mem1D_9_io_output : _T_2953; // @[Mux.scala 31:69:@14633.4]
  assign _T_2927 = RetimeWrapper_104_io_out; // @[package.scala 96:25:@14570.4 package.scala 96:25:@14571.4]
  assign _T_2955 = _T_2927 ? Mem1D_8_io_output : _T_2954; // @[Mux.scala 31:69:@14634.4]
  assign _T_2924 = RetimeWrapper_103_io_out; // @[package.scala 96:25:@14562.4 package.scala 96:25:@14563.4]
  assign _T_2956 = _T_2924 ? Mem1D_7_io_output : _T_2955; // @[Mux.scala 31:69:@14635.4]
  assign _T_2921 = RetimeWrapper_102_io_out; // @[package.scala 96:25:@14554.4 package.scala 96:25:@14555.4]
  assign _T_2957 = _T_2921 ? Mem1D_6_io_output : _T_2956; // @[Mux.scala 31:69:@14636.4]
  assign _T_2918 = RetimeWrapper_101_io_out; // @[package.scala 96:25:@14546.4 package.scala 96:25:@14547.4]
  assign _T_2958 = _T_2918 ? Mem1D_5_io_output : _T_2957; // @[Mux.scala 31:69:@14637.4]
  assign _T_2915 = RetimeWrapper_100_io_out; // @[package.scala 96:25:@14538.4 package.scala 96:25:@14539.4]
  assign _T_2959 = _T_2915 ? Mem1D_4_io_output : _T_2958; // @[Mux.scala 31:69:@14638.4]
  assign _T_2912 = RetimeWrapper_99_io_out; // @[package.scala 96:25:@14530.4 package.scala 96:25:@14531.4]
  assign _T_2960 = _T_2912 ? Mem1D_3_io_output : _T_2959; // @[Mux.scala 31:69:@14639.4]
  assign _T_2909 = RetimeWrapper_98_io_out; // @[package.scala 96:25:@14522.4 package.scala 96:25:@14523.4]
  assign _T_2961 = _T_2909 ? Mem1D_2_io_output : _T_2960; // @[Mux.scala 31:69:@14640.4]
  assign _T_2906 = RetimeWrapper_97_io_out; // @[package.scala 96:25:@14514.4 package.scala 96:25:@14515.4]
  assign _T_2962 = _T_2906 ? Mem1D_1_io_output : _T_2961; // @[Mux.scala 31:69:@14641.4]
  assign _T_2903 = RetimeWrapper_96_io_out; // @[package.scala 96:25:@14506.4 package.scala 96:25:@14507.4]
  assign _T_3088 = RetimeWrapper_126_io_out; // @[package.scala 96:25:@14810.4 package.scala 96:25:@14811.4]
  assign _T_3092 = _T_3088 ? Mem1D_14_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@14820.4]
  assign _T_3085 = RetimeWrapper_125_io_out; // @[package.scala 96:25:@14802.4 package.scala 96:25:@14803.4]
  assign _T_3093 = _T_3085 ? Mem1D_13_io_output : _T_3092; // @[Mux.scala 31:69:@14821.4]
  assign _T_3082 = RetimeWrapper_124_io_out; // @[package.scala 96:25:@14794.4 package.scala 96:25:@14795.4]
  assign _T_3094 = _T_3082 ? Mem1D_12_io_output : _T_3093; // @[Mux.scala 31:69:@14822.4]
  assign _T_3079 = RetimeWrapper_123_io_out; // @[package.scala 96:25:@14786.4 package.scala 96:25:@14787.4]
  assign _T_3095 = _T_3079 ? Mem1D_11_io_output : _T_3094; // @[Mux.scala 31:69:@14823.4]
  assign _T_3076 = RetimeWrapper_122_io_out; // @[package.scala 96:25:@14778.4 package.scala 96:25:@14779.4]
  assign _T_3096 = _T_3076 ? Mem1D_10_io_output : _T_3095; // @[Mux.scala 31:69:@14824.4]
  assign _T_3073 = RetimeWrapper_121_io_out; // @[package.scala 96:25:@14770.4 package.scala 96:25:@14771.4]
  assign _T_3097 = _T_3073 ? Mem1D_9_io_output : _T_3096; // @[Mux.scala 31:69:@14825.4]
  assign _T_3070 = RetimeWrapper_120_io_out; // @[package.scala 96:25:@14762.4 package.scala 96:25:@14763.4]
  assign _T_3098 = _T_3070 ? Mem1D_8_io_output : _T_3097; // @[Mux.scala 31:69:@14826.4]
  assign _T_3067 = RetimeWrapper_119_io_out; // @[package.scala 96:25:@14754.4 package.scala 96:25:@14755.4]
  assign _T_3099 = _T_3067 ? Mem1D_7_io_output : _T_3098; // @[Mux.scala 31:69:@14827.4]
  assign _T_3064 = RetimeWrapper_118_io_out; // @[package.scala 96:25:@14746.4 package.scala 96:25:@14747.4]
  assign _T_3100 = _T_3064 ? Mem1D_6_io_output : _T_3099; // @[Mux.scala 31:69:@14828.4]
  assign _T_3061 = RetimeWrapper_117_io_out; // @[package.scala 96:25:@14738.4 package.scala 96:25:@14739.4]
  assign _T_3101 = _T_3061 ? Mem1D_5_io_output : _T_3100; // @[Mux.scala 31:69:@14829.4]
  assign _T_3058 = RetimeWrapper_116_io_out; // @[package.scala 96:25:@14730.4 package.scala 96:25:@14731.4]
  assign _T_3102 = _T_3058 ? Mem1D_4_io_output : _T_3101; // @[Mux.scala 31:69:@14830.4]
  assign _T_3055 = RetimeWrapper_115_io_out; // @[package.scala 96:25:@14722.4 package.scala 96:25:@14723.4]
  assign _T_3103 = _T_3055 ? Mem1D_3_io_output : _T_3102; // @[Mux.scala 31:69:@14831.4]
  assign _T_3052 = RetimeWrapper_114_io_out; // @[package.scala 96:25:@14714.4 package.scala 96:25:@14715.4]
  assign _T_3104 = _T_3052 ? Mem1D_2_io_output : _T_3103; // @[Mux.scala 31:69:@14832.4]
  assign _T_3049 = RetimeWrapper_113_io_out; // @[package.scala 96:25:@14706.4 package.scala 96:25:@14707.4]
  assign _T_3105 = _T_3049 ? Mem1D_1_io_output : _T_3104; // @[Mux.scala 31:69:@14833.4]
  assign _T_3046 = RetimeWrapper_112_io_out; // @[package.scala 96:25:@14698.4 package.scala 96:25:@14699.4]
  assign _T_3231 = RetimeWrapper_142_io_out; // @[package.scala 96:25:@15002.4 package.scala 96:25:@15003.4]
  assign _T_3235 = _T_3231 ? Mem1D_14_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@15012.4]
  assign _T_3228 = RetimeWrapper_141_io_out; // @[package.scala 96:25:@14994.4 package.scala 96:25:@14995.4]
  assign _T_3236 = _T_3228 ? Mem1D_13_io_output : _T_3235; // @[Mux.scala 31:69:@15013.4]
  assign _T_3225 = RetimeWrapper_140_io_out; // @[package.scala 96:25:@14986.4 package.scala 96:25:@14987.4]
  assign _T_3237 = _T_3225 ? Mem1D_12_io_output : _T_3236; // @[Mux.scala 31:69:@15014.4]
  assign _T_3222 = RetimeWrapper_139_io_out; // @[package.scala 96:25:@14978.4 package.scala 96:25:@14979.4]
  assign _T_3238 = _T_3222 ? Mem1D_11_io_output : _T_3237; // @[Mux.scala 31:69:@15015.4]
  assign _T_3219 = RetimeWrapper_138_io_out; // @[package.scala 96:25:@14970.4 package.scala 96:25:@14971.4]
  assign _T_3239 = _T_3219 ? Mem1D_10_io_output : _T_3238; // @[Mux.scala 31:69:@15016.4]
  assign _T_3216 = RetimeWrapper_137_io_out; // @[package.scala 96:25:@14962.4 package.scala 96:25:@14963.4]
  assign _T_3240 = _T_3216 ? Mem1D_9_io_output : _T_3239; // @[Mux.scala 31:69:@15017.4]
  assign _T_3213 = RetimeWrapper_136_io_out; // @[package.scala 96:25:@14954.4 package.scala 96:25:@14955.4]
  assign _T_3241 = _T_3213 ? Mem1D_8_io_output : _T_3240; // @[Mux.scala 31:69:@15018.4]
  assign _T_3210 = RetimeWrapper_135_io_out; // @[package.scala 96:25:@14946.4 package.scala 96:25:@14947.4]
  assign _T_3242 = _T_3210 ? Mem1D_7_io_output : _T_3241; // @[Mux.scala 31:69:@15019.4]
  assign _T_3207 = RetimeWrapper_134_io_out; // @[package.scala 96:25:@14938.4 package.scala 96:25:@14939.4]
  assign _T_3243 = _T_3207 ? Mem1D_6_io_output : _T_3242; // @[Mux.scala 31:69:@15020.4]
  assign _T_3204 = RetimeWrapper_133_io_out; // @[package.scala 96:25:@14930.4 package.scala 96:25:@14931.4]
  assign _T_3244 = _T_3204 ? Mem1D_5_io_output : _T_3243; // @[Mux.scala 31:69:@15021.4]
  assign _T_3201 = RetimeWrapper_132_io_out; // @[package.scala 96:25:@14922.4 package.scala 96:25:@14923.4]
  assign _T_3245 = _T_3201 ? Mem1D_4_io_output : _T_3244; // @[Mux.scala 31:69:@15022.4]
  assign _T_3198 = RetimeWrapper_131_io_out; // @[package.scala 96:25:@14914.4 package.scala 96:25:@14915.4]
  assign _T_3246 = _T_3198 ? Mem1D_3_io_output : _T_3245; // @[Mux.scala 31:69:@15023.4]
  assign _T_3195 = RetimeWrapper_130_io_out; // @[package.scala 96:25:@14906.4 package.scala 96:25:@14907.4]
  assign _T_3247 = _T_3195 ? Mem1D_2_io_output : _T_3246; // @[Mux.scala 31:69:@15024.4]
  assign _T_3192 = RetimeWrapper_129_io_out; // @[package.scala 96:25:@14898.4 package.scala 96:25:@14899.4]
  assign _T_3248 = _T_3192 ? Mem1D_1_io_output : _T_3247; // @[Mux.scala 31:69:@15025.4]
  assign _T_3189 = RetimeWrapper_128_io_out; // @[package.scala 96:25:@14890.4 package.scala 96:25:@14891.4]
  assign io_rPort_8_output_0 = _T_3189 ? Mem1D_io_output : _T_3248; // @[MemPrimitives.scala 148:13:@15027.4]
  assign io_rPort_7_output_0 = _T_3046 ? Mem1D_io_output : _T_3105; // @[MemPrimitives.scala 148:13:@14835.4]
  assign io_rPort_6_output_0 = _T_2903 ? Mem1D_io_output : _T_2962; // @[MemPrimitives.scala 148:13:@14643.4]
  assign io_rPort_5_output_0 = _T_2760 ? Mem1D_io_output : _T_2819; // @[MemPrimitives.scala 148:13:@14451.4]
  assign io_rPort_4_output_0 = _T_2617 ? Mem1D_io_output : _T_2676; // @[MemPrimitives.scala 148:13:@14259.4]
  assign io_rPort_3_output_0 = _T_2474 ? Mem1D_io_output : _T_2533; // @[MemPrimitives.scala 148:13:@14067.4]
  assign io_rPort_2_output_0 = _T_2331 ? Mem1D_io_output : _T_2390; // @[MemPrimitives.scala 148:13:@13875.4]
  assign io_rPort_1_output_0 = _T_2188 ? Mem1D_io_output : _T_2247; // @[MemPrimitives.scala 148:13:@13683.4]
  assign io_rPort_0_output_0 = _T_2045 ? Mem1D_io_output : _T_2104; // @[MemPrimitives.scala 148:13:@13491.4]
  assign Mem1D_clock = clock; // @[:@11429.4]
  assign Mem1D_reset = reset; // @[:@11430.4]
  assign Mem1D_io_r_ofs_0 = _T_579[0]; // @[MemPrimitives.scala 127:28:@11962.4]
  assign Mem1D_io_r_backpressure = _T_579[1]; // @[MemPrimitives.scala 128:32:@11963.4]
  assign Mem1D_io_w_ofs_0 = _T_322[0]; // @[MemPrimitives.scala 94:28:@11693.4]
  assign Mem1D_io_w_data_0 = _T_322[8:1]; // @[MemPrimitives.scala 95:29:@11694.4]
  assign Mem1D_io_w_en_0 = _T_322[9]; // @[MemPrimitives.scala 96:27:@11695.4]
  assign Mem1D_1_clock = clock; // @[:@11445.4]
  assign Mem1D_1_reset = reset; // @[:@11446.4]
  assign Mem1D_1_io_r_ofs_0 = _T_671[0]; // @[MemPrimitives.scala 127:28:@12051.4]
  assign Mem1D_1_io_r_backpressure = _T_671[1]; // @[MemPrimitives.scala 128:32:@12052.4]
  assign Mem1D_1_io_w_ofs_0 = _T_333[0]; // @[MemPrimitives.scala 94:28:@11705.4]
  assign Mem1D_1_io_w_data_0 = _T_333[8:1]; // @[MemPrimitives.scala 95:29:@11706.4]
  assign Mem1D_1_io_w_en_0 = _T_333[9]; // @[MemPrimitives.scala 96:27:@11707.4]
  assign Mem1D_2_clock = clock; // @[:@11461.4]
  assign Mem1D_2_reset = reset; // @[:@11462.4]
  assign Mem1D_2_io_r_ofs_0 = _T_763[0]; // @[MemPrimitives.scala 127:28:@12140.4]
  assign Mem1D_2_io_r_backpressure = _T_763[1]; // @[MemPrimitives.scala 128:32:@12141.4]
  assign Mem1D_2_io_w_ofs_0 = _T_344[0]; // @[MemPrimitives.scala 94:28:@11717.4]
  assign Mem1D_2_io_w_data_0 = _T_344[8:1]; // @[MemPrimitives.scala 95:29:@11718.4]
  assign Mem1D_2_io_w_en_0 = _T_344[9]; // @[MemPrimitives.scala 96:27:@11719.4]
  assign Mem1D_3_clock = clock; // @[:@11477.4]
  assign Mem1D_3_reset = reset; // @[:@11478.4]
  assign Mem1D_3_io_r_ofs_0 = _T_855[0]; // @[MemPrimitives.scala 127:28:@12229.4]
  assign Mem1D_3_io_r_backpressure = _T_855[1]; // @[MemPrimitives.scala 128:32:@12230.4]
  assign Mem1D_3_io_w_ofs_0 = _T_355[0]; // @[MemPrimitives.scala 94:28:@11729.4]
  assign Mem1D_3_io_w_data_0 = _T_355[8:1]; // @[MemPrimitives.scala 95:29:@11730.4]
  assign Mem1D_3_io_w_en_0 = _T_355[9]; // @[MemPrimitives.scala 96:27:@11731.4]
  assign Mem1D_4_clock = clock; // @[:@11493.4]
  assign Mem1D_4_reset = reset; // @[:@11494.4]
  assign Mem1D_4_io_r_ofs_0 = _T_947[0]; // @[MemPrimitives.scala 127:28:@12318.4]
  assign Mem1D_4_io_r_backpressure = _T_947[1]; // @[MemPrimitives.scala 128:32:@12319.4]
  assign Mem1D_4_io_w_ofs_0 = _T_366[0]; // @[MemPrimitives.scala 94:28:@11741.4]
  assign Mem1D_4_io_w_data_0 = _T_366[8:1]; // @[MemPrimitives.scala 95:29:@11742.4]
  assign Mem1D_4_io_w_en_0 = _T_366[9]; // @[MemPrimitives.scala 96:27:@11743.4]
  assign Mem1D_5_clock = clock; // @[:@11509.4]
  assign Mem1D_5_reset = reset; // @[:@11510.4]
  assign Mem1D_5_io_r_ofs_0 = _T_1039[0]; // @[MemPrimitives.scala 127:28:@12407.4]
  assign Mem1D_5_io_r_backpressure = _T_1039[1]; // @[MemPrimitives.scala 128:32:@12408.4]
  assign Mem1D_5_io_w_ofs_0 = _T_377[0]; // @[MemPrimitives.scala 94:28:@11753.4]
  assign Mem1D_5_io_w_data_0 = _T_377[8:1]; // @[MemPrimitives.scala 95:29:@11754.4]
  assign Mem1D_5_io_w_en_0 = _T_377[9]; // @[MemPrimitives.scala 96:27:@11755.4]
  assign Mem1D_6_clock = clock; // @[:@11525.4]
  assign Mem1D_6_reset = reset; // @[:@11526.4]
  assign Mem1D_6_io_r_ofs_0 = _T_1131[0]; // @[MemPrimitives.scala 127:28:@12496.4]
  assign Mem1D_6_io_r_backpressure = _T_1131[1]; // @[MemPrimitives.scala 128:32:@12497.4]
  assign Mem1D_6_io_w_ofs_0 = _T_388[0]; // @[MemPrimitives.scala 94:28:@11765.4]
  assign Mem1D_6_io_w_data_0 = _T_388[8:1]; // @[MemPrimitives.scala 95:29:@11766.4]
  assign Mem1D_6_io_w_en_0 = _T_388[9]; // @[MemPrimitives.scala 96:27:@11767.4]
  assign Mem1D_7_clock = clock; // @[:@11541.4]
  assign Mem1D_7_reset = reset; // @[:@11542.4]
  assign Mem1D_7_io_r_ofs_0 = _T_1223[0]; // @[MemPrimitives.scala 127:28:@12585.4]
  assign Mem1D_7_io_r_backpressure = _T_1223[1]; // @[MemPrimitives.scala 128:32:@12586.4]
  assign Mem1D_7_io_w_ofs_0 = _T_399[0]; // @[MemPrimitives.scala 94:28:@11777.4]
  assign Mem1D_7_io_w_data_0 = _T_399[8:1]; // @[MemPrimitives.scala 95:29:@11778.4]
  assign Mem1D_7_io_w_en_0 = _T_399[9]; // @[MemPrimitives.scala 96:27:@11779.4]
  assign Mem1D_8_clock = clock; // @[:@11557.4]
  assign Mem1D_8_reset = reset; // @[:@11558.4]
  assign Mem1D_8_io_r_ofs_0 = _T_1315[0]; // @[MemPrimitives.scala 127:28:@12674.4]
  assign Mem1D_8_io_r_backpressure = _T_1315[1]; // @[MemPrimitives.scala 128:32:@12675.4]
  assign Mem1D_8_io_w_ofs_0 = _T_410[0]; // @[MemPrimitives.scala 94:28:@11789.4]
  assign Mem1D_8_io_w_data_0 = _T_410[8:1]; // @[MemPrimitives.scala 95:29:@11790.4]
  assign Mem1D_8_io_w_en_0 = _T_410[9]; // @[MemPrimitives.scala 96:27:@11791.4]
  assign Mem1D_9_clock = clock; // @[:@11573.4]
  assign Mem1D_9_reset = reset; // @[:@11574.4]
  assign Mem1D_9_io_r_ofs_0 = _T_1407[0]; // @[MemPrimitives.scala 127:28:@12763.4]
  assign Mem1D_9_io_r_backpressure = _T_1407[1]; // @[MemPrimitives.scala 128:32:@12764.4]
  assign Mem1D_9_io_w_ofs_0 = _T_421[0]; // @[MemPrimitives.scala 94:28:@11801.4]
  assign Mem1D_9_io_w_data_0 = _T_421[8:1]; // @[MemPrimitives.scala 95:29:@11802.4]
  assign Mem1D_9_io_w_en_0 = _T_421[9]; // @[MemPrimitives.scala 96:27:@11803.4]
  assign Mem1D_10_clock = clock; // @[:@11589.4]
  assign Mem1D_10_reset = reset; // @[:@11590.4]
  assign Mem1D_10_io_r_ofs_0 = _T_1499[0]; // @[MemPrimitives.scala 127:28:@12852.4]
  assign Mem1D_10_io_r_backpressure = _T_1499[1]; // @[MemPrimitives.scala 128:32:@12853.4]
  assign Mem1D_10_io_w_ofs_0 = _T_432[0]; // @[MemPrimitives.scala 94:28:@11813.4]
  assign Mem1D_10_io_w_data_0 = _T_432[8:1]; // @[MemPrimitives.scala 95:29:@11814.4]
  assign Mem1D_10_io_w_en_0 = _T_432[9]; // @[MemPrimitives.scala 96:27:@11815.4]
  assign Mem1D_11_clock = clock; // @[:@11605.4]
  assign Mem1D_11_reset = reset; // @[:@11606.4]
  assign Mem1D_11_io_r_ofs_0 = _T_1591[0]; // @[MemPrimitives.scala 127:28:@12941.4]
  assign Mem1D_11_io_r_backpressure = _T_1591[1]; // @[MemPrimitives.scala 128:32:@12942.4]
  assign Mem1D_11_io_w_ofs_0 = _T_443[0]; // @[MemPrimitives.scala 94:28:@11825.4]
  assign Mem1D_11_io_w_data_0 = _T_443[8:1]; // @[MemPrimitives.scala 95:29:@11826.4]
  assign Mem1D_11_io_w_en_0 = _T_443[9]; // @[MemPrimitives.scala 96:27:@11827.4]
  assign Mem1D_12_clock = clock; // @[:@11621.4]
  assign Mem1D_12_reset = reset; // @[:@11622.4]
  assign Mem1D_12_io_r_ofs_0 = _T_1683[0]; // @[MemPrimitives.scala 127:28:@13030.4]
  assign Mem1D_12_io_r_backpressure = _T_1683[1]; // @[MemPrimitives.scala 128:32:@13031.4]
  assign Mem1D_12_io_w_ofs_0 = _T_454[0]; // @[MemPrimitives.scala 94:28:@11837.4]
  assign Mem1D_12_io_w_data_0 = _T_454[8:1]; // @[MemPrimitives.scala 95:29:@11838.4]
  assign Mem1D_12_io_w_en_0 = _T_454[9]; // @[MemPrimitives.scala 96:27:@11839.4]
  assign Mem1D_13_clock = clock; // @[:@11637.4]
  assign Mem1D_13_reset = reset; // @[:@11638.4]
  assign Mem1D_13_io_r_ofs_0 = _T_1775[0]; // @[MemPrimitives.scala 127:28:@13119.4]
  assign Mem1D_13_io_r_backpressure = _T_1775[1]; // @[MemPrimitives.scala 128:32:@13120.4]
  assign Mem1D_13_io_w_ofs_0 = _T_465[0]; // @[MemPrimitives.scala 94:28:@11849.4]
  assign Mem1D_13_io_w_data_0 = _T_465[8:1]; // @[MemPrimitives.scala 95:29:@11850.4]
  assign Mem1D_13_io_w_en_0 = _T_465[9]; // @[MemPrimitives.scala 96:27:@11851.4]
  assign Mem1D_14_clock = clock; // @[:@11653.4]
  assign Mem1D_14_reset = reset; // @[:@11654.4]
  assign Mem1D_14_io_r_ofs_0 = _T_1867[0]; // @[MemPrimitives.scala 127:28:@13208.4]
  assign Mem1D_14_io_r_backpressure = _T_1867[1]; // @[MemPrimitives.scala 128:32:@13209.4]
  assign Mem1D_14_io_w_ofs_0 = _T_476[0]; // @[MemPrimitives.scala 94:28:@11861.4]
  assign Mem1D_14_io_w_data_0 = _T_476[8:1]; // @[MemPrimitives.scala 95:29:@11862.4]
  assign Mem1D_14_io_w_en_0 = _T_476[9]; // @[MemPrimitives.scala 96:27:@11863.4]
  assign Mem1D_15_clock = clock; // @[:@11669.4]
  assign Mem1D_15_reset = reset; // @[:@11670.4]
  assign Mem1D_15_io_r_ofs_0 = _T_1959[0]; // @[MemPrimitives.scala 127:28:@13297.4]
  assign Mem1D_15_io_r_backpressure = _T_1959[1]; // @[MemPrimitives.scala 128:32:@13298.4]
  assign Mem1D_15_io_w_ofs_0 = _T_487[0]; // @[MemPrimitives.scala 94:28:@11873.4]
  assign Mem1D_15_io_w_data_0 = _T_487[8:1]; // @[MemPrimitives.scala 95:29:@11874.4]
  assign Mem1D_15_io_w_en_0 = _T_487[9]; // @[MemPrimitives.scala 96:27:@11875.4]
  assign StickySelects_clock = clock; // @[:@11913.4]
  assign StickySelects_reset = reset; // @[:@11914.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0 & _T_495; // @[MemPrimitives.scala 122:60:@11915.4]
  assign StickySelects_io_ins_1 = io_rPort_1_en_0 & _T_501; // @[MemPrimitives.scala 122:60:@11916.4]
  assign StickySelects_io_ins_2 = io_rPort_2_en_0 & _T_507; // @[MemPrimitives.scala 122:60:@11917.4]
  assign StickySelects_io_ins_3 = io_rPort_3_en_0 & _T_513; // @[MemPrimitives.scala 122:60:@11918.4]
  assign StickySelects_io_ins_4 = io_rPort_4_en_0 & _T_519; // @[MemPrimitives.scala 122:60:@11919.4]
  assign StickySelects_io_ins_5 = io_rPort_5_en_0 & _T_525; // @[MemPrimitives.scala 122:60:@11920.4]
  assign StickySelects_io_ins_6 = io_rPort_6_en_0 & _T_531; // @[MemPrimitives.scala 122:60:@11921.4]
  assign StickySelects_io_ins_7 = io_rPort_7_en_0 & _T_537; // @[MemPrimitives.scala 122:60:@11922.4]
  assign StickySelects_io_ins_8 = io_rPort_8_en_0 & _T_543; // @[MemPrimitives.scala 122:60:@11923.4]
  assign StickySelects_1_clock = clock; // @[:@12002.4]
  assign StickySelects_1_reset = reset; // @[:@12003.4]
  assign StickySelects_1_io_ins_0 = io_rPort_0_en_0 & _T_587; // @[MemPrimitives.scala 122:60:@12004.4]
  assign StickySelects_1_io_ins_1 = io_rPort_1_en_0 & _T_593; // @[MemPrimitives.scala 122:60:@12005.4]
  assign StickySelects_1_io_ins_2 = io_rPort_2_en_0 & _T_599; // @[MemPrimitives.scala 122:60:@12006.4]
  assign StickySelects_1_io_ins_3 = io_rPort_3_en_0 & _T_605; // @[MemPrimitives.scala 122:60:@12007.4]
  assign StickySelects_1_io_ins_4 = io_rPort_4_en_0 & _T_611; // @[MemPrimitives.scala 122:60:@12008.4]
  assign StickySelects_1_io_ins_5 = io_rPort_5_en_0 & _T_617; // @[MemPrimitives.scala 122:60:@12009.4]
  assign StickySelects_1_io_ins_6 = io_rPort_6_en_0 & _T_623; // @[MemPrimitives.scala 122:60:@12010.4]
  assign StickySelects_1_io_ins_7 = io_rPort_7_en_0 & _T_629; // @[MemPrimitives.scala 122:60:@12011.4]
  assign StickySelects_1_io_ins_8 = io_rPort_8_en_0 & _T_635; // @[MemPrimitives.scala 122:60:@12012.4]
  assign StickySelects_2_clock = clock; // @[:@12091.4]
  assign StickySelects_2_reset = reset; // @[:@12092.4]
  assign StickySelects_2_io_ins_0 = io_rPort_0_en_0 & _T_679; // @[MemPrimitives.scala 122:60:@12093.4]
  assign StickySelects_2_io_ins_1 = io_rPort_1_en_0 & _T_685; // @[MemPrimitives.scala 122:60:@12094.4]
  assign StickySelects_2_io_ins_2 = io_rPort_2_en_0 & _T_691; // @[MemPrimitives.scala 122:60:@12095.4]
  assign StickySelects_2_io_ins_3 = io_rPort_3_en_0 & _T_697; // @[MemPrimitives.scala 122:60:@12096.4]
  assign StickySelects_2_io_ins_4 = io_rPort_4_en_0 & _T_703; // @[MemPrimitives.scala 122:60:@12097.4]
  assign StickySelects_2_io_ins_5 = io_rPort_5_en_0 & _T_709; // @[MemPrimitives.scala 122:60:@12098.4]
  assign StickySelects_2_io_ins_6 = io_rPort_6_en_0 & _T_715; // @[MemPrimitives.scala 122:60:@12099.4]
  assign StickySelects_2_io_ins_7 = io_rPort_7_en_0 & _T_721; // @[MemPrimitives.scala 122:60:@12100.4]
  assign StickySelects_2_io_ins_8 = io_rPort_8_en_0 & _T_727; // @[MemPrimitives.scala 122:60:@12101.4]
  assign StickySelects_3_clock = clock; // @[:@12180.4]
  assign StickySelects_3_reset = reset; // @[:@12181.4]
  assign StickySelects_3_io_ins_0 = io_rPort_0_en_0 & _T_771; // @[MemPrimitives.scala 122:60:@12182.4]
  assign StickySelects_3_io_ins_1 = io_rPort_1_en_0 & _T_777; // @[MemPrimitives.scala 122:60:@12183.4]
  assign StickySelects_3_io_ins_2 = io_rPort_2_en_0 & _T_783; // @[MemPrimitives.scala 122:60:@12184.4]
  assign StickySelects_3_io_ins_3 = io_rPort_3_en_0 & _T_789; // @[MemPrimitives.scala 122:60:@12185.4]
  assign StickySelects_3_io_ins_4 = io_rPort_4_en_0 & _T_795; // @[MemPrimitives.scala 122:60:@12186.4]
  assign StickySelects_3_io_ins_5 = io_rPort_5_en_0 & _T_801; // @[MemPrimitives.scala 122:60:@12187.4]
  assign StickySelects_3_io_ins_6 = io_rPort_6_en_0 & _T_807; // @[MemPrimitives.scala 122:60:@12188.4]
  assign StickySelects_3_io_ins_7 = io_rPort_7_en_0 & _T_813; // @[MemPrimitives.scala 122:60:@12189.4]
  assign StickySelects_3_io_ins_8 = io_rPort_8_en_0 & _T_819; // @[MemPrimitives.scala 122:60:@12190.4]
  assign StickySelects_4_clock = clock; // @[:@12269.4]
  assign StickySelects_4_reset = reset; // @[:@12270.4]
  assign StickySelects_4_io_ins_0 = io_rPort_0_en_0 & _T_863; // @[MemPrimitives.scala 122:60:@12271.4]
  assign StickySelects_4_io_ins_1 = io_rPort_1_en_0 & _T_869; // @[MemPrimitives.scala 122:60:@12272.4]
  assign StickySelects_4_io_ins_2 = io_rPort_2_en_0 & _T_875; // @[MemPrimitives.scala 122:60:@12273.4]
  assign StickySelects_4_io_ins_3 = io_rPort_3_en_0 & _T_881; // @[MemPrimitives.scala 122:60:@12274.4]
  assign StickySelects_4_io_ins_4 = io_rPort_4_en_0 & _T_887; // @[MemPrimitives.scala 122:60:@12275.4]
  assign StickySelects_4_io_ins_5 = io_rPort_5_en_0 & _T_893; // @[MemPrimitives.scala 122:60:@12276.4]
  assign StickySelects_4_io_ins_6 = io_rPort_6_en_0 & _T_899; // @[MemPrimitives.scala 122:60:@12277.4]
  assign StickySelects_4_io_ins_7 = io_rPort_7_en_0 & _T_905; // @[MemPrimitives.scala 122:60:@12278.4]
  assign StickySelects_4_io_ins_8 = io_rPort_8_en_0 & _T_911; // @[MemPrimitives.scala 122:60:@12279.4]
  assign StickySelects_5_clock = clock; // @[:@12358.4]
  assign StickySelects_5_reset = reset; // @[:@12359.4]
  assign StickySelects_5_io_ins_0 = io_rPort_0_en_0 & _T_955; // @[MemPrimitives.scala 122:60:@12360.4]
  assign StickySelects_5_io_ins_1 = io_rPort_1_en_0 & _T_961; // @[MemPrimitives.scala 122:60:@12361.4]
  assign StickySelects_5_io_ins_2 = io_rPort_2_en_0 & _T_967; // @[MemPrimitives.scala 122:60:@12362.4]
  assign StickySelects_5_io_ins_3 = io_rPort_3_en_0 & _T_973; // @[MemPrimitives.scala 122:60:@12363.4]
  assign StickySelects_5_io_ins_4 = io_rPort_4_en_0 & _T_979; // @[MemPrimitives.scala 122:60:@12364.4]
  assign StickySelects_5_io_ins_5 = io_rPort_5_en_0 & _T_985; // @[MemPrimitives.scala 122:60:@12365.4]
  assign StickySelects_5_io_ins_6 = io_rPort_6_en_0 & _T_991; // @[MemPrimitives.scala 122:60:@12366.4]
  assign StickySelects_5_io_ins_7 = io_rPort_7_en_0 & _T_997; // @[MemPrimitives.scala 122:60:@12367.4]
  assign StickySelects_5_io_ins_8 = io_rPort_8_en_0 & _T_1003; // @[MemPrimitives.scala 122:60:@12368.4]
  assign StickySelects_6_clock = clock; // @[:@12447.4]
  assign StickySelects_6_reset = reset; // @[:@12448.4]
  assign StickySelects_6_io_ins_0 = io_rPort_0_en_0 & _T_1047; // @[MemPrimitives.scala 122:60:@12449.4]
  assign StickySelects_6_io_ins_1 = io_rPort_1_en_0 & _T_1053; // @[MemPrimitives.scala 122:60:@12450.4]
  assign StickySelects_6_io_ins_2 = io_rPort_2_en_0 & _T_1059; // @[MemPrimitives.scala 122:60:@12451.4]
  assign StickySelects_6_io_ins_3 = io_rPort_3_en_0 & _T_1065; // @[MemPrimitives.scala 122:60:@12452.4]
  assign StickySelects_6_io_ins_4 = io_rPort_4_en_0 & _T_1071; // @[MemPrimitives.scala 122:60:@12453.4]
  assign StickySelects_6_io_ins_5 = io_rPort_5_en_0 & _T_1077; // @[MemPrimitives.scala 122:60:@12454.4]
  assign StickySelects_6_io_ins_6 = io_rPort_6_en_0 & _T_1083; // @[MemPrimitives.scala 122:60:@12455.4]
  assign StickySelects_6_io_ins_7 = io_rPort_7_en_0 & _T_1089; // @[MemPrimitives.scala 122:60:@12456.4]
  assign StickySelects_6_io_ins_8 = io_rPort_8_en_0 & _T_1095; // @[MemPrimitives.scala 122:60:@12457.4]
  assign StickySelects_7_clock = clock; // @[:@12536.4]
  assign StickySelects_7_reset = reset; // @[:@12537.4]
  assign StickySelects_7_io_ins_0 = io_rPort_0_en_0 & _T_1139; // @[MemPrimitives.scala 122:60:@12538.4]
  assign StickySelects_7_io_ins_1 = io_rPort_1_en_0 & _T_1145; // @[MemPrimitives.scala 122:60:@12539.4]
  assign StickySelects_7_io_ins_2 = io_rPort_2_en_0 & _T_1151; // @[MemPrimitives.scala 122:60:@12540.4]
  assign StickySelects_7_io_ins_3 = io_rPort_3_en_0 & _T_1157; // @[MemPrimitives.scala 122:60:@12541.4]
  assign StickySelects_7_io_ins_4 = io_rPort_4_en_0 & _T_1163; // @[MemPrimitives.scala 122:60:@12542.4]
  assign StickySelects_7_io_ins_5 = io_rPort_5_en_0 & _T_1169; // @[MemPrimitives.scala 122:60:@12543.4]
  assign StickySelects_7_io_ins_6 = io_rPort_6_en_0 & _T_1175; // @[MemPrimitives.scala 122:60:@12544.4]
  assign StickySelects_7_io_ins_7 = io_rPort_7_en_0 & _T_1181; // @[MemPrimitives.scala 122:60:@12545.4]
  assign StickySelects_7_io_ins_8 = io_rPort_8_en_0 & _T_1187; // @[MemPrimitives.scala 122:60:@12546.4]
  assign StickySelects_8_clock = clock; // @[:@12625.4]
  assign StickySelects_8_reset = reset; // @[:@12626.4]
  assign StickySelects_8_io_ins_0 = io_rPort_0_en_0 & _T_1231; // @[MemPrimitives.scala 122:60:@12627.4]
  assign StickySelects_8_io_ins_1 = io_rPort_1_en_0 & _T_1237; // @[MemPrimitives.scala 122:60:@12628.4]
  assign StickySelects_8_io_ins_2 = io_rPort_2_en_0 & _T_1243; // @[MemPrimitives.scala 122:60:@12629.4]
  assign StickySelects_8_io_ins_3 = io_rPort_3_en_0 & _T_1249; // @[MemPrimitives.scala 122:60:@12630.4]
  assign StickySelects_8_io_ins_4 = io_rPort_4_en_0 & _T_1255; // @[MemPrimitives.scala 122:60:@12631.4]
  assign StickySelects_8_io_ins_5 = io_rPort_5_en_0 & _T_1261; // @[MemPrimitives.scala 122:60:@12632.4]
  assign StickySelects_8_io_ins_6 = io_rPort_6_en_0 & _T_1267; // @[MemPrimitives.scala 122:60:@12633.4]
  assign StickySelects_8_io_ins_7 = io_rPort_7_en_0 & _T_1273; // @[MemPrimitives.scala 122:60:@12634.4]
  assign StickySelects_8_io_ins_8 = io_rPort_8_en_0 & _T_1279; // @[MemPrimitives.scala 122:60:@12635.4]
  assign StickySelects_9_clock = clock; // @[:@12714.4]
  assign StickySelects_9_reset = reset; // @[:@12715.4]
  assign StickySelects_9_io_ins_0 = io_rPort_0_en_0 & _T_1323; // @[MemPrimitives.scala 122:60:@12716.4]
  assign StickySelects_9_io_ins_1 = io_rPort_1_en_0 & _T_1329; // @[MemPrimitives.scala 122:60:@12717.4]
  assign StickySelects_9_io_ins_2 = io_rPort_2_en_0 & _T_1335; // @[MemPrimitives.scala 122:60:@12718.4]
  assign StickySelects_9_io_ins_3 = io_rPort_3_en_0 & _T_1341; // @[MemPrimitives.scala 122:60:@12719.4]
  assign StickySelects_9_io_ins_4 = io_rPort_4_en_0 & _T_1347; // @[MemPrimitives.scala 122:60:@12720.4]
  assign StickySelects_9_io_ins_5 = io_rPort_5_en_0 & _T_1353; // @[MemPrimitives.scala 122:60:@12721.4]
  assign StickySelects_9_io_ins_6 = io_rPort_6_en_0 & _T_1359; // @[MemPrimitives.scala 122:60:@12722.4]
  assign StickySelects_9_io_ins_7 = io_rPort_7_en_0 & _T_1365; // @[MemPrimitives.scala 122:60:@12723.4]
  assign StickySelects_9_io_ins_8 = io_rPort_8_en_0 & _T_1371; // @[MemPrimitives.scala 122:60:@12724.4]
  assign StickySelects_10_clock = clock; // @[:@12803.4]
  assign StickySelects_10_reset = reset; // @[:@12804.4]
  assign StickySelects_10_io_ins_0 = io_rPort_0_en_0 & _T_1415; // @[MemPrimitives.scala 122:60:@12805.4]
  assign StickySelects_10_io_ins_1 = io_rPort_1_en_0 & _T_1421; // @[MemPrimitives.scala 122:60:@12806.4]
  assign StickySelects_10_io_ins_2 = io_rPort_2_en_0 & _T_1427; // @[MemPrimitives.scala 122:60:@12807.4]
  assign StickySelects_10_io_ins_3 = io_rPort_3_en_0 & _T_1433; // @[MemPrimitives.scala 122:60:@12808.4]
  assign StickySelects_10_io_ins_4 = io_rPort_4_en_0 & _T_1439; // @[MemPrimitives.scala 122:60:@12809.4]
  assign StickySelects_10_io_ins_5 = io_rPort_5_en_0 & _T_1445; // @[MemPrimitives.scala 122:60:@12810.4]
  assign StickySelects_10_io_ins_6 = io_rPort_6_en_0 & _T_1451; // @[MemPrimitives.scala 122:60:@12811.4]
  assign StickySelects_10_io_ins_7 = io_rPort_7_en_0 & _T_1457; // @[MemPrimitives.scala 122:60:@12812.4]
  assign StickySelects_10_io_ins_8 = io_rPort_8_en_0 & _T_1463; // @[MemPrimitives.scala 122:60:@12813.4]
  assign StickySelects_11_clock = clock; // @[:@12892.4]
  assign StickySelects_11_reset = reset; // @[:@12893.4]
  assign StickySelects_11_io_ins_0 = io_rPort_0_en_0 & _T_1507; // @[MemPrimitives.scala 122:60:@12894.4]
  assign StickySelects_11_io_ins_1 = io_rPort_1_en_0 & _T_1513; // @[MemPrimitives.scala 122:60:@12895.4]
  assign StickySelects_11_io_ins_2 = io_rPort_2_en_0 & _T_1519; // @[MemPrimitives.scala 122:60:@12896.4]
  assign StickySelects_11_io_ins_3 = io_rPort_3_en_0 & _T_1525; // @[MemPrimitives.scala 122:60:@12897.4]
  assign StickySelects_11_io_ins_4 = io_rPort_4_en_0 & _T_1531; // @[MemPrimitives.scala 122:60:@12898.4]
  assign StickySelects_11_io_ins_5 = io_rPort_5_en_0 & _T_1537; // @[MemPrimitives.scala 122:60:@12899.4]
  assign StickySelects_11_io_ins_6 = io_rPort_6_en_0 & _T_1543; // @[MemPrimitives.scala 122:60:@12900.4]
  assign StickySelects_11_io_ins_7 = io_rPort_7_en_0 & _T_1549; // @[MemPrimitives.scala 122:60:@12901.4]
  assign StickySelects_11_io_ins_8 = io_rPort_8_en_0 & _T_1555; // @[MemPrimitives.scala 122:60:@12902.4]
  assign StickySelects_12_clock = clock; // @[:@12981.4]
  assign StickySelects_12_reset = reset; // @[:@12982.4]
  assign StickySelects_12_io_ins_0 = io_rPort_0_en_0 & _T_1599; // @[MemPrimitives.scala 122:60:@12983.4]
  assign StickySelects_12_io_ins_1 = io_rPort_1_en_0 & _T_1605; // @[MemPrimitives.scala 122:60:@12984.4]
  assign StickySelects_12_io_ins_2 = io_rPort_2_en_0 & _T_1611; // @[MemPrimitives.scala 122:60:@12985.4]
  assign StickySelects_12_io_ins_3 = io_rPort_3_en_0 & _T_1617; // @[MemPrimitives.scala 122:60:@12986.4]
  assign StickySelects_12_io_ins_4 = io_rPort_4_en_0 & _T_1623; // @[MemPrimitives.scala 122:60:@12987.4]
  assign StickySelects_12_io_ins_5 = io_rPort_5_en_0 & _T_1629; // @[MemPrimitives.scala 122:60:@12988.4]
  assign StickySelects_12_io_ins_6 = io_rPort_6_en_0 & _T_1635; // @[MemPrimitives.scala 122:60:@12989.4]
  assign StickySelects_12_io_ins_7 = io_rPort_7_en_0 & _T_1641; // @[MemPrimitives.scala 122:60:@12990.4]
  assign StickySelects_12_io_ins_8 = io_rPort_8_en_0 & _T_1647; // @[MemPrimitives.scala 122:60:@12991.4]
  assign StickySelects_13_clock = clock; // @[:@13070.4]
  assign StickySelects_13_reset = reset; // @[:@13071.4]
  assign StickySelects_13_io_ins_0 = io_rPort_0_en_0 & _T_1691; // @[MemPrimitives.scala 122:60:@13072.4]
  assign StickySelects_13_io_ins_1 = io_rPort_1_en_0 & _T_1697; // @[MemPrimitives.scala 122:60:@13073.4]
  assign StickySelects_13_io_ins_2 = io_rPort_2_en_0 & _T_1703; // @[MemPrimitives.scala 122:60:@13074.4]
  assign StickySelects_13_io_ins_3 = io_rPort_3_en_0 & _T_1709; // @[MemPrimitives.scala 122:60:@13075.4]
  assign StickySelects_13_io_ins_4 = io_rPort_4_en_0 & _T_1715; // @[MemPrimitives.scala 122:60:@13076.4]
  assign StickySelects_13_io_ins_5 = io_rPort_5_en_0 & _T_1721; // @[MemPrimitives.scala 122:60:@13077.4]
  assign StickySelects_13_io_ins_6 = io_rPort_6_en_0 & _T_1727; // @[MemPrimitives.scala 122:60:@13078.4]
  assign StickySelects_13_io_ins_7 = io_rPort_7_en_0 & _T_1733; // @[MemPrimitives.scala 122:60:@13079.4]
  assign StickySelects_13_io_ins_8 = io_rPort_8_en_0 & _T_1739; // @[MemPrimitives.scala 122:60:@13080.4]
  assign StickySelects_14_clock = clock; // @[:@13159.4]
  assign StickySelects_14_reset = reset; // @[:@13160.4]
  assign StickySelects_14_io_ins_0 = io_rPort_0_en_0 & _T_1783; // @[MemPrimitives.scala 122:60:@13161.4]
  assign StickySelects_14_io_ins_1 = io_rPort_1_en_0 & _T_1789; // @[MemPrimitives.scala 122:60:@13162.4]
  assign StickySelects_14_io_ins_2 = io_rPort_2_en_0 & _T_1795; // @[MemPrimitives.scala 122:60:@13163.4]
  assign StickySelects_14_io_ins_3 = io_rPort_3_en_0 & _T_1801; // @[MemPrimitives.scala 122:60:@13164.4]
  assign StickySelects_14_io_ins_4 = io_rPort_4_en_0 & _T_1807; // @[MemPrimitives.scala 122:60:@13165.4]
  assign StickySelects_14_io_ins_5 = io_rPort_5_en_0 & _T_1813; // @[MemPrimitives.scala 122:60:@13166.4]
  assign StickySelects_14_io_ins_6 = io_rPort_6_en_0 & _T_1819; // @[MemPrimitives.scala 122:60:@13167.4]
  assign StickySelects_14_io_ins_7 = io_rPort_7_en_0 & _T_1825; // @[MemPrimitives.scala 122:60:@13168.4]
  assign StickySelects_14_io_ins_8 = io_rPort_8_en_0 & _T_1831; // @[MemPrimitives.scala 122:60:@13169.4]
  assign StickySelects_15_clock = clock; // @[:@13248.4]
  assign StickySelects_15_reset = reset; // @[:@13249.4]
  assign StickySelects_15_io_ins_0 = io_rPort_0_en_0 & _T_1875; // @[MemPrimitives.scala 122:60:@13250.4]
  assign StickySelects_15_io_ins_1 = io_rPort_1_en_0 & _T_1881; // @[MemPrimitives.scala 122:60:@13251.4]
  assign StickySelects_15_io_ins_2 = io_rPort_2_en_0 & _T_1887; // @[MemPrimitives.scala 122:60:@13252.4]
  assign StickySelects_15_io_ins_3 = io_rPort_3_en_0 & _T_1893; // @[MemPrimitives.scala 122:60:@13253.4]
  assign StickySelects_15_io_ins_4 = io_rPort_4_en_0 & _T_1899; // @[MemPrimitives.scala 122:60:@13254.4]
  assign StickySelects_15_io_ins_5 = io_rPort_5_en_0 & _T_1905; // @[MemPrimitives.scala 122:60:@13255.4]
  assign StickySelects_15_io_ins_6 = io_rPort_6_en_0 & _T_1911; // @[MemPrimitives.scala 122:60:@13256.4]
  assign StickySelects_15_io_ins_7 = io_rPort_7_en_0 & _T_1917; // @[MemPrimitives.scala 122:60:@13257.4]
  assign StickySelects_15_io_ins_8 = io_rPort_8_en_0 & _T_1923; // @[MemPrimitives.scala 122:60:@13258.4]
  assign RetimeWrapper_clock = clock; // @[:@13350.4]
  assign RetimeWrapper_reset = reset; // @[:@13351.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13353.4]
  assign RetimeWrapper_io_in = _T_495 & io_rPort_0_en_0; // @[package.scala 94:16:@13352.4]
  assign RetimeWrapper_1_clock = clock; // @[:@13358.4]
  assign RetimeWrapper_1_reset = reset; // @[:@13359.4]
  assign RetimeWrapper_1_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13361.4]
  assign RetimeWrapper_1_io_in = _T_587 & io_rPort_0_en_0; // @[package.scala 94:16:@13360.4]
  assign RetimeWrapper_2_clock = clock; // @[:@13366.4]
  assign RetimeWrapper_2_reset = reset; // @[:@13367.4]
  assign RetimeWrapper_2_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13369.4]
  assign RetimeWrapper_2_io_in = _T_679 & io_rPort_0_en_0; // @[package.scala 94:16:@13368.4]
  assign RetimeWrapper_3_clock = clock; // @[:@13374.4]
  assign RetimeWrapper_3_reset = reset; // @[:@13375.4]
  assign RetimeWrapper_3_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13377.4]
  assign RetimeWrapper_3_io_in = _T_771 & io_rPort_0_en_0; // @[package.scala 94:16:@13376.4]
  assign RetimeWrapper_4_clock = clock; // @[:@13382.4]
  assign RetimeWrapper_4_reset = reset; // @[:@13383.4]
  assign RetimeWrapper_4_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13385.4]
  assign RetimeWrapper_4_io_in = _T_863 & io_rPort_0_en_0; // @[package.scala 94:16:@13384.4]
  assign RetimeWrapper_5_clock = clock; // @[:@13390.4]
  assign RetimeWrapper_5_reset = reset; // @[:@13391.4]
  assign RetimeWrapper_5_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13393.4]
  assign RetimeWrapper_5_io_in = _T_955 & io_rPort_0_en_0; // @[package.scala 94:16:@13392.4]
  assign RetimeWrapper_6_clock = clock; // @[:@13398.4]
  assign RetimeWrapper_6_reset = reset; // @[:@13399.4]
  assign RetimeWrapper_6_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13401.4]
  assign RetimeWrapper_6_io_in = _T_1047 & io_rPort_0_en_0; // @[package.scala 94:16:@13400.4]
  assign RetimeWrapper_7_clock = clock; // @[:@13406.4]
  assign RetimeWrapper_7_reset = reset; // @[:@13407.4]
  assign RetimeWrapper_7_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13409.4]
  assign RetimeWrapper_7_io_in = _T_1139 & io_rPort_0_en_0; // @[package.scala 94:16:@13408.4]
  assign RetimeWrapper_8_clock = clock; // @[:@13414.4]
  assign RetimeWrapper_8_reset = reset; // @[:@13415.4]
  assign RetimeWrapper_8_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13417.4]
  assign RetimeWrapper_8_io_in = _T_1231 & io_rPort_0_en_0; // @[package.scala 94:16:@13416.4]
  assign RetimeWrapper_9_clock = clock; // @[:@13422.4]
  assign RetimeWrapper_9_reset = reset; // @[:@13423.4]
  assign RetimeWrapper_9_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13425.4]
  assign RetimeWrapper_9_io_in = _T_1323 & io_rPort_0_en_0; // @[package.scala 94:16:@13424.4]
  assign RetimeWrapper_10_clock = clock; // @[:@13430.4]
  assign RetimeWrapper_10_reset = reset; // @[:@13431.4]
  assign RetimeWrapper_10_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13433.4]
  assign RetimeWrapper_10_io_in = _T_1415 & io_rPort_0_en_0; // @[package.scala 94:16:@13432.4]
  assign RetimeWrapper_11_clock = clock; // @[:@13438.4]
  assign RetimeWrapper_11_reset = reset; // @[:@13439.4]
  assign RetimeWrapper_11_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13441.4]
  assign RetimeWrapper_11_io_in = _T_1507 & io_rPort_0_en_0; // @[package.scala 94:16:@13440.4]
  assign RetimeWrapper_12_clock = clock; // @[:@13446.4]
  assign RetimeWrapper_12_reset = reset; // @[:@13447.4]
  assign RetimeWrapper_12_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13449.4]
  assign RetimeWrapper_12_io_in = _T_1599 & io_rPort_0_en_0; // @[package.scala 94:16:@13448.4]
  assign RetimeWrapper_13_clock = clock; // @[:@13454.4]
  assign RetimeWrapper_13_reset = reset; // @[:@13455.4]
  assign RetimeWrapper_13_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13457.4]
  assign RetimeWrapper_13_io_in = _T_1691 & io_rPort_0_en_0; // @[package.scala 94:16:@13456.4]
  assign RetimeWrapper_14_clock = clock; // @[:@13462.4]
  assign RetimeWrapper_14_reset = reset; // @[:@13463.4]
  assign RetimeWrapper_14_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13465.4]
  assign RetimeWrapper_14_io_in = _T_1783 & io_rPort_0_en_0; // @[package.scala 94:16:@13464.4]
  assign RetimeWrapper_15_clock = clock; // @[:@13470.4]
  assign RetimeWrapper_15_reset = reset; // @[:@13471.4]
  assign RetimeWrapper_15_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13473.4]
  assign RetimeWrapper_15_io_in = _T_1875 & io_rPort_0_en_0; // @[package.scala 94:16:@13472.4]
  assign RetimeWrapper_16_clock = clock; // @[:@13542.4]
  assign RetimeWrapper_16_reset = reset; // @[:@13543.4]
  assign RetimeWrapper_16_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@13545.4]
  assign RetimeWrapper_16_io_in = _T_501 & io_rPort_1_en_0; // @[package.scala 94:16:@13544.4]
  assign RetimeWrapper_17_clock = clock; // @[:@13550.4]
  assign RetimeWrapper_17_reset = reset; // @[:@13551.4]
  assign RetimeWrapper_17_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@13553.4]
  assign RetimeWrapper_17_io_in = _T_593 & io_rPort_1_en_0; // @[package.scala 94:16:@13552.4]
  assign RetimeWrapper_18_clock = clock; // @[:@13558.4]
  assign RetimeWrapper_18_reset = reset; // @[:@13559.4]
  assign RetimeWrapper_18_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@13561.4]
  assign RetimeWrapper_18_io_in = _T_685 & io_rPort_1_en_0; // @[package.scala 94:16:@13560.4]
  assign RetimeWrapper_19_clock = clock; // @[:@13566.4]
  assign RetimeWrapper_19_reset = reset; // @[:@13567.4]
  assign RetimeWrapper_19_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@13569.4]
  assign RetimeWrapper_19_io_in = _T_777 & io_rPort_1_en_0; // @[package.scala 94:16:@13568.4]
  assign RetimeWrapper_20_clock = clock; // @[:@13574.4]
  assign RetimeWrapper_20_reset = reset; // @[:@13575.4]
  assign RetimeWrapper_20_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@13577.4]
  assign RetimeWrapper_20_io_in = _T_869 & io_rPort_1_en_0; // @[package.scala 94:16:@13576.4]
  assign RetimeWrapper_21_clock = clock; // @[:@13582.4]
  assign RetimeWrapper_21_reset = reset; // @[:@13583.4]
  assign RetimeWrapper_21_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@13585.4]
  assign RetimeWrapper_21_io_in = _T_961 & io_rPort_1_en_0; // @[package.scala 94:16:@13584.4]
  assign RetimeWrapper_22_clock = clock; // @[:@13590.4]
  assign RetimeWrapper_22_reset = reset; // @[:@13591.4]
  assign RetimeWrapper_22_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@13593.4]
  assign RetimeWrapper_22_io_in = _T_1053 & io_rPort_1_en_0; // @[package.scala 94:16:@13592.4]
  assign RetimeWrapper_23_clock = clock; // @[:@13598.4]
  assign RetimeWrapper_23_reset = reset; // @[:@13599.4]
  assign RetimeWrapper_23_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@13601.4]
  assign RetimeWrapper_23_io_in = _T_1145 & io_rPort_1_en_0; // @[package.scala 94:16:@13600.4]
  assign RetimeWrapper_24_clock = clock; // @[:@13606.4]
  assign RetimeWrapper_24_reset = reset; // @[:@13607.4]
  assign RetimeWrapper_24_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@13609.4]
  assign RetimeWrapper_24_io_in = _T_1237 & io_rPort_1_en_0; // @[package.scala 94:16:@13608.4]
  assign RetimeWrapper_25_clock = clock; // @[:@13614.4]
  assign RetimeWrapper_25_reset = reset; // @[:@13615.4]
  assign RetimeWrapper_25_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@13617.4]
  assign RetimeWrapper_25_io_in = _T_1329 & io_rPort_1_en_0; // @[package.scala 94:16:@13616.4]
  assign RetimeWrapper_26_clock = clock; // @[:@13622.4]
  assign RetimeWrapper_26_reset = reset; // @[:@13623.4]
  assign RetimeWrapper_26_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@13625.4]
  assign RetimeWrapper_26_io_in = _T_1421 & io_rPort_1_en_0; // @[package.scala 94:16:@13624.4]
  assign RetimeWrapper_27_clock = clock; // @[:@13630.4]
  assign RetimeWrapper_27_reset = reset; // @[:@13631.4]
  assign RetimeWrapper_27_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@13633.4]
  assign RetimeWrapper_27_io_in = _T_1513 & io_rPort_1_en_0; // @[package.scala 94:16:@13632.4]
  assign RetimeWrapper_28_clock = clock; // @[:@13638.4]
  assign RetimeWrapper_28_reset = reset; // @[:@13639.4]
  assign RetimeWrapper_28_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@13641.4]
  assign RetimeWrapper_28_io_in = _T_1605 & io_rPort_1_en_0; // @[package.scala 94:16:@13640.4]
  assign RetimeWrapper_29_clock = clock; // @[:@13646.4]
  assign RetimeWrapper_29_reset = reset; // @[:@13647.4]
  assign RetimeWrapper_29_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@13649.4]
  assign RetimeWrapper_29_io_in = _T_1697 & io_rPort_1_en_0; // @[package.scala 94:16:@13648.4]
  assign RetimeWrapper_30_clock = clock; // @[:@13654.4]
  assign RetimeWrapper_30_reset = reset; // @[:@13655.4]
  assign RetimeWrapper_30_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@13657.4]
  assign RetimeWrapper_30_io_in = _T_1789 & io_rPort_1_en_0; // @[package.scala 94:16:@13656.4]
  assign RetimeWrapper_31_clock = clock; // @[:@13662.4]
  assign RetimeWrapper_31_reset = reset; // @[:@13663.4]
  assign RetimeWrapper_31_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@13665.4]
  assign RetimeWrapper_31_io_in = _T_1881 & io_rPort_1_en_0; // @[package.scala 94:16:@13664.4]
  assign RetimeWrapper_32_clock = clock; // @[:@13734.4]
  assign RetimeWrapper_32_reset = reset; // @[:@13735.4]
  assign RetimeWrapper_32_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@13737.4]
  assign RetimeWrapper_32_io_in = _T_507 & io_rPort_2_en_0; // @[package.scala 94:16:@13736.4]
  assign RetimeWrapper_33_clock = clock; // @[:@13742.4]
  assign RetimeWrapper_33_reset = reset; // @[:@13743.4]
  assign RetimeWrapper_33_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@13745.4]
  assign RetimeWrapper_33_io_in = _T_599 & io_rPort_2_en_0; // @[package.scala 94:16:@13744.4]
  assign RetimeWrapper_34_clock = clock; // @[:@13750.4]
  assign RetimeWrapper_34_reset = reset; // @[:@13751.4]
  assign RetimeWrapper_34_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@13753.4]
  assign RetimeWrapper_34_io_in = _T_691 & io_rPort_2_en_0; // @[package.scala 94:16:@13752.4]
  assign RetimeWrapper_35_clock = clock; // @[:@13758.4]
  assign RetimeWrapper_35_reset = reset; // @[:@13759.4]
  assign RetimeWrapper_35_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@13761.4]
  assign RetimeWrapper_35_io_in = _T_783 & io_rPort_2_en_0; // @[package.scala 94:16:@13760.4]
  assign RetimeWrapper_36_clock = clock; // @[:@13766.4]
  assign RetimeWrapper_36_reset = reset; // @[:@13767.4]
  assign RetimeWrapper_36_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@13769.4]
  assign RetimeWrapper_36_io_in = _T_875 & io_rPort_2_en_0; // @[package.scala 94:16:@13768.4]
  assign RetimeWrapper_37_clock = clock; // @[:@13774.4]
  assign RetimeWrapper_37_reset = reset; // @[:@13775.4]
  assign RetimeWrapper_37_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@13777.4]
  assign RetimeWrapper_37_io_in = _T_967 & io_rPort_2_en_0; // @[package.scala 94:16:@13776.4]
  assign RetimeWrapper_38_clock = clock; // @[:@13782.4]
  assign RetimeWrapper_38_reset = reset; // @[:@13783.4]
  assign RetimeWrapper_38_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@13785.4]
  assign RetimeWrapper_38_io_in = _T_1059 & io_rPort_2_en_0; // @[package.scala 94:16:@13784.4]
  assign RetimeWrapper_39_clock = clock; // @[:@13790.4]
  assign RetimeWrapper_39_reset = reset; // @[:@13791.4]
  assign RetimeWrapper_39_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@13793.4]
  assign RetimeWrapper_39_io_in = _T_1151 & io_rPort_2_en_0; // @[package.scala 94:16:@13792.4]
  assign RetimeWrapper_40_clock = clock; // @[:@13798.4]
  assign RetimeWrapper_40_reset = reset; // @[:@13799.4]
  assign RetimeWrapper_40_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@13801.4]
  assign RetimeWrapper_40_io_in = _T_1243 & io_rPort_2_en_0; // @[package.scala 94:16:@13800.4]
  assign RetimeWrapper_41_clock = clock; // @[:@13806.4]
  assign RetimeWrapper_41_reset = reset; // @[:@13807.4]
  assign RetimeWrapper_41_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@13809.4]
  assign RetimeWrapper_41_io_in = _T_1335 & io_rPort_2_en_0; // @[package.scala 94:16:@13808.4]
  assign RetimeWrapper_42_clock = clock; // @[:@13814.4]
  assign RetimeWrapper_42_reset = reset; // @[:@13815.4]
  assign RetimeWrapper_42_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@13817.4]
  assign RetimeWrapper_42_io_in = _T_1427 & io_rPort_2_en_0; // @[package.scala 94:16:@13816.4]
  assign RetimeWrapper_43_clock = clock; // @[:@13822.4]
  assign RetimeWrapper_43_reset = reset; // @[:@13823.4]
  assign RetimeWrapper_43_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@13825.4]
  assign RetimeWrapper_43_io_in = _T_1519 & io_rPort_2_en_0; // @[package.scala 94:16:@13824.4]
  assign RetimeWrapper_44_clock = clock; // @[:@13830.4]
  assign RetimeWrapper_44_reset = reset; // @[:@13831.4]
  assign RetimeWrapper_44_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@13833.4]
  assign RetimeWrapper_44_io_in = _T_1611 & io_rPort_2_en_0; // @[package.scala 94:16:@13832.4]
  assign RetimeWrapper_45_clock = clock; // @[:@13838.4]
  assign RetimeWrapper_45_reset = reset; // @[:@13839.4]
  assign RetimeWrapper_45_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@13841.4]
  assign RetimeWrapper_45_io_in = _T_1703 & io_rPort_2_en_0; // @[package.scala 94:16:@13840.4]
  assign RetimeWrapper_46_clock = clock; // @[:@13846.4]
  assign RetimeWrapper_46_reset = reset; // @[:@13847.4]
  assign RetimeWrapper_46_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@13849.4]
  assign RetimeWrapper_46_io_in = _T_1795 & io_rPort_2_en_0; // @[package.scala 94:16:@13848.4]
  assign RetimeWrapper_47_clock = clock; // @[:@13854.4]
  assign RetimeWrapper_47_reset = reset; // @[:@13855.4]
  assign RetimeWrapper_47_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@13857.4]
  assign RetimeWrapper_47_io_in = _T_1887 & io_rPort_2_en_0; // @[package.scala 94:16:@13856.4]
  assign RetimeWrapper_48_clock = clock; // @[:@13926.4]
  assign RetimeWrapper_48_reset = reset; // @[:@13927.4]
  assign RetimeWrapper_48_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@13929.4]
  assign RetimeWrapper_48_io_in = _T_513 & io_rPort_3_en_0; // @[package.scala 94:16:@13928.4]
  assign RetimeWrapper_49_clock = clock; // @[:@13934.4]
  assign RetimeWrapper_49_reset = reset; // @[:@13935.4]
  assign RetimeWrapper_49_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@13937.4]
  assign RetimeWrapper_49_io_in = _T_605 & io_rPort_3_en_0; // @[package.scala 94:16:@13936.4]
  assign RetimeWrapper_50_clock = clock; // @[:@13942.4]
  assign RetimeWrapper_50_reset = reset; // @[:@13943.4]
  assign RetimeWrapper_50_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@13945.4]
  assign RetimeWrapper_50_io_in = _T_697 & io_rPort_3_en_0; // @[package.scala 94:16:@13944.4]
  assign RetimeWrapper_51_clock = clock; // @[:@13950.4]
  assign RetimeWrapper_51_reset = reset; // @[:@13951.4]
  assign RetimeWrapper_51_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@13953.4]
  assign RetimeWrapper_51_io_in = _T_789 & io_rPort_3_en_0; // @[package.scala 94:16:@13952.4]
  assign RetimeWrapper_52_clock = clock; // @[:@13958.4]
  assign RetimeWrapper_52_reset = reset; // @[:@13959.4]
  assign RetimeWrapper_52_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@13961.4]
  assign RetimeWrapper_52_io_in = _T_881 & io_rPort_3_en_0; // @[package.scala 94:16:@13960.4]
  assign RetimeWrapper_53_clock = clock; // @[:@13966.4]
  assign RetimeWrapper_53_reset = reset; // @[:@13967.4]
  assign RetimeWrapper_53_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@13969.4]
  assign RetimeWrapper_53_io_in = _T_973 & io_rPort_3_en_0; // @[package.scala 94:16:@13968.4]
  assign RetimeWrapper_54_clock = clock; // @[:@13974.4]
  assign RetimeWrapper_54_reset = reset; // @[:@13975.4]
  assign RetimeWrapper_54_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@13977.4]
  assign RetimeWrapper_54_io_in = _T_1065 & io_rPort_3_en_0; // @[package.scala 94:16:@13976.4]
  assign RetimeWrapper_55_clock = clock; // @[:@13982.4]
  assign RetimeWrapper_55_reset = reset; // @[:@13983.4]
  assign RetimeWrapper_55_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@13985.4]
  assign RetimeWrapper_55_io_in = _T_1157 & io_rPort_3_en_0; // @[package.scala 94:16:@13984.4]
  assign RetimeWrapper_56_clock = clock; // @[:@13990.4]
  assign RetimeWrapper_56_reset = reset; // @[:@13991.4]
  assign RetimeWrapper_56_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@13993.4]
  assign RetimeWrapper_56_io_in = _T_1249 & io_rPort_3_en_0; // @[package.scala 94:16:@13992.4]
  assign RetimeWrapper_57_clock = clock; // @[:@13998.4]
  assign RetimeWrapper_57_reset = reset; // @[:@13999.4]
  assign RetimeWrapper_57_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14001.4]
  assign RetimeWrapper_57_io_in = _T_1341 & io_rPort_3_en_0; // @[package.scala 94:16:@14000.4]
  assign RetimeWrapper_58_clock = clock; // @[:@14006.4]
  assign RetimeWrapper_58_reset = reset; // @[:@14007.4]
  assign RetimeWrapper_58_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14009.4]
  assign RetimeWrapper_58_io_in = _T_1433 & io_rPort_3_en_0; // @[package.scala 94:16:@14008.4]
  assign RetimeWrapper_59_clock = clock; // @[:@14014.4]
  assign RetimeWrapper_59_reset = reset; // @[:@14015.4]
  assign RetimeWrapper_59_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14017.4]
  assign RetimeWrapper_59_io_in = _T_1525 & io_rPort_3_en_0; // @[package.scala 94:16:@14016.4]
  assign RetimeWrapper_60_clock = clock; // @[:@14022.4]
  assign RetimeWrapper_60_reset = reset; // @[:@14023.4]
  assign RetimeWrapper_60_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14025.4]
  assign RetimeWrapper_60_io_in = _T_1617 & io_rPort_3_en_0; // @[package.scala 94:16:@14024.4]
  assign RetimeWrapper_61_clock = clock; // @[:@14030.4]
  assign RetimeWrapper_61_reset = reset; // @[:@14031.4]
  assign RetimeWrapper_61_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14033.4]
  assign RetimeWrapper_61_io_in = _T_1709 & io_rPort_3_en_0; // @[package.scala 94:16:@14032.4]
  assign RetimeWrapper_62_clock = clock; // @[:@14038.4]
  assign RetimeWrapper_62_reset = reset; // @[:@14039.4]
  assign RetimeWrapper_62_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14041.4]
  assign RetimeWrapper_62_io_in = _T_1801 & io_rPort_3_en_0; // @[package.scala 94:16:@14040.4]
  assign RetimeWrapper_63_clock = clock; // @[:@14046.4]
  assign RetimeWrapper_63_reset = reset; // @[:@14047.4]
  assign RetimeWrapper_63_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14049.4]
  assign RetimeWrapper_63_io_in = _T_1893 & io_rPort_3_en_0; // @[package.scala 94:16:@14048.4]
  assign RetimeWrapper_64_clock = clock; // @[:@14118.4]
  assign RetimeWrapper_64_reset = reset; // @[:@14119.4]
  assign RetimeWrapper_64_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14121.4]
  assign RetimeWrapper_64_io_in = _T_519 & io_rPort_4_en_0; // @[package.scala 94:16:@14120.4]
  assign RetimeWrapper_65_clock = clock; // @[:@14126.4]
  assign RetimeWrapper_65_reset = reset; // @[:@14127.4]
  assign RetimeWrapper_65_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14129.4]
  assign RetimeWrapper_65_io_in = _T_611 & io_rPort_4_en_0; // @[package.scala 94:16:@14128.4]
  assign RetimeWrapper_66_clock = clock; // @[:@14134.4]
  assign RetimeWrapper_66_reset = reset; // @[:@14135.4]
  assign RetimeWrapper_66_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14137.4]
  assign RetimeWrapper_66_io_in = _T_703 & io_rPort_4_en_0; // @[package.scala 94:16:@14136.4]
  assign RetimeWrapper_67_clock = clock; // @[:@14142.4]
  assign RetimeWrapper_67_reset = reset; // @[:@14143.4]
  assign RetimeWrapper_67_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14145.4]
  assign RetimeWrapper_67_io_in = _T_795 & io_rPort_4_en_0; // @[package.scala 94:16:@14144.4]
  assign RetimeWrapper_68_clock = clock; // @[:@14150.4]
  assign RetimeWrapper_68_reset = reset; // @[:@14151.4]
  assign RetimeWrapper_68_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14153.4]
  assign RetimeWrapper_68_io_in = _T_887 & io_rPort_4_en_0; // @[package.scala 94:16:@14152.4]
  assign RetimeWrapper_69_clock = clock; // @[:@14158.4]
  assign RetimeWrapper_69_reset = reset; // @[:@14159.4]
  assign RetimeWrapper_69_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14161.4]
  assign RetimeWrapper_69_io_in = _T_979 & io_rPort_4_en_0; // @[package.scala 94:16:@14160.4]
  assign RetimeWrapper_70_clock = clock; // @[:@14166.4]
  assign RetimeWrapper_70_reset = reset; // @[:@14167.4]
  assign RetimeWrapper_70_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14169.4]
  assign RetimeWrapper_70_io_in = _T_1071 & io_rPort_4_en_0; // @[package.scala 94:16:@14168.4]
  assign RetimeWrapper_71_clock = clock; // @[:@14174.4]
  assign RetimeWrapper_71_reset = reset; // @[:@14175.4]
  assign RetimeWrapper_71_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14177.4]
  assign RetimeWrapper_71_io_in = _T_1163 & io_rPort_4_en_0; // @[package.scala 94:16:@14176.4]
  assign RetimeWrapper_72_clock = clock; // @[:@14182.4]
  assign RetimeWrapper_72_reset = reset; // @[:@14183.4]
  assign RetimeWrapper_72_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14185.4]
  assign RetimeWrapper_72_io_in = _T_1255 & io_rPort_4_en_0; // @[package.scala 94:16:@14184.4]
  assign RetimeWrapper_73_clock = clock; // @[:@14190.4]
  assign RetimeWrapper_73_reset = reset; // @[:@14191.4]
  assign RetimeWrapper_73_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14193.4]
  assign RetimeWrapper_73_io_in = _T_1347 & io_rPort_4_en_0; // @[package.scala 94:16:@14192.4]
  assign RetimeWrapper_74_clock = clock; // @[:@14198.4]
  assign RetimeWrapper_74_reset = reset; // @[:@14199.4]
  assign RetimeWrapper_74_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14201.4]
  assign RetimeWrapper_74_io_in = _T_1439 & io_rPort_4_en_0; // @[package.scala 94:16:@14200.4]
  assign RetimeWrapper_75_clock = clock; // @[:@14206.4]
  assign RetimeWrapper_75_reset = reset; // @[:@14207.4]
  assign RetimeWrapper_75_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14209.4]
  assign RetimeWrapper_75_io_in = _T_1531 & io_rPort_4_en_0; // @[package.scala 94:16:@14208.4]
  assign RetimeWrapper_76_clock = clock; // @[:@14214.4]
  assign RetimeWrapper_76_reset = reset; // @[:@14215.4]
  assign RetimeWrapper_76_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14217.4]
  assign RetimeWrapper_76_io_in = _T_1623 & io_rPort_4_en_0; // @[package.scala 94:16:@14216.4]
  assign RetimeWrapper_77_clock = clock; // @[:@14222.4]
  assign RetimeWrapper_77_reset = reset; // @[:@14223.4]
  assign RetimeWrapper_77_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14225.4]
  assign RetimeWrapper_77_io_in = _T_1715 & io_rPort_4_en_0; // @[package.scala 94:16:@14224.4]
  assign RetimeWrapper_78_clock = clock; // @[:@14230.4]
  assign RetimeWrapper_78_reset = reset; // @[:@14231.4]
  assign RetimeWrapper_78_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14233.4]
  assign RetimeWrapper_78_io_in = _T_1807 & io_rPort_4_en_0; // @[package.scala 94:16:@14232.4]
  assign RetimeWrapper_79_clock = clock; // @[:@14238.4]
  assign RetimeWrapper_79_reset = reset; // @[:@14239.4]
  assign RetimeWrapper_79_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14241.4]
  assign RetimeWrapper_79_io_in = _T_1899 & io_rPort_4_en_0; // @[package.scala 94:16:@14240.4]
  assign RetimeWrapper_80_clock = clock; // @[:@14310.4]
  assign RetimeWrapper_80_reset = reset; // @[:@14311.4]
  assign RetimeWrapper_80_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14313.4]
  assign RetimeWrapper_80_io_in = _T_525 & io_rPort_5_en_0; // @[package.scala 94:16:@14312.4]
  assign RetimeWrapper_81_clock = clock; // @[:@14318.4]
  assign RetimeWrapper_81_reset = reset; // @[:@14319.4]
  assign RetimeWrapper_81_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14321.4]
  assign RetimeWrapper_81_io_in = _T_617 & io_rPort_5_en_0; // @[package.scala 94:16:@14320.4]
  assign RetimeWrapper_82_clock = clock; // @[:@14326.4]
  assign RetimeWrapper_82_reset = reset; // @[:@14327.4]
  assign RetimeWrapper_82_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14329.4]
  assign RetimeWrapper_82_io_in = _T_709 & io_rPort_5_en_0; // @[package.scala 94:16:@14328.4]
  assign RetimeWrapper_83_clock = clock; // @[:@14334.4]
  assign RetimeWrapper_83_reset = reset; // @[:@14335.4]
  assign RetimeWrapper_83_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14337.4]
  assign RetimeWrapper_83_io_in = _T_801 & io_rPort_5_en_0; // @[package.scala 94:16:@14336.4]
  assign RetimeWrapper_84_clock = clock; // @[:@14342.4]
  assign RetimeWrapper_84_reset = reset; // @[:@14343.4]
  assign RetimeWrapper_84_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14345.4]
  assign RetimeWrapper_84_io_in = _T_893 & io_rPort_5_en_0; // @[package.scala 94:16:@14344.4]
  assign RetimeWrapper_85_clock = clock; // @[:@14350.4]
  assign RetimeWrapper_85_reset = reset; // @[:@14351.4]
  assign RetimeWrapper_85_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14353.4]
  assign RetimeWrapper_85_io_in = _T_985 & io_rPort_5_en_0; // @[package.scala 94:16:@14352.4]
  assign RetimeWrapper_86_clock = clock; // @[:@14358.4]
  assign RetimeWrapper_86_reset = reset; // @[:@14359.4]
  assign RetimeWrapper_86_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14361.4]
  assign RetimeWrapper_86_io_in = _T_1077 & io_rPort_5_en_0; // @[package.scala 94:16:@14360.4]
  assign RetimeWrapper_87_clock = clock; // @[:@14366.4]
  assign RetimeWrapper_87_reset = reset; // @[:@14367.4]
  assign RetimeWrapper_87_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14369.4]
  assign RetimeWrapper_87_io_in = _T_1169 & io_rPort_5_en_0; // @[package.scala 94:16:@14368.4]
  assign RetimeWrapper_88_clock = clock; // @[:@14374.4]
  assign RetimeWrapper_88_reset = reset; // @[:@14375.4]
  assign RetimeWrapper_88_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14377.4]
  assign RetimeWrapper_88_io_in = _T_1261 & io_rPort_5_en_0; // @[package.scala 94:16:@14376.4]
  assign RetimeWrapper_89_clock = clock; // @[:@14382.4]
  assign RetimeWrapper_89_reset = reset; // @[:@14383.4]
  assign RetimeWrapper_89_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14385.4]
  assign RetimeWrapper_89_io_in = _T_1353 & io_rPort_5_en_0; // @[package.scala 94:16:@14384.4]
  assign RetimeWrapper_90_clock = clock; // @[:@14390.4]
  assign RetimeWrapper_90_reset = reset; // @[:@14391.4]
  assign RetimeWrapper_90_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14393.4]
  assign RetimeWrapper_90_io_in = _T_1445 & io_rPort_5_en_0; // @[package.scala 94:16:@14392.4]
  assign RetimeWrapper_91_clock = clock; // @[:@14398.4]
  assign RetimeWrapper_91_reset = reset; // @[:@14399.4]
  assign RetimeWrapper_91_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14401.4]
  assign RetimeWrapper_91_io_in = _T_1537 & io_rPort_5_en_0; // @[package.scala 94:16:@14400.4]
  assign RetimeWrapper_92_clock = clock; // @[:@14406.4]
  assign RetimeWrapper_92_reset = reset; // @[:@14407.4]
  assign RetimeWrapper_92_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14409.4]
  assign RetimeWrapper_92_io_in = _T_1629 & io_rPort_5_en_0; // @[package.scala 94:16:@14408.4]
  assign RetimeWrapper_93_clock = clock; // @[:@14414.4]
  assign RetimeWrapper_93_reset = reset; // @[:@14415.4]
  assign RetimeWrapper_93_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14417.4]
  assign RetimeWrapper_93_io_in = _T_1721 & io_rPort_5_en_0; // @[package.scala 94:16:@14416.4]
  assign RetimeWrapper_94_clock = clock; // @[:@14422.4]
  assign RetimeWrapper_94_reset = reset; // @[:@14423.4]
  assign RetimeWrapper_94_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14425.4]
  assign RetimeWrapper_94_io_in = _T_1813 & io_rPort_5_en_0; // @[package.scala 94:16:@14424.4]
  assign RetimeWrapper_95_clock = clock; // @[:@14430.4]
  assign RetimeWrapper_95_reset = reset; // @[:@14431.4]
  assign RetimeWrapper_95_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14433.4]
  assign RetimeWrapper_95_io_in = _T_1905 & io_rPort_5_en_0; // @[package.scala 94:16:@14432.4]
  assign RetimeWrapper_96_clock = clock; // @[:@14502.4]
  assign RetimeWrapper_96_reset = reset; // @[:@14503.4]
  assign RetimeWrapper_96_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14505.4]
  assign RetimeWrapper_96_io_in = _T_531 & io_rPort_6_en_0; // @[package.scala 94:16:@14504.4]
  assign RetimeWrapper_97_clock = clock; // @[:@14510.4]
  assign RetimeWrapper_97_reset = reset; // @[:@14511.4]
  assign RetimeWrapper_97_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14513.4]
  assign RetimeWrapper_97_io_in = _T_623 & io_rPort_6_en_0; // @[package.scala 94:16:@14512.4]
  assign RetimeWrapper_98_clock = clock; // @[:@14518.4]
  assign RetimeWrapper_98_reset = reset; // @[:@14519.4]
  assign RetimeWrapper_98_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14521.4]
  assign RetimeWrapper_98_io_in = _T_715 & io_rPort_6_en_0; // @[package.scala 94:16:@14520.4]
  assign RetimeWrapper_99_clock = clock; // @[:@14526.4]
  assign RetimeWrapper_99_reset = reset; // @[:@14527.4]
  assign RetimeWrapper_99_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14529.4]
  assign RetimeWrapper_99_io_in = _T_807 & io_rPort_6_en_0; // @[package.scala 94:16:@14528.4]
  assign RetimeWrapper_100_clock = clock; // @[:@14534.4]
  assign RetimeWrapper_100_reset = reset; // @[:@14535.4]
  assign RetimeWrapper_100_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14537.4]
  assign RetimeWrapper_100_io_in = _T_899 & io_rPort_6_en_0; // @[package.scala 94:16:@14536.4]
  assign RetimeWrapper_101_clock = clock; // @[:@14542.4]
  assign RetimeWrapper_101_reset = reset; // @[:@14543.4]
  assign RetimeWrapper_101_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14545.4]
  assign RetimeWrapper_101_io_in = _T_991 & io_rPort_6_en_0; // @[package.scala 94:16:@14544.4]
  assign RetimeWrapper_102_clock = clock; // @[:@14550.4]
  assign RetimeWrapper_102_reset = reset; // @[:@14551.4]
  assign RetimeWrapper_102_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14553.4]
  assign RetimeWrapper_102_io_in = _T_1083 & io_rPort_6_en_0; // @[package.scala 94:16:@14552.4]
  assign RetimeWrapper_103_clock = clock; // @[:@14558.4]
  assign RetimeWrapper_103_reset = reset; // @[:@14559.4]
  assign RetimeWrapper_103_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14561.4]
  assign RetimeWrapper_103_io_in = _T_1175 & io_rPort_6_en_0; // @[package.scala 94:16:@14560.4]
  assign RetimeWrapper_104_clock = clock; // @[:@14566.4]
  assign RetimeWrapper_104_reset = reset; // @[:@14567.4]
  assign RetimeWrapper_104_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14569.4]
  assign RetimeWrapper_104_io_in = _T_1267 & io_rPort_6_en_0; // @[package.scala 94:16:@14568.4]
  assign RetimeWrapper_105_clock = clock; // @[:@14574.4]
  assign RetimeWrapper_105_reset = reset; // @[:@14575.4]
  assign RetimeWrapper_105_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14577.4]
  assign RetimeWrapper_105_io_in = _T_1359 & io_rPort_6_en_0; // @[package.scala 94:16:@14576.4]
  assign RetimeWrapper_106_clock = clock; // @[:@14582.4]
  assign RetimeWrapper_106_reset = reset; // @[:@14583.4]
  assign RetimeWrapper_106_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14585.4]
  assign RetimeWrapper_106_io_in = _T_1451 & io_rPort_6_en_0; // @[package.scala 94:16:@14584.4]
  assign RetimeWrapper_107_clock = clock; // @[:@14590.4]
  assign RetimeWrapper_107_reset = reset; // @[:@14591.4]
  assign RetimeWrapper_107_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14593.4]
  assign RetimeWrapper_107_io_in = _T_1543 & io_rPort_6_en_0; // @[package.scala 94:16:@14592.4]
  assign RetimeWrapper_108_clock = clock; // @[:@14598.4]
  assign RetimeWrapper_108_reset = reset; // @[:@14599.4]
  assign RetimeWrapper_108_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14601.4]
  assign RetimeWrapper_108_io_in = _T_1635 & io_rPort_6_en_0; // @[package.scala 94:16:@14600.4]
  assign RetimeWrapper_109_clock = clock; // @[:@14606.4]
  assign RetimeWrapper_109_reset = reset; // @[:@14607.4]
  assign RetimeWrapper_109_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14609.4]
  assign RetimeWrapper_109_io_in = _T_1727 & io_rPort_6_en_0; // @[package.scala 94:16:@14608.4]
  assign RetimeWrapper_110_clock = clock; // @[:@14614.4]
  assign RetimeWrapper_110_reset = reset; // @[:@14615.4]
  assign RetimeWrapper_110_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14617.4]
  assign RetimeWrapper_110_io_in = _T_1819 & io_rPort_6_en_0; // @[package.scala 94:16:@14616.4]
  assign RetimeWrapper_111_clock = clock; // @[:@14622.4]
  assign RetimeWrapper_111_reset = reset; // @[:@14623.4]
  assign RetimeWrapper_111_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14625.4]
  assign RetimeWrapper_111_io_in = _T_1911 & io_rPort_6_en_0; // @[package.scala 94:16:@14624.4]
  assign RetimeWrapper_112_clock = clock; // @[:@14694.4]
  assign RetimeWrapper_112_reset = reset; // @[:@14695.4]
  assign RetimeWrapper_112_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14697.4]
  assign RetimeWrapper_112_io_in = _T_537 & io_rPort_7_en_0; // @[package.scala 94:16:@14696.4]
  assign RetimeWrapper_113_clock = clock; // @[:@14702.4]
  assign RetimeWrapper_113_reset = reset; // @[:@14703.4]
  assign RetimeWrapper_113_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14705.4]
  assign RetimeWrapper_113_io_in = _T_629 & io_rPort_7_en_0; // @[package.scala 94:16:@14704.4]
  assign RetimeWrapper_114_clock = clock; // @[:@14710.4]
  assign RetimeWrapper_114_reset = reset; // @[:@14711.4]
  assign RetimeWrapper_114_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14713.4]
  assign RetimeWrapper_114_io_in = _T_721 & io_rPort_7_en_0; // @[package.scala 94:16:@14712.4]
  assign RetimeWrapper_115_clock = clock; // @[:@14718.4]
  assign RetimeWrapper_115_reset = reset; // @[:@14719.4]
  assign RetimeWrapper_115_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14721.4]
  assign RetimeWrapper_115_io_in = _T_813 & io_rPort_7_en_0; // @[package.scala 94:16:@14720.4]
  assign RetimeWrapper_116_clock = clock; // @[:@14726.4]
  assign RetimeWrapper_116_reset = reset; // @[:@14727.4]
  assign RetimeWrapper_116_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14729.4]
  assign RetimeWrapper_116_io_in = _T_905 & io_rPort_7_en_0; // @[package.scala 94:16:@14728.4]
  assign RetimeWrapper_117_clock = clock; // @[:@14734.4]
  assign RetimeWrapper_117_reset = reset; // @[:@14735.4]
  assign RetimeWrapper_117_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14737.4]
  assign RetimeWrapper_117_io_in = _T_997 & io_rPort_7_en_0; // @[package.scala 94:16:@14736.4]
  assign RetimeWrapper_118_clock = clock; // @[:@14742.4]
  assign RetimeWrapper_118_reset = reset; // @[:@14743.4]
  assign RetimeWrapper_118_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14745.4]
  assign RetimeWrapper_118_io_in = _T_1089 & io_rPort_7_en_0; // @[package.scala 94:16:@14744.4]
  assign RetimeWrapper_119_clock = clock; // @[:@14750.4]
  assign RetimeWrapper_119_reset = reset; // @[:@14751.4]
  assign RetimeWrapper_119_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14753.4]
  assign RetimeWrapper_119_io_in = _T_1181 & io_rPort_7_en_0; // @[package.scala 94:16:@14752.4]
  assign RetimeWrapper_120_clock = clock; // @[:@14758.4]
  assign RetimeWrapper_120_reset = reset; // @[:@14759.4]
  assign RetimeWrapper_120_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14761.4]
  assign RetimeWrapper_120_io_in = _T_1273 & io_rPort_7_en_0; // @[package.scala 94:16:@14760.4]
  assign RetimeWrapper_121_clock = clock; // @[:@14766.4]
  assign RetimeWrapper_121_reset = reset; // @[:@14767.4]
  assign RetimeWrapper_121_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14769.4]
  assign RetimeWrapper_121_io_in = _T_1365 & io_rPort_7_en_0; // @[package.scala 94:16:@14768.4]
  assign RetimeWrapper_122_clock = clock; // @[:@14774.4]
  assign RetimeWrapper_122_reset = reset; // @[:@14775.4]
  assign RetimeWrapper_122_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14777.4]
  assign RetimeWrapper_122_io_in = _T_1457 & io_rPort_7_en_0; // @[package.scala 94:16:@14776.4]
  assign RetimeWrapper_123_clock = clock; // @[:@14782.4]
  assign RetimeWrapper_123_reset = reset; // @[:@14783.4]
  assign RetimeWrapper_123_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14785.4]
  assign RetimeWrapper_123_io_in = _T_1549 & io_rPort_7_en_0; // @[package.scala 94:16:@14784.4]
  assign RetimeWrapper_124_clock = clock; // @[:@14790.4]
  assign RetimeWrapper_124_reset = reset; // @[:@14791.4]
  assign RetimeWrapper_124_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14793.4]
  assign RetimeWrapper_124_io_in = _T_1641 & io_rPort_7_en_0; // @[package.scala 94:16:@14792.4]
  assign RetimeWrapper_125_clock = clock; // @[:@14798.4]
  assign RetimeWrapper_125_reset = reset; // @[:@14799.4]
  assign RetimeWrapper_125_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14801.4]
  assign RetimeWrapper_125_io_in = _T_1733 & io_rPort_7_en_0; // @[package.scala 94:16:@14800.4]
  assign RetimeWrapper_126_clock = clock; // @[:@14806.4]
  assign RetimeWrapper_126_reset = reset; // @[:@14807.4]
  assign RetimeWrapper_126_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14809.4]
  assign RetimeWrapper_126_io_in = _T_1825 & io_rPort_7_en_0; // @[package.scala 94:16:@14808.4]
  assign RetimeWrapper_127_clock = clock; // @[:@14814.4]
  assign RetimeWrapper_127_reset = reset; // @[:@14815.4]
  assign RetimeWrapper_127_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14817.4]
  assign RetimeWrapper_127_io_in = _T_1917 & io_rPort_7_en_0; // @[package.scala 94:16:@14816.4]
  assign RetimeWrapper_128_clock = clock; // @[:@14886.4]
  assign RetimeWrapper_128_reset = reset; // @[:@14887.4]
  assign RetimeWrapper_128_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@14889.4]
  assign RetimeWrapper_128_io_in = _T_543 & io_rPort_8_en_0; // @[package.scala 94:16:@14888.4]
  assign RetimeWrapper_129_clock = clock; // @[:@14894.4]
  assign RetimeWrapper_129_reset = reset; // @[:@14895.4]
  assign RetimeWrapper_129_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@14897.4]
  assign RetimeWrapper_129_io_in = _T_635 & io_rPort_8_en_0; // @[package.scala 94:16:@14896.4]
  assign RetimeWrapper_130_clock = clock; // @[:@14902.4]
  assign RetimeWrapper_130_reset = reset; // @[:@14903.4]
  assign RetimeWrapper_130_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@14905.4]
  assign RetimeWrapper_130_io_in = _T_727 & io_rPort_8_en_0; // @[package.scala 94:16:@14904.4]
  assign RetimeWrapper_131_clock = clock; // @[:@14910.4]
  assign RetimeWrapper_131_reset = reset; // @[:@14911.4]
  assign RetimeWrapper_131_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@14913.4]
  assign RetimeWrapper_131_io_in = _T_819 & io_rPort_8_en_0; // @[package.scala 94:16:@14912.4]
  assign RetimeWrapper_132_clock = clock; // @[:@14918.4]
  assign RetimeWrapper_132_reset = reset; // @[:@14919.4]
  assign RetimeWrapper_132_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@14921.4]
  assign RetimeWrapper_132_io_in = _T_911 & io_rPort_8_en_0; // @[package.scala 94:16:@14920.4]
  assign RetimeWrapper_133_clock = clock; // @[:@14926.4]
  assign RetimeWrapper_133_reset = reset; // @[:@14927.4]
  assign RetimeWrapper_133_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@14929.4]
  assign RetimeWrapper_133_io_in = _T_1003 & io_rPort_8_en_0; // @[package.scala 94:16:@14928.4]
  assign RetimeWrapper_134_clock = clock; // @[:@14934.4]
  assign RetimeWrapper_134_reset = reset; // @[:@14935.4]
  assign RetimeWrapper_134_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@14937.4]
  assign RetimeWrapper_134_io_in = _T_1095 & io_rPort_8_en_0; // @[package.scala 94:16:@14936.4]
  assign RetimeWrapper_135_clock = clock; // @[:@14942.4]
  assign RetimeWrapper_135_reset = reset; // @[:@14943.4]
  assign RetimeWrapper_135_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@14945.4]
  assign RetimeWrapper_135_io_in = _T_1187 & io_rPort_8_en_0; // @[package.scala 94:16:@14944.4]
  assign RetimeWrapper_136_clock = clock; // @[:@14950.4]
  assign RetimeWrapper_136_reset = reset; // @[:@14951.4]
  assign RetimeWrapper_136_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@14953.4]
  assign RetimeWrapper_136_io_in = _T_1279 & io_rPort_8_en_0; // @[package.scala 94:16:@14952.4]
  assign RetimeWrapper_137_clock = clock; // @[:@14958.4]
  assign RetimeWrapper_137_reset = reset; // @[:@14959.4]
  assign RetimeWrapper_137_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@14961.4]
  assign RetimeWrapper_137_io_in = _T_1371 & io_rPort_8_en_0; // @[package.scala 94:16:@14960.4]
  assign RetimeWrapper_138_clock = clock; // @[:@14966.4]
  assign RetimeWrapper_138_reset = reset; // @[:@14967.4]
  assign RetimeWrapper_138_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@14969.4]
  assign RetimeWrapper_138_io_in = _T_1463 & io_rPort_8_en_0; // @[package.scala 94:16:@14968.4]
  assign RetimeWrapper_139_clock = clock; // @[:@14974.4]
  assign RetimeWrapper_139_reset = reset; // @[:@14975.4]
  assign RetimeWrapper_139_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@14977.4]
  assign RetimeWrapper_139_io_in = _T_1555 & io_rPort_8_en_0; // @[package.scala 94:16:@14976.4]
  assign RetimeWrapper_140_clock = clock; // @[:@14982.4]
  assign RetimeWrapper_140_reset = reset; // @[:@14983.4]
  assign RetimeWrapper_140_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@14985.4]
  assign RetimeWrapper_140_io_in = _T_1647 & io_rPort_8_en_0; // @[package.scala 94:16:@14984.4]
  assign RetimeWrapper_141_clock = clock; // @[:@14990.4]
  assign RetimeWrapper_141_reset = reset; // @[:@14991.4]
  assign RetimeWrapper_141_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@14993.4]
  assign RetimeWrapper_141_io_in = _T_1739 & io_rPort_8_en_0; // @[package.scala 94:16:@14992.4]
  assign RetimeWrapper_142_clock = clock; // @[:@14998.4]
  assign RetimeWrapper_142_reset = reset; // @[:@14999.4]
  assign RetimeWrapper_142_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15001.4]
  assign RetimeWrapper_142_io_in = _T_1831 & io_rPort_8_en_0; // @[package.scala 94:16:@15000.4]
  assign RetimeWrapper_143_clock = clock; // @[:@15006.4]
  assign RetimeWrapper_143_reset = reset; // @[:@15007.4]
  assign RetimeWrapper_143_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15009.4]
  assign RetimeWrapper_143_io_in = _T_1923 & io_rPort_8_en_0; // @[package.scala 94:16:@15008.4]
endmodule
module SimBlackBoxesfix2fixBox_2( // @[:@15061.2]
  input  [31:0] io_a, // @[:@15064.4]
  output [32:0] io_b // @[:@15064.4]
);
  wire  _T_20; // @[implicits.scala 69:16:@15071.4]
  assign _T_20 = io_a[31]; // @[implicits.scala 69:16:@15071.4]
  assign io_b = {_T_20,io_a}; // @[SimBlackBoxes.scala 99:40:@15076.4]
endmodule
module __2( // @[:@15078.2]
  input  [31:0] io_b, // @[:@15081.4]
  output [32:0] io_result // @[:@15081.4]
);
  wire [31:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@15086.4]
  wire [32:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@15086.4]
  SimBlackBoxesfix2fixBox_2 SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@15086.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@15099.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@15094.4]
endmodule
module RetimeWrapper_197( // @[:@15153.2]
  input         clock, // @[:@15154.4]
  input         reset, // @[:@15155.4]
  input         io_flow, // @[:@15156.4]
  input  [31:0] io_in, // @[:@15156.4]
  output [31:0] io_out // @[:@15156.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@15158.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@15158.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@15158.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@15158.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@15158.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@15158.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@15158.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@15171.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@15170.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@15169.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@15168.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@15167.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@15165.4]
endmodule
module fix2fixBox( // @[:@15173.2]
  input         clock, // @[:@15174.4]
  input         reset, // @[:@15175.4]
  input  [32:0] io_a, // @[:@15176.4]
  input         io_flow, // @[:@15176.4]
  output [31:0] io_b // @[:@15176.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@15186.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@15186.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@15186.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@15186.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@15186.4]
  RetimeWrapper_197 RetimeWrapper ( // @[package.scala 93:22:@15186.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@15193.4]
  assign RetimeWrapper_clock = clock; // @[:@15187.4]
  assign RetimeWrapper_reset = reset; // @[:@15188.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@15190.4]
  assign RetimeWrapper_io_in = io_a[31:0]; // @[package.scala 94:16:@15189.4]
endmodule
module x297_sum( // @[:@15195.2]
  input         clock, // @[:@15196.4]
  input         reset, // @[:@15197.4]
  input  [31:0] io_a, // @[:@15198.4]
  input  [31:0] io_b, // @[:@15198.4]
  input         io_flow, // @[:@15198.4]
  output [31:0] io_result // @[:@15198.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@15206.4]
  wire [32:0] __io_result; // @[Math.scala 709:24:@15206.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@15213.4]
  wire [32:0] __1_io_result; // @[Math.scala 709:24:@15213.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@15231.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@15231.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@15231.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@15231.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@15231.4]
  wire [32:0] a_upcast_number; // @[Math.scala 712:22:@15211.4 Math.scala 713:14:@15212.4]
  wire [32:0] b_upcast_number; // @[Math.scala 712:22:@15218.4 Math.scala 713:14:@15219.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@15220.4]
  __2 _ ( // @[Math.scala 709:24:@15206.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 709:24:@15213.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox fix2fixBox ( // @[Math.scala 141:30:@15231.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@15211.4 Math.scala 713:14:@15212.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@15218.4 Math.scala 713:14:@15219.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@15220.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@15239.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@15209.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@15216.4]
  assign fix2fixBox_clock = clock; // @[:@15232.4]
  assign fix2fixBox_reset = reset; // @[:@15233.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@15234.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@15237.4]
endmodule
module RetimeWrapper_203( // @[:@15413.2]
  input         clock, // @[:@15414.4]
  input         reset, // @[:@15415.4]
  input         io_flow, // @[:@15416.4]
  input  [31:0] io_in, // @[:@15416.4]
  output [31:0] io_out // @[:@15416.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@15418.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@15418.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@15418.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@15418.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@15418.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@15418.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@15418.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@15431.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@15430.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@15429.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@15428.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@15427.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@15425.4]
endmodule
module RetimeWrapper_208( // @[:@15721.2]
  input         clock, // @[:@15722.4]
  input         reset, // @[:@15723.4]
  input         io_flow, // @[:@15724.4]
  input  [31:0] io_in, // @[:@15724.4]
  output [31:0] io_out // @[:@15724.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@15726.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@15726.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@15726.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@15726.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@15726.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@15726.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(5)) sr ( // @[RetimeShiftRegister.scala 15:20:@15726.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@15739.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@15738.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@15737.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@15736.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@15735.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@15733.4]
endmodule
module RetimeWrapper_210( // @[:@15785.2]
  input         clock, // @[:@15786.4]
  input         reset, // @[:@15787.4]
  input         io_flow, // @[:@15788.4]
  input  [31:0] io_in, // @[:@15788.4]
  output [31:0] io_out // @[:@15788.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@15790.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@15790.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@15790.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@15790.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@15790.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@15790.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@15790.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@15803.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@15802.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@15801.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@15800.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@15799.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@15797.4]
endmodule
module RetimeWrapper_211( // @[:@15817.2]
  input   clock, // @[:@15818.4]
  input   reset, // @[:@15819.4]
  input   io_flow, // @[:@15820.4]
  input   io_in, // @[:@15820.4]
  output  io_out // @[:@15820.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@15822.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@15822.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@15822.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@15822.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@15822.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@15822.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(5)) sr ( // @[RetimeShiftRegister.scala 15:20:@15822.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@15835.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@15834.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@15833.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@15832.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@15831.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@15829.4]
endmodule
module RetimeWrapper_212( // @[:@15849.2]
  input   clock, // @[:@15850.4]
  input   reset, // @[:@15851.4]
  input   io_flow, // @[:@15852.4]
  input   io_in, // @[:@15852.4]
  output  io_out // @[:@15852.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@15854.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@15854.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@15854.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@15854.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@15854.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@15854.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(4)) sr ( // @[RetimeShiftRegister.scala 15:20:@15854.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@15867.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@15866.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@15865.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@15864.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@15863.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@15861.4]
endmodule
module x323_rdcol( // @[:@16003.2]
  input         clock, // @[:@16004.4]
  input         reset, // @[:@16005.4]
  input  [31:0] io_a, // @[:@16006.4]
  input  [31:0] io_b, // @[:@16006.4]
  input         io_flow, // @[:@16006.4]
  output [31:0] io_result // @[:@16006.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@16014.4]
  wire [32:0] __io_result; // @[Math.scala 709:24:@16014.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@16021.4]
  wire [32:0] __1_io_result; // @[Math.scala 709:24:@16021.4]
  wire  fix2fixBox_clock; // @[Math.scala 182:30:@16040.4]
  wire  fix2fixBox_reset; // @[Math.scala 182:30:@16040.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 182:30:@16040.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 182:30:@16040.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 182:30:@16040.4]
  wire [32:0] a_upcast_number; // @[Math.scala 712:22:@16019.4 Math.scala 713:14:@16020.4]
  wire [32:0] b_upcast_number; // @[Math.scala 712:22:@16026.4 Math.scala 713:14:@16027.4]
  wire [33:0] _T_21; // @[Math.scala 177:37:@16028.4]
  wire [33:0] _T_22; // @[Math.scala 177:37:@16029.4]
  __2 _ ( // @[Math.scala 709:24:@16014.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 709:24:@16021.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox fix2fixBox ( // @[Math.scala 182:30:@16040.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@16019.4 Math.scala 713:14:@16020.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@16026.4 Math.scala 713:14:@16027.4]
  assign _T_21 = a_upcast_number - b_upcast_number; // @[Math.scala 177:37:@16028.4]
  assign _T_22 = $unsigned(_T_21); // @[Math.scala 177:37:@16029.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 188:17:@16048.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@16017.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@16024.4]
  assign fix2fixBox_clock = clock; // @[:@16041.4]
  assign fix2fixBox_reset = reset; // @[:@16042.4]
  assign fix2fixBox_io_a = _T_22[32:0]; // @[Math.scala 183:23:@16043.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 186:26:@16046.4]
endmodule
module RetimeWrapper_220( // @[:@16402.2]
  input   clock, // @[:@16403.4]
  input   reset, // @[:@16404.4]
  input   io_flow, // @[:@16405.4]
  input   io_in, // @[:@16405.4]
  output  io_out // @[:@16405.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@16407.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@16407.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@16407.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@16407.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@16407.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@16407.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@16407.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@16420.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@16419.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@16418.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@16417.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@16416.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@16414.4]
endmodule
module RetimeWrapper_229( // @[:@17136.2]
  input         clock, // @[:@17137.4]
  input         reset, // @[:@17138.4]
  input         io_flow, // @[:@17139.4]
  input  [31:0] io_in, // @[:@17139.4]
  output [31:0] io_out // @[:@17139.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@17141.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@17141.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@17141.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@17141.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@17141.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@17141.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(4)) sr ( // @[RetimeShiftRegister.scala 15:20:@17141.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@17154.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@17153.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@17152.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@17151.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@17150.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@17148.4]
endmodule
module SimBlackBoxesfix2fixBox_30( // @[:@19249.2]
  input  [7:0] io_a, // @[:@19252.4]
  output [8:0] io_b // @[:@19252.4]
);
  assign io_b = {1'h0,io_a}; // @[SimBlackBoxes.scala 99:40:@19263.4]
endmodule
module __30( // @[:@19265.2]
  input  [7:0] io_b, // @[:@19268.4]
  output [8:0] io_result // @[:@19268.4]
);
  wire [7:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@19273.4]
  wire [8:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@19273.4]
  SimBlackBoxesfix2fixBox_30 SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@19273.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@19286.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@19281.4]
endmodule
module fix2fixBox_14( // @[:@19327.2]
  input  [8:0] io_a, // @[:@19330.4]
  output [7:0] io_b // @[:@19330.4]
);
  assign io_b = io_a[7:0]; // @[Converter.scala 95:38:@19340.4]
endmodule
module x472_x11( // @[:@19342.2]
  input  [7:0] io_a, // @[:@19345.4]
  input  [7:0] io_b, // @[:@19345.4]
  output [7:0] io_result // @[:@19345.4]
);
  wire [7:0] __io_b; // @[Math.scala 709:24:@19353.4]
  wire [8:0] __io_result; // @[Math.scala 709:24:@19353.4]
  wire [7:0] __1_io_b; // @[Math.scala 709:24:@19360.4]
  wire [8:0] __1_io_result; // @[Math.scala 709:24:@19360.4]
  wire [8:0] fix2fixBox_io_a; // @[Math.scala 141:30:@19370.4]
  wire [7:0] fix2fixBox_io_b; // @[Math.scala 141:30:@19370.4]
  wire [8:0] a_upcast_number; // @[Math.scala 712:22:@19358.4 Math.scala 713:14:@19359.4]
  wire [8:0] b_upcast_number; // @[Math.scala 712:22:@19365.4 Math.scala 713:14:@19366.4]
  wire [9:0] _T_21; // @[Math.scala 136:37:@19367.4]
  __30 _ ( // @[Math.scala 709:24:@19353.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __30 __1 ( // @[Math.scala 709:24:@19360.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_14 fix2fixBox ( // @[Math.scala 141:30:@19370.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@19358.4 Math.scala 713:14:@19359.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@19365.4 Math.scala 713:14:@19366.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@19367.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@19378.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@19356.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@19363.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@19373.4]
endmodule
module fix2fixBox_20( // @[:@20209.2]
  input        clock, // @[:@20210.4]
  input        reset, // @[:@20211.4]
  input  [8:0] io_a, // @[:@20212.4]
  input        io_flow, // @[:@20212.4]
  output [7:0] io_b // @[:@20212.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@20222.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@20222.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@20222.4]
  wire [7:0] RetimeWrapper_io_in; // @[package.scala 93:22:@20222.4]
  wire [7:0] RetimeWrapper_io_out; // @[package.scala 93:22:@20222.4]
  RetimeWrapper_21 RetimeWrapper ( // @[package.scala 93:22:@20222.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@20229.4]
  assign RetimeWrapper_clock = clock; // @[:@20223.4]
  assign RetimeWrapper_reset = reset; // @[:@20224.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@20226.4]
  assign RetimeWrapper_io_in = io_a[7:0]; // @[package.scala 94:16:@20225.4]
endmodule
module x478_x11( // @[:@20231.2]
  input        clock, // @[:@20232.4]
  input        reset, // @[:@20233.4]
  input  [7:0] io_a, // @[:@20234.4]
  input  [7:0] io_b, // @[:@20234.4]
  input        io_flow, // @[:@20234.4]
  output [7:0] io_result // @[:@20234.4]
);
  wire [7:0] __io_b; // @[Math.scala 709:24:@20242.4]
  wire [8:0] __io_result; // @[Math.scala 709:24:@20242.4]
  wire [7:0] __1_io_b; // @[Math.scala 709:24:@20249.4]
  wire [8:0] __1_io_result; // @[Math.scala 709:24:@20249.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@20259.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@20259.4]
  wire [8:0] fix2fixBox_io_a; // @[Math.scala 141:30:@20259.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@20259.4]
  wire [7:0] fix2fixBox_io_b; // @[Math.scala 141:30:@20259.4]
  wire [8:0] a_upcast_number; // @[Math.scala 712:22:@20247.4 Math.scala 713:14:@20248.4]
  wire [8:0] b_upcast_number; // @[Math.scala 712:22:@20254.4 Math.scala 713:14:@20255.4]
  wire [9:0] _T_21; // @[Math.scala 136:37:@20256.4]
  __30 _ ( // @[Math.scala 709:24:@20242.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __30 __1 ( // @[Math.scala 709:24:@20249.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_20 fix2fixBox ( // @[Math.scala 141:30:@20259.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@20247.4 Math.scala 713:14:@20248.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@20254.4 Math.scala 713:14:@20255.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@20256.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@20267.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@20245.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@20252.4]
  assign fix2fixBox_clock = clock; // @[:@20260.4]
  assign fix2fixBox_reset = reset; // @[:@20261.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@20262.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@20265.4]
endmodule
module RetimeWrapper_266( // @[:@20281.2]
  input        clock, // @[:@20282.4]
  input        reset, // @[:@20283.4]
  input        io_flow, // @[:@20284.4]
  input  [7:0] io_in, // @[:@20284.4]
  output [7:0] io_out // @[:@20284.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@20286.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@20286.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@20286.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@20286.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@20286.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@20286.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@20286.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@20299.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@20298.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@20297.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@20296.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@20295.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@20293.4]
endmodule
module RetimeWrapper_267( // @[:@20444.2]
  input        clock, // @[:@20445.4]
  input        reset, // @[:@20446.4]
  input        io_flow, // @[:@20447.4]
  input  [7:0] io_in, // @[:@20447.4]
  output [7:0] io_out // @[:@20447.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@20449.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@20449.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@20449.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@20449.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@20449.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@20449.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@20449.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@20462.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@20461.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@20460.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@20459.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@20458.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@20456.4]
endmodule
module x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1( // @[:@20560.2]
  input          clock, // @[:@20561.4]
  input          reset, // @[:@20562.4]
  output         io_in_x270_TREADY, // @[:@20563.4]
  input  [255:0] io_in_x270_TDATA, // @[:@20563.4]
  input  [7:0]   io_in_x270_TID, // @[:@20563.4]
  input  [7:0]   io_in_x270_TDEST, // @[:@20563.4]
  output         io_in_x271_TVALID, // @[:@20563.4]
  input          io_in_x271_TREADY, // @[:@20563.4]
  output [255:0] io_in_x271_TDATA, // @[:@20563.4]
  input          io_sigsIn_backpressure, // @[:@20563.4]
  input          io_sigsIn_datapathEn, // @[:@20563.4]
  input          io_sigsIn_break, // @[:@20563.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_1, // @[:@20563.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_0, // @[:@20563.4]
  input          io_sigsIn_cchainOutputs_0_oobs_0, // @[:@20563.4]
  input          io_sigsIn_cchainOutputs_0_oobs_1, // @[:@20563.4]
  input          io_rr // @[:@20563.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@20577.4]
  wire [31:0] __io_result; // @[Math.scala 709:24:@20577.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@20589.4]
  wire [31:0] __1_io_result; // @[Math.scala 709:24:@20589.4]
  wire  x283_lb_0_clock; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire  x283_lb_0_reset; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire [2:0] x283_lb_0_io_rPort_8_banks_1; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire [2:0] x283_lb_0_io_rPort_8_banks_0; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire  x283_lb_0_io_rPort_8_ofs_0; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire  x283_lb_0_io_rPort_8_en_0; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire  x283_lb_0_io_rPort_8_backpressure; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire [7:0] x283_lb_0_io_rPort_8_output_0; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire [2:0] x283_lb_0_io_rPort_7_banks_1; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire [2:0] x283_lb_0_io_rPort_7_banks_0; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire  x283_lb_0_io_rPort_7_ofs_0; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire  x283_lb_0_io_rPort_7_en_0; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire  x283_lb_0_io_rPort_7_backpressure; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire [7:0] x283_lb_0_io_rPort_7_output_0; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire [2:0] x283_lb_0_io_rPort_6_banks_1; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire [2:0] x283_lb_0_io_rPort_6_banks_0; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire  x283_lb_0_io_rPort_6_ofs_0; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire  x283_lb_0_io_rPort_6_en_0; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire  x283_lb_0_io_rPort_6_backpressure; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire [7:0] x283_lb_0_io_rPort_6_output_0; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire [2:0] x283_lb_0_io_rPort_5_banks_1; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire [2:0] x283_lb_0_io_rPort_5_banks_0; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire  x283_lb_0_io_rPort_5_ofs_0; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire  x283_lb_0_io_rPort_5_en_0; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire  x283_lb_0_io_rPort_5_backpressure; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire [7:0] x283_lb_0_io_rPort_5_output_0; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire [2:0] x283_lb_0_io_rPort_4_banks_1; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire [2:0] x283_lb_0_io_rPort_4_banks_0; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire  x283_lb_0_io_rPort_4_ofs_0; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire  x283_lb_0_io_rPort_4_en_0; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire  x283_lb_0_io_rPort_4_backpressure; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire [7:0] x283_lb_0_io_rPort_4_output_0; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire [2:0] x283_lb_0_io_rPort_3_banks_1; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire [2:0] x283_lb_0_io_rPort_3_banks_0; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire  x283_lb_0_io_rPort_3_ofs_0; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire  x283_lb_0_io_rPort_3_en_0; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire  x283_lb_0_io_rPort_3_backpressure; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire [7:0] x283_lb_0_io_rPort_3_output_0; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire [2:0] x283_lb_0_io_rPort_2_banks_1; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire [2:0] x283_lb_0_io_rPort_2_banks_0; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire  x283_lb_0_io_rPort_2_ofs_0; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire  x283_lb_0_io_rPort_2_en_0; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire  x283_lb_0_io_rPort_2_backpressure; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire [7:0] x283_lb_0_io_rPort_2_output_0; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire [2:0] x283_lb_0_io_rPort_1_banks_1; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire [2:0] x283_lb_0_io_rPort_1_banks_0; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire  x283_lb_0_io_rPort_1_ofs_0; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire  x283_lb_0_io_rPort_1_en_0; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire  x283_lb_0_io_rPort_1_backpressure; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire [7:0] x283_lb_0_io_rPort_1_output_0; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire [2:0] x283_lb_0_io_rPort_0_banks_1; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire [2:0] x283_lb_0_io_rPort_0_banks_0; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire  x283_lb_0_io_rPort_0_ofs_0; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire  x283_lb_0_io_rPort_0_en_0; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire  x283_lb_0_io_rPort_0_backpressure; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire [7:0] x283_lb_0_io_rPort_0_output_0; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire [2:0] x283_lb_0_io_wPort_0_banks_1; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire [2:0] x283_lb_0_io_wPort_0_banks_0; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire  x283_lb_0_io_wPort_0_ofs_0; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire [7:0] x283_lb_0_io_wPort_0_data_0; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire  x283_lb_0_io_wPort_0_en_0; // @[m_x283_lb_0.scala 35:17:@20599.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@20679.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@20679.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@20679.4]
  wire [7:0] RetimeWrapper_io_in; // @[package.scala 93:22:@20679.4]
  wire [7:0] RetimeWrapper_io_out; // @[package.scala 93:22:@20679.4]
  wire  x297_sum_1_clock; // @[Math.scala 150:24:@20784.4]
  wire  x297_sum_1_reset; // @[Math.scala 150:24:@20784.4]
  wire [31:0] x297_sum_1_io_a; // @[Math.scala 150:24:@20784.4]
  wire [31:0] x297_sum_1_io_b; // @[Math.scala 150:24:@20784.4]
  wire  x297_sum_1_io_flow; // @[Math.scala 150:24:@20784.4]
  wire [31:0] x297_sum_1_io_result; // @[Math.scala 150:24:@20784.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@20794.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@20794.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@20794.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@20794.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@20794.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@20803.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@20803.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@20803.4]
  wire [31:0] RetimeWrapper_2_io_in; // @[package.scala 93:22:@20803.4]
  wire [31:0] RetimeWrapper_2_io_out; // @[package.scala 93:22:@20803.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@20812.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@20812.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@20812.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@20812.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@20812.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@20821.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@20821.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@20821.4]
  wire [31:0] RetimeWrapper_4_io_in; // @[package.scala 93:22:@20821.4]
  wire [31:0] RetimeWrapper_4_io_out; // @[package.scala 93:22:@20821.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@20832.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@20832.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@20832.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@20832.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@20832.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@20853.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@20853.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@20853.4]
  wire [31:0] RetimeWrapper_6_io_in; // @[package.scala 93:22:@20853.4]
  wire [31:0] RetimeWrapper_6_io_out; // @[package.scala 93:22:@20853.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@20869.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@20869.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@20869.4]
  wire [31:0] RetimeWrapper_7_io_in; // @[package.scala 93:22:@20869.4]
  wire [31:0] RetimeWrapper_7_io_out; // @[package.scala 93:22:@20869.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@20922.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@20922.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@20922.4]
  wire [31:0] RetimeWrapper_8_io_in; // @[package.scala 93:22:@20922.4]
  wire [31:0] RetimeWrapper_8_io_out; // @[package.scala 93:22:@20922.4]
  wire  x314_sum_1_clock; // @[Math.scala 150:24:@20931.4]
  wire  x314_sum_1_reset; // @[Math.scala 150:24:@20931.4]
  wire [31:0] x314_sum_1_io_a; // @[Math.scala 150:24:@20931.4]
  wire [31:0] x314_sum_1_io_b; // @[Math.scala 150:24:@20931.4]
  wire  x314_sum_1_io_flow; // @[Math.scala 150:24:@20931.4]
  wire [31:0] x314_sum_1_io_result; // @[Math.scala 150:24:@20931.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@20941.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@20941.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@20941.4]
  wire [31:0] RetimeWrapper_9_io_in; // @[package.scala 93:22:@20941.4]
  wire [31:0] RetimeWrapper_9_io_out; // @[package.scala 93:22:@20941.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@20950.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@20950.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@20950.4]
  wire [31:0] RetimeWrapper_10_io_in; // @[package.scala 93:22:@20950.4]
  wire [31:0] RetimeWrapper_10_io_out; // @[package.scala 93:22:@20950.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@20959.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@20959.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@20959.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@20959.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@20959.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@20968.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@20968.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@20968.4]
  wire [31:0] RetimeWrapper_12_io_in; // @[package.scala 93:22:@20968.4]
  wire [31:0] RetimeWrapper_12_io_out; // @[package.scala 93:22:@20968.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@20980.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@20980.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@20980.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@20980.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@20980.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@20999.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@20999.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@20999.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@20999.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@20999.4]
  wire  x323_rdcol_1_clock; // @[Math.scala 191:24:@21015.4]
  wire  x323_rdcol_1_reset; // @[Math.scala 191:24:@21015.4]
  wire [31:0] x323_rdcol_1_io_a; // @[Math.scala 191:24:@21015.4]
  wire [31:0] x323_rdcol_1_io_b; // @[Math.scala 191:24:@21015.4]
  wire  x323_rdcol_1_io_flow; // @[Math.scala 191:24:@21015.4]
  wire [31:0] x323_rdcol_1_io_result; // @[Math.scala 191:24:@21015.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@21032.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@21032.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@21032.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@21032.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@21032.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@21067.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@21067.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@21067.4]
  wire [31:0] RetimeWrapper_16_io_in; // @[package.scala 93:22:@21067.4]
  wire [31:0] RetimeWrapper_16_io_out; // @[package.scala 93:22:@21067.4]
  wire  x333_sum_1_clock; // @[Math.scala 150:24:@21078.4]
  wire  x333_sum_1_reset; // @[Math.scala 150:24:@21078.4]
  wire [31:0] x333_sum_1_io_a; // @[Math.scala 150:24:@21078.4]
  wire [31:0] x333_sum_1_io_b; // @[Math.scala 150:24:@21078.4]
  wire  x333_sum_1_io_flow; // @[Math.scala 150:24:@21078.4]
  wire [31:0] x333_sum_1_io_result; // @[Math.scala 150:24:@21078.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@21088.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@21088.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@21088.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@21088.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@21088.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@21097.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@21097.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@21097.4]
  wire [31:0] RetimeWrapper_18_io_in; // @[package.scala 93:22:@21097.4]
  wire [31:0] RetimeWrapper_18_io_out; // @[package.scala 93:22:@21097.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@21109.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@21109.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@21109.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@21109.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@21109.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@21128.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@21128.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@21128.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@21128.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@21128.4]
  wire  x342_rdcol_1_clock; // @[Math.scala 191:24:@21144.4]
  wire  x342_rdcol_1_reset; // @[Math.scala 191:24:@21144.4]
  wire [31:0] x342_rdcol_1_io_a; // @[Math.scala 191:24:@21144.4]
  wire [31:0] x342_rdcol_1_io_b; // @[Math.scala 191:24:@21144.4]
  wire  x342_rdcol_1_io_flow; // @[Math.scala 191:24:@21144.4]
  wire [31:0] x342_rdcol_1_io_result; // @[Math.scala 191:24:@21144.4]
  wire  x352_sum_1_clock; // @[Math.scala 150:24:@21187.4]
  wire  x352_sum_1_reset; // @[Math.scala 150:24:@21187.4]
  wire [31:0] x352_sum_1_io_a; // @[Math.scala 150:24:@21187.4]
  wire [31:0] x352_sum_1_io_b; // @[Math.scala 150:24:@21187.4]
  wire  x352_sum_1_io_flow; // @[Math.scala 150:24:@21187.4]
  wire [31:0] x352_sum_1_io_result; // @[Math.scala 150:24:@21187.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@21197.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@21197.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@21197.4]
  wire [31:0] RetimeWrapper_21_io_in; // @[package.scala 93:22:@21197.4]
  wire [31:0] RetimeWrapper_21_io_out; // @[package.scala 93:22:@21197.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@21206.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@21206.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@21206.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@21206.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@21206.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@21218.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@21218.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@21218.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@21218.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@21218.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@21237.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@21237.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@21237.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@21237.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@21237.4]
  wire  x361_rdrow_1_clock; // @[Math.scala 191:24:@21253.4]
  wire  x361_rdrow_1_reset; // @[Math.scala 191:24:@21253.4]
  wire [31:0] x361_rdrow_1_io_a; // @[Math.scala 191:24:@21253.4]
  wire [31:0] x361_rdrow_1_io_b; // @[Math.scala 191:24:@21253.4]
  wire  x361_rdrow_1_io_flow; // @[Math.scala 191:24:@21253.4]
  wire [31:0] x361_rdrow_1_io_result; // @[Math.scala 191:24:@21253.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@21270.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@21270.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@21270.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@21270.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@21270.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@21316.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@21316.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@21316.4]
  wire [31:0] RetimeWrapper_26_io_in; // @[package.scala 93:22:@21316.4]
  wire [31:0] RetimeWrapper_26_io_out; // @[package.scala 93:22:@21316.4]
  wire  x371_sum_1_clock; // @[Math.scala 150:24:@21325.4]
  wire  x371_sum_1_reset; // @[Math.scala 150:24:@21325.4]
  wire [31:0] x371_sum_1_io_a; // @[Math.scala 150:24:@21325.4]
  wire [31:0] x371_sum_1_io_b; // @[Math.scala 150:24:@21325.4]
  wire  x371_sum_1_io_flow; // @[Math.scala 150:24:@21325.4]
  wire [31:0] x371_sum_1_io_result; // @[Math.scala 150:24:@21325.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@21335.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@21335.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@21335.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@21335.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@21335.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@21344.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@21344.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@21344.4]
  wire [31:0] RetimeWrapper_28_io_in; // @[package.scala 93:22:@21344.4]
  wire [31:0] RetimeWrapper_28_io_out; // @[package.scala 93:22:@21344.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@21356.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@21356.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@21356.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@21356.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@21356.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@21375.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@21375.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@21375.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@21375.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@21375.4]
  wire  x388_sum_1_clock; // @[Math.scala 150:24:@21395.4]
  wire  x388_sum_1_reset; // @[Math.scala 150:24:@21395.4]
  wire [31:0] x388_sum_1_io_a; // @[Math.scala 150:24:@21395.4]
  wire [31:0] x388_sum_1_io_b; // @[Math.scala 150:24:@21395.4]
  wire  x388_sum_1_io_flow; // @[Math.scala 150:24:@21395.4]
  wire [31:0] x388_sum_1_io_result; // @[Math.scala 150:24:@21395.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@21405.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@21405.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@21405.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@21405.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@21405.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@21417.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@21417.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@21417.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@21417.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@21417.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@21436.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@21436.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@21436.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@21436.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@21436.4]
  wire  x405_sum_1_clock; // @[Math.scala 150:24:@21456.4]
  wire  x405_sum_1_reset; // @[Math.scala 150:24:@21456.4]
  wire [31:0] x405_sum_1_io_a; // @[Math.scala 150:24:@21456.4]
  wire [31:0] x405_sum_1_io_b; // @[Math.scala 150:24:@21456.4]
  wire  x405_sum_1_io_flow; // @[Math.scala 150:24:@21456.4]
  wire [31:0] x405_sum_1_io_result; // @[Math.scala 150:24:@21456.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@21466.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@21466.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@21466.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@21466.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@21466.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@21478.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@21478.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@21478.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@21478.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@21478.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@21497.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@21497.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@21497.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@21497.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@21497.4]
  wire  x414_rdrow_1_clock; // @[Math.scala 191:24:@21515.4]
  wire  x414_rdrow_1_reset; // @[Math.scala 191:24:@21515.4]
  wire [31:0] x414_rdrow_1_io_a; // @[Math.scala 191:24:@21515.4]
  wire [31:0] x414_rdrow_1_io_b; // @[Math.scala 191:24:@21515.4]
  wire  x414_rdrow_1_io_flow; // @[Math.scala 191:24:@21515.4]
  wire [31:0] x414_rdrow_1_io_result; // @[Math.scala 191:24:@21515.4]
  wire  x424_sum_1_clock; // @[Math.scala 150:24:@21569.4]
  wire  x424_sum_1_reset; // @[Math.scala 150:24:@21569.4]
  wire [31:0] x424_sum_1_io_a; // @[Math.scala 150:24:@21569.4]
  wire [31:0] x424_sum_1_io_b; // @[Math.scala 150:24:@21569.4]
  wire  x424_sum_1_io_flow; // @[Math.scala 150:24:@21569.4]
  wire [31:0] x424_sum_1_io_result; // @[Math.scala 150:24:@21569.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@21579.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@21579.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@21579.4]
  wire [31:0] RetimeWrapper_37_io_in; // @[package.scala 93:22:@21579.4]
  wire [31:0] RetimeWrapper_37_io_out; // @[package.scala 93:22:@21579.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@21588.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@21588.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@21588.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@21588.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@21588.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@21600.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@21600.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@21600.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@21600.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@21600.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@21619.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@21619.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@21619.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@21619.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@21619.4]
  wire  x441_sum_1_clock; // @[Math.scala 150:24:@21639.4]
  wire  x441_sum_1_reset; // @[Math.scala 150:24:@21639.4]
  wire [31:0] x441_sum_1_io_a; // @[Math.scala 150:24:@21639.4]
  wire [31:0] x441_sum_1_io_b; // @[Math.scala 150:24:@21639.4]
  wire  x441_sum_1_io_flow; // @[Math.scala 150:24:@21639.4]
  wire [31:0] x441_sum_1_io_result; // @[Math.scala 150:24:@21639.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@21649.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@21649.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@21649.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@21649.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@21649.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@21661.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@21661.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@21661.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@21661.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@21661.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@21680.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@21680.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@21680.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@21680.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@21680.4]
  wire  x458_sum_1_clock; // @[Math.scala 150:24:@21700.4]
  wire  x458_sum_1_reset; // @[Math.scala 150:24:@21700.4]
  wire [31:0] x458_sum_1_io_a; // @[Math.scala 150:24:@21700.4]
  wire [31:0] x458_sum_1_io_b; // @[Math.scala 150:24:@21700.4]
  wire  x458_sum_1_io_flow; // @[Math.scala 150:24:@21700.4]
  wire [31:0] x458_sum_1_io_result; // @[Math.scala 150:24:@21700.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@21710.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@21710.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@21710.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@21710.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@21710.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@21722.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@21722.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@21722.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@21722.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@21722.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@21741.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@21741.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@21741.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@21741.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@21741.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@21755.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@21755.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@21755.4]
  wire [7:0] RetimeWrapper_47_io_in; // @[package.scala 93:22:@21755.4]
  wire [7:0] RetimeWrapper_47_io_out; // @[package.scala 93:22:@21755.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@21769.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@21769.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@21769.4]
  wire [7:0] RetimeWrapper_48_io_in; // @[package.scala 93:22:@21769.4]
  wire [7:0] RetimeWrapper_48_io_out; // @[package.scala 93:22:@21769.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@21783.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@21783.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@21783.4]
  wire [7:0] RetimeWrapper_49_io_in; // @[package.scala 93:22:@21783.4]
  wire [7:0] RetimeWrapper_49_io_out; // @[package.scala 93:22:@21783.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@21797.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@21797.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@21797.4]
  wire [7:0] RetimeWrapper_50_io_in; // @[package.scala 93:22:@21797.4]
  wire [7:0] RetimeWrapper_50_io_out; // @[package.scala 93:22:@21797.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@21811.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@21811.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@21811.4]
  wire [7:0] RetimeWrapper_51_io_in; // @[package.scala 93:22:@21811.4]
  wire [7:0] RetimeWrapper_51_io_out; // @[package.scala 93:22:@21811.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@21825.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@21825.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@21825.4]
  wire [7:0] RetimeWrapper_52_io_in; // @[package.scala 93:22:@21825.4]
  wire [7:0] RetimeWrapper_52_io_out; // @[package.scala 93:22:@21825.4]
  wire [7:0] x472_x11_1_io_a; // @[Math.scala 150:24:@21834.4]
  wire [7:0] x472_x11_1_io_b; // @[Math.scala 150:24:@21834.4]
  wire [7:0] x472_x11_1_io_result; // @[Math.scala 150:24:@21834.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@21844.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@21844.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@21844.4]
  wire [7:0] RetimeWrapper_53_io_in; // @[package.scala 93:22:@21844.4]
  wire [7:0] RetimeWrapper_53_io_out; // @[package.scala 93:22:@21844.4]
  wire [7:0] x473_x12_1_io_a; // @[Math.scala 150:24:@21853.4]
  wire [7:0] x473_x12_1_io_b; // @[Math.scala 150:24:@21853.4]
  wire [7:0] x473_x12_1_io_result; // @[Math.scala 150:24:@21853.4]
  wire [7:0] x474_x11_1_io_a; // @[Math.scala 150:24:@21863.4]
  wire [7:0] x474_x11_1_io_b; // @[Math.scala 150:24:@21863.4]
  wire [7:0] x474_x11_1_io_result; // @[Math.scala 150:24:@21863.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@21873.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@21873.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@21873.4]
  wire [7:0] RetimeWrapper_54_io_in; // @[package.scala 93:22:@21873.4]
  wire [7:0] RetimeWrapper_54_io_out; // @[package.scala 93:22:@21873.4]
  wire [7:0] x475_x12_1_io_a; // @[Math.scala 150:24:@21884.4]
  wire [7:0] x475_x12_1_io_b; // @[Math.scala 150:24:@21884.4]
  wire [7:0] x475_x12_1_io_result; // @[Math.scala 150:24:@21884.4]
  wire [7:0] x476_x11_1_io_a; // @[Math.scala 150:24:@21894.4]
  wire [7:0] x476_x11_1_io_b; // @[Math.scala 150:24:@21894.4]
  wire [7:0] x476_x11_1_io_result; // @[Math.scala 150:24:@21894.4]
  wire [7:0] x477_x12_1_io_a; // @[Math.scala 150:24:@21904.4]
  wire [7:0] x477_x12_1_io_b; // @[Math.scala 150:24:@21904.4]
  wire [7:0] x477_x12_1_io_result; // @[Math.scala 150:24:@21904.4]
  wire  x478_x11_1_clock; // @[Math.scala 150:24:@21914.4]
  wire  x478_x11_1_reset; // @[Math.scala 150:24:@21914.4]
  wire [7:0] x478_x11_1_io_a; // @[Math.scala 150:24:@21914.4]
  wire [7:0] x478_x11_1_io_b; // @[Math.scala 150:24:@21914.4]
  wire  x478_x11_1_io_flow; // @[Math.scala 150:24:@21914.4]
  wire [7:0] x478_x11_1_io_result; // @[Math.scala 150:24:@21914.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@21924.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@21924.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@21924.4]
  wire [7:0] RetimeWrapper_55_io_in; // @[package.scala 93:22:@21924.4]
  wire [7:0] RetimeWrapper_55_io_out; // @[package.scala 93:22:@21924.4]
  wire [7:0] x479_sum_1_io_a; // @[Math.scala 150:24:@21933.4]
  wire [7:0] x479_sum_1_io_b; // @[Math.scala 150:24:@21933.4]
  wire [7:0] x479_sum_1_io_result; // @[Math.scala 150:24:@21933.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@21954.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@21954.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@21954.4]
  wire [7:0] RetimeWrapper_56_io_in; // @[package.scala 93:22:@21954.4]
  wire [7:0] RetimeWrapper_56_io_out; // @[package.scala 93:22:@21954.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@21963.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@21963.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@21963.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@21963.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@21963.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@21972.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@21972.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@21972.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@21972.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@21972.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@21981.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@21981.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@21981.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@21981.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@21981.4]
  wire  b281; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 62:18:@20597.4]
  wire  b282; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 63:18:@20598.4]
  wire  _T_206; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 68:30:@20667.4]
  wire  _T_207; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 68:37:@20668.4]
  wire  _T_211; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 70:76:@20673.4]
  wire  _T_212; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 70:62:@20674.4]
  wire  _T_214; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 70:101:@20675.4]
  wire [31:0] b279_number; // @[Math.scala 712:22:@20582.4 Math.scala 713:14:@20583.4]
  wire [31:0] _T_240; // @[Math.scala 499:52:@20698.4]
  wire  x288; // @[Math.scala 499:44:@20706.4]
  wire  x289; // @[Math.scala 499:44:@20713.4]
  wire  x290; // @[Math.scala 499:44:@20720.4]
  wire [31:0] _T_287; // @[Mux.scala 19:72:@20732.4]
  wire [31:0] _T_289; // @[Mux.scala 19:72:@20733.4]
  wire [31:0] _T_291; // @[Mux.scala 19:72:@20734.4]
  wire [31:0] _T_293; // @[Mux.scala 19:72:@20736.4]
  wire [31:0] x291_number; // @[Mux.scala 19:72:@20737.4]
  wire [31:0] _T_305; // @[Math.scala 406:49:@20747.4]
  wire [31:0] _T_307; // @[Math.scala 406:56:@20749.4]
  wire [31:0] _T_308; // @[Math.scala 406:56:@20750.4]
  wire [31:0] b280_number; // @[Math.scala 712:22:@20594.4 Math.scala 713:14:@20595.4]
  wire [31:0] _T_317; // @[Math.scala 406:49:@20758.4]
  wire [31:0] _T_319; // @[Math.scala 406:56:@20760.4]
  wire [31:0] _T_320; // @[Math.scala 406:56:@20761.4]
  wire  _T_325; // @[FixedPoint.scala 50:25:@20767.4]
  wire [1:0] _T_329; // @[Bitwise.scala 72:12:@20769.4]
  wire [29:0] _T_330; // @[FixedPoint.scala 18:52:@20770.4]
  wire  _T_335; // @[FixedPoint.scala 50:25:@20776.4]
  wire [1:0] _T_339; // @[Bitwise.scala 72:12:@20778.4]
  wire [29:0] _T_340; // @[FixedPoint.scala 18:52:@20779.4]
  wire  _T_358; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 113:101:@20829.4]
  wire  _T_362; // @[package.scala 96:25:@20837.4 package.scala 96:25:@20838.4]
  wire  _T_364; // @[implicits.scala 55:10:@20839.4]
  wire  _T_365; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 113:118:@20840.4]
  wire  _T_367; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 113:205:@20842.4]
  wire  _T_368; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 113:224:@20843.4]
  wire  x588_b281_D1; // @[package.scala 96:25:@20817.4 package.scala 96:25:@20818.4]
  wire  _T_369; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 113:250:@20844.4]
  wire  x586_b282_D1; // @[package.scala 96:25:@20799.4 package.scala 96:25:@20800.4]
  wire [31:0] x590_b279_D3_number; // @[package.scala 96:25:@20858.4 package.scala 96:25:@20859.4]
  wire [31:0] _T_379; // @[Math.scala 465:37:@20864.4]
  wire  x304; // @[Math.scala 465:44:@20866.4]
  wire [31:0] x591_b280_D3_number; // @[package.scala 96:25:@20874.4 package.scala 96:25:@20875.4]
  wire [31:0] _T_390; // @[Math.scala 465:37:@20880.4]
  wire  x305; // @[Math.scala 465:44:@20882.4]
  wire  x306; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 124:24:@20885.4]
  wire [31:0] _T_406; // @[Math.scala 406:56:@20896.4]
  wire [31:0] _T_407; // @[Math.scala 406:56:@20897.4]
  wire [31:0] x549_number; // @[implicits.scala 133:21:@20898.4]
  wire [31:0] _T_416; // @[Math.scala 406:49:@20905.4]
  wire [31:0] _T_418; // @[Math.scala 406:56:@20907.4]
  wire [31:0] _T_419; // @[Math.scala 406:56:@20908.4]
  wire  _T_424; // @[FixedPoint.scala 50:25:@20914.4]
  wire [1:0] _T_428; // @[Bitwise.scala 72:12:@20916.4]
  wire [29:0] _T_429; // @[FixedPoint.scala 18:52:@20917.4]
  wire  _T_460; // @[package.scala 96:25:@20985.4 package.scala 96:25:@20986.4]
  wire  _T_462; // @[implicits.scala 55:10:@20987.4]
  wire  _T_463; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 149:146:@20988.4]
  wire  x595_x307_D2; // @[package.scala 96:25:@20964.4 package.scala 96:25:@20965.4]
  wire  x597_x306_D4; // @[package.scala 96:25:@21004.4 package.scala 96:25:@21005.4]
  wire [7:0] x319_rd_0_number; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 145:29:@20976.4 sm_x485_inr_Foreach_SAMPLER_BOX.scala 149:274:@20995.4]
  wire [31:0] x323_rdcol_number; // @[Math.scala 195:22:@21021.4 Math.scala 196:14:@21022.4]
  wire [31:0] _T_487; // @[Math.scala 465:37:@21027.4]
  wire  x324; // @[Math.scala 465:44:@21029.4]
  wire  x598_x304_D1; // @[package.scala 96:25:@21037.4 package.scala 96:25:@21038.4]
  wire  x325; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 163:24:@21041.4]
  wire [31:0] _T_506; // @[Math.scala 406:56:@21052.4]
  wire [31:0] _T_507; // @[Math.scala 406:56:@21053.4]
  wire  _T_512; // @[FixedPoint.scala 50:25:@21059.4]
  wire [1:0] _T_516; // @[Bitwise.scala 72:12:@21061.4]
  wire [29:0] _T_517; // @[FixedPoint.scala 18:52:@21062.4]
  wire  _T_544; // @[package.scala 96:25:@21114.4 package.scala 96:25:@21115.4]
  wire  _T_546; // @[implicits.scala 55:10:@21116.4]
  wire  _T_547; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 190:194:@21117.4]
  wire  x600_x326_D1; // @[package.scala 96:25:@21093.4 package.scala 96:25:@21094.4]
  wire  x602_x325_D3; // @[package.scala 96:25:@21133.4 package.scala 96:25:@21134.4]
  wire [7:0] x338_rd_0_number; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 186:29:@21105.4 sm_x485_inr_Foreach_SAMPLER_BOX.scala 190:322:@21124.4]
  wire [31:0] x342_rdcol_number; // @[Math.scala 195:22:@21150.4 Math.scala 196:14:@21151.4]
  wire [31:0] _T_571; // @[Math.scala 465:37:@21156.4]
  wire  x343; // @[Math.scala 465:44:@21158.4]
  wire  x344; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 202:59:@21161.4]
  wire [31:0] _T_587; // @[Math.scala 406:56:@21172.4]
  wire [31:0] _T_588; // @[Math.scala 406:56:@21173.4]
  wire  _T_593; // @[FixedPoint.scala 50:25:@21179.4]
  wire [1:0] _T_597; // @[Bitwise.scala 72:12:@21181.4]
  wire [29:0] _T_598; // @[FixedPoint.scala 18:52:@21182.4]
  wire  _T_620; // @[package.scala 96:25:@21223.4 package.scala 96:25:@21224.4]
  wire  _T_622; // @[implicits.scala 55:10:@21225.4]
  wire  _T_623; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 219:194:@21226.4]
  wire  x604_x345_D1; // @[package.scala 96:25:@21211.4 package.scala 96:25:@21212.4]
  wire  x605_x344_D3; // @[package.scala 96:25:@21242.4 package.scala 96:25:@21243.4]
  wire [7:0] x357_rd_0_number; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 215:29:@21214.4 sm_x485_inr_Foreach_SAMPLER_BOX.scala 219:322:@21233.4]
  wire [31:0] x361_rdrow_number; // @[Math.scala 195:22:@21259.4 Math.scala 196:14:@21260.4]
  wire [31:0] _T_647; // @[Math.scala 465:37:@21265.4]
  wire  x362; // @[Math.scala 465:44:@21267.4]
  wire  x606_x305_D1; // @[package.scala 96:25:@21275.4 package.scala 96:25:@21276.4]
  wire  x363; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 233:24:@21279.4]
  wire [31:0] _T_666; // @[Math.scala 406:56:@21290.4]
  wire [31:0] _T_667; // @[Math.scala 406:56:@21291.4]
  wire [31:0] x558_number; // @[implicits.scala 133:21:@21292.4]
  wire [31:0] _T_676; // @[Math.scala 406:49:@21299.4]
  wire [31:0] _T_678; // @[Math.scala 406:56:@21301.4]
  wire [31:0] _T_679; // @[Math.scala 406:56:@21302.4]
  wire  _T_684; // @[FixedPoint.scala 50:25:@21308.4]
  wire [1:0] _T_688; // @[Bitwise.scala 72:12:@21310.4]
  wire [29:0] _T_689; // @[FixedPoint.scala 18:52:@21311.4]
  wire  _T_714; // @[package.scala 96:25:@21361.4 package.scala 96:25:@21362.4]
  wire  _T_716; // @[implicits.scala 55:10:@21363.4]
  wire  _T_717; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 254:194:@21364.4]
  wire  x608_x364_D1; // @[package.scala 96:25:@21340.4 package.scala 96:25:@21341.4]
  wire  x610_x363_D3; // @[package.scala 96:25:@21380.4 package.scala 96:25:@21381.4]
  wire [7:0] x376_rd_0_number; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 250:29:@21352.4 sm_x485_inr_Foreach_SAMPLER_BOX.scala 254:322:@21371.4]
  wire  x380; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 262:24:@21389.4]
  wire  _T_750; // @[package.scala 96:25:@21422.4 package.scala 96:25:@21423.4]
  wire  _T_752; // @[implicits.scala 55:10:@21424.4]
  wire  _T_753; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 273:194:@21425.4]
  wire  x611_x381_D1; // @[package.scala 96:25:@21410.4 package.scala 96:25:@21411.4]
  wire  x612_x380_D3; // @[package.scala 96:25:@21441.4 package.scala 96:25:@21442.4]
  wire [7:0] x393_rd_0_number; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 269:29:@21413.4 sm_x485_inr_Foreach_SAMPLER_BOX.scala 273:322:@21432.4]
  wire  x397; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 281:24:@21450.4]
  wire  _T_786; // @[package.scala 96:25:@21483.4 package.scala 96:25:@21484.4]
  wire  _T_788; // @[implicits.scala 55:10:@21485.4]
  wire  _T_789; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 292:194:@21486.4]
  wire  x613_x398_D1; // @[package.scala 96:25:@21471.4 package.scala 96:25:@21472.4]
  wire  x614_x397_D3; // @[package.scala 96:25:@21502.4 package.scala 96:25:@21503.4]
  wire [7:0] x410_rd_0_number; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 288:29:@21474.4 sm_x485_inr_Foreach_SAMPLER_BOX.scala 292:322:@21493.4]
  wire [31:0] x414_rdrow_number; // @[Math.scala 195:22:@21521.4 Math.scala 196:14:@21522.4]
  wire [31:0] _T_815; // @[Math.scala 465:37:@21527.4]
  wire  x415; // @[Math.scala 465:44:@21529.4]
  wire  x416; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 312:24:@21532.4]
  wire [31:0] _T_831; // @[Math.scala 406:56:@21543.4]
  wire [31:0] _T_832; // @[Math.scala 406:56:@21544.4]
  wire [31:0] x567_number; // @[implicits.scala 133:21:@21545.4]
  wire [31:0] _T_841; // @[Math.scala 406:49:@21552.4]
  wire [31:0] _T_843; // @[Math.scala 406:56:@21554.4]
  wire [31:0] _T_844; // @[Math.scala 406:56:@21555.4]
  wire  _T_849; // @[FixedPoint.scala 50:25:@21561.4]
  wire [1:0] _T_853; // @[Bitwise.scala 72:12:@21563.4]
  wire [29:0] _T_854; // @[FixedPoint.scala 18:52:@21564.4]
  wire  _T_876; // @[package.scala 96:25:@21605.4 package.scala 96:25:@21606.4]
  wire  _T_878; // @[implicits.scala 55:10:@21607.4]
  wire  _T_879; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 331:194:@21608.4]
  wire  x616_x417_D1; // @[package.scala 96:25:@21593.4 package.scala 96:25:@21594.4]
  wire  x617_x416_D3; // @[package.scala 96:25:@21624.4 package.scala 96:25:@21625.4]
  wire [7:0] x429_rd_0_number; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 327:29:@21596.4 sm_x485_inr_Foreach_SAMPLER_BOX.scala 331:322:@21615.4]
  wire  x433; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 339:24:@21633.4]
  wire  _T_912; // @[package.scala 96:25:@21666.4 package.scala 96:25:@21667.4]
  wire  _T_914; // @[implicits.scala 55:10:@21668.4]
  wire  _T_915; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 350:194:@21669.4]
  wire  x618_x434_D1; // @[package.scala 96:25:@21654.4 package.scala 96:25:@21655.4]
  wire  x619_x433_D3; // @[package.scala 96:25:@21685.4 package.scala 96:25:@21686.4]
  wire [7:0] x446_rd_0_number; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 346:29:@21657.4 sm_x485_inr_Foreach_SAMPLER_BOX.scala 350:322:@21676.4]
  wire  x450; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 358:24:@21694.4]
  wire  _T_948; // @[package.scala 96:25:@21727.4 package.scala 96:25:@21728.4]
  wire  _T_950; // @[implicits.scala 55:10:@21729.4]
  wire  _T_951; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 369:194:@21730.4]
  wire  x620_x451_D1; // @[package.scala 96:25:@21715.4 package.scala 96:25:@21716.4]
  wire  x621_x450_D3; // @[package.scala 96:25:@21746.4 package.scala 96:25:@21747.4]
  wire [7:0] x463_rd_0_number; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 365:29:@21718.4 sm_x485_inr_Foreach_SAMPLER_BOX.scala 369:322:@21737.4]
  wire [7:0] x622_x577_D1_number; // @[package.scala 96:25:@21760.4 package.scala 96:25:@21761.4]
  wire [8:0] _GEN_0; // @[Math.scala 450:32:@21765.4]
  wire [8:0] _T_969; // @[Math.scala 450:32:@21765.4]
  wire [7:0] x623_x579_D1_number; // @[package.scala 96:25:@21774.4 package.scala 96:25:@21775.4]
  wire [8:0] _GEN_1; // @[Math.scala 450:32:@21779.4]
  wire [8:0] _T_976; // @[Math.scala 450:32:@21779.4]
  wire [7:0] x624_x580_D1_number; // @[package.scala 96:25:@21788.4 package.scala 96:25:@21789.4]
  wire [9:0] _GEN_2; // @[Math.scala 450:32:@21793.4]
  wire [9:0] _T_983; // @[Math.scala 450:32:@21793.4]
  wire [7:0] x625_x581_D1_number; // @[package.scala 96:25:@21802.4 package.scala 96:25:@21803.4]
  wire [8:0] _GEN_3; // @[Math.scala 450:32:@21807.4]
  wire [8:0] _T_990; // @[Math.scala 450:32:@21807.4]
  wire [7:0] x626_x583_D1_number; // @[package.scala 96:25:@21816.4 package.scala 96:25:@21817.4]
  wire [8:0] _GEN_4; // @[Math.scala 450:32:@21821.4]
  wire [8:0] _T_997; // @[Math.scala 450:32:@21821.4]
  wire [7:0] x479_sum_number; // @[Math.scala 154:22:@21939.4 Math.scala 155:14:@21940.4]
  wire [3:0] _T_1044; // @[FixedPoint.scala 18:52:@21945.4]
  wire  _T_1065; // @[package.scala 96:25:@21986.4 package.scala 96:25:@21987.4]
  wire  _T_1067; // @[implicits.scala 55:10:@21988.4]
  wire  x632_b281_D12; // @[package.scala 96:25:@21977.4 package.scala 96:25:@21978.4]
  wire  _T_1068; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 439:116:@21989.4]
  wire  x631_b282_D12; // @[package.scala 96:25:@21968.4 package.scala 96:25:@21969.4]
  wire  _T_1069; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 439:122:@21990.4]
  wire [31:0] x297_sum_number; // @[Math.scala 154:22:@20790.4 Math.scala 155:14:@20791.4]
  wire [31:0] x587_x548_D1_number; // @[package.scala 96:25:@20808.4 package.scala 96:25:@20809.4]
  wire [31:0] x589_x547_D1_number; // @[package.scala 96:25:@20826.4 package.scala 96:25:@20827.4]
  wire [31:0] x593_x314_sum_D1_number; // @[package.scala 96:25:@20946.4 package.scala 96:25:@20947.4]
  wire [31:0] x594_x548_D5_number; // @[package.scala 96:25:@20955.4 package.scala 96:25:@20956.4]
  wire [31:0] x596_x550_D2_number; // @[package.scala 96:25:@20973.4 package.scala 96:25:@20974.4]
  wire [31:0] x333_sum_number; // @[Math.scala 154:22:@21084.4 Math.scala 155:14:@21085.4]
  wire [31:0] x601_x554_D1_number; // @[package.scala 96:25:@21102.4 package.scala 96:25:@21103.4]
  wire [31:0] x352_sum_number; // @[Math.scala 154:22:@21193.4 Math.scala 155:14:@21194.4]
  wire [31:0] x603_x557_D1_number; // @[package.scala 96:25:@21202.4 package.scala 96:25:@21203.4]
  wire [31:0] x371_sum_number; // @[Math.scala 154:22:@21331.4 Math.scala 155:14:@21332.4]
  wire [31:0] x609_x559_D1_number; // @[package.scala 96:25:@21349.4 package.scala 96:25:@21350.4]
  wire [31:0] x388_sum_number; // @[Math.scala 154:22:@21401.4 Math.scala 155:14:@21402.4]
  wire [31:0] x405_sum_number; // @[Math.scala 154:22:@21462.4 Math.scala 155:14:@21463.4]
  wire [31:0] x424_sum_number; // @[Math.scala 154:22:@21575.4 Math.scala 155:14:@21576.4]
  wire [31:0] x615_x568_D1_number; // @[package.scala 96:25:@21584.4 package.scala 96:25:@21585.4]
  wire [31:0] x441_sum_number; // @[Math.scala 154:22:@21645.4 Math.scala 155:14:@21646.4]
  wire [31:0] x458_sum_number; // @[Math.scala 154:22:@21706.4 Math.scala 155:14:@21707.4]
  _ _ ( // @[Math.scala 709:24:@20577.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 709:24:@20589.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  x283_lb_0 x283_lb_0 ( // @[m_x283_lb_0.scala 35:17:@20599.4]
    .clock(x283_lb_0_clock),
    .reset(x283_lb_0_reset),
    .io_rPort_8_banks_1(x283_lb_0_io_rPort_8_banks_1),
    .io_rPort_8_banks_0(x283_lb_0_io_rPort_8_banks_0),
    .io_rPort_8_ofs_0(x283_lb_0_io_rPort_8_ofs_0),
    .io_rPort_8_en_0(x283_lb_0_io_rPort_8_en_0),
    .io_rPort_8_backpressure(x283_lb_0_io_rPort_8_backpressure),
    .io_rPort_8_output_0(x283_lb_0_io_rPort_8_output_0),
    .io_rPort_7_banks_1(x283_lb_0_io_rPort_7_banks_1),
    .io_rPort_7_banks_0(x283_lb_0_io_rPort_7_banks_0),
    .io_rPort_7_ofs_0(x283_lb_0_io_rPort_7_ofs_0),
    .io_rPort_7_en_0(x283_lb_0_io_rPort_7_en_0),
    .io_rPort_7_backpressure(x283_lb_0_io_rPort_7_backpressure),
    .io_rPort_7_output_0(x283_lb_0_io_rPort_7_output_0),
    .io_rPort_6_banks_1(x283_lb_0_io_rPort_6_banks_1),
    .io_rPort_6_banks_0(x283_lb_0_io_rPort_6_banks_0),
    .io_rPort_6_ofs_0(x283_lb_0_io_rPort_6_ofs_0),
    .io_rPort_6_en_0(x283_lb_0_io_rPort_6_en_0),
    .io_rPort_6_backpressure(x283_lb_0_io_rPort_6_backpressure),
    .io_rPort_6_output_0(x283_lb_0_io_rPort_6_output_0),
    .io_rPort_5_banks_1(x283_lb_0_io_rPort_5_banks_1),
    .io_rPort_5_banks_0(x283_lb_0_io_rPort_5_banks_0),
    .io_rPort_5_ofs_0(x283_lb_0_io_rPort_5_ofs_0),
    .io_rPort_5_en_0(x283_lb_0_io_rPort_5_en_0),
    .io_rPort_5_backpressure(x283_lb_0_io_rPort_5_backpressure),
    .io_rPort_5_output_0(x283_lb_0_io_rPort_5_output_0),
    .io_rPort_4_banks_1(x283_lb_0_io_rPort_4_banks_1),
    .io_rPort_4_banks_0(x283_lb_0_io_rPort_4_banks_0),
    .io_rPort_4_ofs_0(x283_lb_0_io_rPort_4_ofs_0),
    .io_rPort_4_en_0(x283_lb_0_io_rPort_4_en_0),
    .io_rPort_4_backpressure(x283_lb_0_io_rPort_4_backpressure),
    .io_rPort_4_output_0(x283_lb_0_io_rPort_4_output_0),
    .io_rPort_3_banks_1(x283_lb_0_io_rPort_3_banks_1),
    .io_rPort_3_banks_0(x283_lb_0_io_rPort_3_banks_0),
    .io_rPort_3_ofs_0(x283_lb_0_io_rPort_3_ofs_0),
    .io_rPort_3_en_0(x283_lb_0_io_rPort_3_en_0),
    .io_rPort_3_backpressure(x283_lb_0_io_rPort_3_backpressure),
    .io_rPort_3_output_0(x283_lb_0_io_rPort_3_output_0),
    .io_rPort_2_banks_1(x283_lb_0_io_rPort_2_banks_1),
    .io_rPort_2_banks_0(x283_lb_0_io_rPort_2_banks_0),
    .io_rPort_2_ofs_0(x283_lb_0_io_rPort_2_ofs_0),
    .io_rPort_2_en_0(x283_lb_0_io_rPort_2_en_0),
    .io_rPort_2_backpressure(x283_lb_0_io_rPort_2_backpressure),
    .io_rPort_2_output_0(x283_lb_0_io_rPort_2_output_0),
    .io_rPort_1_banks_1(x283_lb_0_io_rPort_1_banks_1),
    .io_rPort_1_banks_0(x283_lb_0_io_rPort_1_banks_0),
    .io_rPort_1_ofs_0(x283_lb_0_io_rPort_1_ofs_0),
    .io_rPort_1_en_0(x283_lb_0_io_rPort_1_en_0),
    .io_rPort_1_backpressure(x283_lb_0_io_rPort_1_backpressure),
    .io_rPort_1_output_0(x283_lb_0_io_rPort_1_output_0),
    .io_rPort_0_banks_1(x283_lb_0_io_rPort_0_banks_1),
    .io_rPort_0_banks_0(x283_lb_0_io_rPort_0_banks_0),
    .io_rPort_0_ofs_0(x283_lb_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x283_lb_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x283_lb_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x283_lb_0_io_rPort_0_output_0),
    .io_wPort_0_banks_1(x283_lb_0_io_wPort_0_banks_1),
    .io_wPort_0_banks_0(x283_lb_0_io_wPort_0_banks_0),
    .io_wPort_0_ofs_0(x283_lb_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x283_lb_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x283_lb_0_io_wPort_0_en_0)
  );
  RetimeWrapper_21 RetimeWrapper ( // @[package.scala 93:22:@20679.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x297_sum x297_sum_1 ( // @[Math.scala 150:24:@20784.4]
    .clock(x297_sum_1_clock),
    .reset(x297_sum_1_reset),
    .io_a(x297_sum_1_io_a),
    .io_b(x297_sum_1_io_b),
    .io_flow(x297_sum_1_io_flow),
    .io_result(x297_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@20794.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_197 RetimeWrapper_2 ( // @[package.scala 93:22:@20803.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@20812.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_197 RetimeWrapper_4 ( // @[package.scala 93:22:@20821.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@20832.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_203 RetimeWrapper_6 ( // @[package.scala 93:22:@20853.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_203 RetimeWrapper_7 ( // @[package.scala 93:22:@20869.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_203 RetimeWrapper_8 ( // @[package.scala 93:22:@20922.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  x297_sum x314_sum_1 ( // @[Math.scala 150:24:@20931.4]
    .clock(x314_sum_1_clock),
    .reset(x314_sum_1_reset),
    .io_a(x314_sum_1_io_a),
    .io_b(x314_sum_1_io_b),
    .io_flow(x314_sum_1_io_flow),
    .io_result(x314_sum_1_io_result)
  );
  RetimeWrapper_197 RetimeWrapper_9 ( // @[package.scala 93:22:@20941.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_208 RetimeWrapper_10 ( // @[package.scala 93:22:@20950.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_11 ( // @[package.scala 93:22:@20959.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_210 RetimeWrapper_12 ( // @[package.scala 93:22:@20968.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_211 RetimeWrapper_13 ( // @[package.scala 93:22:@20980.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_212 RetimeWrapper_14 ( // @[package.scala 93:22:@20999.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  x323_rdcol x323_rdcol_1 ( // @[Math.scala 191:24:@21015.4]
    .clock(x323_rdcol_1_clock),
    .reset(x323_rdcol_1_reset),
    .io_a(x323_rdcol_1_io_a),
    .io_b(x323_rdcol_1_io_b),
    .io_flow(x323_rdcol_1_io_flow),
    .io_result(x323_rdcol_1_io_result)
  );
  RetimeWrapper RetimeWrapper_15 ( // @[package.scala 93:22:@21032.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_197 RetimeWrapper_16 ( // @[package.scala 93:22:@21067.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  x297_sum x333_sum_1 ( // @[Math.scala 150:24:@21078.4]
    .clock(x333_sum_1_clock),
    .reset(x333_sum_1_reset),
    .io_a(x333_sum_1_io_a),
    .io_b(x333_sum_1_io_b),
    .io_flow(x333_sum_1_io_flow),
    .io_result(x333_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_17 ( // @[package.scala 93:22:@21088.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_197 RetimeWrapper_18 ( // @[package.scala 93:22:@21097.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_211 RetimeWrapper_19 ( // @[package.scala 93:22:@21109.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_220 RetimeWrapper_20 ( // @[package.scala 93:22:@21128.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  x323_rdcol x342_rdcol_1 ( // @[Math.scala 191:24:@21144.4]
    .clock(x342_rdcol_1_clock),
    .reset(x342_rdcol_1_reset),
    .io_a(x342_rdcol_1_io_a),
    .io_b(x342_rdcol_1_io_b),
    .io_flow(x342_rdcol_1_io_flow),
    .io_result(x342_rdcol_1_io_result)
  );
  x297_sum x352_sum_1 ( // @[Math.scala 150:24:@21187.4]
    .clock(x352_sum_1_clock),
    .reset(x352_sum_1_reset),
    .io_a(x352_sum_1_io_a),
    .io_b(x352_sum_1_io_b),
    .io_flow(x352_sum_1_io_flow),
    .io_result(x352_sum_1_io_result)
  );
  RetimeWrapper_197 RetimeWrapper_21 ( // @[package.scala 93:22:@21197.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper RetimeWrapper_22 ( // @[package.scala 93:22:@21206.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_211 RetimeWrapper_23 ( // @[package.scala 93:22:@21218.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_220 RetimeWrapper_24 ( // @[package.scala 93:22:@21237.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  x323_rdcol x361_rdrow_1 ( // @[Math.scala 191:24:@21253.4]
    .clock(x361_rdrow_1_clock),
    .reset(x361_rdrow_1_reset),
    .io_a(x361_rdrow_1_io_a),
    .io_b(x361_rdrow_1_io_b),
    .io_flow(x361_rdrow_1_io_flow),
    .io_result(x361_rdrow_1_io_result)
  );
  RetimeWrapper RetimeWrapper_25 ( // @[package.scala 93:22:@21270.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_229 RetimeWrapper_26 ( // @[package.scala 93:22:@21316.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  x297_sum x371_sum_1 ( // @[Math.scala 150:24:@21325.4]
    .clock(x371_sum_1_clock),
    .reset(x371_sum_1_reset),
    .io_a(x371_sum_1_io_a),
    .io_b(x371_sum_1_io_b),
    .io_flow(x371_sum_1_io_flow),
    .io_result(x371_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_27 ( // @[package.scala 93:22:@21335.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_197 RetimeWrapper_28 ( // @[package.scala 93:22:@21344.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_211 RetimeWrapper_29 ( // @[package.scala 93:22:@21356.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_220 RetimeWrapper_30 ( // @[package.scala 93:22:@21375.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  x297_sum x388_sum_1 ( // @[Math.scala 150:24:@21395.4]
    .clock(x388_sum_1_clock),
    .reset(x388_sum_1_reset),
    .io_a(x388_sum_1_io_a),
    .io_b(x388_sum_1_io_b),
    .io_flow(x388_sum_1_io_flow),
    .io_result(x388_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_31 ( // @[package.scala 93:22:@21405.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_211 RetimeWrapper_32 ( // @[package.scala 93:22:@21417.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_220 RetimeWrapper_33 ( // @[package.scala 93:22:@21436.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  x297_sum x405_sum_1 ( // @[Math.scala 150:24:@21456.4]
    .clock(x405_sum_1_clock),
    .reset(x405_sum_1_reset),
    .io_a(x405_sum_1_io_a),
    .io_b(x405_sum_1_io_b),
    .io_flow(x405_sum_1_io_flow),
    .io_result(x405_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_34 ( // @[package.scala 93:22:@21466.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_211 RetimeWrapper_35 ( // @[package.scala 93:22:@21478.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_220 RetimeWrapper_36 ( // @[package.scala 93:22:@21497.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  x323_rdcol x414_rdrow_1 ( // @[Math.scala 191:24:@21515.4]
    .clock(x414_rdrow_1_clock),
    .reset(x414_rdrow_1_reset),
    .io_a(x414_rdrow_1_io_a),
    .io_b(x414_rdrow_1_io_b),
    .io_flow(x414_rdrow_1_io_flow),
    .io_result(x414_rdrow_1_io_result)
  );
  x297_sum x424_sum_1 ( // @[Math.scala 150:24:@21569.4]
    .clock(x424_sum_1_clock),
    .reset(x424_sum_1_reset),
    .io_a(x424_sum_1_io_a),
    .io_b(x424_sum_1_io_b),
    .io_flow(x424_sum_1_io_flow),
    .io_result(x424_sum_1_io_result)
  );
  RetimeWrapper_197 RetimeWrapper_37 ( // @[package.scala 93:22:@21579.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper RetimeWrapper_38 ( // @[package.scala 93:22:@21588.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_211 RetimeWrapper_39 ( // @[package.scala 93:22:@21600.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_220 RetimeWrapper_40 ( // @[package.scala 93:22:@21619.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  x297_sum x441_sum_1 ( // @[Math.scala 150:24:@21639.4]
    .clock(x441_sum_1_clock),
    .reset(x441_sum_1_reset),
    .io_a(x441_sum_1_io_a),
    .io_b(x441_sum_1_io_b),
    .io_flow(x441_sum_1_io_flow),
    .io_result(x441_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_41 ( // @[package.scala 93:22:@21649.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_211 RetimeWrapper_42 ( // @[package.scala 93:22:@21661.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_220 RetimeWrapper_43 ( // @[package.scala 93:22:@21680.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  x297_sum x458_sum_1 ( // @[Math.scala 150:24:@21700.4]
    .clock(x458_sum_1_clock),
    .reset(x458_sum_1_reset),
    .io_a(x458_sum_1_io_a),
    .io_b(x458_sum_1_io_b),
    .io_flow(x458_sum_1_io_flow),
    .io_result(x458_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_44 ( // @[package.scala 93:22:@21710.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_211 RetimeWrapper_45 ( // @[package.scala 93:22:@21722.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_220 RetimeWrapper_46 ( // @[package.scala 93:22:@21741.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_47 ( // @[package.scala 93:22:@21755.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_48 ( // @[package.scala 93:22:@21769.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_49 ( // @[package.scala 93:22:@21783.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_50 ( // @[package.scala 93:22:@21797.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_51 ( // @[package.scala 93:22:@21811.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_52 ( // @[package.scala 93:22:@21825.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  x472_x11 x472_x11_1 ( // @[Math.scala 150:24:@21834.4]
    .io_a(x472_x11_1_io_a),
    .io_b(x472_x11_1_io_b),
    .io_result(x472_x11_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_53 ( // @[package.scala 93:22:@21844.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  x472_x11 x473_x12_1 ( // @[Math.scala 150:24:@21853.4]
    .io_a(x473_x12_1_io_a),
    .io_b(x473_x12_1_io_b),
    .io_result(x473_x12_1_io_result)
  );
  x472_x11 x474_x11_1 ( // @[Math.scala 150:24:@21863.4]
    .io_a(x474_x11_1_io_a),
    .io_b(x474_x11_1_io_b),
    .io_result(x474_x11_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_54 ( // @[package.scala 93:22:@21873.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  x472_x11 x475_x12_1 ( // @[Math.scala 150:24:@21884.4]
    .io_a(x475_x12_1_io_a),
    .io_b(x475_x12_1_io_b),
    .io_result(x475_x12_1_io_result)
  );
  x472_x11 x476_x11_1 ( // @[Math.scala 150:24:@21894.4]
    .io_a(x476_x11_1_io_a),
    .io_b(x476_x11_1_io_b),
    .io_result(x476_x11_1_io_result)
  );
  x472_x11 x477_x12_1 ( // @[Math.scala 150:24:@21904.4]
    .io_a(x477_x12_1_io_a),
    .io_b(x477_x12_1_io_b),
    .io_result(x477_x12_1_io_result)
  );
  x478_x11 x478_x11_1 ( // @[Math.scala 150:24:@21914.4]
    .clock(x478_x11_1_clock),
    .reset(x478_x11_1_reset),
    .io_a(x478_x11_1_io_a),
    .io_b(x478_x11_1_io_b),
    .io_flow(x478_x11_1_io_flow),
    .io_result(x478_x11_1_io_result)
  );
  RetimeWrapper_266 RetimeWrapper_55 ( // @[package.scala 93:22:@21924.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  x472_x11 x479_sum_1 ( // @[Math.scala 150:24:@21933.4]
    .io_a(x479_sum_1_io_a),
    .io_b(x479_sum_1_io_b),
    .io_result(x479_sum_1_io_result)
  );
  RetimeWrapper_267 RetimeWrapper_56 ( // @[package.scala 93:22:@21954.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper_12 RetimeWrapper_57 ( // @[package.scala 93:22:@21963.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper_12 RetimeWrapper_58 ( // @[package.scala 93:22:@21972.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_12 RetimeWrapper_59 ( // @[package.scala 93:22:@21981.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  assign b281 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 62:18:@20597.4]
  assign b282 = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 63:18:@20598.4]
  assign _T_206 = b281 & b282; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 68:30:@20667.4]
  assign _T_207 = _T_206 & io_sigsIn_datapathEn; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 68:37:@20668.4]
  assign _T_211 = io_in_x270_TID == 8'h0; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 70:76:@20673.4]
  assign _T_212 = _T_207 & _T_211; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 70:62:@20674.4]
  assign _T_214 = io_in_x270_TDEST == 8'h0; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 70:101:@20675.4]
  assign b279_number = __io_result; // @[Math.scala 712:22:@20582.4 Math.scala 713:14:@20583.4]
  assign _T_240 = $signed(b279_number); // @[Math.scala 499:52:@20698.4]
  assign x288 = $signed(32'sh1) == $signed(_T_240); // @[Math.scala 499:44:@20706.4]
  assign x289 = $signed(32'sh2) == $signed(_T_240); // @[Math.scala 499:44:@20713.4]
  assign x290 = $signed(32'sh3) == $signed(_T_240); // @[Math.scala 499:44:@20720.4]
  assign _T_287 = x288 ? 32'h1 : 32'h0; // @[Mux.scala 19:72:@20732.4]
  assign _T_289 = x289 ? 32'h2 : 32'h0; // @[Mux.scala 19:72:@20733.4]
  assign _T_291 = x290 ? 32'h3 : 32'h0; // @[Mux.scala 19:72:@20734.4]
  assign _T_293 = _T_287 | _T_289; // @[Mux.scala 19:72:@20736.4]
  assign x291_number = _T_293 | _T_291; // @[Mux.scala 19:72:@20737.4]
  assign _T_305 = $signed(x291_number); // @[Math.scala 406:49:@20747.4]
  assign _T_307 = $signed(_T_305) & $signed(32'sh3); // @[Math.scala 406:56:@20749.4]
  assign _T_308 = $signed(_T_307); // @[Math.scala 406:56:@20750.4]
  assign b280_number = __1_io_result; // @[Math.scala 712:22:@20594.4 Math.scala 713:14:@20595.4]
  assign _T_317 = $signed(b280_number); // @[Math.scala 406:49:@20758.4]
  assign _T_319 = $signed(_T_317) & $signed(32'sh3); // @[Math.scala 406:56:@20760.4]
  assign _T_320 = $signed(_T_319); // @[Math.scala 406:56:@20761.4]
  assign _T_325 = x291_number[31]; // @[FixedPoint.scala 50:25:@20767.4]
  assign _T_329 = _T_325 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@20769.4]
  assign _T_330 = x291_number[31:2]; // @[FixedPoint.scala 18:52:@20770.4]
  assign _T_335 = b280_number[31]; // @[FixedPoint.scala 50:25:@20776.4]
  assign _T_339 = _T_335 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@20778.4]
  assign _T_340 = b280_number[31:2]; // @[FixedPoint.scala 18:52:@20779.4]
  assign _T_358 = ~ io_sigsIn_break; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 113:101:@20829.4]
  assign _T_362 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@20837.4 package.scala 96:25:@20838.4]
  assign _T_364 = io_rr ? _T_362 : 1'h0; // @[implicits.scala 55:10:@20839.4]
  assign _T_365 = _T_358 & _T_364; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 113:118:@20840.4]
  assign _T_367 = _T_365 & _T_358; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 113:205:@20842.4]
  assign _T_368 = _T_367 & io_sigsIn_backpressure; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 113:224:@20843.4]
  assign x588_b281_D1 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@20817.4 package.scala 96:25:@20818.4]
  assign _T_369 = _T_368 & x588_b281_D1; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 113:250:@20844.4]
  assign x586_b282_D1 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@20799.4 package.scala 96:25:@20800.4]
  assign x590_b279_D3_number = RetimeWrapper_6_io_out; // @[package.scala 96:25:@20858.4 package.scala 96:25:@20859.4]
  assign _T_379 = $signed(x590_b279_D3_number); // @[Math.scala 465:37:@20864.4]
  assign x304 = $signed(_T_379) < $signed(32'sh0); // @[Math.scala 465:44:@20866.4]
  assign x591_b280_D3_number = RetimeWrapper_7_io_out; // @[package.scala 96:25:@20874.4 package.scala 96:25:@20875.4]
  assign _T_390 = $signed(x591_b280_D3_number); // @[Math.scala 465:37:@20880.4]
  assign x305 = $signed(_T_390) < $signed(32'sh0); // @[Math.scala 465:44:@20882.4]
  assign x306 = x304 | x305; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 124:24:@20885.4]
  assign _T_406 = $signed(_T_379) & $signed(32'sh3); // @[Math.scala 406:56:@20896.4]
  assign _T_407 = $signed(_T_406); // @[Math.scala 406:56:@20897.4]
  assign x549_number = $unsigned(_T_407); // @[implicits.scala 133:21:@20898.4]
  assign _T_416 = $signed(x549_number); // @[Math.scala 406:49:@20905.4]
  assign _T_418 = $signed(_T_416) & $signed(32'sh3); // @[Math.scala 406:56:@20907.4]
  assign _T_419 = $signed(_T_418); // @[Math.scala 406:56:@20908.4]
  assign _T_424 = x549_number[31]; // @[FixedPoint.scala 50:25:@20914.4]
  assign _T_428 = _T_424 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@20916.4]
  assign _T_429 = x549_number[31:2]; // @[FixedPoint.scala 18:52:@20917.4]
  assign _T_460 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@20985.4 package.scala 96:25:@20986.4]
  assign _T_462 = io_rr ? _T_460 : 1'h0; // @[implicits.scala 55:10:@20987.4]
  assign _T_463 = _T_358 & _T_462; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 149:146:@20988.4]
  assign x595_x307_D2 = RetimeWrapper_11_io_out; // @[package.scala 96:25:@20964.4 package.scala 96:25:@20965.4]
  assign x597_x306_D4 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@21004.4 package.scala 96:25:@21005.4]
  assign x319_rd_0_number = x283_lb_0_io_rPort_7_output_0; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 145:29:@20976.4 sm_x485_inr_Foreach_SAMPLER_BOX.scala 149:274:@20995.4]
  assign x323_rdcol_number = x323_rdcol_1_io_result; // @[Math.scala 195:22:@21021.4 Math.scala 196:14:@21022.4]
  assign _T_487 = $signed(x323_rdcol_number); // @[Math.scala 465:37:@21027.4]
  assign x324 = $signed(_T_487) < $signed(32'sh0); // @[Math.scala 465:44:@21029.4]
  assign x598_x304_D1 = RetimeWrapper_15_io_out; // @[package.scala 96:25:@21037.4 package.scala 96:25:@21038.4]
  assign x325 = x598_x304_D1 | x324; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 163:24:@21041.4]
  assign _T_506 = $signed(_T_487) & $signed(32'sh3); // @[Math.scala 406:56:@21052.4]
  assign _T_507 = $signed(_T_506); // @[Math.scala 406:56:@21053.4]
  assign _T_512 = x323_rdcol_number[31]; // @[FixedPoint.scala 50:25:@21059.4]
  assign _T_516 = _T_512 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@21061.4]
  assign _T_517 = x323_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@21062.4]
  assign _T_544 = RetimeWrapper_19_io_out; // @[package.scala 96:25:@21114.4 package.scala 96:25:@21115.4]
  assign _T_546 = io_rr ? _T_544 : 1'h0; // @[implicits.scala 55:10:@21116.4]
  assign _T_547 = _T_358 & _T_546; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 190:194:@21117.4]
  assign x600_x326_D1 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@21093.4 package.scala 96:25:@21094.4]
  assign x602_x325_D3 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@21133.4 package.scala 96:25:@21134.4]
  assign x338_rd_0_number = x283_lb_0_io_rPort_5_output_0; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 186:29:@21105.4 sm_x485_inr_Foreach_SAMPLER_BOX.scala 190:322:@21124.4]
  assign x342_rdcol_number = x342_rdcol_1_io_result; // @[Math.scala 195:22:@21150.4 Math.scala 196:14:@21151.4]
  assign _T_571 = $signed(x342_rdcol_number); // @[Math.scala 465:37:@21156.4]
  assign x343 = $signed(_T_571) < $signed(32'sh0); // @[Math.scala 465:44:@21158.4]
  assign x344 = x598_x304_D1 | x343; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 202:59:@21161.4]
  assign _T_587 = $signed(_T_571) & $signed(32'sh3); // @[Math.scala 406:56:@21172.4]
  assign _T_588 = $signed(_T_587); // @[Math.scala 406:56:@21173.4]
  assign _T_593 = x342_rdcol_number[31]; // @[FixedPoint.scala 50:25:@21179.4]
  assign _T_597 = _T_593 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@21181.4]
  assign _T_598 = x342_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@21182.4]
  assign _T_620 = RetimeWrapper_23_io_out; // @[package.scala 96:25:@21223.4 package.scala 96:25:@21224.4]
  assign _T_622 = io_rr ? _T_620 : 1'h0; // @[implicits.scala 55:10:@21225.4]
  assign _T_623 = _T_358 & _T_622; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 219:194:@21226.4]
  assign x604_x345_D1 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@21211.4 package.scala 96:25:@21212.4]
  assign x605_x344_D3 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@21242.4 package.scala 96:25:@21243.4]
  assign x357_rd_0_number = x283_lb_0_io_rPort_0_output_0; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 215:29:@21214.4 sm_x485_inr_Foreach_SAMPLER_BOX.scala 219:322:@21233.4]
  assign x361_rdrow_number = x361_rdrow_1_io_result; // @[Math.scala 195:22:@21259.4 Math.scala 196:14:@21260.4]
  assign _T_647 = $signed(x361_rdrow_number); // @[Math.scala 465:37:@21265.4]
  assign x362 = $signed(_T_647) < $signed(32'sh0); // @[Math.scala 465:44:@21267.4]
  assign x606_x305_D1 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@21275.4 package.scala 96:25:@21276.4]
  assign x363 = x362 | x606_x305_D1; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 233:24:@21279.4]
  assign _T_666 = $signed(_T_647) & $signed(32'sh3); // @[Math.scala 406:56:@21290.4]
  assign _T_667 = $signed(_T_666); // @[Math.scala 406:56:@21291.4]
  assign x558_number = $unsigned(_T_667); // @[implicits.scala 133:21:@21292.4]
  assign _T_676 = $signed(x558_number); // @[Math.scala 406:49:@21299.4]
  assign _T_678 = $signed(_T_676) & $signed(32'sh3); // @[Math.scala 406:56:@21301.4]
  assign _T_679 = $signed(_T_678); // @[Math.scala 406:56:@21302.4]
  assign _T_684 = x558_number[31]; // @[FixedPoint.scala 50:25:@21308.4]
  assign _T_688 = _T_684 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@21310.4]
  assign _T_689 = x558_number[31:2]; // @[FixedPoint.scala 18:52:@21311.4]
  assign _T_714 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@21361.4 package.scala 96:25:@21362.4]
  assign _T_716 = io_rr ? _T_714 : 1'h0; // @[implicits.scala 55:10:@21363.4]
  assign _T_717 = _T_358 & _T_716; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 254:194:@21364.4]
  assign x608_x364_D1 = RetimeWrapper_27_io_out; // @[package.scala 96:25:@21340.4 package.scala 96:25:@21341.4]
  assign x610_x363_D3 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@21380.4 package.scala 96:25:@21381.4]
  assign x376_rd_0_number = x283_lb_0_io_rPort_1_output_0; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 250:29:@21352.4 sm_x485_inr_Foreach_SAMPLER_BOX.scala 254:322:@21371.4]
  assign x380 = x362 | x324; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 262:24:@21389.4]
  assign _T_750 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@21422.4 package.scala 96:25:@21423.4]
  assign _T_752 = io_rr ? _T_750 : 1'h0; // @[implicits.scala 55:10:@21424.4]
  assign _T_753 = _T_358 & _T_752; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 273:194:@21425.4]
  assign x611_x381_D1 = RetimeWrapper_31_io_out; // @[package.scala 96:25:@21410.4 package.scala 96:25:@21411.4]
  assign x612_x380_D3 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@21441.4 package.scala 96:25:@21442.4]
  assign x393_rd_0_number = x283_lb_0_io_rPort_3_output_0; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 269:29:@21413.4 sm_x485_inr_Foreach_SAMPLER_BOX.scala 273:322:@21432.4]
  assign x397 = x362 | x343; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 281:24:@21450.4]
  assign _T_786 = RetimeWrapper_35_io_out; // @[package.scala 96:25:@21483.4 package.scala 96:25:@21484.4]
  assign _T_788 = io_rr ? _T_786 : 1'h0; // @[implicits.scala 55:10:@21485.4]
  assign _T_789 = _T_358 & _T_788; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 292:194:@21486.4]
  assign x613_x398_D1 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@21471.4 package.scala 96:25:@21472.4]
  assign x614_x397_D3 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@21502.4 package.scala 96:25:@21503.4]
  assign x410_rd_0_number = x283_lb_0_io_rPort_8_output_0; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 288:29:@21474.4 sm_x485_inr_Foreach_SAMPLER_BOX.scala 292:322:@21493.4]
  assign x414_rdrow_number = x414_rdrow_1_io_result; // @[Math.scala 195:22:@21521.4 Math.scala 196:14:@21522.4]
  assign _T_815 = $signed(x414_rdrow_number); // @[Math.scala 465:37:@21527.4]
  assign x415 = $signed(_T_815) < $signed(32'sh0); // @[Math.scala 465:44:@21529.4]
  assign x416 = x415 | x606_x305_D1; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 312:24:@21532.4]
  assign _T_831 = $signed(_T_815) & $signed(32'sh3); // @[Math.scala 406:56:@21543.4]
  assign _T_832 = $signed(_T_831); // @[Math.scala 406:56:@21544.4]
  assign x567_number = $unsigned(_T_832); // @[implicits.scala 133:21:@21545.4]
  assign _T_841 = $signed(x567_number); // @[Math.scala 406:49:@21552.4]
  assign _T_843 = $signed(_T_841) & $signed(32'sh3); // @[Math.scala 406:56:@21554.4]
  assign _T_844 = $signed(_T_843); // @[Math.scala 406:56:@21555.4]
  assign _T_849 = x567_number[31]; // @[FixedPoint.scala 50:25:@21561.4]
  assign _T_853 = _T_849 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@21563.4]
  assign _T_854 = x567_number[31:2]; // @[FixedPoint.scala 18:52:@21564.4]
  assign _T_876 = RetimeWrapper_39_io_out; // @[package.scala 96:25:@21605.4 package.scala 96:25:@21606.4]
  assign _T_878 = io_rr ? _T_876 : 1'h0; // @[implicits.scala 55:10:@21607.4]
  assign _T_879 = _T_358 & _T_878; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 331:194:@21608.4]
  assign x616_x417_D1 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@21593.4 package.scala 96:25:@21594.4]
  assign x617_x416_D3 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@21624.4 package.scala 96:25:@21625.4]
  assign x429_rd_0_number = x283_lb_0_io_rPort_2_output_0; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 327:29:@21596.4 sm_x485_inr_Foreach_SAMPLER_BOX.scala 331:322:@21615.4]
  assign x433 = x415 | x324; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 339:24:@21633.4]
  assign _T_912 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@21666.4 package.scala 96:25:@21667.4]
  assign _T_914 = io_rr ? _T_912 : 1'h0; // @[implicits.scala 55:10:@21668.4]
  assign _T_915 = _T_358 & _T_914; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 350:194:@21669.4]
  assign x618_x434_D1 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@21654.4 package.scala 96:25:@21655.4]
  assign x619_x433_D3 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@21685.4 package.scala 96:25:@21686.4]
  assign x446_rd_0_number = x283_lb_0_io_rPort_6_output_0; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 346:29:@21657.4 sm_x485_inr_Foreach_SAMPLER_BOX.scala 350:322:@21676.4]
  assign x450 = x415 | x343; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 358:24:@21694.4]
  assign _T_948 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@21727.4 package.scala 96:25:@21728.4]
  assign _T_950 = io_rr ? _T_948 : 1'h0; // @[implicits.scala 55:10:@21729.4]
  assign _T_951 = _T_358 & _T_950; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 369:194:@21730.4]
  assign x620_x451_D1 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@21715.4 package.scala 96:25:@21716.4]
  assign x621_x450_D3 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@21746.4 package.scala 96:25:@21747.4]
  assign x463_rd_0_number = x283_lb_0_io_rPort_4_output_0; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 365:29:@21718.4 sm_x485_inr_Foreach_SAMPLER_BOX.scala 369:322:@21737.4]
  assign x622_x577_D1_number = RetimeWrapper_47_io_out; // @[package.scala 96:25:@21760.4 package.scala 96:25:@21761.4]
  assign _GEN_0 = {{1'd0}, x622_x577_D1_number}; // @[Math.scala 450:32:@21765.4]
  assign _T_969 = _GEN_0 << 1; // @[Math.scala 450:32:@21765.4]
  assign x623_x579_D1_number = RetimeWrapper_48_io_out; // @[package.scala 96:25:@21774.4 package.scala 96:25:@21775.4]
  assign _GEN_1 = {{1'd0}, x623_x579_D1_number}; // @[Math.scala 450:32:@21779.4]
  assign _T_976 = _GEN_1 << 1; // @[Math.scala 450:32:@21779.4]
  assign x624_x580_D1_number = RetimeWrapper_49_io_out; // @[package.scala 96:25:@21788.4 package.scala 96:25:@21789.4]
  assign _GEN_2 = {{2'd0}, x624_x580_D1_number}; // @[Math.scala 450:32:@21793.4]
  assign _T_983 = _GEN_2 << 2; // @[Math.scala 450:32:@21793.4]
  assign x625_x581_D1_number = RetimeWrapper_50_io_out; // @[package.scala 96:25:@21802.4 package.scala 96:25:@21803.4]
  assign _GEN_3 = {{1'd0}, x625_x581_D1_number}; // @[Math.scala 450:32:@21807.4]
  assign _T_990 = _GEN_3 << 1; // @[Math.scala 450:32:@21807.4]
  assign x626_x583_D1_number = RetimeWrapper_51_io_out; // @[package.scala 96:25:@21816.4 package.scala 96:25:@21817.4]
  assign _GEN_4 = {{1'd0}, x626_x583_D1_number}; // @[Math.scala 450:32:@21821.4]
  assign _T_997 = _GEN_4 << 1; // @[Math.scala 450:32:@21821.4]
  assign x479_sum_number = x479_sum_1_io_result; // @[Math.scala 154:22:@21939.4 Math.scala 155:14:@21940.4]
  assign _T_1044 = x479_sum_number[7:4]; // @[FixedPoint.scala 18:52:@21945.4]
  assign _T_1065 = RetimeWrapper_59_io_out; // @[package.scala 96:25:@21986.4 package.scala 96:25:@21987.4]
  assign _T_1067 = io_rr ? _T_1065 : 1'h0; // @[implicits.scala 55:10:@21988.4]
  assign x632_b281_D12 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@21977.4 package.scala 96:25:@21978.4]
  assign _T_1068 = _T_1067 & x632_b281_D12; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 439:116:@21989.4]
  assign x631_b282_D12 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@21968.4 package.scala 96:25:@21969.4]
  assign _T_1069 = _T_1068 & x631_b282_D12; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 439:122:@21990.4]
  assign x297_sum_number = x297_sum_1_io_result; // @[Math.scala 154:22:@20790.4 Math.scala 155:14:@20791.4]
  assign x587_x548_D1_number = RetimeWrapper_2_io_out; // @[package.scala 96:25:@20808.4 package.scala 96:25:@20809.4]
  assign x589_x547_D1_number = RetimeWrapper_4_io_out; // @[package.scala 96:25:@20826.4 package.scala 96:25:@20827.4]
  assign x593_x314_sum_D1_number = RetimeWrapper_9_io_out; // @[package.scala 96:25:@20946.4 package.scala 96:25:@20947.4]
  assign x594_x548_D5_number = RetimeWrapper_10_io_out; // @[package.scala 96:25:@20955.4 package.scala 96:25:@20956.4]
  assign x596_x550_D2_number = RetimeWrapper_12_io_out; // @[package.scala 96:25:@20973.4 package.scala 96:25:@20974.4]
  assign x333_sum_number = x333_sum_1_io_result; // @[Math.scala 154:22:@21084.4 Math.scala 155:14:@21085.4]
  assign x601_x554_D1_number = RetimeWrapper_18_io_out; // @[package.scala 96:25:@21102.4 package.scala 96:25:@21103.4]
  assign x352_sum_number = x352_sum_1_io_result; // @[Math.scala 154:22:@21193.4 Math.scala 155:14:@21194.4]
  assign x603_x557_D1_number = RetimeWrapper_21_io_out; // @[package.scala 96:25:@21202.4 package.scala 96:25:@21203.4]
  assign x371_sum_number = x371_sum_1_io_result; // @[Math.scala 154:22:@21331.4 Math.scala 155:14:@21332.4]
  assign x609_x559_D1_number = RetimeWrapper_28_io_out; // @[package.scala 96:25:@21349.4 package.scala 96:25:@21350.4]
  assign x388_sum_number = x388_sum_1_io_result; // @[Math.scala 154:22:@21401.4 Math.scala 155:14:@21402.4]
  assign x405_sum_number = x405_sum_1_io_result; // @[Math.scala 154:22:@21462.4 Math.scala 155:14:@21463.4]
  assign x424_sum_number = x424_sum_1_io_result; // @[Math.scala 154:22:@21575.4 Math.scala 155:14:@21576.4]
  assign x615_x568_D1_number = RetimeWrapper_37_io_out; // @[package.scala 96:25:@21584.4 package.scala 96:25:@21585.4]
  assign x441_sum_number = x441_sum_1_io_result; // @[Math.scala 154:22:@21645.4 Math.scala 155:14:@21646.4]
  assign x458_sum_number = x458_sum_1_io_result; // @[Math.scala 154:22:@21706.4 Math.scala 155:14:@21707.4]
  assign io_in_x270_TREADY = _T_212 & _T_214; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 68:22:@20669.4 sm_x485_inr_Foreach_SAMPLER_BOX.scala 70:22:@20677.4]
  assign io_in_x271_TVALID = _T_1069 & io_sigsIn_backpressure; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 439:22:@21992.4]
  assign io_in_x271_TDATA = {{248'd0}, RetimeWrapper_56_io_out}; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 440:24:@21993.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 710:17:@20580.4]
  assign __1_io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_1); // @[Math.scala 710:17:@20592.4]
  assign x283_lb_0_clock = clock; // @[:@20600.4]
  assign x283_lb_0_reset = reset; // @[:@20601.4]
  assign x283_lb_0_io_rPort_8_banks_1 = x603_x557_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@21489.4]
  assign x283_lb_0_io_rPort_8_banks_0 = x609_x559_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@21488.4]
  assign x283_lb_0_io_rPort_8_ofs_0 = x405_sum_number[0]; // @[MemInterfaceType.scala 107:54:@21490.4]
  assign x283_lb_0_io_rPort_8_en_0 = _T_789 & x613_x398_D1; // @[MemInterfaceType.scala 110:79:@21492.4]
  assign x283_lb_0_io_rPort_8_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@21491.4]
  assign x283_lb_0_io_rPort_7_banks_1 = x594_x548_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@20991.4]
  assign x283_lb_0_io_rPort_7_banks_0 = x596_x550_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@20990.4]
  assign x283_lb_0_io_rPort_7_ofs_0 = x593_x314_sum_D1_number[0]; // @[MemInterfaceType.scala 107:54:@20992.4]
  assign x283_lb_0_io_rPort_7_en_0 = _T_463 & x595_x307_D2; // @[MemInterfaceType.scala 110:79:@20994.4]
  assign x283_lb_0_io_rPort_7_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@20993.4]
  assign x283_lb_0_io_rPort_6_banks_1 = x601_x554_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@21672.4]
  assign x283_lb_0_io_rPort_6_banks_0 = x615_x568_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@21671.4]
  assign x283_lb_0_io_rPort_6_ofs_0 = x441_sum_number[0]; // @[MemInterfaceType.scala 107:54:@21673.4]
  assign x283_lb_0_io_rPort_6_en_0 = _T_915 & x618_x434_D1; // @[MemInterfaceType.scala 110:79:@21675.4]
  assign x283_lb_0_io_rPort_6_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@21674.4]
  assign x283_lb_0_io_rPort_5_banks_1 = x601_x554_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@21120.4]
  assign x283_lb_0_io_rPort_5_banks_0 = x596_x550_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@21119.4]
  assign x283_lb_0_io_rPort_5_ofs_0 = x333_sum_number[0]; // @[MemInterfaceType.scala 107:54:@21121.4]
  assign x283_lb_0_io_rPort_5_en_0 = _T_547 & x600_x326_D1; // @[MemInterfaceType.scala 110:79:@21123.4]
  assign x283_lb_0_io_rPort_5_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@21122.4]
  assign x283_lb_0_io_rPort_4_banks_1 = x603_x557_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@21733.4]
  assign x283_lb_0_io_rPort_4_banks_0 = x615_x568_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@21732.4]
  assign x283_lb_0_io_rPort_4_ofs_0 = x458_sum_number[0]; // @[MemInterfaceType.scala 107:54:@21734.4]
  assign x283_lb_0_io_rPort_4_en_0 = _T_951 & x620_x451_D1; // @[MemInterfaceType.scala 110:79:@21736.4]
  assign x283_lb_0_io_rPort_4_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@21735.4]
  assign x283_lb_0_io_rPort_3_banks_1 = x601_x554_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@21428.4]
  assign x283_lb_0_io_rPort_3_banks_0 = x609_x559_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@21427.4]
  assign x283_lb_0_io_rPort_3_ofs_0 = x388_sum_number[0]; // @[MemInterfaceType.scala 107:54:@21429.4]
  assign x283_lb_0_io_rPort_3_en_0 = _T_753 & x611_x381_D1; // @[MemInterfaceType.scala 110:79:@21431.4]
  assign x283_lb_0_io_rPort_3_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@21430.4]
  assign x283_lb_0_io_rPort_2_banks_1 = x594_x548_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@21611.4]
  assign x283_lb_0_io_rPort_2_banks_0 = x615_x568_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@21610.4]
  assign x283_lb_0_io_rPort_2_ofs_0 = x424_sum_number[0]; // @[MemInterfaceType.scala 107:54:@21612.4]
  assign x283_lb_0_io_rPort_2_en_0 = _T_879 & x616_x417_D1; // @[MemInterfaceType.scala 110:79:@21614.4]
  assign x283_lb_0_io_rPort_2_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@21613.4]
  assign x283_lb_0_io_rPort_1_banks_1 = x594_x548_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@21367.4]
  assign x283_lb_0_io_rPort_1_banks_0 = x609_x559_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@21366.4]
  assign x283_lb_0_io_rPort_1_ofs_0 = x371_sum_number[0]; // @[MemInterfaceType.scala 107:54:@21368.4]
  assign x283_lb_0_io_rPort_1_en_0 = _T_717 & x608_x364_D1; // @[MemInterfaceType.scala 110:79:@21370.4]
  assign x283_lb_0_io_rPort_1_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@21369.4]
  assign x283_lb_0_io_rPort_0_banks_1 = x603_x557_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@21229.4]
  assign x283_lb_0_io_rPort_0_banks_0 = x596_x550_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@21228.4]
  assign x283_lb_0_io_rPort_0_ofs_0 = x352_sum_number[0]; // @[MemInterfaceType.scala 107:54:@21230.4]
  assign x283_lb_0_io_rPort_0_en_0 = _T_623 & x604_x345_D1; // @[MemInterfaceType.scala 110:79:@21232.4]
  assign x283_lb_0_io_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@21231.4]
  assign x283_lb_0_io_wPort_0_banks_1 = x587_x548_D1_number[2:0]; // @[MemInterfaceType.scala 88:58:@20847.4]
  assign x283_lb_0_io_wPort_0_banks_0 = x589_x547_D1_number[2:0]; // @[MemInterfaceType.scala 88:58:@20846.4]
  assign x283_lb_0_io_wPort_0_ofs_0 = x297_sum_number[0]; // @[MemInterfaceType.scala 89:54:@20848.4]
  assign x283_lb_0_io_wPort_0_data_0 = RetimeWrapper_io_out; // @[MemInterfaceType.scala 90:56:@20849.4]
  assign x283_lb_0_io_wPort_0_en_0 = _T_369 & x586_b282_D1; // @[MemInterfaceType.scala 93:57:@20851.4]
  assign RetimeWrapper_clock = clock; // @[:@20680.4]
  assign RetimeWrapper_reset = reset; // @[:@20681.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@20683.4]
  assign RetimeWrapper_io_in = io_in_x270_TDATA[7:0]; // @[package.scala 94:16:@20682.4]
  assign x297_sum_1_clock = clock; // @[:@20785.4]
  assign x297_sum_1_reset = reset; // @[:@20786.4]
  assign x297_sum_1_io_a = {_T_329,_T_330}; // @[Math.scala 151:17:@20787.4]
  assign x297_sum_1_io_b = {_T_339,_T_340}; // @[Math.scala 152:17:@20788.4]
  assign x297_sum_1_io_flow = io_in_x271_TREADY; // @[Math.scala 153:20:@20789.4]
  assign RetimeWrapper_1_clock = clock; // @[:@20795.4]
  assign RetimeWrapper_1_reset = reset; // @[:@20796.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@20798.4]
  assign RetimeWrapper_1_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@20797.4]
  assign RetimeWrapper_2_clock = clock; // @[:@20804.4]
  assign RetimeWrapper_2_reset = reset; // @[:@20805.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@20807.4]
  assign RetimeWrapper_2_io_in = $unsigned(_T_320); // @[package.scala 94:16:@20806.4]
  assign RetimeWrapper_3_clock = clock; // @[:@20813.4]
  assign RetimeWrapper_3_reset = reset; // @[:@20814.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@20816.4]
  assign RetimeWrapper_3_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@20815.4]
  assign RetimeWrapper_4_clock = clock; // @[:@20822.4]
  assign RetimeWrapper_4_reset = reset; // @[:@20823.4]
  assign RetimeWrapper_4_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@20825.4]
  assign RetimeWrapper_4_io_in = $unsigned(_T_308); // @[package.scala 94:16:@20824.4]
  assign RetimeWrapper_5_clock = clock; // @[:@20833.4]
  assign RetimeWrapper_5_reset = reset; // @[:@20834.4]
  assign RetimeWrapper_5_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@20836.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@20835.4]
  assign RetimeWrapper_6_clock = clock; // @[:@20854.4]
  assign RetimeWrapper_6_reset = reset; // @[:@20855.4]
  assign RetimeWrapper_6_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@20857.4]
  assign RetimeWrapper_6_io_in = __io_result; // @[package.scala 94:16:@20856.4]
  assign RetimeWrapper_7_clock = clock; // @[:@20870.4]
  assign RetimeWrapper_7_reset = reset; // @[:@20871.4]
  assign RetimeWrapper_7_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@20873.4]
  assign RetimeWrapper_7_io_in = __1_io_result; // @[package.scala 94:16:@20872.4]
  assign RetimeWrapper_8_clock = clock; // @[:@20923.4]
  assign RetimeWrapper_8_reset = reset; // @[:@20924.4]
  assign RetimeWrapper_8_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@20926.4]
  assign RetimeWrapper_8_io_in = {_T_339,_T_340}; // @[package.scala 94:16:@20925.4]
  assign x314_sum_1_clock = clock; // @[:@20932.4]
  assign x314_sum_1_reset = reset; // @[:@20933.4]
  assign x314_sum_1_io_a = {_T_428,_T_429}; // @[Math.scala 151:17:@20934.4]
  assign x314_sum_1_io_b = RetimeWrapper_8_io_out; // @[Math.scala 152:17:@20935.4]
  assign x314_sum_1_io_flow = io_in_x271_TREADY; // @[Math.scala 153:20:@20936.4]
  assign RetimeWrapper_9_clock = clock; // @[:@20942.4]
  assign RetimeWrapper_9_reset = reset; // @[:@20943.4]
  assign RetimeWrapper_9_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@20945.4]
  assign RetimeWrapper_9_io_in = x314_sum_1_io_result; // @[package.scala 94:16:@20944.4]
  assign RetimeWrapper_10_clock = clock; // @[:@20951.4]
  assign RetimeWrapper_10_reset = reset; // @[:@20952.4]
  assign RetimeWrapper_10_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@20954.4]
  assign RetimeWrapper_10_io_in = $unsigned(_T_320); // @[package.scala 94:16:@20953.4]
  assign RetimeWrapper_11_clock = clock; // @[:@20960.4]
  assign RetimeWrapper_11_reset = reset; // @[:@20961.4]
  assign RetimeWrapper_11_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@20963.4]
  assign RetimeWrapper_11_io_in = ~ x306; // @[package.scala 94:16:@20962.4]
  assign RetimeWrapper_12_clock = clock; // @[:@20969.4]
  assign RetimeWrapper_12_reset = reset; // @[:@20970.4]
  assign RetimeWrapper_12_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@20972.4]
  assign RetimeWrapper_12_io_in = $unsigned(_T_419); // @[package.scala 94:16:@20971.4]
  assign RetimeWrapper_13_clock = clock; // @[:@20981.4]
  assign RetimeWrapper_13_reset = reset; // @[:@20982.4]
  assign RetimeWrapper_13_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@20984.4]
  assign RetimeWrapper_13_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@20983.4]
  assign RetimeWrapper_14_clock = clock; // @[:@21000.4]
  assign RetimeWrapper_14_reset = reset; // @[:@21001.4]
  assign RetimeWrapper_14_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21003.4]
  assign RetimeWrapper_14_io_in = x304 | x305; // @[package.scala 94:16:@21002.4]
  assign x323_rdcol_1_clock = clock; // @[:@21016.4]
  assign x323_rdcol_1_reset = reset; // @[:@21017.4]
  assign x323_rdcol_1_io_a = RetimeWrapper_7_io_out; // @[Math.scala 192:17:@21018.4]
  assign x323_rdcol_1_io_b = 32'h1; // @[Math.scala 193:17:@21019.4]
  assign x323_rdcol_1_io_flow = io_in_x271_TREADY; // @[Math.scala 194:20:@21020.4]
  assign RetimeWrapper_15_clock = clock; // @[:@21033.4]
  assign RetimeWrapper_15_reset = reset; // @[:@21034.4]
  assign RetimeWrapper_15_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21036.4]
  assign RetimeWrapper_15_io_in = $signed(_T_379) < $signed(32'sh0); // @[package.scala 94:16:@21035.4]
  assign RetimeWrapper_16_clock = clock; // @[:@21068.4]
  assign RetimeWrapper_16_reset = reset; // @[:@21069.4]
  assign RetimeWrapper_16_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21071.4]
  assign RetimeWrapper_16_io_in = {_T_428,_T_429}; // @[package.scala 94:16:@21070.4]
  assign x333_sum_1_clock = clock; // @[:@21079.4]
  assign x333_sum_1_reset = reset; // @[:@21080.4]
  assign x333_sum_1_io_a = RetimeWrapper_16_io_out; // @[Math.scala 151:17:@21081.4]
  assign x333_sum_1_io_b = {_T_516,_T_517}; // @[Math.scala 152:17:@21082.4]
  assign x333_sum_1_io_flow = io_in_x271_TREADY; // @[Math.scala 153:20:@21083.4]
  assign RetimeWrapper_17_clock = clock; // @[:@21089.4]
  assign RetimeWrapper_17_reset = reset; // @[:@21090.4]
  assign RetimeWrapper_17_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21092.4]
  assign RetimeWrapper_17_io_in = ~ x325; // @[package.scala 94:16:@21091.4]
  assign RetimeWrapper_18_clock = clock; // @[:@21098.4]
  assign RetimeWrapper_18_reset = reset; // @[:@21099.4]
  assign RetimeWrapper_18_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21101.4]
  assign RetimeWrapper_18_io_in = $unsigned(_T_507); // @[package.scala 94:16:@21100.4]
  assign RetimeWrapper_19_clock = clock; // @[:@21110.4]
  assign RetimeWrapper_19_reset = reset; // @[:@21111.4]
  assign RetimeWrapper_19_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21113.4]
  assign RetimeWrapper_19_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@21112.4]
  assign RetimeWrapper_20_clock = clock; // @[:@21129.4]
  assign RetimeWrapper_20_reset = reset; // @[:@21130.4]
  assign RetimeWrapper_20_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21132.4]
  assign RetimeWrapper_20_io_in = x598_x304_D1 | x324; // @[package.scala 94:16:@21131.4]
  assign x342_rdcol_1_clock = clock; // @[:@21145.4]
  assign x342_rdcol_1_reset = reset; // @[:@21146.4]
  assign x342_rdcol_1_io_a = RetimeWrapper_7_io_out; // @[Math.scala 192:17:@21147.4]
  assign x342_rdcol_1_io_b = 32'h2; // @[Math.scala 193:17:@21148.4]
  assign x342_rdcol_1_io_flow = io_in_x271_TREADY; // @[Math.scala 194:20:@21149.4]
  assign x352_sum_1_clock = clock; // @[:@21188.4]
  assign x352_sum_1_reset = reset; // @[:@21189.4]
  assign x352_sum_1_io_a = RetimeWrapper_16_io_out; // @[Math.scala 151:17:@21190.4]
  assign x352_sum_1_io_b = {_T_597,_T_598}; // @[Math.scala 152:17:@21191.4]
  assign x352_sum_1_io_flow = io_in_x271_TREADY; // @[Math.scala 153:20:@21192.4]
  assign RetimeWrapper_21_clock = clock; // @[:@21198.4]
  assign RetimeWrapper_21_reset = reset; // @[:@21199.4]
  assign RetimeWrapper_21_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21201.4]
  assign RetimeWrapper_21_io_in = $unsigned(_T_588); // @[package.scala 94:16:@21200.4]
  assign RetimeWrapper_22_clock = clock; // @[:@21207.4]
  assign RetimeWrapper_22_reset = reset; // @[:@21208.4]
  assign RetimeWrapper_22_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21210.4]
  assign RetimeWrapper_22_io_in = ~ x344; // @[package.scala 94:16:@21209.4]
  assign RetimeWrapper_23_clock = clock; // @[:@21219.4]
  assign RetimeWrapper_23_reset = reset; // @[:@21220.4]
  assign RetimeWrapper_23_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21222.4]
  assign RetimeWrapper_23_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@21221.4]
  assign RetimeWrapper_24_clock = clock; // @[:@21238.4]
  assign RetimeWrapper_24_reset = reset; // @[:@21239.4]
  assign RetimeWrapper_24_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21241.4]
  assign RetimeWrapper_24_io_in = x598_x304_D1 | x343; // @[package.scala 94:16:@21240.4]
  assign x361_rdrow_1_clock = clock; // @[:@21254.4]
  assign x361_rdrow_1_reset = reset; // @[:@21255.4]
  assign x361_rdrow_1_io_a = RetimeWrapper_6_io_out; // @[Math.scala 192:17:@21256.4]
  assign x361_rdrow_1_io_b = 32'h1; // @[Math.scala 193:17:@21257.4]
  assign x361_rdrow_1_io_flow = io_in_x271_TREADY; // @[Math.scala 194:20:@21258.4]
  assign RetimeWrapper_25_clock = clock; // @[:@21271.4]
  assign RetimeWrapper_25_reset = reset; // @[:@21272.4]
  assign RetimeWrapper_25_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21274.4]
  assign RetimeWrapper_25_io_in = $signed(_T_390) < $signed(32'sh0); // @[package.scala 94:16:@21273.4]
  assign RetimeWrapper_26_clock = clock; // @[:@21317.4]
  assign RetimeWrapper_26_reset = reset; // @[:@21318.4]
  assign RetimeWrapper_26_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21320.4]
  assign RetimeWrapper_26_io_in = {_T_339,_T_340}; // @[package.scala 94:16:@21319.4]
  assign x371_sum_1_clock = clock; // @[:@21326.4]
  assign x371_sum_1_reset = reset; // @[:@21327.4]
  assign x371_sum_1_io_a = {_T_688,_T_689}; // @[Math.scala 151:17:@21328.4]
  assign x371_sum_1_io_b = RetimeWrapper_26_io_out; // @[Math.scala 152:17:@21329.4]
  assign x371_sum_1_io_flow = io_in_x271_TREADY; // @[Math.scala 153:20:@21330.4]
  assign RetimeWrapper_27_clock = clock; // @[:@21336.4]
  assign RetimeWrapper_27_reset = reset; // @[:@21337.4]
  assign RetimeWrapper_27_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21339.4]
  assign RetimeWrapper_27_io_in = ~ x363; // @[package.scala 94:16:@21338.4]
  assign RetimeWrapper_28_clock = clock; // @[:@21345.4]
  assign RetimeWrapper_28_reset = reset; // @[:@21346.4]
  assign RetimeWrapper_28_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21348.4]
  assign RetimeWrapper_28_io_in = $unsigned(_T_679); // @[package.scala 94:16:@21347.4]
  assign RetimeWrapper_29_clock = clock; // @[:@21357.4]
  assign RetimeWrapper_29_reset = reset; // @[:@21358.4]
  assign RetimeWrapper_29_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21360.4]
  assign RetimeWrapper_29_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@21359.4]
  assign RetimeWrapper_30_clock = clock; // @[:@21376.4]
  assign RetimeWrapper_30_reset = reset; // @[:@21377.4]
  assign RetimeWrapper_30_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21379.4]
  assign RetimeWrapper_30_io_in = x362 | x606_x305_D1; // @[package.scala 94:16:@21378.4]
  assign x388_sum_1_clock = clock; // @[:@21396.4]
  assign x388_sum_1_reset = reset; // @[:@21397.4]
  assign x388_sum_1_io_a = {_T_688,_T_689}; // @[Math.scala 151:17:@21398.4]
  assign x388_sum_1_io_b = {_T_516,_T_517}; // @[Math.scala 152:17:@21399.4]
  assign x388_sum_1_io_flow = io_in_x271_TREADY; // @[Math.scala 153:20:@21400.4]
  assign RetimeWrapper_31_clock = clock; // @[:@21406.4]
  assign RetimeWrapper_31_reset = reset; // @[:@21407.4]
  assign RetimeWrapper_31_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21409.4]
  assign RetimeWrapper_31_io_in = ~ x380; // @[package.scala 94:16:@21408.4]
  assign RetimeWrapper_32_clock = clock; // @[:@21418.4]
  assign RetimeWrapper_32_reset = reset; // @[:@21419.4]
  assign RetimeWrapper_32_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21421.4]
  assign RetimeWrapper_32_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@21420.4]
  assign RetimeWrapper_33_clock = clock; // @[:@21437.4]
  assign RetimeWrapper_33_reset = reset; // @[:@21438.4]
  assign RetimeWrapper_33_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21440.4]
  assign RetimeWrapper_33_io_in = x362 | x324; // @[package.scala 94:16:@21439.4]
  assign x405_sum_1_clock = clock; // @[:@21457.4]
  assign x405_sum_1_reset = reset; // @[:@21458.4]
  assign x405_sum_1_io_a = {_T_688,_T_689}; // @[Math.scala 151:17:@21459.4]
  assign x405_sum_1_io_b = {_T_597,_T_598}; // @[Math.scala 152:17:@21460.4]
  assign x405_sum_1_io_flow = io_in_x271_TREADY; // @[Math.scala 153:20:@21461.4]
  assign RetimeWrapper_34_clock = clock; // @[:@21467.4]
  assign RetimeWrapper_34_reset = reset; // @[:@21468.4]
  assign RetimeWrapper_34_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21470.4]
  assign RetimeWrapper_34_io_in = ~ x397; // @[package.scala 94:16:@21469.4]
  assign RetimeWrapper_35_clock = clock; // @[:@21479.4]
  assign RetimeWrapper_35_reset = reset; // @[:@21480.4]
  assign RetimeWrapper_35_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21482.4]
  assign RetimeWrapper_35_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@21481.4]
  assign RetimeWrapper_36_clock = clock; // @[:@21498.4]
  assign RetimeWrapper_36_reset = reset; // @[:@21499.4]
  assign RetimeWrapper_36_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21501.4]
  assign RetimeWrapper_36_io_in = x362 | x343; // @[package.scala 94:16:@21500.4]
  assign x414_rdrow_1_clock = clock; // @[:@21516.4]
  assign x414_rdrow_1_reset = reset; // @[:@21517.4]
  assign x414_rdrow_1_io_a = RetimeWrapper_6_io_out; // @[Math.scala 192:17:@21518.4]
  assign x414_rdrow_1_io_b = 32'h2; // @[Math.scala 193:17:@21519.4]
  assign x414_rdrow_1_io_flow = io_in_x271_TREADY; // @[Math.scala 194:20:@21520.4]
  assign x424_sum_1_clock = clock; // @[:@21570.4]
  assign x424_sum_1_reset = reset; // @[:@21571.4]
  assign x424_sum_1_io_a = {_T_853,_T_854}; // @[Math.scala 151:17:@21572.4]
  assign x424_sum_1_io_b = RetimeWrapper_26_io_out; // @[Math.scala 152:17:@21573.4]
  assign x424_sum_1_io_flow = io_in_x271_TREADY; // @[Math.scala 153:20:@21574.4]
  assign RetimeWrapper_37_clock = clock; // @[:@21580.4]
  assign RetimeWrapper_37_reset = reset; // @[:@21581.4]
  assign RetimeWrapper_37_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21583.4]
  assign RetimeWrapper_37_io_in = $unsigned(_T_844); // @[package.scala 94:16:@21582.4]
  assign RetimeWrapper_38_clock = clock; // @[:@21589.4]
  assign RetimeWrapper_38_reset = reset; // @[:@21590.4]
  assign RetimeWrapper_38_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21592.4]
  assign RetimeWrapper_38_io_in = ~ x416; // @[package.scala 94:16:@21591.4]
  assign RetimeWrapper_39_clock = clock; // @[:@21601.4]
  assign RetimeWrapper_39_reset = reset; // @[:@21602.4]
  assign RetimeWrapper_39_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21604.4]
  assign RetimeWrapper_39_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@21603.4]
  assign RetimeWrapper_40_clock = clock; // @[:@21620.4]
  assign RetimeWrapper_40_reset = reset; // @[:@21621.4]
  assign RetimeWrapper_40_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21623.4]
  assign RetimeWrapper_40_io_in = x415 | x606_x305_D1; // @[package.scala 94:16:@21622.4]
  assign x441_sum_1_clock = clock; // @[:@21640.4]
  assign x441_sum_1_reset = reset; // @[:@21641.4]
  assign x441_sum_1_io_a = {_T_853,_T_854}; // @[Math.scala 151:17:@21642.4]
  assign x441_sum_1_io_b = {_T_516,_T_517}; // @[Math.scala 152:17:@21643.4]
  assign x441_sum_1_io_flow = io_in_x271_TREADY; // @[Math.scala 153:20:@21644.4]
  assign RetimeWrapper_41_clock = clock; // @[:@21650.4]
  assign RetimeWrapper_41_reset = reset; // @[:@21651.4]
  assign RetimeWrapper_41_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21653.4]
  assign RetimeWrapper_41_io_in = ~ x433; // @[package.scala 94:16:@21652.4]
  assign RetimeWrapper_42_clock = clock; // @[:@21662.4]
  assign RetimeWrapper_42_reset = reset; // @[:@21663.4]
  assign RetimeWrapper_42_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21665.4]
  assign RetimeWrapper_42_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@21664.4]
  assign RetimeWrapper_43_clock = clock; // @[:@21681.4]
  assign RetimeWrapper_43_reset = reset; // @[:@21682.4]
  assign RetimeWrapper_43_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21684.4]
  assign RetimeWrapper_43_io_in = x415 | x324; // @[package.scala 94:16:@21683.4]
  assign x458_sum_1_clock = clock; // @[:@21701.4]
  assign x458_sum_1_reset = reset; // @[:@21702.4]
  assign x458_sum_1_io_a = {_T_853,_T_854}; // @[Math.scala 151:17:@21703.4]
  assign x458_sum_1_io_b = {_T_597,_T_598}; // @[Math.scala 152:17:@21704.4]
  assign x458_sum_1_io_flow = io_in_x271_TREADY; // @[Math.scala 153:20:@21705.4]
  assign RetimeWrapper_44_clock = clock; // @[:@21711.4]
  assign RetimeWrapper_44_reset = reset; // @[:@21712.4]
  assign RetimeWrapper_44_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21714.4]
  assign RetimeWrapper_44_io_in = ~ x450; // @[package.scala 94:16:@21713.4]
  assign RetimeWrapper_45_clock = clock; // @[:@21723.4]
  assign RetimeWrapper_45_reset = reset; // @[:@21724.4]
  assign RetimeWrapper_45_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21726.4]
  assign RetimeWrapper_45_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@21725.4]
  assign RetimeWrapper_46_clock = clock; // @[:@21742.4]
  assign RetimeWrapper_46_reset = reset; // @[:@21743.4]
  assign RetimeWrapper_46_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21745.4]
  assign RetimeWrapper_46_io_in = x415 | x343; // @[package.scala 94:16:@21744.4]
  assign RetimeWrapper_47_clock = clock; // @[:@21756.4]
  assign RetimeWrapper_47_reset = reset; // @[:@21757.4]
  assign RetimeWrapper_47_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21759.4]
  assign RetimeWrapper_47_io_in = x602_x325_D3 ? 8'h0 : x338_rd_0_number; // @[package.scala 94:16:@21758.4]
  assign RetimeWrapper_48_clock = clock; // @[:@21770.4]
  assign RetimeWrapper_48_reset = reset; // @[:@21771.4]
  assign RetimeWrapper_48_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21773.4]
  assign RetimeWrapper_48_io_in = x610_x363_D3 ? 8'h0 : x376_rd_0_number; // @[package.scala 94:16:@21772.4]
  assign RetimeWrapper_49_clock = clock; // @[:@21784.4]
  assign RetimeWrapper_49_reset = reset; // @[:@21785.4]
  assign RetimeWrapper_49_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21787.4]
  assign RetimeWrapper_49_io_in = x612_x380_D3 ? 8'h0 : x393_rd_0_number; // @[package.scala 94:16:@21786.4]
  assign RetimeWrapper_50_clock = clock; // @[:@21798.4]
  assign RetimeWrapper_50_reset = reset; // @[:@21799.4]
  assign RetimeWrapper_50_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21801.4]
  assign RetimeWrapper_50_io_in = x614_x397_D3 ? 8'h0 : x410_rd_0_number; // @[package.scala 94:16:@21800.4]
  assign RetimeWrapper_51_clock = clock; // @[:@21812.4]
  assign RetimeWrapper_51_reset = reset; // @[:@21813.4]
  assign RetimeWrapper_51_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21815.4]
  assign RetimeWrapper_51_io_in = x619_x433_D3 ? 8'h0 : x446_rd_0_number; // @[package.scala 94:16:@21814.4]
  assign RetimeWrapper_52_clock = clock; // @[:@21826.4]
  assign RetimeWrapper_52_reset = reset; // @[:@21827.4]
  assign RetimeWrapper_52_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21829.4]
  assign RetimeWrapper_52_io_in = x597_x306_D4 ? 8'h0 : x319_rd_0_number; // @[package.scala 94:16:@21828.4]
  assign x472_x11_1_io_a = RetimeWrapper_52_io_out; // @[Math.scala 151:17:@21837.4]
  assign x472_x11_1_io_b = _T_969[7:0]; // @[Math.scala 152:17:@21838.4]
  assign RetimeWrapper_53_clock = clock; // @[:@21845.4]
  assign RetimeWrapper_53_reset = reset; // @[:@21846.4]
  assign RetimeWrapper_53_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21848.4]
  assign RetimeWrapper_53_io_in = x605_x344_D3 ? 8'h0 : x357_rd_0_number; // @[package.scala 94:16:@21847.4]
  assign x473_x12_1_io_a = RetimeWrapper_53_io_out; // @[Math.scala 151:17:@21856.4]
  assign x473_x12_1_io_b = _T_976[7:0]; // @[Math.scala 152:17:@21857.4]
  assign x474_x11_1_io_a = _T_983[7:0]; // @[Math.scala 151:17:@21866.4]
  assign x474_x11_1_io_b = _T_990[7:0]; // @[Math.scala 152:17:@21867.4]
  assign RetimeWrapper_54_clock = clock; // @[:@21874.4]
  assign RetimeWrapper_54_reset = reset; // @[:@21875.4]
  assign RetimeWrapper_54_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21877.4]
  assign RetimeWrapper_54_io_in = x617_x416_D3 ? 8'h0 : x429_rd_0_number; // @[package.scala 94:16:@21876.4]
  assign x475_x12_1_io_a = RetimeWrapper_54_io_out; // @[Math.scala 151:17:@21887.4]
  assign x475_x12_1_io_b = _T_997[7:0]; // @[Math.scala 152:17:@21888.4]
  assign x476_x11_1_io_a = x472_x11_1_io_result; // @[Math.scala 151:17:@21897.4]
  assign x476_x11_1_io_b = x473_x12_1_io_result; // @[Math.scala 152:17:@21898.4]
  assign x477_x12_1_io_a = x474_x11_1_io_result; // @[Math.scala 151:17:@21907.4]
  assign x477_x12_1_io_b = x475_x12_1_io_result; // @[Math.scala 152:17:@21908.4]
  assign x478_x11_1_clock = clock; // @[:@21915.4]
  assign x478_x11_1_reset = reset; // @[:@21916.4]
  assign x478_x11_1_io_a = x476_x11_1_io_result; // @[Math.scala 151:17:@21917.4]
  assign x478_x11_1_io_b = x477_x12_1_io_result; // @[Math.scala 152:17:@21918.4]
  assign x478_x11_1_io_flow = io_in_x271_TREADY; // @[Math.scala 153:20:@21919.4]
  assign RetimeWrapper_55_clock = clock; // @[:@21925.4]
  assign RetimeWrapper_55_reset = reset; // @[:@21926.4]
  assign RetimeWrapper_55_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21928.4]
  assign RetimeWrapper_55_io_in = x621_x450_D3 ? 8'h0 : x463_rd_0_number; // @[package.scala 94:16:@21927.4]
  assign x479_sum_1_io_a = x478_x11_1_io_result; // @[Math.scala 151:17:@21936.4]
  assign x479_sum_1_io_b = RetimeWrapper_55_io_out; // @[Math.scala 152:17:@21937.4]
  assign RetimeWrapper_56_clock = clock; // @[:@21955.4]
  assign RetimeWrapper_56_reset = reset; // @[:@21956.4]
  assign RetimeWrapper_56_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21958.4]
  assign RetimeWrapper_56_io_in = {4'h0,_T_1044}; // @[package.scala 94:16:@21957.4]
  assign RetimeWrapper_57_clock = clock; // @[:@21964.4]
  assign RetimeWrapper_57_reset = reset; // @[:@21965.4]
  assign RetimeWrapper_57_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21967.4]
  assign RetimeWrapper_57_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@21966.4]
  assign RetimeWrapper_58_clock = clock; // @[:@21973.4]
  assign RetimeWrapper_58_reset = reset; // @[:@21974.4]
  assign RetimeWrapper_58_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21976.4]
  assign RetimeWrapper_58_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@21975.4]
  assign RetimeWrapper_59_clock = clock; // @[:@21982.4]
  assign RetimeWrapper_59_reset = reset; // @[:@21983.4]
  assign RetimeWrapper_59_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21985.4]
  assign RetimeWrapper_59_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@21984.4]
endmodule
module x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1( // @[:@22003.2]
  input          clock, // @[:@22004.4]
  input          reset, // @[:@22005.4]
  input          io_in_x270_TVALID, // @[:@22006.4]
  output         io_in_x270_TREADY, // @[:@22006.4]
  input  [255:0] io_in_x270_TDATA, // @[:@22006.4]
  input  [7:0]   io_in_x270_TID, // @[:@22006.4]
  input  [7:0]   io_in_x270_TDEST, // @[:@22006.4]
  output         io_in_x271_TVALID, // @[:@22006.4]
  input          io_in_x271_TREADY, // @[:@22006.4]
  output [255:0] io_in_x271_TDATA, // @[:@22006.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@22006.4]
  input          io_sigsIn_smChildAcks_0, // @[:@22006.4]
  output         io_sigsOut_smDoneIn_0, // @[:@22006.4]
  output         io_sigsOut_smCtrCopyDone_0, // @[:@22006.4]
  input          io_rr // @[:@22006.4]
);
  wire  x278_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@22016.4]
  wire  x278_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@22016.4]
  wire  x278_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@22016.4]
  wire  x278_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@22016.4]
  wire [31:0] x278_ctrchain_io_output_counts_1; // @[SpatialBlocks.scala 37:22:@22016.4]
  wire [31:0] x278_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@22016.4]
  wire  x278_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@22016.4]
  wire  x278_ctrchain_io_output_oobs_1; // @[SpatialBlocks.scala 37:22:@22016.4]
  wire  x278_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@22016.4]
  wire  x485_inr_Foreach_SAMPLER_BOX_sm_clock; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 32:18:@22075.4]
  wire  x485_inr_Foreach_SAMPLER_BOX_sm_reset; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 32:18:@22075.4]
  wire  x485_inr_Foreach_SAMPLER_BOX_sm_io_enable; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 32:18:@22075.4]
  wire  x485_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 32:18:@22075.4]
  wire  x485_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 32:18:@22075.4]
  wire  x485_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 32:18:@22075.4]
  wire  x485_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 32:18:@22075.4]
  wire  x485_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 32:18:@22075.4]
  wire  x485_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 32:18:@22075.4]
  wire  x485_inr_Foreach_SAMPLER_BOX_sm_io_parentAck; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 32:18:@22075.4]
  wire  x485_inr_Foreach_SAMPLER_BOX_sm_io_backpressure; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 32:18:@22075.4]
  wire  x485_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 32:18:@22075.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@22103.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@22103.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@22103.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@22103.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@22103.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@22145.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@22145.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@22145.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@22145.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@22145.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@22153.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@22153.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@22153.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@22153.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@22153.4]
  wire  x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_clock; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 452:24:@22185.4]
  wire  x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_reset; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 452:24:@22185.4]
  wire  x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x270_TREADY; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 452:24:@22185.4]
  wire [255:0] x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x270_TDATA; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 452:24:@22185.4]
  wire [7:0] x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x270_TID; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 452:24:@22185.4]
  wire [7:0] x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x270_TDEST; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 452:24:@22185.4]
  wire  x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x271_TVALID; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 452:24:@22185.4]
  wire  x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x271_TREADY; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 452:24:@22185.4]
  wire [255:0] x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x271_TDATA; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 452:24:@22185.4]
  wire  x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 452:24:@22185.4]
  wire  x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 452:24:@22185.4]
  wire  x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 452:24:@22185.4]
  wire [31:0] x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 452:24:@22185.4]
  wire [31:0] x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 452:24:@22185.4]
  wire  x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 452:24:@22185.4]
  wire  x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 452:24:@22185.4]
  wire  x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_rr; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 452:24:@22185.4]
  wire  _T_239; // @[package.scala 96:25:@22108.4 package.scala 96:25:@22109.4]
  wire  x485_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[sm_x486_outr_UnitPipe.scala 68:66:@22114.4]
  wire  _T_252; // @[package.scala 96:25:@22150.4 package.scala 96:25:@22151.4]
  wire  _T_258; // @[package.scala 96:25:@22158.4 package.scala 96:25:@22159.4]
  wire  _T_261; // @[SpatialBlocks.scala 110:93:@22161.4]
  wire  x485_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn; // @[SpatialBlocks.scala 110:90:@22162.4]
  wire  _T_263; // @[SpatialBlocks.scala 128:36:@22170.4]
  wire  _T_264; // @[SpatialBlocks.scala 128:78:@22171.4]
  wire  _T_269; // @[SpatialBlocks.scala 130:61:@22180.4]
  x278_ctrchain x278_ctrchain ( // @[SpatialBlocks.scala 37:22:@22016.4]
    .clock(x278_ctrchain_clock),
    .reset(x278_ctrchain_reset),
    .io_input_reset(x278_ctrchain_io_input_reset),
    .io_input_enable(x278_ctrchain_io_input_enable),
    .io_output_counts_1(x278_ctrchain_io_output_counts_1),
    .io_output_counts_0(x278_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x278_ctrchain_io_output_oobs_0),
    .io_output_oobs_1(x278_ctrchain_io_output_oobs_1),
    .io_output_done(x278_ctrchain_io_output_done)
  );
  x485_inr_Foreach_SAMPLER_BOX_sm x485_inr_Foreach_SAMPLER_BOX_sm ( // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 32:18:@22075.4]
    .clock(x485_inr_Foreach_SAMPLER_BOX_sm_clock),
    .reset(x485_inr_Foreach_SAMPLER_BOX_sm_reset),
    .io_enable(x485_inr_Foreach_SAMPLER_BOX_sm_io_enable),
    .io_done(x485_inr_Foreach_SAMPLER_BOX_sm_io_done),
    .io_doneLatch(x485_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch),
    .io_ctrDone(x485_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone),
    .io_datapathEn(x485_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn),
    .io_ctrInc(x485_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc),
    .io_ctrRst(x485_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst),
    .io_parentAck(x485_inr_Foreach_SAMPLER_BOX_sm_io_parentAck),
    .io_backpressure(x485_inr_Foreach_SAMPLER_BOX_sm_io_backpressure),
    .io_break(x485_inr_Foreach_SAMPLER_BOX_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@22103.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@22145.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@22153.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1 x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1 ( // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 452:24:@22185.4]
    .clock(x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_clock),
    .reset(x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_reset),
    .io_in_x270_TREADY(x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x270_TREADY),
    .io_in_x270_TDATA(x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x270_TDATA),
    .io_in_x270_TID(x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x270_TID),
    .io_in_x270_TDEST(x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x270_TDEST),
    .io_in_x271_TVALID(x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x271_TVALID),
    .io_in_x271_TREADY(x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x271_TREADY),
    .io_in_x271_TDATA(x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x271_TDATA),
    .io_sigsIn_backpressure(x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_1(x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsIn_cchainOutputs_0_oobs_1(x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1),
    .io_rr(x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_rr)
  );
  assign _T_239 = RetimeWrapper_io_out; // @[package.scala 96:25:@22108.4 package.scala 96:25:@22109.4]
  assign x485_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure = io_in_x270_TVALID | x485_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x486_outr_UnitPipe.scala 68:66:@22114.4]
  assign _T_252 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@22150.4 package.scala 96:25:@22151.4]
  assign _T_258 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@22158.4 package.scala 96:25:@22159.4]
  assign _T_261 = ~ _T_258; // @[SpatialBlocks.scala 110:93:@22161.4]
  assign x485_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn = _T_252 & _T_261; // @[SpatialBlocks.scala 110:90:@22162.4]
  assign _T_263 = x485_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[SpatialBlocks.scala 128:36:@22170.4]
  assign _T_264 = ~ x485_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[SpatialBlocks.scala 128:78:@22171.4]
  assign _T_269 = x485_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[SpatialBlocks.scala 130:61:@22180.4]
  assign io_in_x270_TREADY = x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x270_TREADY; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 48:23:@22242.4]
  assign io_in_x271_TVALID = x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x271_TVALID; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 49:23:@22252.4]
  assign io_in_x271_TDATA = x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x271_TDATA; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 49:23:@22250.4]
  assign io_sigsOut_smDoneIn_0 = x485_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[SpatialBlocks.scala 127:53:@22168.4]
  assign io_sigsOut_smCtrCopyDone_0 = x485_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[SpatialBlocks.scala 139:125:@22184.4]
  assign x278_ctrchain_clock = clock; // @[:@22017.4]
  assign x278_ctrchain_reset = reset; // @[:@22018.4]
  assign x278_ctrchain_io_input_reset = x485_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[SpatialBlocks.scala 130:103:@22183.4]
  assign x278_ctrchain_io_input_enable = _T_269 & x485_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 104:75:@22138.4 SpatialBlocks.scala 130:45:@22182.4]
  assign x485_inr_Foreach_SAMPLER_BOX_sm_clock = clock; // @[:@22076.4]
  assign x485_inr_Foreach_SAMPLER_BOX_sm_reset = reset; // @[:@22077.4]
  assign x485_inr_Foreach_SAMPLER_BOX_sm_io_enable = x485_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn & x485_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 112:18:@22165.4]
  assign x485_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone = io_rr ? _T_239 : 1'h0; // @[sm_x486_outr_UnitPipe.scala 66:50:@22111.4]
  assign x485_inr_Foreach_SAMPLER_BOX_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 114:21:@22167.4]
  assign x485_inr_Foreach_SAMPLER_BOX_sm_io_backpressure = io_in_x271_TREADY | x485_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[SpatialBlocks.scala 105:24:@22139.4]
  assign x485_inr_Foreach_SAMPLER_BOX_sm_io_break = 1'h0; // @[sm_x486_outr_UnitPipe.scala 70:48:@22117.4]
  assign RetimeWrapper_clock = clock; // @[:@22104.4]
  assign RetimeWrapper_reset = reset; // @[:@22105.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@22107.4]
  assign RetimeWrapper_io_in = x278_ctrchain_io_output_done; // @[package.scala 94:16:@22106.4]
  assign RetimeWrapper_1_clock = clock; // @[:@22146.4]
  assign RetimeWrapper_1_reset = reset; // @[:@22147.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@22149.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@22148.4]
  assign RetimeWrapper_2_clock = clock; // @[:@22154.4]
  assign RetimeWrapper_2_reset = reset; // @[:@22155.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@22157.4]
  assign RetimeWrapper_2_io_in = x485_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[package.scala 94:16:@22156.4]
  assign x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_clock = clock; // @[:@22186.4]
  assign x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_reset = reset; // @[:@22187.4]
  assign x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x270_TDATA = io_in_x270_TDATA; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 48:23:@22241.4]
  assign x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x270_TID = io_in_x270_TID; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 48:23:@22237.4]
  assign x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x270_TDEST = io_in_x270_TDEST; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 48:23:@22236.4]
  assign x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x271_TREADY = io_in_x271_TREADY; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 49:23:@22251.4]
  assign x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure = io_in_x271_TREADY | x485_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 456:22:@22269.4]
  assign x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn = _T_263 & _T_264; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 456:22:@22267.4]
  assign x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break = x485_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 456:22:@22265.4]
  assign x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1 = x278_ctrchain_io_output_counts_1; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 456:22:@22260.4]
  assign x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = x278_ctrchain_io_output_counts_0; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 456:22:@22259.4]
  assign x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x278_ctrchain_io_output_oobs_0; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 456:22:@22257.4]
  assign x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1 = x278_ctrchain_io_output_oobs_1; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 456:22:@22258.4]
  assign x485_inr_Foreach_SAMPLER_BOX_kernelx485_inr_Foreach_SAMPLER_BOX_concrete1_io_rr = io_rr; // @[sm_x485_inr_Foreach_SAMPLER_BOX.scala 455:18:@22253.4]
endmodule
module RootController_kernelRootController_concrete1( // @[:@22282.2]
  input          clock, // @[:@22283.4]
  input          reset, // @[:@22284.4]
  input          io_in_x270_TVALID, // @[:@22285.4]
  output         io_in_x270_TREADY, // @[:@22285.4]
  input  [255:0] io_in_x270_TDATA, // @[:@22285.4]
  input  [7:0]   io_in_x270_TID, // @[:@22285.4]
  input  [7:0]   io_in_x270_TDEST, // @[:@22285.4]
  output         io_in_x271_TVALID, // @[:@22285.4]
  input          io_in_x271_TREADY, // @[:@22285.4]
  output [255:0] io_in_x271_TDATA, // @[:@22285.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@22285.4]
  input          io_sigsIn_smChildAcks_0, // @[:@22285.4]
  output         io_sigsOut_smDoneIn_0, // @[:@22285.4]
  input          io_rr // @[:@22285.4]
);
  wire  x486_outr_UnitPipe_sm_clock; // @[sm_x486_outr_UnitPipe.scala 32:18:@22426.4]
  wire  x486_outr_UnitPipe_sm_reset; // @[sm_x486_outr_UnitPipe.scala 32:18:@22426.4]
  wire  x486_outr_UnitPipe_sm_io_enable; // @[sm_x486_outr_UnitPipe.scala 32:18:@22426.4]
  wire  x486_outr_UnitPipe_sm_io_done; // @[sm_x486_outr_UnitPipe.scala 32:18:@22426.4]
  wire  x486_outr_UnitPipe_sm_io_parentAck; // @[sm_x486_outr_UnitPipe.scala 32:18:@22426.4]
  wire  x486_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x486_outr_UnitPipe.scala 32:18:@22426.4]
  wire  x486_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x486_outr_UnitPipe.scala 32:18:@22426.4]
  wire  x486_outr_UnitPipe_sm_io_childAck_0; // @[sm_x486_outr_UnitPipe.scala 32:18:@22426.4]
  wire  x486_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x486_outr_UnitPipe.scala 32:18:@22426.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@22478.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@22478.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@22478.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@22478.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@22478.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@22486.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@22486.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@22486.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@22486.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@22486.4]
  wire  x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_clock; // @[sm_x486_outr_UnitPipe.scala 75:24:@22513.4]
  wire  x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_reset; // @[sm_x486_outr_UnitPipe.scala 75:24:@22513.4]
  wire  x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_io_in_x270_TVALID; // @[sm_x486_outr_UnitPipe.scala 75:24:@22513.4]
  wire  x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_io_in_x270_TREADY; // @[sm_x486_outr_UnitPipe.scala 75:24:@22513.4]
  wire [255:0] x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_io_in_x270_TDATA; // @[sm_x486_outr_UnitPipe.scala 75:24:@22513.4]
  wire [7:0] x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_io_in_x270_TID; // @[sm_x486_outr_UnitPipe.scala 75:24:@22513.4]
  wire [7:0] x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_io_in_x270_TDEST; // @[sm_x486_outr_UnitPipe.scala 75:24:@22513.4]
  wire  x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_io_in_x271_TVALID; // @[sm_x486_outr_UnitPipe.scala 75:24:@22513.4]
  wire  x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_io_in_x271_TREADY; // @[sm_x486_outr_UnitPipe.scala 75:24:@22513.4]
  wire [255:0] x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_io_in_x271_TDATA; // @[sm_x486_outr_UnitPipe.scala 75:24:@22513.4]
  wire  x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x486_outr_UnitPipe.scala 75:24:@22513.4]
  wire  x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x486_outr_UnitPipe.scala 75:24:@22513.4]
  wire  x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x486_outr_UnitPipe.scala 75:24:@22513.4]
  wire  x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x486_outr_UnitPipe.scala 75:24:@22513.4]
  wire  x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_io_rr; // @[sm_x486_outr_UnitPipe.scala 75:24:@22513.4]
  wire  _T_246; // @[package.scala 96:25:@22483.4 package.scala 96:25:@22484.4]
  wire  _T_252; // @[package.scala 96:25:@22491.4 package.scala 96:25:@22492.4]
  wire  _T_255; // @[SpatialBlocks.scala 110:93:@22494.4]
  x486_outr_UnitPipe_sm x486_outr_UnitPipe_sm ( // @[sm_x486_outr_UnitPipe.scala 32:18:@22426.4]
    .clock(x486_outr_UnitPipe_sm_clock),
    .reset(x486_outr_UnitPipe_sm_reset),
    .io_enable(x486_outr_UnitPipe_sm_io_enable),
    .io_done(x486_outr_UnitPipe_sm_io_done),
    .io_parentAck(x486_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x486_outr_UnitPipe_sm_io_doneIn_0),
    .io_enableOut_0(x486_outr_UnitPipe_sm_io_enableOut_0),
    .io_childAck_0(x486_outr_UnitPipe_sm_io_childAck_0),
    .io_ctrCopyDone_0(x486_outr_UnitPipe_sm_io_ctrCopyDone_0)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@22478.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@22486.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1 x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1 ( // @[sm_x486_outr_UnitPipe.scala 75:24:@22513.4]
    .clock(x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_clock),
    .reset(x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_reset),
    .io_in_x270_TVALID(x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_io_in_x270_TVALID),
    .io_in_x270_TREADY(x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_io_in_x270_TREADY),
    .io_in_x270_TDATA(x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_io_in_x270_TDATA),
    .io_in_x270_TID(x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_io_in_x270_TID),
    .io_in_x270_TDEST(x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_io_in_x270_TDEST),
    .io_in_x271_TVALID(x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_io_in_x271_TVALID),
    .io_in_x271_TREADY(x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_io_in_x271_TREADY),
    .io_in_x271_TDATA(x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_io_in_x271_TDATA),
    .io_sigsIn_smEnableOuts_0(x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smCtrCopyDone_0(x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_rr(x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_246 = RetimeWrapper_io_out; // @[package.scala 96:25:@22483.4 package.scala 96:25:@22484.4]
  assign _T_252 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@22491.4 package.scala 96:25:@22492.4]
  assign _T_255 = ~ _T_252; // @[SpatialBlocks.scala 110:93:@22494.4]
  assign io_in_x270_TREADY = x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_io_in_x270_TREADY; // @[sm_x486_outr_UnitPipe.scala 48:23:@22568.4]
  assign io_in_x271_TVALID = x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_io_in_x271_TVALID; // @[sm_x486_outr_UnitPipe.scala 49:23:@22578.4]
  assign io_in_x271_TDATA = x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_io_in_x271_TDATA; // @[sm_x486_outr_UnitPipe.scala 49:23:@22576.4]
  assign io_sigsOut_smDoneIn_0 = x486_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 127:53:@22501.4]
  assign x486_outr_UnitPipe_sm_clock = clock; // @[:@22427.4]
  assign x486_outr_UnitPipe_sm_reset = reset; // @[:@22428.4]
  assign x486_outr_UnitPipe_sm_io_enable = _T_246 & _T_255; // @[SpatialBlocks.scala 112:18:@22498.4]
  assign x486_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 114:21:@22500.4]
  assign x486_outr_UnitPipe_sm_io_doneIn_0 = x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 102:67:@22470.4]
  assign x486_outr_UnitPipe_sm_io_ctrCopyDone_0 = x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 132:80:@22512.4]
  assign RetimeWrapper_clock = clock; // @[:@22479.4]
  assign RetimeWrapper_reset = reset; // @[:@22480.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@22482.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@22481.4]
  assign RetimeWrapper_1_clock = clock; // @[:@22487.4]
  assign RetimeWrapper_1_reset = reset; // @[:@22488.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@22490.4]
  assign RetimeWrapper_1_io_in = x486_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@22489.4]
  assign x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_clock = clock; // @[:@22514.4]
  assign x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_reset = reset; // @[:@22515.4]
  assign x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_io_in_x270_TVALID = io_in_x270_TVALID; // @[sm_x486_outr_UnitPipe.scala 48:23:@22569.4]
  assign x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_io_in_x270_TDATA = io_in_x270_TDATA; // @[sm_x486_outr_UnitPipe.scala 48:23:@22567.4]
  assign x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_io_in_x270_TID = io_in_x270_TID; // @[sm_x486_outr_UnitPipe.scala 48:23:@22563.4]
  assign x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_io_in_x270_TDEST = io_in_x270_TDEST; // @[sm_x486_outr_UnitPipe.scala 48:23:@22562.4]
  assign x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_io_in_x271_TREADY = io_in_x271_TREADY; // @[sm_x486_outr_UnitPipe.scala 49:23:@22577.4]
  assign x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x486_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x486_outr_UnitPipe.scala 79:22:@22587.4]
  assign x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x486_outr_UnitPipe_sm_io_childAck_0; // @[sm_x486_outr_UnitPipe.scala 79:22:@22585.4]
  assign x486_outr_UnitPipe_kernelx486_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x486_outr_UnitPipe.scala 78:18:@22579.4]
endmodule
module AccelUnit( // @[:@22606.2]
  input          clock, // @[:@22607.4]
  input          reset, // @[:@22608.4]
  input          io_enable, // @[:@22609.4]
  output         io_done, // @[:@22609.4]
  input          io_reset, // @[:@22609.4]
  input          io_memStreams_loads_0_cmd_ready, // @[:@22609.4]
  output         io_memStreams_loads_0_cmd_valid, // @[:@22609.4]
  output [63:0]  io_memStreams_loads_0_cmd_bits_addr, // @[:@22609.4]
  output [31:0]  io_memStreams_loads_0_cmd_bits_size, // @[:@22609.4]
  output         io_memStreams_loads_0_data_ready, // @[:@22609.4]
  input          io_memStreams_loads_0_data_valid, // @[:@22609.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_0, // @[:@22609.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_1, // @[:@22609.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_2, // @[:@22609.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_3, // @[:@22609.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_4, // @[:@22609.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_5, // @[:@22609.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_6, // @[:@22609.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_7, // @[:@22609.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_8, // @[:@22609.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_9, // @[:@22609.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_10, // @[:@22609.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_11, // @[:@22609.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_12, // @[:@22609.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_13, // @[:@22609.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_14, // @[:@22609.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_15, // @[:@22609.4]
  input          io_memStreams_stores_0_cmd_ready, // @[:@22609.4]
  output         io_memStreams_stores_0_cmd_valid, // @[:@22609.4]
  output [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@22609.4]
  output [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@22609.4]
  input          io_memStreams_stores_0_data_ready, // @[:@22609.4]
  output         io_memStreams_stores_0_data_valid, // @[:@22609.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_0, // @[:@22609.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_1, // @[:@22609.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_2, // @[:@22609.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_3, // @[:@22609.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_4, // @[:@22609.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_5, // @[:@22609.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_6, // @[:@22609.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_7, // @[:@22609.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_8, // @[:@22609.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_9, // @[:@22609.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_10, // @[:@22609.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_11, // @[:@22609.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_12, // @[:@22609.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_13, // @[:@22609.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_14, // @[:@22609.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_15, // @[:@22609.4]
  output [15:0]  io_memStreams_stores_0_data_bits_wstrb, // @[:@22609.4]
  output         io_memStreams_stores_0_wresp_ready, // @[:@22609.4]
  input          io_memStreams_stores_0_wresp_valid, // @[:@22609.4]
  input          io_memStreams_stores_0_wresp_bits, // @[:@22609.4]
  input          io_memStreams_gathers_0_cmd_ready, // @[:@22609.4]
  output         io_memStreams_gathers_0_cmd_valid, // @[:@22609.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_0, // @[:@22609.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_1, // @[:@22609.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_2, // @[:@22609.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_3, // @[:@22609.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_4, // @[:@22609.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_5, // @[:@22609.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_6, // @[:@22609.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_7, // @[:@22609.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_8, // @[:@22609.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_9, // @[:@22609.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_10, // @[:@22609.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_11, // @[:@22609.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_12, // @[:@22609.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_13, // @[:@22609.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_14, // @[:@22609.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_15, // @[:@22609.4]
  output         io_memStreams_gathers_0_data_ready, // @[:@22609.4]
  input          io_memStreams_gathers_0_data_valid, // @[:@22609.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_0, // @[:@22609.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_1, // @[:@22609.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_2, // @[:@22609.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_3, // @[:@22609.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_4, // @[:@22609.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_5, // @[:@22609.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_6, // @[:@22609.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_7, // @[:@22609.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_8, // @[:@22609.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_9, // @[:@22609.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_10, // @[:@22609.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_11, // @[:@22609.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_12, // @[:@22609.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_13, // @[:@22609.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_14, // @[:@22609.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_15, // @[:@22609.4]
  input          io_memStreams_scatters_0_cmd_ready, // @[:@22609.4]
  output         io_memStreams_scatters_0_cmd_valid, // @[:@22609.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_0, // @[:@22609.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_1, // @[:@22609.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_2, // @[:@22609.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_3, // @[:@22609.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_4, // @[:@22609.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_5, // @[:@22609.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_6, // @[:@22609.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_7, // @[:@22609.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_8, // @[:@22609.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_9, // @[:@22609.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_10, // @[:@22609.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_11, // @[:@22609.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_12, // @[:@22609.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_13, // @[:@22609.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_14, // @[:@22609.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_15, // @[:@22609.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_0, // @[:@22609.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_1, // @[:@22609.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_2, // @[:@22609.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_3, // @[:@22609.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_4, // @[:@22609.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_5, // @[:@22609.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_6, // @[:@22609.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_7, // @[:@22609.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_8, // @[:@22609.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_9, // @[:@22609.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_10, // @[:@22609.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_11, // @[:@22609.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_12, // @[:@22609.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_13, // @[:@22609.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_14, // @[:@22609.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_15, // @[:@22609.4]
  output         io_memStreams_scatters_0_wresp_ready, // @[:@22609.4]
  input          io_memStreams_scatters_0_wresp_valid, // @[:@22609.4]
  input          io_memStreams_scatters_0_wresp_bits, // @[:@22609.4]
  input          io_axiStreamsIn_0_TVALID, // @[:@22609.4]
  output         io_axiStreamsIn_0_TREADY, // @[:@22609.4]
  input  [255:0] io_axiStreamsIn_0_TDATA, // @[:@22609.4]
  input  [31:0]  io_axiStreamsIn_0_TSTRB, // @[:@22609.4]
  input  [31:0]  io_axiStreamsIn_0_TKEEP, // @[:@22609.4]
  input          io_axiStreamsIn_0_TLAST, // @[:@22609.4]
  input  [7:0]   io_axiStreamsIn_0_TID, // @[:@22609.4]
  input  [7:0]   io_axiStreamsIn_0_TDEST, // @[:@22609.4]
  input  [31:0]  io_axiStreamsIn_0_TUSER, // @[:@22609.4]
  output         io_axiStreamsOut_0_TVALID, // @[:@22609.4]
  input          io_axiStreamsOut_0_TREADY, // @[:@22609.4]
  output [255:0] io_axiStreamsOut_0_TDATA, // @[:@22609.4]
  output [31:0]  io_axiStreamsOut_0_TSTRB, // @[:@22609.4]
  output [31:0]  io_axiStreamsOut_0_TKEEP, // @[:@22609.4]
  output         io_axiStreamsOut_0_TLAST, // @[:@22609.4]
  output [7:0]   io_axiStreamsOut_0_TID, // @[:@22609.4]
  output [7:0]   io_axiStreamsOut_0_TDEST, // @[:@22609.4]
  output [31:0]  io_axiStreamsOut_0_TUSER, // @[:@22609.4]
  output         io_heap_0_req_valid, // @[:@22609.4]
  output         io_heap_0_req_bits_allocDealloc, // @[:@22609.4]
  output [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@22609.4]
  input          io_heap_0_resp_valid, // @[:@22609.4]
  input          io_heap_0_resp_bits_allocDealloc, // @[:@22609.4]
  input  [63:0]  io_heap_0_resp_bits_sizeAddr, // @[:@22609.4]
  input  [63:0]  io_argIns_0, // @[:@22609.4]
  input  [63:0]  io_argIns_1, // @[:@22609.4]
  input          io_argOuts_0_port_ready, // @[:@22609.4]
  output         io_argOuts_0_port_valid, // @[:@22609.4]
  output [63:0]  io_argOuts_0_port_bits, // @[:@22609.4]
  input  [63:0]  io_argOuts_0_echo // @[:@22609.4]
);
  wire  SingleCounter_clock; // @[Main.scala 35:32:@22772.4]
  wire  SingleCounter_reset; // @[Main.scala 35:32:@22772.4]
  wire  SingleCounter_io_input_reset; // @[Main.scala 35:32:@22772.4]
  wire  SingleCounter_io_output_done; // @[Main.scala 35:32:@22772.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@22790.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@22790.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@22790.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@22790.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@22790.4]
  wire  SRFF_clock; // @[Main.scala 39:28:@22799.4]
  wire  SRFF_reset; // @[Main.scala 39:28:@22799.4]
  wire  SRFF_io_input_set; // @[Main.scala 39:28:@22799.4]
  wire  SRFF_io_input_reset; // @[Main.scala 39:28:@22799.4]
  wire  SRFF_io_input_asyn_reset; // @[Main.scala 39:28:@22799.4]
  wire  SRFF_io_output; // @[Main.scala 39:28:@22799.4]
  wire  RootController_sm_clock; // @[sm_RootController.scala 32:18:@22837.4]
  wire  RootController_sm_reset; // @[sm_RootController.scala 32:18:@22837.4]
  wire  RootController_sm_io_enable; // @[sm_RootController.scala 32:18:@22837.4]
  wire  RootController_sm_io_done; // @[sm_RootController.scala 32:18:@22837.4]
  wire  RootController_sm_io_rst; // @[sm_RootController.scala 32:18:@22837.4]
  wire  RootController_sm_io_ctrDone; // @[sm_RootController.scala 32:18:@22837.4]
  wire  RootController_sm_io_ctrInc; // @[sm_RootController.scala 32:18:@22837.4]
  wire  RootController_sm_io_doneIn_0; // @[sm_RootController.scala 32:18:@22837.4]
  wire  RootController_sm_io_enableOut_0; // @[sm_RootController.scala 32:18:@22837.4]
  wire  RootController_sm_io_childAck_0; // @[sm_RootController.scala 32:18:@22837.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@22869.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@22869.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@22869.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@22869.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@22869.4]
  wire  RootController_kernelRootController_concrete1_clock; // @[sm_RootController.scala 73:24:@22928.4]
  wire  RootController_kernelRootController_concrete1_reset; // @[sm_RootController.scala 73:24:@22928.4]
  wire  RootController_kernelRootController_concrete1_io_in_x270_TVALID; // @[sm_RootController.scala 73:24:@22928.4]
  wire  RootController_kernelRootController_concrete1_io_in_x270_TREADY; // @[sm_RootController.scala 73:24:@22928.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x270_TDATA; // @[sm_RootController.scala 73:24:@22928.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x270_TID; // @[sm_RootController.scala 73:24:@22928.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x270_TDEST; // @[sm_RootController.scala 73:24:@22928.4]
  wire  RootController_kernelRootController_concrete1_io_in_x271_TVALID; // @[sm_RootController.scala 73:24:@22928.4]
  wire  RootController_kernelRootController_concrete1_io_in_x271_TREADY; // @[sm_RootController.scala 73:24:@22928.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x271_TDATA; // @[sm_RootController.scala 73:24:@22928.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_RootController.scala 73:24:@22928.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0; // @[sm_RootController.scala 73:24:@22928.4]
  wire  RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[sm_RootController.scala 73:24:@22928.4]
  wire  RootController_kernelRootController_concrete1_io_rr; // @[sm_RootController.scala 73:24:@22928.4]
  wire  _T_599; // @[package.scala 96:25:@22795.4 package.scala 96:25:@22796.4]
  wire  _T_664; // @[Main.scala 41:50:@22865.4]
  wire  _T_665; // @[Main.scala 41:59:@22866.4]
  wire  _T_677; // @[package.scala 100:49:@22886.4]
  reg  _T_680; // @[package.scala 48:56:@22887.4]
  reg [31:0] _RAND_0;
  SingleCounter SingleCounter ( // @[Main.scala 35:32:@22772.4]
    .clock(SingleCounter_clock),
    .reset(SingleCounter_reset),
    .io_input_reset(SingleCounter_io_input_reset),
    .io_output_done(SingleCounter_io_output_done)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@22790.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  SRFF SRFF ( // @[Main.scala 39:28:@22799.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  RootController_sm RootController_sm ( // @[sm_RootController.scala 32:18:@22837.4]
    .clock(RootController_sm_clock),
    .reset(RootController_sm_reset),
    .io_enable(RootController_sm_io_enable),
    .io_done(RootController_sm_io_done),
    .io_rst(RootController_sm_io_rst),
    .io_ctrDone(RootController_sm_io_ctrDone),
    .io_ctrInc(RootController_sm_io_ctrInc),
    .io_doneIn_0(RootController_sm_io_doneIn_0),
    .io_enableOut_0(RootController_sm_io_enableOut_0),
    .io_childAck_0(RootController_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@22869.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RootController_kernelRootController_concrete1 RootController_kernelRootController_concrete1 ( // @[sm_RootController.scala 73:24:@22928.4]
    .clock(RootController_kernelRootController_concrete1_clock),
    .reset(RootController_kernelRootController_concrete1_reset),
    .io_in_x270_TVALID(RootController_kernelRootController_concrete1_io_in_x270_TVALID),
    .io_in_x270_TREADY(RootController_kernelRootController_concrete1_io_in_x270_TREADY),
    .io_in_x270_TDATA(RootController_kernelRootController_concrete1_io_in_x270_TDATA),
    .io_in_x270_TID(RootController_kernelRootController_concrete1_io_in_x270_TID),
    .io_in_x270_TDEST(RootController_kernelRootController_concrete1_io_in_x270_TDEST),
    .io_in_x271_TVALID(RootController_kernelRootController_concrete1_io_in_x271_TVALID),
    .io_in_x271_TREADY(RootController_kernelRootController_concrete1_io_in_x271_TREADY),
    .io_in_x271_TDATA(RootController_kernelRootController_concrete1_io_in_x271_TDATA),
    .io_sigsIn_smEnableOuts_0(RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(RootController_kernelRootController_concrete1_io_rr)
  );
  assign _T_599 = RetimeWrapper_io_out; // @[package.scala 96:25:@22795.4 package.scala 96:25:@22796.4]
  assign _T_664 = io_enable & _T_599; // @[Main.scala 41:50:@22865.4]
  assign _T_665 = ~ SRFF_io_output; // @[Main.scala 41:59:@22866.4]
  assign _T_677 = RootController_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@22886.4]
  assign io_done = SRFF_io_output; // @[Main.scala 48:23:@22885.4]
  assign io_memStreams_loads_0_cmd_valid = 1'h0;
  assign io_memStreams_loads_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_loads_0_cmd_bits_size = 32'h0;
  assign io_memStreams_loads_0_data_ready = 1'h0;
  assign io_memStreams_stores_0_cmd_valid = 1'h0;
  assign io_memStreams_stores_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_stores_0_cmd_bits_size = 32'h0;
  assign io_memStreams_stores_0_data_valid = 1'h0;
  assign io_memStreams_stores_0_data_bits_wdata_0 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_1 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_2 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_3 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_4 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_5 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_6 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_7 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_8 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_9 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_10 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_11 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_12 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_13 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_14 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_15 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wstrb = 16'h0;
  assign io_memStreams_stores_0_wresp_ready = 1'h0;
  assign io_memStreams_gathers_0_cmd_valid = 1'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_0 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_1 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_2 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_3 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_4 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_5 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_6 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_7 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_8 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_9 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_10 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_11 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_12 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_13 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_14 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_15 = 64'h0;
  assign io_memStreams_gathers_0_data_ready = 1'h0;
  assign io_memStreams_scatters_0_cmd_valid = 1'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_0 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_1 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_2 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_3 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_4 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_5 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_6 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_7 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_8 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_9 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_10 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_11 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_12 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_13 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_14 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_15 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_0 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_1 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_2 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_3 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_4 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_5 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_6 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_7 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_8 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_9 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_10 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_11 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_12 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_13 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_14 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_15 = 32'h0;
  assign io_memStreams_scatters_0_wresp_ready = 1'h0;
  assign io_axiStreamsIn_0_TREADY = RootController_kernelRootController_concrete1_io_in_x270_TREADY; // @[sm_RootController.scala 48:23:@22983.4]
  assign io_axiStreamsOut_0_TVALID = RootController_kernelRootController_concrete1_io_in_x271_TVALID; // @[sm_RootController.scala 49:23:@22993.4]
  assign io_axiStreamsOut_0_TDATA = RootController_kernelRootController_concrete1_io_in_x271_TDATA; // @[sm_RootController.scala 49:23:@22991.4]
  assign io_axiStreamsOut_0_TSTRB = 32'hffffffff; // @[sm_RootController.scala 49:23:@22990.4]
  assign io_axiStreamsOut_0_TKEEP = 32'hffffffff; // @[sm_RootController.scala 49:23:@22989.4]
  assign io_axiStreamsOut_0_TLAST = 1'h0; // @[sm_RootController.scala 49:23:@22988.4]
  assign io_axiStreamsOut_0_TID = 8'h0; // @[sm_RootController.scala 49:23:@22987.4]
  assign io_axiStreamsOut_0_TDEST = 8'h0; // @[sm_RootController.scala 49:23:@22986.4]
  assign io_axiStreamsOut_0_TUSER = 32'h4; // @[sm_RootController.scala 49:23:@22985.4]
  assign io_heap_0_req_valid = 1'h0;
  assign io_heap_0_req_bits_allocDealloc = 1'h0;
  assign io_heap_0_req_bits_sizeAddr = 64'h0;
  assign io_argOuts_0_port_valid = 1'h0;
  assign io_argOuts_0_port_bits = 64'h0;
  assign SingleCounter_clock = clock; // @[:@22773.4]
  assign SingleCounter_reset = reset; // @[:@22774.4]
  assign SingleCounter_io_input_reset = reset; // @[Main.scala 36:79:@22788.4]
  assign RetimeWrapper_clock = clock; // @[:@22791.4]
  assign RetimeWrapper_reset = reset; // @[:@22792.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@22794.4]
  assign RetimeWrapper_io_in = SingleCounter_io_output_done; // @[package.scala 94:16:@22793.4]
  assign SRFF_clock = clock; // @[:@22800.4]
  assign SRFF_reset = reset; // @[:@22801.4]
  assign SRFF_io_input_set = RootController_sm_io_done; // @[Main.scala 57:29:@23020.4]
  assign SRFF_io_input_reset = RetimeWrapper_1_io_out; // @[Main.scala 46:31:@22883.4]
  assign SRFF_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[Main.scala 47:36:@22884.4]
  assign RootController_sm_clock = clock; // @[:@22838.4]
  assign RootController_sm_reset = reset; // @[:@22839.4]
  assign RootController_sm_io_enable = _T_664 & _T_665; // @[Main.scala 45:33:@22882.4 SpatialBlocks.scala 112:18:@22916.4]
  assign RootController_sm_io_rst = RetimeWrapper_1_io_out; // @[SpatialBlocks.scala 106:15:@22910.4]
  assign RootController_sm_io_ctrDone = RootController_sm_io_ctrInc & _T_680; // @[Main.scala 49:34:@22890.4]
  assign RootController_sm_io_doneIn_0 = RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 102:67:@22907.4]
  assign RetimeWrapper_1_clock = clock; // @[:@22870.4]
  assign RetimeWrapper_1_reset = reset; // @[:@22871.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@22873.4]
  assign RetimeWrapper_1_io_in = reset | io_reset; // @[package.scala 94:16:@22872.4]
  assign RootController_kernelRootController_concrete1_clock = clock; // @[:@22929.4]
  assign RootController_kernelRootController_concrete1_reset = reset; // @[:@22930.4]
  assign RootController_kernelRootController_concrete1_io_in_x270_TVALID = io_axiStreamsIn_0_TVALID; // @[sm_RootController.scala 48:23:@22984.4]
  assign RootController_kernelRootController_concrete1_io_in_x270_TDATA = io_axiStreamsIn_0_TDATA; // @[sm_RootController.scala 48:23:@22982.4]
  assign RootController_kernelRootController_concrete1_io_in_x270_TID = io_axiStreamsIn_0_TID; // @[sm_RootController.scala 48:23:@22978.4]
  assign RootController_kernelRootController_concrete1_io_in_x270_TDEST = io_axiStreamsIn_0_TDEST; // @[sm_RootController.scala 48:23:@22977.4]
  assign RootController_kernelRootController_concrete1_io_in_x271_TREADY = io_axiStreamsOut_0_TREADY; // @[sm_RootController.scala 49:23:@22992.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0 = RootController_sm_io_enableOut_0; // @[sm_RootController.scala 77:22:@23002.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0 = RootController_sm_io_childAck_0; // @[sm_RootController.scala 77:22:@23000.4]
  assign RootController_kernelRootController_concrete1_io_rr = RetimeWrapper_io_out; // @[sm_RootController.scala 76:18:@22994.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_680 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_680 <= 1'h0;
    end else begin
      _T_680 <= _T_677;
    end
  end
endmodule
module SpatialIP( // @[:@23022.2]
  input         clock, // @[:@23023.4]
  input         reset, // @[:@23024.4]
  input  [31:0] io_raddr, // @[:@23025.4]
  input         io_wen, // @[:@23025.4]
  input  [31:0] io_waddr, // @[:@23025.4]
  input  [63:0] io_wdata, // @[:@23025.4]
  output [63:0] io_rdata // @[:@23025.4]
);
  wire  accel_clock; // @[Instantiator.scala 53:44:@23027.4]
  wire  accel_reset; // @[Instantiator.scala 53:44:@23027.4]
  wire  accel_io_enable; // @[Instantiator.scala 53:44:@23027.4]
  wire  accel_io_done; // @[Instantiator.scala 53:44:@23027.4]
  wire  accel_io_reset; // @[Instantiator.scala 53:44:@23027.4]
  wire  accel_io_memStreams_loads_0_cmd_ready; // @[Instantiator.scala 53:44:@23027.4]
  wire  accel_io_memStreams_loads_0_cmd_valid; // @[Instantiator.scala 53:44:@23027.4]
  wire [63:0] accel_io_memStreams_loads_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_loads_0_cmd_bits_size; // @[Instantiator.scala 53:44:@23027.4]
  wire  accel_io_memStreams_loads_0_data_ready; // @[Instantiator.scala 53:44:@23027.4]
  wire  accel_io_memStreams_loads_0_data_valid; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_0; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_1; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_2; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_3; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_4; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_5; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_6; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_7; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_8; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_9; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_10; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_11; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_12; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_13; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_14; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_15; // @[Instantiator.scala 53:44:@23027.4]
  wire  accel_io_memStreams_stores_0_cmd_ready; // @[Instantiator.scala 53:44:@23027.4]
  wire  accel_io_memStreams_stores_0_cmd_valid; // @[Instantiator.scala 53:44:@23027.4]
  wire [63:0] accel_io_memStreams_stores_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_stores_0_cmd_bits_size; // @[Instantiator.scala 53:44:@23027.4]
  wire  accel_io_memStreams_stores_0_data_ready; // @[Instantiator.scala 53:44:@23027.4]
  wire  accel_io_memStreams_stores_0_data_valid; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_1; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_2; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_3; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_4; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_5; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_6; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_7; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_8; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_9; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_10; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_11; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_12; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_13; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_14; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_15; // @[Instantiator.scala 53:44:@23027.4]
  wire [15:0] accel_io_memStreams_stores_0_data_bits_wstrb; // @[Instantiator.scala 53:44:@23027.4]
  wire  accel_io_memStreams_stores_0_wresp_ready; // @[Instantiator.scala 53:44:@23027.4]
  wire  accel_io_memStreams_stores_0_wresp_valid; // @[Instantiator.scala 53:44:@23027.4]
  wire  accel_io_memStreams_stores_0_wresp_bits; // @[Instantiator.scala 53:44:@23027.4]
  wire  accel_io_memStreams_gathers_0_cmd_ready; // @[Instantiator.scala 53:44:@23027.4]
  wire  accel_io_memStreams_gathers_0_cmd_valid; // @[Instantiator.scala 53:44:@23027.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_0; // @[Instantiator.scala 53:44:@23027.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_1; // @[Instantiator.scala 53:44:@23027.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_2; // @[Instantiator.scala 53:44:@23027.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_3; // @[Instantiator.scala 53:44:@23027.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_4; // @[Instantiator.scala 53:44:@23027.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_5; // @[Instantiator.scala 53:44:@23027.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_6; // @[Instantiator.scala 53:44:@23027.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_7; // @[Instantiator.scala 53:44:@23027.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_8; // @[Instantiator.scala 53:44:@23027.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_9; // @[Instantiator.scala 53:44:@23027.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_10; // @[Instantiator.scala 53:44:@23027.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_11; // @[Instantiator.scala 53:44:@23027.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_12; // @[Instantiator.scala 53:44:@23027.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_13; // @[Instantiator.scala 53:44:@23027.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_14; // @[Instantiator.scala 53:44:@23027.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_15; // @[Instantiator.scala 53:44:@23027.4]
  wire  accel_io_memStreams_gathers_0_data_ready; // @[Instantiator.scala 53:44:@23027.4]
  wire  accel_io_memStreams_gathers_0_data_valid; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_0; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_1; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_2; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_3; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_4; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_5; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_6; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_7; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_8; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_9; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_10; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_11; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_12; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_13; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_14; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_15; // @[Instantiator.scala 53:44:@23027.4]
  wire  accel_io_memStreams_scatters_0_cmd_ready; // @[Instantiator.scala 53:44:@23027.4]
  wire  accel_io_memStreams_scatters_0_cmd_valid; // @[Instantiator.scala 53:44:@23027.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0; // @[Instantiator.scala 53:44:@23027.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1; // @[Instantiator.scala 53:44:@23027.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2; // @[Instantiator.scala 53:44:@23027.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3; // @[Instantiator.scala 53:44:@23027.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4; // @[Instantiator.scala 53:44:@23027.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5; // @[Instantiator.scala 53:44:@23027.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6; // @[Instantiator.scala 53:44:@23027.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7; // @[Instantiator.scala 53:44:@23027.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8; // @[Instantiator.scala 53:44:@23027.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9; // @[Instantiator.scala 53:44:@23027.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10; // @[Instantiator.scala 53:44:@23027.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11; // @[Instantiator.scala 53:44:@23027.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12; // @[Instantiator.scala 53:44:@23027.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13; // @[Instantiator.scala 53:44:@23027.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14; // @[Instantiator.scala 53:44:@23027.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_0; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_1; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_2; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_3; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_4; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_5; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_6; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_7; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_8; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_9; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_10; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_11; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_12; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_13; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_14; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_15; // @[Instantiator.scala 53:44:@23027.4]
  wire  accel_io_memStreams_scatters_0_wresp_ready; // @[Instantiator.scala 53:44:@23027.4]
  wire  accel_io_memStreams_scatters_0_wresp_valid; // @[Instantiator.scala 53:44:@23027.4]
  wire  accel_io_memStreams_scatters_0_wresp_bits; // @[Instantiator.scala 53:44:@23027.4]
  wire  accel_io_axiStreamsIn_0_TVALID; // @[Instantiator.scala 53:44:@23027.4]
  wire  accel_io_axiStreamsIn_0_TREADY; // @[Instantiator.scala 53:44:@23027.4]
  wire [255:0] accel_io_axiStreamsIn_0_TDATA; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_axiStreamsIn_0_TSTRB; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_axiStreamsIn_0_TKEEP; // @[Instantiator.scala 53:44:@23027.4]
  wire  accel_io_axiStreamsIn_0_TLAST; // @[Instantiator.scala 53:44:@23027.4]
  wire [7:0] accel_io_axiStreamsIn_0_TID; // @[Instantiator.scala 53:44:@23027.4]
  wire [7:0] accel_io_axiStreamsIn_0_TDEST; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_axiStreamsIn_0_TUSER; // @[Instantiator.scala 53:44:@23027.4]
  wire  accel_io_axiStreamsOut_0_TVALID; // @[Instantiator.scala 53:44:@23027.4]
  wire  accel_io_axiStreamsOut_0_TREADY; // @[Instantiator.scala 53:44:@23027.4]
  wire [255:0] accel_io_axiStreamsOut_0_TDATA; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_axiStreamsOut_0_TSTRB; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_axiStreamsOut_0_TKEEP; // @[Instantiator.scala 53:44:@23027.4]
  wire  accel_io_axiStreamsOut_0_TLAST; // @[Instantiator.scala 53:44:@23027.4]
  wire [7:0] accel_io_axiStreamsOut_0_TID; // @[Instantiator.scala 53:44:@23027.4]
  wire [7:0] accel_io_axiStreamsOut_0_TDEST; // @[Instantiator.scala 53:44:@23027.4]
  wire [31:0] accel_io_axiStreamsOut_0_TUSER; // @[Instantiator.scala 53:44:@23027.4]
  wire  accel_io_heap_0_req_valid; // @[Instantiator.scala 53:44:@23027.4]
  wire  accel_io_heap_0_req_bits_allocDealloc; // @[Instantiator.scala 53:44:@23027.4]
  wire [63:0] accel_io_heap_0_req_bits_sizeAddr; // @[Instantiator.scala 53:44:@23027.4]
  wire  accel_io_heap_0_resp_valid; // @[Instantiator.scala 53:44:@23027.4]
  wire  accel_io_heap_0_resp_bits_allocDealloc; // @[Instantiator.scala 53:44:@23027.4]
  wire [63:0] accel_io_heap_0_resp_bits_sizeAddr; // @[Instantiator.scala 53:44:@23027.4]
  wire [63:0] accel_io_argIns_0; // @[Instantiator.scala 53:44:@23027.4]
  wire [63:0] accel_io_argIns_1; // @[Instantiator.scala 53:44:@23027.4]
  wire  accel_io_argOuts_0_port_ready; // @[Instantiator.scala 53:44:@23027.4]
  wire  accel_io_argOuts_0_port_valid; // @[Instantiator.scala 53:44:@23027.4]
  wire [63:0] accel_io_argOuts_0_port_bits; // @[Instantiator.scala 53:44:@23027.4]
  wire [63:0] accel_io_argOuts_0_echo; // @[Instantiator.scala 53:44:@23027.4]
  AccelUnit accel ( // @[Instantiator.scala 53:44:@23027.4]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_enable(accel_io_enable),
    .io_done(accel_io_done),
    .io_reset(accel_io_reset),
    .io_memStreams_loads_0_cmd_ready(accel_io_memStreams_loads_0_cmd_ready),
    .io_memStreams_loads_0_cmd_valid(accel_io_memStreams_loads_0_cmd_valid),
    .io_memStreams_loads_0_cmd_bits_addr(accel_io_memStreams_loads_0_cmd_bits_addr),
    .io_memStreams_loads_0_cmd_bits_size(accel_io_memStreams_loads_0_cmd_bits_size),
    .io_memStreams_loads_0_data_ready(accel_io_memStreams_loads_0_data_ready),
    .io_memStreams_loads_0_data_valid(accel_io_memStreams_loads_0_data_valid),
    .io_memStreams_loads_0_data_bits_rdata_0(accel_io_memStreams_loads_0_data_bits_rdata_0),
    .io_memStreams_loads_0_data_bits_rdata_1(accel_io_memStreams_loads_0_data_bits_rdata_1),
    .io_memStreams_loads_0_data_bits_rdata_2(accel_io_memStreams_loads_0_data_bits_rdata_2),
    .io_memStreams_loads_0_data_bits_rdata_3(accel_io_memStreams_loads_0_data_bits_rdata_3),
    .io_memStreams_loads_0_data_bits_rdata_4(accel_io_memStreams_loads_0_data_bits_rdata_4),
    .io_memStreams_loads_0_data_bits_rdata_5(accel_io_memStreams_loads_0_data_bits_rdata_5),
    .io_memStreams_loads_0_data_bits_rdata_6(accel_io_memStreams_loads_0_data_bits_rdata_6),
    .io_memStreams_loads_0_data_bits_rdata_7(accel_io_memStreams_loads_0_data_bits_rdata_7),
    .io_memStreams_loads_0_data_bits_rdata_8(accel_io_memStreams_loads_0_data_bits_rdata_8),
    .io_memStreams_loads_0_data_bits_rdata_9(accel_io_memStreams_loads_0_data_bits_rdata_9),
    .io_memStreams_loads_0_data_bits_rdata_10(accel_io_memStreams_loads_0_data_bits_rdata_10),
    .io_memStreams_loads_0_data_bits_rdata_11(accel_io_memStreams_loads_0_data_bits_rdata_11),
    .io_memStreams_loads_0_data_bits_rdata_12(accel_io_memStreams_loads_0_data_bits_rdata_12),
    .io_memStreams_loads_0_data_bits_rdata_13(accel_io_memStreams_loads_0_data_bits_rdata_13),
    .io_memStreams_loads_0_data_bits_rdata_14(accel_io_memStreams_loads_0_data_bits_rdata_14),
    .io_memStreams_loads_0_data_bits_rdata_15(accel_io_memStreams_loads_0_data_bits_rdata_15),
    .io_memStreams_stores_0_cmd_ready(accel_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(accel_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(accel_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(accel_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(accel_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(accel_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(accel_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wdata_1(accel_io_memStreams_stores_0_data_bits_wdata_1),
    .io_memStreams_stores_0_data_bits_wdata_2(accel_io_memStreams_stores_0_data_bits_wdata_2),
    .io_memStreams_stores_0_data_bits_wdata_3(accel_io_memStreams_stores_0_data_bits_wdata_3),
    .io_memStreams_stores_0_data_bits_wdata_4(accel_io_memStreams_stores_0_data_bits_wdata_4),
    .io_memStreams_stores_0_data_bits_wdata_5(accel_io_memStreams_stores_0_data_bits_wdata_5),
    .io_memStreams_stores_0_data_bits_wdata_6(accel_io_memStreams_stores_0_data_bits_wdata_6),
    .io_memStreams_stores_0_data_bits_wdata_7(accel_io_memStreams_stores_0_data_bits_wdata_7),
    .io_memStreams_stores_0_data_bits_wdata_8(accel_io_memStreams_stores_0_data_bits_wdata_8),
    .io_memStreams_stores_0_data_bits_wdata_9(accel_io_memStreams_stores_0_data_bits_wdata_9),
    .io_memStreams_stores_0_data_bits_wdata_10(accel_io_memStreams_stores_0_data_bits_wdata_10),
    .io_memStreams_stores_0_data_bits_wdata_11(accel_io_memStreams_stores_0_data_bits_wdata_11),
    .io_memStreams_stores_0_data_bits_wdata_12(accel_io_memStreams_stores_0_data_bits_wdata_12),
    .io_memStreams_stores_0_data_bits_wdata_13(accel_io_memStreams_stores_0_data_bits_wdata_13),
    .io_memStreams_stores_0_data_bits_wdata_14(accel_io_memStreams_stores_0_data_bits_wdata_14),
    .io_memStreams_stores_0_data_bits_wdata_15(accel_io_memStreams_stores_0_data_bits_wdata_15),
    .io_memStreams_stores_0_data_bits_wstrb(accel_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(accel_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(accel_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(accel_io_memStreams_stores_0_wresp_bits),
    .io_memStreams_gathers_0_cmd_ready(accel_io_memStreams_gathers_0_cmd_ready),
    .io_memStreams_gathers_0_cmd_valid(accel_io_memStreams_gathers_0_cmd_valid),
    .io_memStreams_gathers_0_cmd_bits_addr_0(accel_io_memStreams_gathers_0_cmd_bits_addr_0),
    .io_memStreams_gathers_0_cmd_bits_addr_1(accel_io_memStreams_gathers_0_cmd_bits_addr_1),
    .io_memStreams_gathers_0_cmd_bits_addr_2(accel_io_memStreams_gathers_0_cmd_bits_addr_2),
    .io_memStreams_gathers_0_cmd_bits_addr_3(accel_io_memStreams_gathers_0_cmd_bits_addr_3),
    .io_memStreams_gathers_0_cmd_bits_addr_4(accel_io_memStreams_gathers_0_cmd_bits_addr_4),
    .io_memStreams_gathers_0_cmd_bits_addr_5(accel_io_memStreams_gathers_0_cmd_bits_addr_5),
    .io_memStreams_gathers_0_cmd_bits_addr_6(accel_io_memStreams_gathers_0_cmd_bits_addr_6),
    .io_memStreams_gathers_0_cmd_bits_addr_7(accel_io_memStreams_gathers_0_cmd_bits_addr_7),
    .io_memStreams_gathers_0_cmd_bits_addr_8(accel_io_memStreams_gathers_0_cmd_bits_addr_8),
    .io_memStreams_gathers_0_cmd_bits_addr_9(accel_io_memStreams_gathers_0_cmd_bits_addr_9),
    .io_memStreams_gathers_0_cmd_bits_addr_10(accel_io_memStreams_gathers_0_cmd_bits_addr_10),
    .io_memStreams_gathers_0_cmd_bits_addr_11(accel_io_memStreams_gathers_0_cmd_bits_addr_11),
    .io_memStreams_gathers_0_cmd_bits_addr_12(accel_io_memStreams_gathers_0_cmd_bits_addr_12),
    .io_memStreams_gathers_0_cmd_bits_addr_13(accel_io_memStreams_gathers_0_cmd_bits_addr_13),
    .io_memStreams_gathers_0_cmd_bits_addr_14(accel_io_memStreams_gathers_0_cmd_bits_addr_14),
    .io_memStreams_gathers_0_cmd_bits_addr_15(accel_io_memStreams_gathers_0_cmd_bits_addr_15),
    .io_memStreams_gathers_0_data_ready(accel_io_memStreams_gathers_0_data_ready),
    .io_memStreams_gathers_0_data_valid(accel_io_memStreams_gathers_0_data_valid),
    .io_memStreams_gathers_0_data_bits_0(accel_io_memStreams_gathers_0_data_bits_0),
    .io_memStreams_gathers_0_data_bits_1(accel_io_memStreams_gathers_0_data_bits_1),
    .io_memStreams_gathers_0_data_bits_2(accel_io_memStreams_gathers_0_data_bits_2),
    .io_memStreams_gathers_0_data_bits_3(accel_io_memStreams_gathers_0_data_bits_3),
    .io_memStreams_gathers_0_data_bits_4(accel_io_memStreams_gathers_0_data_bits_4),
    .io_memStreams_gathers_0_data_bits_5(accel_io_memStreams_gathers_0_data_bits_5),
    .io_memStreams_gathers_0_data_bits_6(accel_io_memStreams_gathers_0_data_bits_6),
    .io_memStreams_gathers_0_data_bits_7(accel_io_memStreams_gathers_0_data_bits_7),
    .io_memStreams_gathers_0_data_bits_8(accel_io_memStreams_gathers_0_data_bits_8),
    .io_memStreams_gathers_0_data_bits_9(accel_io_memStreams_gathers_0_data_bits_9),
    .io_memStreams_gathers_0_data_bits_10(accel_io_memStreams_gathers_0_data_bits_10),
    .io_memStreams_gathers_0_data_bits_11(accel_io_memStreams_gathers_0_data_bits_11),
    .io_memStreams_gathers_0_data_bits_12(accel_io_memStreams_gathers_0_data_bits_12),
    .io_memStreams_gathers_0_data_bits_13(accel_io_memStreams_gathers_0_data_bits_13),
    .io_memStreams_gathers_0_data_bits_14(accel_io_memStreams_gathers_0_data_bits_14),
    .io_memStreams_gathers_0_data_bits_15(accel_io_memStreams_gathers_0_data_bits_15),
    .io_memStreams_scatters_0_cmd_ready(accel_io_memStreams_scatters_0_cmd_ready),
    .io_memStreams_scatters_0_cmd_valid(accel_io_memStreams_scatters_0_cmd_valid),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_0(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_1(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_2(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_3(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_4(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_5(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_6(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_7(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_8(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_9(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_10(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_11(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_12(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_13(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_14(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_15(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15),
    .io_memStreams_scatters_0_cmd_bits_wdata_0(accel_io_memStreams_scatters_0_cmd_bits_wdata_0),
    .io_memStreams_scatters_0_cmd_bits_wdata_1(accel_io_memStreams_scatters_0_cmd_bits_wdata_1),
    .io_memStreams_scatters_0_cmd_bits_wdata_2(accel_io_memStreams_scatters_0_cmd_bits_wdata_2),
    .io_memStreams_scatters_0_cmd_bits_wdata_3(accel_io_memStreams_scatters_0_cmd_bits_wdata_3),
    .io_memStreams_scatters_0_cmd_bits_wdata_4(accel_io_memStreams_scatters_0_cmd_bits_wdata_4),
    .io_memStreams_scatters_0_cmd_bits_wdata_5(accel_io_memStreams_scatters_0_cmd_bits_wdata_5),
    .io_memStreams_scatters_0_cmd_bits_wdata_6(accel_io_memStreams_scatters_0_cmd_bits_wdata_6),
    .io_memStreams_scatters_0_cmd_bits_wdata_7(accel_io_memStreams_scatters_0_cmd_bits_wdata_7),
    .io_memStreams_scatters_0_cmd_bits_wdata_8(accel_io_memStreams_scatters_0_cmd_bits_wdata_8),
    .io_memStreams_scatters_0_cmd_bits_wdata_9(accel_io_memStreams_scatters_0_cmd_bits_wdata_9),
    .io_memStreams_scatters_0_cmd_bits_wdata_10(accel_io_memStreams_scatters_0_cmd_bits_wdata_10),
    .io_memStreams_scatters_0_cmd_bits_wdata_11(accel_io_memStreams_scatters_0_cmd_bits_wdata_11),
    .io_memStreams_scatters_0_cmd_bits_wdata_12(accel_io_memStreams_scatters_0_cmd_bits_wdata_12),
    .io_memStreams_scatters_0_cmd_bits_wdata_13(accel_io_memStreams_scatters_0_cmd_bits_wdata_13),
    .io_memStreams_scatters_0_cmd_bits_wdata_14(accel_io_memStreams_scatters_0_cmd_bits_wdata_14),
    .io_memStreams_scatters_0_cmd_bits_wdata_15(accel_io_memStreams_scatters_0_cmd_bits_wdata_15),
    .io_memStreams_scatters_0_wresp_ready(accel_io_memStreams_scatters_0_wresp_ready),
    .io_memStreams_scatters_0_wresp_valid(accel_io_memStreams_scatters_0_wresp_valid),
    .io_memStreams_scatters_0_wresp_bits(accel_io_memStreams_scatters_0_wresp_bits),
    .io_axiStreamsIn_0_TVALID(accel_io_axiStreamsIn_0_TVALID),
    .io_axiStreamsIn_0_TREADY(accel_io_axiStreamsIn_0_TREADY),
    .io_axiStreamsIn_0_TDATA(accel_io_axiStreamsIn_0_TDATA),
    .io_axiStreamsIn_0_TSTRB(accel_io_axiStreamsIn_0_TSTRB),
    .io_axiStreamsIn_0_TKEEP(accel_io_axiStreamsIn_0_TKEEP),
    .io_axiStreamsIn_0_TLAST(accel_io_axiStreamsIn_0_TLAST),
    .io_axiStreamsIn_0_TID(accel_io_axiStreamsIn_0_TID),
    .io_axiStreamsIn_0_TDEST(accel_io_axiStreamsIn_0_TDEST),
    .io_axiStreamsIn_0_TUSER(accel_io_axiStreamsIn_0_TUSER),
    .io_axiStreamsOut_0_TVALID(accel_io_axiStreamsOut_0_TVALID),
    .io_axiStreamsOut_0_TREADY(accel_io_axiStreamsOut_0_TREADY),
    .io_axiStreamsOut_0_TDATA(accel_io_axiStreamsOut_0_TDATA),
    .io_axiStreamsOut_0_TSTRB(accel_io_axiStreamsOut_0_TSTRB),
    .io_axiStreamsOut_0_TKEEP(accel_io_axiStreamsOut_0_TKEEP),
    .io_axiStreamsOut_0_TLAST(accel_io_axiStreamsOut_0_TLAST),
    .io_axiStreamsOut_0_TID(accel_io_axiStreamsOut_0_TID),
    .io_axiStreamsOut_0_TDEST(accel_io_axiStreamsOut_0_TDEST),
    .io_axiStreamsOut_0_TUSER(accel_io_axiStreamsOut_0_TUSER),
    .io_heap_0_req_valid(accel_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(accel_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(accel_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(accel_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(accel_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(accel_io_heap_0_resp_bits_sizeAddr),
    .io_argIns_0(accel_io_argIns_0),
    .io_argIns_1(accel_io_argIns_1),
    .io_argOuts_0_port_ready(accel_io_argOuts_0_port_ready),
    .io_argOuts_0_port_valid(accel_io_argOuts_0_port_valid),
    .io_argOuts_0_port_bits(accel_io_argOuts_0_port_bits),
    .io_argOuts_0_echo(accel_io_argOuts_0_echo)
  );
  assign io_rdata = 64'h0;
  assign accel_clock = clock; // @[:@23028.4]
  assign accel_reset = reset; // @[:@23029.4]
  assign accel_io_enable = 1'h0;
  assign accel_io_reset = 1'h0;
  assign accel_io_memStreams_loads_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_loads_0_data_valid = 1'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_0 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_1 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_2 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_3 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_4 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_5 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_6 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_7 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_8 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_9 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_10 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_11 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_12 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_13 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_14 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_15 = 32'h0;
  assign accel_io_memStreams_stores_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_stores_0_data_ready = 1'h0;
  assign accel_io_memStreams_stores_0_wresp_valid = 1'h0;
  assign accel_io_memStreams_stores_0_wresp_bits = 1'h0;
  assign accel_io_memStreams_gathers_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_gathers_0_data_valid = 1'h0;
  assign accel_io_memStreams_gathers_0_data_bits_0 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_1 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_2 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_3 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_4 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_5 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_6 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_7 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_8 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_9 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_10 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_11 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_12 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_13 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_14 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_15 = 32'h0;
  assign accel_io_memStreams_scatters_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_scatters_0_wresp_valid = 1'h0;
  assign accel_io_memStreams_scatters_0_wresp_bits = 1'h0;
  assign accel_io_axiStreamsIn_0_TVALID = 1'h0;
  assign accel_io_axiStreamsIn_0_TDATA = 256'h0;
  assign accel_io_axiStreamsIn_0_TSTRB = 32'h0;
  assign accel_io_axiStreamsIn_0_TKEEP = 32'h0;
  assign accel_io_axiStreamsIn_0_TLAST = 1'h0;
  assign accel_io_axiStreamsIn_0_TID = 8'h0;
  assign accel_io_axiStreamsIn_0_TDEST = 8'h0;
  assign accel_io_axiStreamsIn_0_TUSER = 32'h0;
  assign accel_io_axiStreamsOut_0_TREADY = 1'h0;
  assign accel_io_heap_0_resp_valid = 1'h0;
  assign accel_io_heap_0_resp_bits_allocDealloc = 1'h0;
  assign accel_io_heap_0_resp_bits_sizeAddr = 64'h0;
  assign accel_io_argIns_0 = 64'h0;
  assign accel_io_argIns_1 = 64'h0;
  assign accel_io_argOuts_0_port_ready = 1'h0;
  assign accel_io_argOuts_0_echo = 64'h0;
endmodule
