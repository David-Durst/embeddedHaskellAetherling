// Latency = 4
module top(
  input CLK/*verilator public*/, 
  input [7:0] I_0_0_0/*verilator public*/, 
  output [7:0] O_0_0_0/*verilator public*/, 
  input [7:0] I_1_0_0/*verilator public*/, 
  output [7:0] O_1_0_0/*verilator public*/, 
  output valid_down/*verilator public*/, 
  input valid_up/*verilator public*/
);
  wire dontcare;
  wire [31:0] io_output_counts_1;
  wire [31:0] io_output_counts_0;

  x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1 sampler_box ( // @[m_x55_ctr_0.scala 26:17:@1721.4]
    .clock(CLK), // @[:@1296.4]
    .reset('b0), // @[:@1297.4]
    .io_in_x270_TREADY(dontcare), // @[:@1298.4]
    .io_in_x270_TDATA({I_0_0_0,I_1_0_0}), // @[:@1298.4]
    .io_in_x270_TID(8'h0),
    .io_in_x270_TDEST(8'h0),
    .io_in_x271_TVALID(valid_down), // @[:@1298.4]
    .io_in_x271_TDATA({O_0_0_0,O_1_0_0}), // @[:@1298.4]
    .io_in_x271_TREADY(1'b1), // @[:@1298.4]
    .io_sigsIn_datapathEn(valid_up), // @[:@1298.4]
    .io_sigsIn_backpressure(1'b1), // @[:@20563.4]
    .io_sigsIn_break(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_1(io_output_counts_1), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_0(io_output_counts_0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_0(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_1(1'b0), // @[:@20563.4]
    .io_rr('b1) // @[:@1298.4]
  );

  wire dontcare2;

  wire io_output_oobs_0;
  wire io_output_oobs_1;
  x278_ctrchain cchain ( // @[:@2879.2]
    .clock(CLK), // @[:@2880.4]
    .reset(1'b0), // @[:@2881.4]
    .io_input_reset(1'b0), // @[:@2882.4]
    .io_input_enable(valid_up), // @[:@2882.4]
    .io_output_counts_1(io_output_counts_1), // @[:@2882.4]
    .io_output_counts_0(io_output_counts_0), // @[:@2882.4]
    .io_output_oobs_0(io_output_oobs_0), // @[:@2882.4]
    .io_output_oobs_1(io_output_oobs_1), // @[:@2882.4]
    .io_output_done(dontcare2) // @[:@2882.4]
  );

endmodule

module RetimeShiftRegister
#(
    parameter WIDTH = 1,
    parameter STAGES = 1)
(
    input clock,
    input reset,
    input flow,
    input [WIDTH-1:0] init,
    input [WIDTH-1:0] in,
    output reg [WIDTH-1:0] out
);
  integer i;
  reg [WIDTH-1:0] sr[STAGES:0]; // Create 'STAGES' number of register, each 'WIDTH' bits wide

   /* synopsys dc_tcl_script_begin
    set_ungroup [current_design] true
    set_flatten true -effort high -phase true -design [current_design]
    set_dont_retime [current_design] false
    set_optimize_registers true -design [current_design]
    */
  always @(posedge clock) begin
    if (reset) begin
      for(i=0; i<STAGES; i=i+1) begin
        sr[i] <= init;
      end
    end else begin
      if (flow) begin 
        sr[0] <= in;
        for(i=1; i<STAGES; i=i+1) begin
          sr[i] <= sr[i-1];
        end
      end
    end
  end

  always @(*) begin
    out = sr[STAGES-1];
  end
endmodule
module FF( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  output [31:0] io_rPort_0_output_0, // @[:@6.4]
  input  [31:0] io_wPort_0_data_0, // @[:@6.4]
  input         io_wPort_0_reset, // @[:@6.4]
  input         io_wPort_0_en_0 // @[:@6.4]
);
  reg [31:0] ff; // @[MemPrimitives.scala 173:19:@21.4]
  reg [31:0] _RAND_0;
  wire [31:0] _T_68; // @[MemPrimitives.scala 177:32:@23.4]
  wire [31:0] _T_69; // @[MemPrimitives.scala 177:12:@24.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 177:32:@23.4]
  assign _T_69 = io_wPort_0_reset ? 32'h0 : _T_68; // @[MemPrimitives.scala 177:12:@24.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 178:34:@26.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 32'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 32'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SRFF( // @[:@28.2]
  input   clock, // @[:@29.4]
  input   reset, // @[:@30.4]
  input   io_input_set, // @[:@31.4]
  input   io_input_reset, // @[:@31.4]
  input   io_input_asyn_reset, // @[:@31.4]
  output  io_output // @[:@31.4]
);
  reg  _T_15; // @[SRFF.scala 20:21:@33.4]
  reg [31:0] _RAND_0;
  wire  _T_19; // @[SRFF.scala 21:74:@34.4]
  wire  _T_20; // @[SRFF.scala 21:48:@35.4]
  wire  _T_21; // @[SRFF.scala 21:14:@36.4]
  assign _T_19 = io_input_reset ? 1'h0 : _T_15; // @[SRFF.scala 21:74:@34.4]
  assign _T_20 = io_input_set ? 1'h1 : _T_19; // @[SRFF.scala 21:48:@35.4]
  assign _T_21 = io_input_asyn_reset ? 1'h0 : _T_20; // @[SRFF.scala 21:14:@36.4]
  assign io_output = io_input_asyn_reset ? 1'h0 : _T_15; // @[SRFF.scala 22:15:@39.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_15 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_15 <= 1'h0;
    end else begin
      if (io_input_asyn_reset) begin
        _T_15 <= 1'h0;
      end else begin
        if (io_input_set) begin
          _T_15 <= 1'h1;
        end else begin
          if (io_input_reset) begin
            _T_15 <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module SingleCounter( // @[:@41.2]
  input   clock, // @[:@42.4]
  input   reset, // @[:@43.4]
  input   io_input_reset, // @[:@44.4]
  output  io_output_done // @[:@44.4]
);
  wire  bases_0_clock; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_reset; // @[Counter.scala 253:53:@57.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 253:53:@57.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 253:53:@57.4]
  wire  SRFF_clock; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_set; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_output; // @[Counter.scala 255:22:@73.4]
  wire [31:0] _T_48; // @[Counter.scala 279:52:@101.4]
  wire [32:0] _T_50; // @[Counter.scala 283:33:@102.4]
  wire [31:0] _T_51; // @[Counter.scala 283:33:@103.4]
  wire [31:0] _T_52; // @[Counter.scala 283:33:@104.4]
  wire  _T_57; // @[Counter.scala 285:18:@106.4]
  wire [31:0] _T_68; // @[Counter.scala 291:115:@114.4]
  wire [31:0] _T_71; // @[Counter.scala 291:152:@117.4]
  wire [31:0] _T_72; // @[Counter.scala 291:74:@118.4]
  FF bases_0 ( // @[Counter.scala 253:53:@57.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 255:22:@73.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 279:52:@101.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@102.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@103.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 283:33:@104.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh13); // @[Counter.scala 285:18:@106.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 291:115:@114.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 291:152:@117.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 291:74:@118.4]
  assign io_output_done = $signed(_T_52) >= $signed(32'sh13); // @[Counter.scala 325:20:@127.4]
  assign bases_0_clock = clock; // @[:@58.4]
  assign bases_0_reset = reset; // @[:@59.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 291:31:@120.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 273:27:@99.4]
  assign bases_0_io_wPort_0_en_0 = 1'h1; // @[Counter.scala 276:29:@100.4]
  assign SRFF_clock = clock; // @[:@74.4]
  assign SRFF_reset = reset; // @[:@75.4]
  assign SRFF_io_input_set = io_input_reset == 1'h0; // @[Counter.scala 256:23:@78.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 257:25:@80.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 258:30:@81.4]
endmodule
module RetimeWrapper( // @[:@144.2]
  input   clock, // @[:@145.4]
  input   reset, // @[:@146.4]
  input   io_flow, // @[:@147.4]
  input   io_in, // @[:@147.4]
  output  io_out // @[:@147.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@149.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@149.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@162.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@161.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@160.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@159.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@158.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@156.4]
endmodule
module RootController_sm( // @[:@312.2]
  input   clock, // @[:@313.4]
  input   reset, // @[:@314.4]
  input   io_enable, // @[:@315.4]
  output  io_done, // @[:@315.4]
  input   io_rst, // @[:@315.4]
  input   io_ctrDone, // @[:@315.4]
  output  io_ctrInc, // @[:@315.4]
  input   io_doneIn_0, // @[:@315.4]
  output  io_enableOut_0, // @[:@315.4]
  output  io_childAck_0 // @[:@315.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@318.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@321.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@338.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@433.4]
  wire  finished; // @[Controllers.scala 81:26:@324.4]
  wire  synchronize; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  wire  _T_122; // @[Controllers.scala 128:33:@371.4]
  wire  _T_124; // @[Controllers.scala 128:54:@372.4]
  wire  _T_125; // @[Controllers.scala 128:52:@373.4]
  wire  _T_126; // @[Controllers.scala 128:66:@374.4]
  wire  _T_128; // @[Controllers.scala 128:98:@376.4]
  wire  _T_129; // @[Controllers.scala 128:96:@377.4]
  wire  _T_131; // @[Controllers.scala 128:123:@378.4]
  wire  _T_133; // @[Controllers.scala 129:48:@381.4]
  wire  _T_138; // @[Controllers.scala 130:52:@386.4]
  wire  _T_139; // @[Controllers.scala 130:50:@387.4]
  wire  _T_147; // @[Controllers.scala 130:129:@393.4]
  wire  _T_150; // @[Controllers.scala 131:45:@396.4]
  wire  _T_154; // @[Controllers.scala 213:68:@402.4]
  wire  _T_156; // @[Controllers.scala 213:90:@404.4]
  wire  _T_158; // @[Controllers.scala 213:132:@406.4]
  wire  _T_159; // @[Controllers.scala 213:130:@407.4]
  wire  _T_160; // @[Controllers.scala 213:156:@408.4]
  reg  _T_166; // @[package.scala 48:56:@412.4]
  reg [31:0] _RAND_0;
  reg  _T_180; // @[package.scala 48:56:@430.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@318.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@321.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@338.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@357.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@416.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@433.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  assign finished = done_0_io_output | io_done; // @[Controllers.scala 81:26:@324.4]
  assign synchronize = RetimeWrapper_io_out; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  assign _T_122 = done_0_io_output == 1'h0; // @[Controllers.scala 128:33:@371.4]
  assign _T_124 = io_ctrDone == 1'h0; // @[Controllers.scala 128:54:@372.4]
  assign _T_125 = _T_122 & _T_124; // @[Controllers.scala 128:52:@373.4]
  assign _T_126 = _T_125 & io_enable; // @[Controllers.scala 128:66:@374.4]
  assign _T_128 = ~ iterDone_0_io_output; // @[Controllers.scala 128:98:@376.4]
  assign _T_129 = _T_126 & _T_128; // @[Controllers.scala 128:96:@377.4]
  assign _T_131 = io_doneIn_0 == 1'h0; // @[Controllers.scala 128:123:@378.4]
  assign _T_133 = io_doneIn_0 | io_rst; // @[Controllers.scala 129:48:@381.4]
  assign _T_138 = synchronize == 1'h0; // @[Controllers.scala 130:52:@386.4]
  assign _T_139 = io_doneIn_0 & _T_138; // @[Controllers.scala 130:50:@387.4]
  assign _T_147 = finished == 1'h0; // @[Controllers.scala 130:129:@393.4]
  assign _T_150 = io_rst == 1'h0; // @[Controllers.scala 131:45:@396.4]
  assign _T_154 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@402.4]
  assign _T_156 = _T_154 & _T_128; // @[Controllers.scala 213:90:@404.4]
  assign _T_158 = ~ done_0_io_output; // @[Controllers.scala 213:132:@406.4]
  assign _T_159 = _T_156 & _T_158; // @[Controllers.scala 213:130:@407.4]
  assign _T_160 = ~ io_ctrDone; // @[Controllers.scala 213:156:@408.4]
  assign io_done = RetimeWrapper_2_io_out; // @[Controllers.scala 245:13:@440.4]
  assign io_ctrInc = io_doneIn_0; // @[Controllers.scala 122:17:@356.4]
  assign io_enableOut_0 = _T_159 & _T_160; // @[Controllers.scala 213:55:@410.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@401.4]
  assign active_0_clock = clock; // @[:@319.4]
  assign active_0_reset = reset; // @[:@320.4]
  assign active_0_io_input_set = _T_129 & _T_131; // @[Controllers.scala 128:30:@380.4]
  assign active_0_io_input_reset = _T_133 | done_0_io_output; // @[Controllers.scala 129:32:@385.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@326.4]
  assign done_0_clock = clock; // @[:@322.4]
  assign done_0_reset = reset; // @[:@323.4]
  assign done_0_io_input_set = io_ctrDone & _T_150; // @[Controllers.scala 131:28:@399.4]
  assign done_0_io_input_reset = io_rst | done_0_io_output; // @[Controllers.scala 86:33:@336.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@327.4]
  assign iterDone_0_clock = clock; // @[:@339.4]
  assign iterDone_0_reset = reset; // @[:@340.4]
  assign iterDone_0_io_input_set = _T_139 & _T_147; // @[Controllers.scala 130:32:@395.4]
  assign iterDone_0_io_input_reset = synchronize | io_rst; // @[Controllers.scala 92:37:@350.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@341.4]
  assign RetimeWrapper_clock = clock; // @[:@358.4]
  assign RetimeWrapper_reset = reset; // @[:@359.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@361.4]
  assign RetimeWrapper_io_in = io_doneIn_0; // @[package.scala 94:16:@360.4]
  assign RetimeWrapper_1_clock = clock; // @[:@417.4]
  assign RetimeWrapper_1_reset = reset; // @[:@418.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@420.4]
  assign RetimeWrapper_1_io_in = done_0_io_output & _T_166; // @[package.scala 94:16:@419.4]
  assign RetimeWrapper_2_clock = clock; // @[:@434.4]
  assign RetimeWrapper_2_reset = reset; // @[:@435.4]
  assign RetimeWrapper_2_io_flow = io_enable; // @[package.scala 95:18:@437.4]
  assign RetimeWrapper_2_io_in = done_0_io_output & _T_180; // @[package.scala 94:16:@436.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_166 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_180 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_166 <= 1'h0;
    end else begin
      _T_166 <= _T_122;
    end
    if (reset) begin
      _T_180 <= 1'h0;
    end else begin
      _T_180 <= _T_122;
    end
  end
endmodule
module x473_outr_UnitPipe_sm( // @[:@2389.2]
  input   clock, // @[:@2390.4]
  input   reset, // @[:@2391.4]
  input   io_enable, // @[:@2392.4]
  output  io_done, // @[:@2392.4]
  input   io_parentAck, // @[:@2392.4]
  input   io_doneIn_0, // @[:@2392.4]
  output  io_enableOut_0, // @[:@2392.4]
  output  io_childAck_0, // @[:@2392.4]
  input   io_ctrCopyDone_0 // @[:@2392.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@2395.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@2395.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@2395.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@2395.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@2395.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@2395.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@2398.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@2398.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@2398.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@2398.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@2398.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@2398.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@2415.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@2415.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@2415.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@2415.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@2415.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@2415.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@2446.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@2446.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@2446.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@2446.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@2446.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@2460.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@2460.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@2460.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@2460.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@2460.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@2478.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@2478.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@2478.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@2478.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@2478.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@2515.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@2515.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@2515.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@2515.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@2515.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@2532.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@2532.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@2532.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@2532.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@2532.4]
  wire  _T_105; // @[Controllers.scala 165:35:@2430.4]
  wire  _T_107; // @[Controllers.scala 165:60:@2431.4]
  wire  _T_108; // @[Controllers.scala 165:58:@2432.4]
  wire  _T_110; // @[Controllers.scala 165:76:@2433.4]
  wire  _T_111; // @[Controllers.scala 165:74:@2434.4]
  wire  _T_115; // @[Controllers.scala 165:109:@2437.4]
  wire  _T_118; // @[Controllers.scala 165:141:@2439.4]
  wire  _T_126; // @[package.scala 96:25:@2451.4 package.scala 96:25:@2452.4]
  wire  _T_130; // @[Controllers.scala 167:54:@2454.4]
  wire  _T_131; // @[Controllers.scala 167:52:@2455.4]
  wire  _T_138; // @[package.scala 96:25:@2465.4 package.scala 96:25:@2466.4]
  wire  _T_156; // @[package.scala 96:25:@2483.4 package.scala 96:25:@2484.4]
  wire  _T_160; // @[Controllers.scala 169:67:@2486.4]
  wire  _T_161; // @[Controllers.scala 169:86:@2487.4]
  wire  _T_174; // @[Controllers.scala 213:68:@2501.4]
  wire  _T_176; // @[Controllers.scala 213:90:@2503.4]
  wire  _T_178; // @[Controllers.scala 213:132:@2505.4]
  reg  _T_186; // @[package.scala 48:56:@2511.4]
  reg [31:0] _RAND_0;
  wire  _T_187; // @[package.scala 100:41:@2513.4]
  reg  _T_200; // @[package.scala 48:56:@2529.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@2395.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@2398.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@2415.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@2446.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@2460.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@2478.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@2515.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@2532.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_105 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@2430.4]
  assign _T_107 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@2431.4]
  assign _T_108 = _T_105 & _T_107; // @[Controllers.scala 165:58:@2432.4]
  assign _T_110 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@2433.4]
  assign _T_111 = _T_108 & _T_110; // @[Controllers.scala 165:74:@2434.4]
  assign _T_115 = _T_111 & io_enable; // @[Controllers.scala 165:109:@2437.4]
  assign _T_118 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@2439.4]
  assign _T_126 = RetimeWrapper_io_out; // @[package.scala 96:25:@2451.4 package.scala 96:25:@2452.4]
  assign _T_130 = _T_126 == 1'h0; // @[Controllers.scala 167:54:@2454.4]
  assign _T_131 = io_doneIn_0 | _T_130; // @[Controllers.scala 167:52:@2455.4]
  assign _T_138 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@2465.4 package.scala 96:25:@2466.4]
  assign _T_156 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@2483.4 package.scala 96:25:@2484.4]
  assign _T_160 = _T_156 == 1'h0; // @[Controllers.scala 169:67:@2486.4]
  assign _T_161 = _T_160 & io_enable; // @[Controllers.scala 169:86:@2487.4]
  assign _T_174 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@2501.4]
  assign _T_176 = _T_174 & _T_105; // @[Controllers.scala 213:90:@2503.4]
  assign _T_178 = ~ done_0_io_output; // @[Controllers.scala 213:132:@2505.4]
  assign _T_187 = done_0_io_output & _T_186; // @[package.scala 100:41:@2513.4]
  assign io_done = RetimeWrapper_4_io_out; // @[Controllers.scala 245:13:@2539.4]
  assign io_enableOut_0 = _T_176 & _T_178; // @[Controllers.scala 213:55:@2509.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@2500.4]
  assign active_0_clock = clock; // @[:@2396.4]
  assign active_0_reset = reset; // @[:@2397.4]
  assign active_0_io_input_set = _T_115 & _T_118; // @[Controllers.scala 165:32:@2441.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@2445.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@2403.4]
  assign done_0_clock = clock; // @[:@2399.4]
  assign done_0_reset = reset; // @[:@2400.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_161; // @[Controllers.scala 169:30:@2491.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@2413.4 Controllers.scala 170:32:@2498.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@2404.4]
  assign iterDone_0_clock = clock; // @[:@2416.4]
  assign iterDone_0_reset = reset; // @[:@2417.4]
  assign iterDone_0_io_input_set = _T_131 & io_enable; // @[Controllers.scala 167:34:@2459.4]
  assign iterDone_0_io_input_reset = _T_138 | io_parentAck; // @[Controllers.scala 92:37:@2427.4 Controllers.scala 168:36:@2475.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@2418.4]
  assign RetimeWrapper_clock = clock; // @[:@2447.4]
  assign RetimeWrapper_reset = reset; // @[:@2448.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@2450.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@2449.4]
  assign RetimeWrapper_1_clock = clock; // @[:@2461.4]
  assign RetimeWrapper_1_reset = reset; // @[:@2462.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@2464.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@2463.4]
  assign RetimeWrapper_2_clock = clock; // @[:@2479.4]
  assign RetimeWrapper_2_reset = reset; // @[:@2480.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@2482.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@2481.4]
  assign RetimeWrapper_3_clock = clock; // @[:@2516.4]
  assign RetimeWrapper_3_reset = reset; // @[:@2517.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@2519.4]
  assign RetimeWrapper_3_io_in = _T_187 | io_parentAck; // @[package.scala 94:16:@2518.4]
  assign RetimeWrapper_4_clock = clock; // @[:@2533.4]
  assign RetimeWrapper_4_reset = reset; // @[:@2534.4]
  assign RetimeWrapper_4_io_flow = io_enable; // @[package.scala 95:18:@2536.4]
  assign RetimeWrapper_4_io_in = done_0_io_output & _T_200; // @[package.scala 94:16:@2535.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_186 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_200 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_186 <= 1'h0;
    end else begin
      _T_186 <= _T_110;
    end
    if (reset) begin
      _T_200 <= 1'h0;
    end else begin
      _T_200 <= _T_110;
    end
  end
endmodule
module SingleCounter_1( // @[:@2659.2]
  input         clock, // @[:@2660.4]
  input         reset, // @[:@2661.4]
  input         io_input_reset, // @[:@2662.4]
  input         io_input_enable, // @[:@2662.4]
  output [31:0] io_output_count_0, // @[:@2662.4]
  output        io_output_oobs_0, // @[:@2662.4]
  output        io_output_done, // @[:@2662.4]
  output        io_output_saturated // @[:@2662.4]
);
  wire  bases_0_clock; // @[Counter.scala 253:53:@2675.4]
  wire  bases_0_reset; // @[Counter.scala 253:53:@2675.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 253:53:@2675.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 253:53:@2675.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 253:53:@2675.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 253:53:@2675.4]
  wire  SRFF_clock; // @[Counter.scala 255:22:@2691.4]
  wire  SRFF_reset; // @[Counter.scala 255:22:@2691.4]
  wire  SRFF_io_input_set; // @[Counter.scala 255:22:@2691.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 255:22:@2691.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 255:22:@2691.4]
  wire  SRFF_io_output; // @[Counter.scala 255:22:@2691.4]
  wire  _T_36; // @[Counter.scala 256:45:@2694.4]
  wire [31:0] _T_48; // @[Counter.scala 279:52:@2719.4]
  wire [32:0] _T_50; // @[Counter.scala 283:33:@2720.4]
  wire [31:0] _T_51; // @[Counter.scala 283:33:@2721.4]
  wire [31:0] _T_52; // @[Counter.scala 283:33:@2722.4]
  wire  _T_57; // @[Counter.scala 285:18:@2724.4]
  wire [31:0] _T_68; // @[Counter.scala 291:115:@2732.4]
  wire [31:0] _T_71; // @[Counter.scala 291:152:@2735.4]
  wire [31:0] _T_72; // @[Counter.scala 291:74:@2736.4]
  wire  _T_75; // @[Counter.scala 314:102:@2740.4]
  wire  _T_77; // @[Counter.scala 314:130:@2741.4]
  FF bases_0 ( // @[Counter.scala 253:53:@2675.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 255:22:@2691.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 256:45:@2694.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 279:52:@2719.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@2720.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@2721.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 283:33:@2722.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh4); // @[Counter.scala 285:18:@2724.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 291:115:@2732.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 291:152:@2735.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 291:74:@2736.4]
  assign _T_75 = $signed(_T_48) < $signed(32'sh0); // @[Counter.scala 314:102:@2740.4]
  assign _T_77 = $signed(_T_48) >= $signed(32'sh4); // @[Counter.scala 314:130:@2741.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 296:28:@2739.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 314:60:@2743.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 325:20:@2745.4]
  assign io_output_saturated = $signed(_T_52) >= $signed(32'sh4); // @[Counter.scala 332:25:@2748.4]
  assign bases_0_clock = clock; // @[:@2676.4]
  assign bases_0_reset = reset; // @[:@2677.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 291:31:@2738.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 273:27:@2717.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 276:29:@2718.4]
  assign SRFF_clock = clock; // @[:@2692.4]
  assign SRFF_reset = reset; // @[:@2693.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 256:23:@2696.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 257:25:@2698.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 258:30:@2699.4]
endmodule
module SingleCounter_2( // @[:@2788.2]
  input         clock, // @[:@2789.4]
  input         reset, // @[:@2790.4]
  input         io_setup_saturate, // @[:@2791.4]
  input         io_input_reset, // @[:@2791.4]
  input         io_input_enable, // @[:@2791.4]
  output [31:0] io_output_count_0, // @[:@2791.4]
  output        io_output_oobs_0, // @[:@2791.4]
  output        io_output_done // @[:@2791.4]
);
  wire  bases_0_clock; // @[Counter.scala 253:53:@2804.4]
  wire  bases_0_reset; // @[Counter.scala 253:53:@2804.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 253:53:@2804.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 253:53:@2804.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 253:53:@2804.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 253:53:@2804.4]
  wire  SRFF_clock; // @[Counter.scala 255:22:@2820.4]
  wire  SRFF_reset; // @[Counter.scala 255:22:@2820.4]
  wire  SRFF_io_input_set; // @[Counter.scala 255:22:@2820.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 255:22:@2820.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 255:22:@2820.4]
  wire  SRFF_io_output; // @[Counter.scala 255:22:@2820.4]
  wire  _T_36; // @[Counter.scala 256:45:@2823.4]
  wire [31:0] _T_48; // @[Counter.scala 279:52:@2848.4]
  wire [32:0] _T_50; // @[Counter.scala 283:33:@2849.4]
  wire [31:0] _T_51; // @[Counter.scala 283:33:@2850.4]
  wire [31:0] _T_52; // @[Counter.scala 283:33:@2851.4]
  wire  _T_57; // @[Counter.scala 285:18:@2853.4]
  wire [31:0] _T_68; // @[Counter.scala 291:115:@2861.4]
  wire [31:0] _T_70; // @[Counter.scala 291:85:@2863.4]
  wire [31:0] _T_71; // @[Counter.scala 291:152:@2864.4]
  wire [31:0] _T_72; // @[Counter.scala 291:74:@2865.4]
  wire  _T_75; // @[Counter.scala 314:102:@2869.4]
  wire  _T_77; // @[Counter.scala 314:130:@2870.4]
  FF bases_0 ( // @[Counter.scala 253:53:@2804.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 255:22:@2820.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 256:45:@2823.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 279:52:@2848.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh2); // @[Counter.scala 283:33:@2849.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh2); // @[Counter.scala 283:33:@2850.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 283:33:@2851.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh4); // @[Counter.scala 285:18:@2853.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 291:115:@2861.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 32'h0; // @[Counter.scala 291:85:@2863.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 291:152:@2864.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 291:74:@2865.4]
  assign _T_75 = $signed(_T_48) < $signed(32'sh0); // @[Counter.scala 314:102:@2869.4]
  assign _T_77 = $signed(_T_48) >= $signed(32'sh4); // @[Counter.scala 314:130:@2870.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 296:28:@2868.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 314:60:@2872.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 325:20:@2874.4]
  assign bases_0_clock = clock; // @[:@2805.4]
  assign bases_0_reset = reset; // @[:@2806.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 291:31:@2867.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 273:27:@2846.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 276:29:@2847.4]
  assign SRFF_clock = clock; // @[:@2821.4]
  assign SRFF_reset = reset; // @[:@2822.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 256:23:@2825.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 257:25:@2827.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 258:30:@2828.4]
endmodule
module x278_ctrchain( // @[:@2879.2]
  input         clock, // @[:@2880.4]
  input         reset, // @[:@2881.4]
  input         io_input_reset, // @[:@2882.4]
  input         io_input_enable, // @[:@2882.4]
  output [31:0] io_output_counts_1, // @[:@2882.4]
  output [31:0] io_output_counts_0, // @[:@2882.4]
  output        io_output_oobs_0, // @[:@2882.4]
  output        io_output_oobs_1, // @[:@2882.4]
  output        io_output_done // @[:@2882.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_reset; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 505:46:@2884.4]
  wire [31:0] ctrs_0_io_output_count_0; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_io_output_saturated; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_1_clock; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_reset; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_io_setup_saturate; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_io_input_reset; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_io_input_enable; // @[Counter.scala 505:46:@2887.4]
  wire [31:0] ctrs_1_io_output_count_0; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_io_output_oobs_0; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_io_output_done; // @[Counter.scala 505:46:@2887.4]
  wire  isDone; // @[Counter.scala 533:51:@2904.4]
  reg  wasDone; // @[Counter.scala 534:24:@2905.4]
  reg [31:0] _RAND_0;
  wire  _T_64; // @[Counter.scala 538:69:@2913.4]
  wire  _T_66; // @[Counter.scala 538:80:@2914.4]
  reg  doneLatch; // @[Counter.scala 542:26:@2919.4]
  reg [31:0] _RAND_1;
  wire  _T_73; // @[Counter.scala 543:48:@2920.4]
  wire  _T_74; // @[Counter.scala 543:19:@2921.4]
  SingleCounter_1 ctrs_0 ( // @[Counter.scala 505:46:@2884.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done),
    .io_output_saturated(ctrs_0_io_output_saturated)
  );
  SingleCounter_2 ctrs_1 ( // @[Counter.scala 505:46:@2887.4]
    .clock(ctrs_1_clock),
    .reset(ctrs_1_reset),
    .io_setup_saturate(ctrs_1_io_setup_saturate),
    .io_input_reset(ctrs_1_io_input_reset),
    .io_input_enable(ctrs_1_io_input_enable),
    .io_output_count_0(ctrs_1_io_output_count_0),
    .io_output_oobs_0(ctrs_1_io_output_oobs_0),
    .io_output_done(ctrs_1_io_output_done)
  );
  assign isDone = ctrs_0_io_output_done & ctrs_1_io_output_done; // @[Counter.scala 533:51:@2904.4]
  assign _T_64 = io_input_enable & isDone; // @[Counter.scala 538:69:@2913.4]
  assign _T_66 = wasDone == 1'h0; // @[Counter.scala 538:80:@2914.4]
  assign _T_73 = isDone ? 1'h1 : doneLatch; // @[Counter.scala 543:48:@2920.4]
  assign _T_74 = io_input_reset ? 1'h0 : _T_73; // @[Counter.scala 543:19:@2921.4]
  assign io_output_counts_1 = ctrs_1_io_output_count_0; // @[Counter.scala 549:32:@2926.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 549:32:@2923.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 550:30:@2925.4]
  assign io_output_oobs_1 = ctrs_1_io_output_oobs_0 | doneLatch; // @[Counter.scala 550:30:@2928.4]
  assign io_output_done = _T_64 & _T_66; // @[Counter.scala 538:18:@2916.4]
  assign ctrs_0_clock = clock; // @[:@2885.4]
  assign ctrs_0_reset = reset; // @[:@2886.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 512:24:@2893.4]
  assign ctrs_0_io_input_enable = ctrs_1_io_output_done & io_input_enable; // @[Counter.scala 518:29:@2900.4]
  assign ctrs_1_clock = clock; // @[:@2888.4]
  assign ctrs_1_reset = reset; // @[:@2889.4]
  assign ctrs_1_io_setup_saturate = ctrs_0_io_output_saturated; // @[Counter.scala 524:31:@2903.4]
  assign ctrs_1_io_input_reset = io_input_reset; // @[Counter.scala 512:24:@2897.4]
  assign ctrs_1_io_input_enable = io_input_enable; // @[Counter.scala 516:33:@2898.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= isDone;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (isDone) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module RetimeWrapper_12( // @[:@2968.2]
  input   clock, // @[:@2969.4]
  input   reset, // @[:@2970.4]
  input   io_flow, // @[:@2971.4]
  input   io_in, // @[:@2971.4]
  output  io_out // @[:@2971.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(20)) sr ( // @[RetimeShiftRegister.scala 15:20:@2973.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@2986.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@2985.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@2984.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@2983.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@2982.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@2980.4]
endmodule
module RetimeWrapper_16( // @[:@3096.2]
  input   clock, // @[:@3097.4]
  input   reset, // @[:@3098.4]
  input   io_flow, // @[:@3099.4]
  input   io_in, // @[:@3099.4]
  output  io_out // @[:@3099.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(19)) sr ( // @[RetimeShiftRegister.scala 15:20:@3101.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3114.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3113.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3112.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3111.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3110.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3108.4]
endmodule
module x472_inr_Foreach_SAMPLER_BOX_sm( // @[:@3116.2]
  input   clock, // @[:@3117.4]
  input   reset, // @[:@3118.4]
  input   io_enable, // @[:@3119.4]
  output  io_done, // @[:@3119.4]
  output  io_doneLatch, // @[:@3119.4]
  input   io_ctrDone, // @[:@3119.4]
  output  io_datapathEn, // @[:@3119.4]
  output  io_ctrInc, // @[:@3119.4]
  output  io_ctrRst, // @[:@3119.4]
  input   io_parentAck, // @[:@3119.4]
  input   io_backpressure, // @[:@3119.4]
  input   io_break // @[:@3119.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@3121.4]
  wire  active_reset; // @[Controllers.scala 261:22:@3121.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@3121.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@3121.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@3121.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@3121.4]
  wire  done_clock; // @[Controllers.scala 262:20:@3124.4]
  wire  done_reset; // @[Controllers.scala 262:20:@3124.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@3124.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@3124.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@3124.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@3124.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3158.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3158.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3158.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@3158.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@3158.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@3180.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@3180.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@3180.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@3180.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@3180.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@3192.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@3192.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@3192.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@3192.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@3192.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@3200.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@3200.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@3200.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@3200.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@3200.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@3216.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@3216.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@3216.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@3216.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@3216.4]
  wire  _T_80; // @[Controllers.scala 264:48:@3129.4]
  wire  _T_81; // @[Controllers.scala 264:46:@3130.4]
  wire  _T_82; // @[Controllers.scala 264:62:@3131.4]
  wire  _T_83; // @[Controllers.scala 264:60:@3132.4]
  wire  _T_100; // @[package.scala 100:49:@3149.4]
  reg  _T_103; // @[package.scala 48:56:@3150.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@3163.4 package.scala 96:25:@3164.4]
  wire  _T_110; // @[package.scala 100:49:@3165.4]
  reg  _T_113; // @[package.scala 48:56:@3166.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@3168.4]
  wire  _T_118; // @[Controllers.scala 283:41:@3173.4]
  wire  _T_119; // @[Controllers.scala 283:59:@3174.4]
  wire  _T_121; // @[Controllers.scala 284:37:@3177.4]
  wire  _T_124; // @[package.scala 96:25:@3185.4 package.scala 96:25:@3186.4]
  wire  _T_126; // @[package.scala 100:49:@3187.4]
  reg  _T_129; // @[package.scala 48:56:@3188.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@3210.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@3212.4]
  reg  _T_153; // @[package.scala 48:56:@3213.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@3221.4 package.scala 96:25:@3222.4]
  wire  _T_158; // @[Controllers.scala 292:61:@3223.4]
  wire  _T_159; // @[Controllers.scala 292:24:@3224.4]
  SRFF active ( // @[Controllers.scala 261:22:@3121.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@3124.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_12 RetimeWrapper ( // @[package.scala 93:22:@3158.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_12 RetimeWrapper_1 ( // @[package.scala 93:22:@3180.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@3192.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@3200.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_16 RetimeWrapper_4 ( // @[package.scala 93:22:@3216.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@3129.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@3130.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@3131.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@3132.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@3149.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@3163.4 package.scala 96:25:@3164.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@3165.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@3168.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@3173.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@3174.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@3177.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@3185.4 package.scala 96:25:@3186.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@3187.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@3212.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@3221.4 package.scala 96:25:@3222.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@3223.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@3224.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@3191.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@3226.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@3176.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@3179.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@3171.4]
  assign active_clock = clock; // @[:@3122.4]
  assign active_reset = reset; // @[:@3123.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@3134.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@3138.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@3139.4]
  assign done_clock = clock; // @[:@3125.4]
  assign done_reset = reset; // @[:@3126.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@3154.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@3147.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@3148.4]
  assign RetimeWrapper_clock = clock; // @[:@3159.4]
  assign RetimeWrapper_reset = reset; // @[:@3160.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@3162.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@3161.4]
  assign RetimeWrapper_1_clock = clock; // @[:@3181.4]
  assign RetimeWrapper_1_reset = reset; // @[:@3182.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@3184.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@3183.4]
  assign RetimeWrapper_2_clock = clock; // @[:@3193.4]
  assign RetimeWrapper_2_reset = reset; // @[:@3194.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@3196.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@3195.4]
  assign RetimeWrapper_3_clock = clock; // @[:@3201.4]
  assign RetimeWrapper_3_reset = reset; // @[:@3202.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@3204.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@3203.4]
  assign RetimeWrapper_4_clock = clock; // @[:@3217.4]
  assign RetimeWrapper_4_reset = reset; // @[:@3218.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@3220.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@3219.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module SimBlackBoxesfix2fixBox( // @[:@3332.2]
  input  [31:0] io_a, // @[:@3335.4]
  output [31:0] io_b // @[:@3335.4]
);
  assign io_b = io_a; // @[SimBlackBoxes.scala 99:40:@3345.4]
endmodule
module _( // @[:@3347.2]
  input  [31:0] io_b, // @[:@3350.4]
  output [31:0] io_result // @[:@3350.4]
);
  wire [31:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@3355.4]
  wire [31:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@3355.4]
  SimBlackBoxesfix2fixBox SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@3355.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@3368.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@3363.4]
endmodule
module RetimeWrapper_21( // @[:@3452.2]
  input        clock, // @[:@3453.4]
  input        reset, // @[:@3454.4]
  input        io_flow, // @[:@3455.4]
  input  [7:0] io_in, // @[:@3455.4]
  output [7:0] io_out // @[:@3455.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@3457.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3470.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3469.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@3468.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3467.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3466.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3464.4]
endmodule
module Mem1D_4( // @[:@3472.2]
  input        clock, // @[:@3473.4]
  input        reset, // @[:@3474.4]
  input        io_r_ofs_0, // @[:@3475.4]
  input        io_r_backpressure, // @[:@3475.4]
  input        io_w_ofs_0, // @[:@3475.4]
  input  [7:0] io_w_data_0, // @[:@3475.4]
  input        io_w_en_0, // @[:@3475.4]
  output [7:0] io_output // @[:@3475.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3485.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3485.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3485.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@3485.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@3485.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@3494.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@3494.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@3494.4]
  wire [7:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@3494.4]
  wire [7:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@3494.4]
  reg [7:0] _T_127; // @[MemPrimitives.scala 560:26:@3479.4]
  reg [31:0] _RAND_0;
  wire  _T_130; // @[MemPrimitives.scala 561:61:@3481.4]
  wire  _T_131; // @[MemPrimitives.scala 561:44:@3482.4]
  wire [7:0] _T_132; // @[MemPrimitives.scala 561:19:@3483.4]
  wire  _T_135; // @[package.scala 96:25:@3490.4 package.scala 96:25:@3491.4]
  wire  _T_137; // @[Mux.scala 46:19:@3492.4]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@3485.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_1 ( // @[package.scala 93:22:@3494.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign _T_130 = io_w_ofs_0 == 1'h0; // @[MemPrimitives.scala 561:61:@3481.4]
  assign _T_131 = io_w_en_0 & _T_130; // @[MemPrimitives.scala 561:44:@3482.4]
  assign _T_132 = _T_131 ? io_w_data_0 : _T_127; // @[MemPrimitives.scala 561:19:@3483.4]
  assign _T_135 = RetimeWrapper_io_out; // @[package.scala 96:25:@3490.4 package.scala 96:25:@3491.4]
  assign _T_137 = 1'h0 == _T_135; // @[Mux.scala 46:19:@3492.4]
  assign io_output = RetimeWrapper_1_io_out; // @[MemPrimitives.scala 565:17:@3501.4]
  assign RetimeWrapper_clock = clock; // @[:@3486.4]
  assign RetimeWrapper_reset = reset; // @[:@3487.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@3489.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@3488.4]
  assign RetimeWrapper_1_clock = clock; // @[:@3495.4]
  assign RetimeWrapper_1_reset = reset; // @[:@3496.4]
  assign RetimeWrapper_1_io_flow = io_r_backpressure; // @[package.scala 95:18:@3498.4]
  assign RetimeWrapper_1_io_in = _T_137 ? _T_127 : 8'h0; // @[package.scala 94:16:@3497.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_127 = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_127 <= 8'h0;
    end else begin
      if (_T_131) begin
        _T_127 <= io_w_data_0;
      end
    end
  end
endmodule
module StickySelects( // @[:@4928.2]
  input   clock, // @[:@4929.4]
  input   reset, // @[:@4930.4]
  input   io_ins_0, // @[:@4931.4]
  input   io_ins_1, // @[:@4931.4]
  input   io_ins_2, // @[:@4931.4]
  input   io_ins_3, // @[:@4931.4]
  input   io_ins_4, // @[:@4931.4]
  input   io_ins_5, // @[:@4931.4]
  output  io_outs_0, // @[:@4931.4]
  output  io_outs_1, // @[:@4931.4]
  output  io_outs_2, // @[:@4931.4]
  output  io_outs_3, // @[:@4931.4]
  output  io_outs_4, // @[:@4931.4]
  output  io_outs_5 // @[:@4931.4]
);
  reg  _T_19; // @[StickySelects.scala 21:22:@4933.4]
  reg [31:0] _RAND_0;
  wire  _T_20; // @[StickySelects.scala 22:54:@4934.4]
  wire  _T_21; // @[StickySelects.scala 22:54:@4935.4]
  wire  _T_22; // @[StickySelects.scala 22:54:@4936.4]
  wire  _T_23; // @[StickySelects.scala 22:54:@4937.4]
  wire  _T_25; // @[StickySelects.scala 24:52:@4938.4]
  wire  _T_26; // @[StickySelects.scala 24:21:@4939.4]
  reg  _T_29; // @[StickySelects.scala 21:22:@4941.4]
  reg [31:0] _RAND_1;
  wire  _T_30; // @[StickySelects.scala 22:54:@4942.4]
  wire  _T_31; // @[StickySelects.scala 22:54:@4943.4]
  wire  _T_32; // @[StickySelects.scala 22:54:@4944.4]
  wire  _T_33; // @[StickySelects.scala 22:54:@4945.4]
  wire  _T_35; // @[StickySelects.scala 24:52:@4946.4]
  wire  _T_36; // @[StickySelects.scala 24:21:@4947.4]
  reg  _T_39; // @[StickySelects.scala 21:22:@4949.4]
  reg [31:0] _RAND_2;
  wire  _T_40; // @[StickySelects.scala 22:54:@4950.4]
  wire  _T_41; // @[StickySelects.scala 22:54:@4951.4]
  wire  _T_42; // @[StickySelects.scala 22:54:@4952.4]
  wire  _T_43; // @[StickySelects.scala 22:54:@4953.4]
  wire  _T_45; // @[StickySelects.scala 24:52:@4954.4]
  wire  _T_46; // @[StickySelects.scala 24:21:@4955.4]
  reg  _T_49; // @[StickySelects.scala 21:22:@4957.4]
  reg [31:0] _RAND_3;
  wire  _T_51; // @[StickySelects.scala 22:54:@4959.4]
  wire  _T_52; // @[StickySelects.scala 22:54:@4960.4]
  wire  _T_53; // @[StickySelects.scala 22:54:@4961.4]
  wire  _T_55; // @[StickySelects.scala 24:52:@4962.4]
  wire  _T_56; // @[StickySelects.scala 24:21:@4963.4]
  reg  _T_59; // @[StickySelects.scala 21:22:@4965.4]
  reg [31:0] _RAND_4;
  wire  _T_62; // @[StickySelects.scala 22:54:@4968.4]
  wire  _T_63; // @[StickySelects.scala 22:54:@4969.4]
  wire  _T_65; // @[StickySelects.scala 24:52:@4970.4]
  wire  _T_66; // @[StickySelects.scala 24:21:@4971.4]
  reg  _T_69; // @[StickySelects.scala 21:22:@4973.4]
  reg [31:0] _RAND_5;
  wire  _T_73; // @[StickySelects.scala 22:54:@4977.4]
  wire  _T_75; // @[StickySelects.scala 24:52:@4978.4]
  wire  _T_76; // @[StickySelects.scala 24:21:@4979.4]
  assign _T_20 = io_ins_1 | io_ins_2; // @[StickySelects.scala 22:54:@4934.4]
  assign _T_21 = _T_20 | io_ins_3; // @[StickySelects.scala 22:54:@4935.4]
  assign _T_22 = _T_21 | io_ins_4; // @[StickySelects.scala 22:54:@4936.4]
  assign _T_23 = _T_22 | io_ins_5; // @[StickySelects.scala 22:54:@4937.4]
  assign _T_25 = io_ins_0 | _T_19; // @[StickySelects.scala 24:52:@4938.4]
  assign _T_26 = _T_23 ? 1'h0 : _T_25; // @[StickySelects.scala 24:21:@4939.4]
  assign _T_30 = io_ins_0 | io_ins_2; // @[StickySelects.scala 22:54:@4942.4]
  assign _T_31 = _T_30 | io_ins_3; // @[StickySelects.scala 22:54:@4943.4]
  assign _T_32 = _T_31 | io_ins_4; // @[StickySelects.scala 22:54:@4944.4]
  assign _T_33 = _T_32 | io_ins_5; // @[StickySelects.scala 22:54:@4945.4]
  assign _T_35 = io_ins_1 | _T_29; // @[StickySelects.scala 24:52:@4946.4]
  assign _T_36 = _T_33 ? 1'h0 : _T_35; // @[StickySelects.scala 24:21:@4947.4]
  assign _T_40 = io_ins_0 | io_ins_1; // @[StickySelects.scala 22:54:@4950.4]
  assign _T_41 = _T_40 | io_ins_3; // @[StickySelects.scala 22:54:@4951.4]
  assign _T_42 = _T_41 | io_ins_4; // @[StickySelects.scala 22:54:@4952.4]
  assign _T_43 = _T_42 | io_ins_5; // @[StickySelects.scala 22:54:@4953.4]
  assign _T_45 = io_ins_2 | _T_39; // @[StickySelects.scala 24:52:@4954.4]
  assign _T_46 = _T_43 ? 1'h0 : _T_45; // @[StickySelects.scala 24:21:@4955.4]
  assign _T_51 = _T_40 | io_ins_2; // @[StickySelects.scala 22:54:@4959.4]
  assign _T_52 = _T_51 | io_ins_4; // @[StickySelects.scala 22:54:@4960.4]
  assign _T_53 = _T_52 | io_ins_5; // @[StickySelects.scala 22:54:@4961.4]
  assign _T_55 = io_ins_3 | _T_49; // @[StickySelects.scala 24:52:@4962.4]
  assign _T_56 = _T_53 ? 1'h0 : _T_55; // @[StickySelects.scala 24:21:@4963.4]
  assign _T_62 = _T_51 | io_ins_3; // @[StickySelects.scala 22:54:@4968.4]
  assign _T_63 = _T_62 | io_ins_5; // @[StickySelects.scala 22:54:@4969.4]
  assign _T_65 = io_ins_4 | _T_59; // @[StickySelects.scala 24:52:@4970.4]
  assign _T_66 = _T_63 ? 1'h0 : _T_65; // @[StickySelects.scala 24:21:@4971.4]
  assign _T_73 = _T_62 | io_ins_4; // @[StickySelects.scala 22:54:@4977.4]
  assign _T_75 = io_ins_5 | _T_69; // @[StickySelects.scala 24:52:@4978.4]
  assign _T_76 = _T_73 ? 1'h0 : _T_75; // @[StickySelects.scala 24:21:@4979.4]
  assign io_outs_0 = _T_23 ? 1'h0 : _T_25; // @[StickySelects.scala 28:52:@4981.4]
  assign io_outs_1 = _T_33 ? 1'h0 : _T_35; // @[StickySelects.scala 28:52:@4982.4]
  assign io_outs_2 = _T_43 ? 1'h0 : _T_45; // @[StickySelects.scala 28:52:@4983.4]
  assign io_outs_3 = _T_53 ? 1'h0 : _T_55; // @[StickySelects.scala 28:52:@4984.4]
  assign io_outs_4 = _T_63 ? 1'h0 : _T_65; // @[StickySelects.scala 28:52:@4985.4]
  assign io_outs_5 = _T_73 ? 1'h0 : _T_75; // @[StickySelects.scala 28:52:@4986.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_29 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_39 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_49 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_59 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_69 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (_T_23) begin
        _T_19 <= 1'h0;
      end else begin
        _T_19 <= _T_25;
      end
    end
    if (reset) begin
      _T_29 <= 1'h0;
    end else begin
      if (_T_33) begin
        _T_29 <= 1'h0;
      end else begin
        _T_29 <= _T_35;
      end
    end
    if (reset) begin
      _T_39 <= 1'h0;
    end else begin
      if (_T_43) begin
        _T_39 <= 1'h0;
      end else begin
        _T_39 <= _T_45;
      end
    end
    if (reset) begin
      _T_49 <= 1'h0;
    end else begin
      if (_T_53) begin
        _T_49 <= 1'h0;
      end else begin
        _T_49 <= _T_55;
      end
    end
    if (reset) begin
      _T_59 <= 1'h0;
    end else begin
      if (_T_63) begin
        _T_59 <= 1'h0;
      end else begin
        _T_59 <= _T_65;
      end
    end
    if (reset) begin
      _T_69 <= 1'h0;
    end else begin
      if (_T_73) begin
        _T_69 <= 1'h0;
      end else begin
        _T_69 <= _T_75;
      end
    end
  end
endmodule
module RetimeWrapper_52( // @[:@5900.2]
  input   clock, // @[:@5901.4]
  input   reset, // @[:@5902.4]
  input   io_flow, // @[:@5903.4]
  input   io_in, // @[:@5903.4]
  output  io_out // @[:@5903.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@5905.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@5905.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@5905.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@5905.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@5905.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@5905.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@5905.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@5918.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@5917.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@5916.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@5915.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@5914.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@5912.4]
endmodule
module x283_lb_0( // @[:@8960.2]
  input        clock, // @[:@8961.4]
  input        reset, // @[:@8962.4]
  input  [2:0] io_rPort_11_banks_1, // @[:@8963.4]
  input  [2:0] io_rPort_11_banks_0, // @[:@8963.4]
  input        io_rPort_11_ofs_0, // @[:@8963.4]
  input        io_rPort_11_en_0, // @[:@8963.4]
  input        io_rPort_11_backpressure, // @[:@8963.4]
  output [7:0] io_rPort_11_output_0, // @[:@8963.4]
  input  [2:0] io_rPort_10_banks_1, // @[:@8963.4]
  input  [2:0] io_rPort_10_banks_0, // @[:@8963.4]
  input        io_rPort_10_ofs_0, // @[:@8963.4]
  input        io_rPort_10_en_0, // @[:@8963.4]
  input        io_rPort_10_backpressure, // @[:@8963.4]
  output [7:0] io_rPort_10_output_0, // @[:@8963.4]
  input  [2:0] io_rPort_9_banks_1, // @[:@8963.4]
  input  [2:0] io_rPort_9_banks_0, // @[:@8963.4]
  input        io_rPort_9_ofs_0, // @[:@8963.4]
  input        io_rPort_9_en_0, // @[:@8963.4]
  input        io_rPort_9_backpressure, // @[:@8963.4]
  output [7:0] io_rPort_9_output_0, // @[:@8963.4]
  input  [2:0] io_rPort_8_banks_1, // @[:@8963.4]
  input  [2:0] io_rPort_8_banks_0, // @[:@8963.4]
  input        io_rPort_8_ofs_0, // @[:@8963.4]
  input        io_rPort_8_en_0, // @[:@8963.4]
  input        io_rPort_8_backpressure, // @[:@8963.4]
  output [7:0] io_rPort_8_output_0, // @[:@8963.4]
  input  [2:0] io_rPort_7_banks_1, // @[:@8963.4]
  input  [2:0] io_rPort_7_banks_0, // @[:@8963.4]
  input        io_rPort_7_ofs_0, // @[:@8963.4]
  input        io_rPort_7_en_0, // @[:@8963.4]
  input        io_rPort_7_backpressure, // @[:@8963.4]
  output [7:0] io_rPort_7_output_0, // @[:@8963.4]
  input  [2:0] io_rPort_6_banks_1, // @[:@8963.4]
  input  [2:0] io_rPort_6_banks_0, // @[:@8963.4]
  input        io_rPort_6_ofs_0, // @[:@8963.4]
  input        io_rPort_6_en_0, // @[:@8963.4]
  input        io_rPort_6_backpressure, // @[:@8963.4]
  output [7:0] io_rPort_6_output_0, // @[:@8963.4]
  input  [2:0] io_rPort_5_banks_1, // @[:@8963.4]
  input  [2:0] io_rPort_5_banks_0, // @[:@8963.4]
  input        io_rPort_5_ofs_0, // @[:@8963.4]
  input        io_rPort_5_en_0, // @[:@8963.4]
  input        io_rPort_5_backpressure, // @[:@8963.4]
  output [7:0] io_rPort_5_output_0, // @[:@8963.4]
  input  [2:0] io_rPort_4_banks_1, // @[:@8963.4]
  input  [2:0] io_rPort_4_banks_0, // @[:@8963.4]
  input        io_rPort_4_ofs_0, // @[:@8963.4]
  input        io_rPort_4_en_0, // @[:@8963.4]
  input        io_rPort_4_backpressure, // @[:@8963.4]
  output [7:0] io_rPort_4_output_0, // @[:@8963.4]
  input  [2:0] io_rPort_3_banks_1, // @[:@8963.4]
  input  [2:0] io_rPort_3_banks_0, // @[:@8963.4]
  input        io_rPort_3_ofs_0, // @[:@8963.4]
  input        io_rPort_3_en_0, // @[:@8963.4]
  input        io_rPort_3_backpressure, // @[:@8963.4]
  output [7:0] io_rPort_3_output_0, // @[:@8963.4]
  input  [2:0] io_rPort_2_banks_1, // @[:@8963.4]
  input  [2:0] io_rPort_2_banks_0, // @[:@8963.4]
  input        io_rPort_2_ofs_0, // @[:@8963.4]
  input        io_rPort_2_en_0, // @[:@8963.4]
  input        io_rPort_2_backpressure, // @[:@8963.4]
  output [7:0] io_rPort_2_output_0, // @[:@8963.4]
  input  [2:0] io_rPort_1_banks_1, // @[:@8963.4]
  input  [2:0] io_rPort_1_banks_0, // @[:@8963.4]
  input        io_rPort_1_ofs_0, // @[:@8963.4]
  input        io_rPort_1_en_0, // @[:@8963.4]
  input        io_rPort_1_backpressure, // @[:@8963.4]
  output [7:0] io_rPort_1_output_0, // @[:@8963.4]
  input  [2:0] io_rPort_0_banks_1, // @[:@8963.4]
  input  [2:0] io_rPort_0_banks_0, // @[:@8963.4]
  input        io_rPort_0_ofs_0, // @[:@8963.4]
  input        io_rPort_0_en_0, // @[:@8963.4]
  input        io_rPort_0_backpressure, // @[:@8963.4]
  output [7:0] io_rPort_0_output_0, // @[:@8963.4]
  input  [2:0] io_wPort_1_banks_1, // @[:@8963.4]
  input  [2:0] io_wPort_1_banks_0, // @[:@8963.4]
  input        io_wPort_1_ofs_0, // @[:@8963.4]
  input  [7:0] io_wPort_1_data_0, // @[:@8963.4]
  input        io_wPort_1_en_0, // @[:@8963.4]
  input  [2:0] io_wPort_0_banks_1, // @[:@8963.4]
  input  [2:0] io_wPort_0_banks_0, // @[:@8963.4]
  input        io_wPort_0_ofs_0, // @[:@8963.4]
  input  [7:0] io_wPort_0_data_0, // @[:@8963.4]
  input        io_wPort_0_en_0 // @[:@8963.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@9054.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@9054.4]
  wire  Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9054.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9054.4]
  wire  Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9054.4]
  wire [7:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@9054.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@9054.4]
  wire [7:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@9054.4]
  wire  Mem1D_1_clock; // @[MemPrimitives.scala 64:21:@9070.4]
  wire  Mem1D_1_reset; // @[MemPrimitives.scala 64:21:@9070.4]
  wire  Mem1D_1_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9070.4]
  wire  Mem1D_1_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9070.4]
  wire  Mem1D_1_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9070.4]
  wire [7:0] Mem1D_1_io_w_data_0; // @[MemPrimitives.scala 64:21:@9070.4]
  wire  Mem1D_1_io_w_en_0; // @[MemPrimitives.scala 64:21:@9070.4]
  wire [7:0] Mem1D_1_io_output; // @[MemPrimitives.scala 64:21:@9070.4]
  wire  Mem1D_2_clock; // @[MemPrimitives.scala 64:21:@9086.4]
  wire  Mem1D_2_reset; // @[MemPrimitives.scala 64:21:@9086.4]
  wire  Mem1D_2_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9086.4]
  wire  Mem1D_2_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9086.4]
  wire  Mem1D_2_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9086.4]
  wire [7:0] Mem1D_2_io_w_data_0; // @[MemPrimitives.scala 64:21:@9086.4]
  wire  Mem1D_2_io_w_en_0; // @[MemPrimitives.scala 64:21:@9086.4]
  wire [7:0] Mem1D_2_io_output; // @[MemPrimitives.scala 64:21:@9086.4]
  wire  Mem1D_3_clock; // @[MemPrimitives.scala 64:21:@9102.4]
  wire  Mem1D_3_reset; // @[MemPrimitives.scala 64:21:@9102.4]
  wire  Mem1D_3_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9102.4]
  wire  Mem1D_3_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9102.4]
  wire  Mem1D_3_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9102.4]
  wire [7:0] Mem1D_3_io_w_data_0; // @[MemPrimitives.scala 64:21:@9102.4]
  wire  Mem1D_3_io_w_en_0; // @[MemPrimitives.scala 64:21:@9102.4]
  wire [7:0] Mem1D_3_io_output; // @[MemPrimitives.scala 64:21:@9102.4]
  wire  Mem1D_4_clock; // @[MemPrimitives.scala 64:21:@9118.4]
  wire  Mem1D_4_reset; // @[MemPrimitives.scala 64:21:@9118.4]
  wire  Mem1D_4_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9118.4]
  wire  Mem1D_4_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9118.4]
  wire  Mem1D_4_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9118.4]
  wire [7:0] Mem1D_4_io_w_data_0; // @[MemPrimitives.scala 64:21:@9118.4]
  wire  Mem1D_4_io_w_en_0; // @[MemPrimitives.scala 64:21:@9118.4]
  wire [7:0] Mem1D_4_io_output; // @[MemPrimitives.scala 64:21:@9118.4]
  wire  Mem1D_5_clock; // @[MemPrimitives.scala 64:21:@9134.4]
  wire  Mem1D_5_reset; // @[MemPrimitives.scala 64:21:@9134.4]
  wire  Mem1D_5_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9134.4]
  wire  Mem1D_5_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9134.4]
  wire  Mem1D_5_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9134.4]
  wire [7:0] Mem1D_5_io_w_data_0; // @[MemPrimitives.scala 64:21:@9134.4]
  wire  Mem1D_5_io_w_en_0; // @[MemPrimitives.scala 64:21:@9134.4]
  wire [7:0] Mem1D_5_io_output; // @[MemPrimitives.scala 64:21:@9134.4]
  wire  Mem1D_6_clock; // @[MemPrimitives.scala 64:21:@9150.4]
  wire  Mem1D_6_reset; // @[MemPrimitives.scala 64:21:@9150.4]
  wire  Mem1D_6_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9150.4]
  wire  Mem1D_6_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9150.4]
  wire  Mem1D_6_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9150.4]
  wire [7:0] Mem1D_6_io_w_data_0; // @[MemPrimitives.scala 64:21:@9150.4]
  wire  Mem1D_6_io_w_en_0; // @[MemPrimitives.scala 64:21:@9150.4]
  wire [7:0] Mem1D_6_io_output; // @[MemPrimitives.scala 64:21:@9150.4]
  wire  Mem1D_7_clock; // @[MemPrimitives.scala 64:21:@9166.4]
  wire  Mem1D_7_reset; // @[MemPrimitives.scala 64:21:@9166.4]
  wire  Mem1D_7_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9166.4]
  wire  Mem1D_7_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9166.4]
  wire  Mem1D_7_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9166.4]
  wire [7:0] Mem1D_7_io_w_data_0; // @[MemPrimitives.scala 64:21:@9166.4]
  wire  Mem1D_7_io_w_en_0; // @[MemPrimitives.scala 64:21:@9166.4]
  wire [7:0] Mem1D_7_io_output; // @[MemPrimitives.scala 64:21:@9166.4]
  wire  Mem1D_8_clock; // @[MemPrimitives.scala 64:21:@9182.4]
  wire  Mem1D_8_reset; // @[MemPrimitives.scala 64:21:@9182.4]
  wire  Mem1D_8_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9182.4]
  wire  Mem1D_8_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9182.4]
  wire  Mem1D_8_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9182.4]
  wire [7:0] Mem1D_8_io_w_data_0; // @[MemPrimitives.scala 64:21:@9182.4]
  wire  Mem1D_8_io_w_en_0; // @[MemPrimitives.scala 64:21:@9182.4]
  wire [7:0] Mem1D_8_io_output; // @[MemPrimitives.scala 64:21:@9182.4]
  wire  Mem1D_9_clock; // @[MemPrimitives.scala 64:21:@9198.4]
  wire  Mem1D_9_reset; // @[MemPrimitives.scala 64:21:@9198.4]
  wire  Mem1D_9_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9198.4]
  wire  Mem1D_9_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9198.4]
  wire  Mem1D_9_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9198.4]
  wire [7:0] Mem1D_9_io_w_data_0; // @[MemPrimitives.scala 64:21:@9198.4]
  wire  Mem1D_9_io_w_en_0; // @[MemPrimitives.scala 64:21:@9198.4]
  wire [7:0] Mem1D_9_io_output; // @[MemPrimitives.scala 64:21:@9198.4]
  wire  Mem1D_10_clock; // @[MemPrimitives.scala 64:21:@9214.4]
  wire  Mem1D_10_reset; // @[MemPrimitives.scala 64:21:@9214.4]
  wire  Mem1D_10_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9214.4]
  wire  Mem1D_10_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9214.4]
  wire  Mem1D_10_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9214.4]
  wire [7:0] Mem1D_10_io_w_data_0; // @[MemPrimitives.scala 64:21:@9214.4]
  wire  Mem1D_10_io_w_en_0; // @[MemPrimitives.scala 64:21:@9214.4]
  wire [7:0] Mem1D_10_io_output; // @[MemPrimitives.scala 64:21:@9214.4]
  wire  Mem1D_11_clock; // @[MemPrimitives.scala 64:21:@9230.4]
  wire  Mem1D_11_reset; // @[MemPrimitives.scala 64:21:@9230.4]
  wire  Mem1D_11_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9230.4]
  wire  Mem1D_11_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9230.4]
  wire  Mem1D_11_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9230.4]
  wire [7:0] Mem1D_11_io_w_data_0; // @[MemPrimitives.scala 64:21:@9230.4]
  wire  Mem1D_11_io_w_en_0; // @[MemPrimitives.scala 64:21:@9230.4]
  wire [7:0] Mem1D_11_io_output; // @[MemPrimitives.scala 64:21:@9230.4]
  wire  Mem1D_12_clock; // @[MemPrimitives.scala 64:21:@9246.4]
  wire  Mem1D_12_reset; // @[MemPrimitives.scala 64:21:@9246.4]
  wire  Mem1D_12_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9246.4]
  wire  Mem1D_12_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9246.4]
  wire  Mem1D_12_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9246.4]
  wire [7:0] Mem1D_12_io_w_data_0; // @[MemPrimitives.scala 64:21:@9246.4]
  wire  Mem1D_12_io_w_en_0; // @[MemPrimitives.scala 64:21:@9246.4]
  wire [7:0] Mem1D_12_io_output; // @[MemPrimitives.scala 64:21:@9246.4]
  wire  Mem1D_13_clock; // @[MemPrimitives.scala 64:21:@9262.4]
  wire  Mem1D_13_reset; // @[MemPrimitives.scala 64:21:@9262.4]
  wire  Mem1D_13_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9262.4]
  wire  Mem1D_13_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9262.4]
  wire  Mem1D_13_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9262.4]
  wire [7:0] Mem1D_13_io_w_data_0; // @[MemPrimitives.scala 64:21:@9262.4]
  wire  Mem1D_13_io_w_en_0; // @[MemPrimitives.scala 64:21:@9262.4]
  wire [7:0] Mem1D_13_io_output; // @[MemPrimitives.scala 64:21:@9262.4]
  wire  Mem1D_14_clock; // @[MemPrimitives.scala 64:21:@9278.4]
  wire  Mem1D_14_reset; // @[MemPrimitives.scala 64:21:@9278.4]
  wire  Mem1D_14_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9278.4]
  wire  Mem1D_14_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9278.4]
  wire  Mem1D_14_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9278.4]
  wire [7:0] Mem1D_14_io_w_data_0; // @[MemPrimitives.scala 64:21:@9278.4]
  wire  Mem1D_14_io_w_en_0; // @[MemPrimitives.scala 64:21:@9278.4]
  wire [7:0] Mem1D_14_io_output; // @[MemPrimitives.scala 64:21:@9278.4]
  wire  Mem1D_15_clock; // @[MemPrimitives.scala 64:21:@9294.4]
  wire  Mem1D_15_reset; // @[MemPrimitives.scala 64:21:@9294.4]
  wire  Mem1D_15_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9294.4]
  wire  Mem1D_15_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9294.4]
  wire  Mem1D_15_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9294.4]
  wire [7:0] Mem1D_15_io_w_data_0; // @[MemPrimitives.scala 64:21:@9294.4]
  wire  Mem1D_15_io_w_en_0; // @[MemPrimitives.scala 64:21:@9294.4]
  wire [7:0] Mem1D_15_io_output; // @[MemPrimitives.scala 64:21:@9294.4]
  wire  StickySelects_clock; // @[MemPrimitives.scala 121:29:@9526.4]
  wire  StickySelects_reset; // @[MemPrimitives.scala 121:29:@9526.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 121:29:@9526.4]
  wire  StickySelects_io_ins_1; // @[MemPrimitives.scala 121:29:@9526.4]
  wire  StickySelects_io_ins_2; // @[MemPrimitives.scala 121:29:@9526.4]
  wire  StickySelects_io_ins_3; // @[MemPrimitives.scala 121:29:@9526.4]
  wire  StickySelects_io_ins_4; // @[MemPrimitives.scala 121:29:@9526.4]
  wire  StickySelects_io_ins_5; // @[MemPrimitives.scala 121:29:@9526.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 121:29:@9526.4]
  wire  StickySelects_io_outs_1; // @[MemPrimitives.scala 121:29:@9526.4]
  wire  StickySelects_io_outs_2; // @[MemPrimitives.scala 121:29:@9526.4]
  wire  StickySelects_io_outs_3; // @[MemPrimitives.scala 121:29:@9526.4]
  wire  StickySelects_io_outs_4; // @[MemPrimitives.scala 121:29:@9526.4]
  wire  StickySelects_io_outs_5; // @[MemPrimitives.scala 121:29:@9526.4]
  wire  StickySelects_1_clock; // @[MemPrimitives.scala 121:29:@9588.4]
  wire  StickySelects_1_reset; // @[MemPrimitives.scala 121:29:@9588.4]
  wire  StickySelects_1_io_ins_0; // @[MemPrimitives.scala 121:29:@9588.4]
  wire  StickySelects_1_io_ins_1; // @[MemPrimitives.scala 121:29:@9588.4]
  wire  StickySelects_1_io_ins_2; // @[MemPrimitives.scala 121:29:@9588.4]
  wire  StickySelects_1_io_ins_3; // @[MemPrimitives.scala 121:29:@9588.4]
  wire  StickySelects_1_io_ins_4; // @[MemPrimitives.scala 121:29:@9588.4]
  wire  StickySelects_1_io_ins_5; // @[MemPrimitives.scala 121:29:@9588.4]
  wire  StickySelects_1_io_outs_0; // @[MemPrimitives.scala 121:29:@9588.4]
  wire  StickySelects_1_io_outs_1; // @[MemPrimitives.scala 121:29:@9588.4]
  wire  StickySelects_1_io_outs_2; // @[MemPrimitives.scala 121:29:@9588.4]
  wire  StickySelects_1_io_outs_3; // @[MemPrimitives.scala 121:29:@9588.4]
  wire  StickySelects_1_io_outs_4; // @[MemPrimitives.scala 121:29:@9588.4]
  wire  StickySelects_1_io_outs_5; // @[MemPrimitives.scala 121:29:@9588.4]
  wire  StickySelects_2_clock; // @[MemPrimitives.scala 121:29:@9650.4]
  wire  StickySelects_2_reset; // @[MemPrimitives.scala 121:29:@9650.4]
  wire  StickySelects_2_io_ins_0; // @[MemPrimitives.scala 121:29:@9650.4]
  wire  StickySelects_2_io_ins_1; // @[MemPrimitives.scala 121:29:@9650.4]
  wire  StickySelects_2_io_ins_2; // @[MemPrimitives.scala 121:29:@9650.4]
  wire  StickySelects_2_io_ins_3; // @[MemPrimitives.scala 121:29:@9650.4]
  wire  StickySelects_2_io_ins_4; // @[MemPrimitives.scala 121:29:@9650.4]
  wire  StickySelects_2_io_ins_5; // @[MemPrimitives.scala 121:29:@9650.4]
  wire  StickySelects_2_io_outs_0; // @[MemPrimitives.scala 121:29:@9650.4]
  wire  StickySelects_2_io_outs_1; // @[MemPrimitives.scala 121:29:@9650.4]
  wire  StickySelects_2_io_outs_2; // @[MemPrimitives.scala 121:29:@9650.4]
  wire  StickySelects_2_io_outs_3; // @[MemPrimitives.scala 121:29:@9650.4]
  wire  StickySelects_2_io_outs_4; // @[MemPrimitives.scala 121:29:@9650.4]
  wire  StickySelects_2_io_outs_5; // @[MemPrimitives.scala 121:29:@9650.4]
  wire  StickySelects_3_clock; // @[MemPrimitives.scala 121:29:@9712.4]
  wire  StickySelects_3_reset; // @[MemPrimitives.scala 121:29:@9712.4]
  wire  StickySelects_3_io_ins_0; // @[MemPrimitives.scala 121:29:@9712.4]
  wire  StickySelects_3_io_ins_1; // @[MemPrimitives.scala 121:29:@9712.4]
  wire  StickySelects_3_io_ins_2; // @[MemPrimitives.scala 121:29:@9712.4]
  wire  StickySelects_3_io_ins_3; // @[MemPrimitives.scala 121:29:@9712.4]
  wire  StickySelects_3_io_ins_4; // @[MemPrimitives.scala 121:29:@9712.4]
  wire  StickySelects_3_io_ins_5; // @[MemPrimitives.scala 121:29:@9712.4]
  wire  StickySelects_3_io_outs_0; // @[MemPrimitives.scala 121:29:@9712.4]
  wire  StickySelects_3_io_outs_1; // @[MemPrimitives.scala 121:29:@9712.4]
  wire  StickySelects_3_io_outs_2; // @[MemPrimitives.scala 121:29:@9712.4]
  wire  StickySelects_3_io_outs_3; // @[MemPrimitives.scala 121:29:@9712.4]
  wire  StickySelects_3_io_outs_4; // @[MemPrimitives.scala 121:29:@9712.4]
  wire  StickySelects_3_io_outs_5; // @[MemPrimitives.scala 121:29:@9712.4]
  wire  StickySelects_4_clock; // @[MemPrimitives.scala 121:29:@9774.4]
  wire  StickySelects_4_reset; // @[MemPrimitives.scala 121:29:@9774.4]
  wire  StickySelects_4_io_ins_0; // @[MemPrimitives.scala 121:29:@9774.4]
  wire  StickySelects_4_io_ins_1; // @[MemPrimitives.scala 121:29:@9774.4]
  wire  StickySelects_4_io_ins_2; // @[MemPrimitives.scala 121:29:@9774.4]
  wire  StickySelects_4_io_ins_3; // @[MemPrimitives.scala 121:29:@9774.4]
  wire  StickySelects_4_io_ins_4; // @[MemPrimitives.scala 121:29:@9774.4]
  wire  StickySelects_4_io_ins_5; // @[MemPrimitives.scala 121:29:@9774.4]
  wire  StickySelects_4_io_outs_0; // @[MemPrimitives.scala 121:29:@9774.4]
  wire  StickySelects_4_io_outs_1; // @[MemPrimitives.scala 121:29:@9774.4]
  wire  StickySelects_4_io_outs_2; // @[MemPrimitives.scala 121:29:@9774.4]
  wire  StickySelects_4_io_outs_3; // @[MemPrimitives.scala 121:29:@9774.4]
  wire  StickySelects_4_io_outs_4; // @[MemPrimitives.scala 121:29:@9774.4]
  wire  StickySelects_4_io_outs_5; // @[MemPrimitives.scala 121:29:@9774.4]
  wire  StickySelects_5_clock; // @[MemPrimitives.scala 121:29:@9836.4]
  wire  StickySelects_5_reset; // @[MemPrimitives.scala 121:29:@9836.4]
  wire  StickySelects_5_io_ins_0; // @[MemPrimitives.scala 121:29:@9836.4]
  wire  StickySelects_5_io_ins_1; // @[MemPrimitives.scala 121:29:@9836.4]
  wire  StickySelects_5_io_ins_2; // @[MemPrimitives.scala 121:29:@9836.4]
  wire  StickySelects_5_io_ins_3; // @[MemPrimitives.scala 121:29:@9836.4]
  wire  StickySelects_5_io_ins_4; // @[MemPrimitives.scala 121:29:@9836.4]
  wire  StickySelects_5_io_ins_5; // @[MemPrimitives.scala 121:29:@9836.4]
  wire  StickySelects_5_io_outs_0; // @[MemPrimitives.scala 121:29:@9836.4]
  wire  StickySelects_5_io_outs_1; // @[MemPrimitives.scala 121:29:@9836.4]
  wire  StickySelects_5_io_outs_2; // @[MemPrimitives.scala 121:29:@9836.4]
  wire  StickySelects_5_io_outs_3; // @[MemPrimitives.scala 121:29:@9836.4]
  wire  StickySelects_5_io_outs_4; // @[MemPrimitives.scala 121:29:@9836.4]
  wire  StickySelects_5_io_outs_5; // @[MemPrimitives.scala 121:29:@9836.4]
  wire  StickySelects_6_clock; // @[MemPrimitives.scala 121:29:@9898.4]
  wire  StickySelects_6_reset; // @[MemPrimitives.scala 121:29:@9898.4]
  wire  StickySelects_6_io_ins_0; // @[MemPrimitives.scala 121:29:@9898.4]
  wire  StickySelects_6_io_ins_1; // @[MemPrimitives.scala 121:29:@9898.4]
  wire  StickySelects_6_io_ins_2; // @[MemPrimitives.scala 121:29:@9898.4]
  wire  StickySelects_6_io_ins_3; // @[MemPrimitives.scala 121:29:@9898.4]
  wire  StickySelects_6_io_ins_4; // @[MemPrimitives.scala 121:29:@9898.4]
  wire  StickySelects_6_io_ins_5; // @[MemPrimitives.scala 121:29:@9898.4]
  wire  StickySelects_6_io_outs_0; // @[MemPrimitives.scala 121:29:@9898.4]
  wire  StickySelects_6_io_outs_1; // @[MemPrimitives.scala 121:29:@9898.4]
  wire  StickySelects_6_io_outs_2; // @[MemPrimitives.scala 121:29:@9898.4]
  wire  StickySelects_6_io_outs_3; // @[MemPrimitives.scala 121:29:@9898.4]
  wire  StickySelects_6_io_outs_4; // @[MemPrimitives.scala 121:29:@9898.4]
  wire  StickySelects_6_io_outs_5; // @[MemPrimitives.scala 121:29:@9898.4]
  wire  StickySelects_7_clock; // @[MemPrimitives.scala 121:29:@9960.4]
  wire  StickySelects_7_reset; // @[MemPrimitives.scala 121:29:@9960.4]
  wire  StickySelects_7_io_ins_0; // @[MemPrimitives.scala 121:29:@9960.4]
  wire  StickySelects_7_io_ins_1; // @[MemPrimitives.scala 121:29:@9960.4]
  wire  StickySelects_7_io_ins_2; // @[MemPrimitives.scala 121:29:@9960.4]
  wire  StickySelects_7_io_ins_3; // @[MemPrimitives.scala 121:29:@9960.4]
  wire  StickySelects_7_io_ins_4; // @[MemPrimitives.scala 121:29:@9960.4]
  wire  StickySelects_7_io_ins_5; // @[MemPrimitives.scala 121:29:@9960.4]
  wire  StickySelects_7_io_outs_0; // @[MemPrimitives.scala 121:29:@9960.4]
  wire  StickySelects_7_io_outs_1; // @[MemPrimitives.scala 121:29:@9960.4]
  wire  StickySelects_7_io_outs_2; // @[MemPrimitives.scala 121:29:@9960.4]
  wire  StickySelects_7_io_outs_3; // @[MemPrimitives.scala 121:29:@9960.4]
  wire  StickySelects_7_io_outs_4; // @[MemPrimitives.scala 121:29:@9960.4]
  wire  StickySelects_7_io_outs_5; // @[MemPrimitives.scala 121:29:@9960.4]
  wire  StickySelects_8_clock; // @[MemPrimitives.scala 121:29:@10022.4]
  wire  StickySelects_8_reset; // @[MemPrimitives.scala 121:29:@10022.4]
  wire  StickySelects_8_io_ins_0; // @[MemPrimitives.scala 121:29:@10022.4]
  wire  StickySelects_8_io_ins_1; // @[MemPrimitives.scala 121:29:@10022.4]
  wire  StickySelects_8_io_ins_2; // @[MemPrimitives.scala 121:29:@10022.4]
  wire  StickySelects_8_io_ins_3; // @[MemPrimitives.scala 121:29:@10022.4]
  wire  StickySelects_8_io_ins_4; // @[MemPrimitives.scala 121:29:@10022.4]
  wire  StickySelects_8_io_ins_5; // @[MemPrimitives.scala 121:29:@10022.4]
  wire  StickySelects_8_io_outs_0; // @[MemPrimitives.scala 121:29:@10022.4]
  wire  StickySelects_8_io_outs_1; // @[MemPrimitives.scala 121:29:@10022.4]
  wire  StickySelects_8_io_outs_2; // @[MemPrimitives.scala 121:29:@10022.4]
  wire  StickySelects_8_io_outs_3; // @[MemPrimitives.scala 121:29:@10022.4]
  wire  StickySelects_8_io_outs_4; // @[MemPrimitives.scala 121:29:@10022.4]
  wire  StickySelects_8_io_outs_5; // @[MemPrimitives.scala 121:29:@10022.4]
  wire  StickySelects_9_clock; // @[MemPrimitives.scala 121:29:@10084.4]
  wire  StickySelects_9_reset; // @[MemPrimitives.scala 121:29:@10084.4]
  wire  StickySelects_9_io_ins_0; // @[MemPrimitives.scala 121:29:@10084.4]
  wire  StickySelects_9_io_ins_1; // @[MemPrimitives.scala 121:29:@10084.4]
  wire  StickySelects_9_io_ins_2; // @[MemPrimitives.scala 121:29:@10084.4]
  wire  StickySelects_9_io_ins_3; // @[MemPrimitives.scala 121:29:@10084.4]
  wire  StickySelects_9_io_ins_4; // @[MemPrimitives.scala 121:29:@10084.4]
  wire  StickySelects_9_io_ins_5; // @[MemPrimitives.scala 121:29:@10084.4]
  wire  StickySelects_9_io_outs_0; // @[MemPrimitives.scala 121:29:@10084.4]
  wire  StickySelects_9_io_outs_1; // @[MemPrimitives.scala 121:29:@10084.4]
  wire  StickySelects_9_io_outs_2; // @[MemPrimitives.scala 121:29:@10084.4]
  wire  StickySelects_9_io_outs_3; // @[MemPrimitives.scala 121:29:@10084.4]
  wire  StickySelects_9_io_outs_4; // @[MemPrimitives.scala 121:29:@10084.4]
  wire  StickySelects_9_io_outs_5; // @[MemPrimitives.scala 121:29:@10084.4]
  wire  StickySelects_10_clock; // @[MemPrimitives.scala 121:29:@10146.4]
  wire  StickySelects_10_reset; // @[MemPrimitives.scala 121:29:@10146.4]
  wire  StickySelects_10_io_ins_0; // @[MemPrimitives.scala 121:29:@10146.4]
  wire  StickySelects_10_io_ins_1; // @[MemPrimitives.scala 121:29:@10146.4]
  wire  StickySelects_10_io_ins_2; // @[MemPrimitives.scala 121:29:@10146.4]
  wire  StickySelects_10_io_ins_3; // @[MemPrimitives.scala 121:29:@10146.4]
  wire  StickySelects_10_io_ins_4; // @[MemPrimitives.scala 121:29:@10146.4]
  wire  StickySelects_10_io_ins_5; // @[MemPrimitives.scala 121:29:@10146.4]
  wire  StickySelects_10_io_outs_0; // @[MemPrimitives.scala 121:29:@10146.4]
  wire  StickySelects_10_io_outs_1; // @[MemPrimitives.scala 121:29:@10146.4]
  wire  StickySelects_10_io_outs_2; // @[MemPrimitives.scala 121:29:@10146.4]
  wire  StickySelects_10_io_outs_3; // @[MemPrimitives.scala 121:29:@10146.4]
  wire  StickySelects_10_io_outs_4; // @[MemPrimitives.scala 121:29:@10146.4]
  wire  StickySelects_10_io_outs_5; // @[MemPrimitives.scala 121:29:@10146.4]
  wire  StickySelects_11_clock; // @[MemPrimitives.scala 121:29:@10208.4]
  wire  StickySelects_11_reset; // @[MemPrimitives.scala 121:29:@10208.4]
  wire  StickySelects_11_io_ins_0; // @[MemPrimitives.scala 121:29:@10208.4]
  wire  StickySelects_11_io_ins_1; // @[MemPrimitives.scala 121:29:@10208.4]
  wire  StickySelects_11_io_ins_2; // @[MemPrimitives.scala 121:29:@10208.4]
  wire  StickySelects_11_io_ins_3; // @[MemPrimitives.scala 121:29:@10208.4]
  wire  StickySelects_11_io_ins_4; // @[MemPrimitives.scala 121:29:@10208.4]
  wire  StickySelects_11_io_ins_5; // @[MemPrimitives.scala 121:29:@10208.4]
  wire  StickySelects_11_io_outs_0; // @[MemPrimitives.scala 121:29:@10208.4]
  wire  StickySelects_11_io_outs_1; // @[MemPrimitives.scala 121:29:@10208.4]
  wire  StickySelects_11_io_outs_2; // @[MemPrimitives.scala 121:29:@10208.4]
  wire  StickySelects_11_io_outs_3; // @[MemPrimitives.scala 121:29:@10208.4]
  wire  StickySelects_11_io_outs_4; // @[MemPrimitives.scala 121:29:@10208.4]
  wire  StickySelects_11_io_outs_5; // @[MemPrimitives.scala 121:29:@10208.4]
  wire  StickySelects_12_clock; // @[MemPrimitives.scala 121:29:@10270.4]
  wire  StickySelects_12_reset; // @[MemPrimitives.scala 121:29:@10270.4]
  wire  StickySelects_12_io_ins_0; // @[MemPrimitives.scala 121:29:@10270.4]
  wire  StickySelects_12_io_ins_1; // @[MemPrimitives.scala 121:29:@10270.4]
  wire  StickySelects_12_io_ins_2; // @[MemPrimitives.scala 121:29:@10270.4]
  wire  StickySelects_12_io_ins_3; // @[MemPrimitives.scala 121:29:@10270.4]
  wire  StickySelects_12_io_ins_4; // @[MemPrimitives.scala 121:29:@10270.4]
  wire  StickySelects_12_io_ins_5; // @[MemPrimitives.scala 121:29:@10270.4]
  wire  StickySelects_12_io_outs_0; // @[MemPrimitives.scala 121:29:@10270.4]
  wire  StickySelects_12_io_outs_1; // @[MemPrimitives.scala 121:29:@10270.4]
  wire  StickySelects_12_io_outs_2; // @[MemPrimitives.scala 121:29:@10270.4]
  wire  StickySelects_12_io_outs_3; // @[MemPrimitives.scala 121:29:@10270.4]
  wire  StickySelects_12_io_outs_4; // @[MemPrimitives.scala 121:29:@10270.4]
  wire  StickySelects_12_io_outs_5; // @[MemPrimitives.scala 121:29:@10270.4]
  wire  StickySelects_13_clock; // @[MemPrimitives.scala 121:29:@10332.4]
  wire  StickySelects_13_reset; // @[MemPrimitives.scala 121:29:@10332.4]
  wire  StickySelects_13_io_ins_0; // @[MemPrimitives.scala 121:29:@10332.4]
  wire  StickySelects_13_io_ins_1; // @[MemPrimitives.scala 121:29:@10332.4]
  wire  StickySelects_13_io_ins_2; // @[MemPrimitives.scala 121:29:@10332.4]
  wire  StickySelects_13_io_ins_3; // @[MemPrimitives.scala 121:29:@10332.4]
  wire  StickySelects_13_io_ins_4; // @[MemPrimitives.scala 121:29:@10332.4]
  wire  StickySelects_13_io_ins_5; // @[MemPrimitives.scala 121:29:@10332.4]
  wire  StickySelects_13_io_outs_0; // @[MemPrimitives.scala 121:29:@10332.4]
  wire  StickySelects_13_io_outs_1; // @[MemPrimitives.scala 121:29:@10332.4]
  wire  StickySelects_13_io_outs_2; // @[MemPrimitives.scala 121:29:@10332.4]
  wire  StickySelects_13_io_outs_3; // @[MemPrimitives.scala 121:29:@10332.4]
  wire  StickySelects_13_io_outs_4; // @[MemPrimitives.scala 121:29:@10332.4]
  wire  StickySelects_13_io_outs_5; // @[MemPrimitives.scala 121:29:@10332.4]
  wire  StickySelects_14_clock; // @[MemPrimitives.scala 121:29:@10394.4]
  wire  StickySelects_14_reset; // @[MemPrimitives.scala 121:29:@10394.4]
  wire  StickySelects_14_io_ins_0; // @[MemPrimitives.scala 121:29:@10394.4]
  wire  StickySelects_14_io_ins_1; // @[MemPrimitives.scala 121:29:@10394.4]
  wire  StickySelects_14_io_ins_2; // @[MemPrimitives.scala 121:29:@10394.4]
  wire  StickySelects_14_io_ins_3; // @[MemPrimitives.scala 121:29:@10394.4]
  wire  StickySelects_14_io_ins_4; // @[MemPrimitives.scala 121:29:@10394.4]
  wire  StickySelects_14_io_ins_5; // @[MemPrimitives.scala 121:29:@10394.4]
  wire  StickySelects_14_io_outs_0; // @[MemPrimitives.scala 121:29:@10394.4]
  wire  StickySelects_14_io_outs_1; // @[MemPrimitives.scala 121:29:@10394.4]
  wire  StickySelects_14_io_outs_2; // @[MemPrimitives.scala 121:29:@10394.4]
  wire  StickySelects_14_io_outs_3; // @[MemPrimitives.scala 121:29:@10394.4]
  wire  StickySelects_14_io_outs_4; // @[MemPrimitives.scala 121:29:@10394.4]
  wire  StickySelects_14_io_outs_5; // @[MemPrimitives.scala 121:29:@10394.4]
  wire  StickySelects_15_clock; // @[MemPrimitives.scala 121:29:@10456.4]
  wire  StickySelects_15_reset; // @[MemPrimitives.scala 121:29:@10456.4]
  wire  StickySelects_15_io_ins_0; // @[MemPrimitives.scala 121:29:@10456.4]
  wire  StickySelects_15_io_ins_1; // @[MemPrimitives.scala 121:29:@10456.4]
  wire  StickySelects_15_io_ins_2; // @[MemPrimitives.scala 121:29:@10456.4]
  wire  StickySelects_15_io_ins_3; // @[MemPrimitives.scala 121:29:@10456.4]
  wire  StickySelects_15_io_ins_4; // @[MemPrimitives.scala 121:29:@10456.4]
  wire  StickySelects_15_io_ins_5; // @[MemPrimitives.scala 121:29:@10456.4]
  wire  StickySelects_15_io_outs_0; // @[MemPrimitives.scala 121:29:@10456.4]
  wire  StickySelects_15_io_outs_1; // @[MemPrimitives.scala 121:29:@10456.4]
  wire  StickySelects_15_io_outs_2; // @[MemPrimitives.scala 121:29:@10456.4]
  wire  StickySelects_15_io_outs_3; // @[MemPrimitives.scala 121:29:@10456.4]
  wire  StickySelects_15_io_outs_4; // @[MemPrimitives.scala 121:29:@10456.4]
  wire  StickySelects_15_io_outs_5; // @[MemPrimitives.scala 121:29:@10456.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@10519.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@10519.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@10519.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@10519.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@10519.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@10527.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@10527.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@10527.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@10527.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@10527.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@10535.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@10535.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@10535.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@10535.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@10535.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@10543.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@10543.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@10543.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@10543.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@10543.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@10551.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@10551.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@10551.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@10551.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@10551.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@10559.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@10559.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@10559.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@10559.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@10559.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@10567.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@10567.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@10567.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@10567.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@10567.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@10575.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@10575.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@10575.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@10575.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@10575.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@10615.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@10615.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@10615.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@10615.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@10615.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@10623.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@10623.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@10623.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@10623.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@10623.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@10631.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@10631.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@10631.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@10631.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@10631.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@10639.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@10639.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@10639.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@10639.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@10639.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@10647.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@10647.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@10647.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@10647.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@10647.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@10655.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@10655.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@10655.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@10655.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@10655.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@10663.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@10663.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@10663.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@10663.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@10663.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@10671.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@10671.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@10671.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@10671.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@10671.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@10711.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@10711.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@10711.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@10711.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@10711.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@10719.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@10719.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@10719.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@10719.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@10719.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@10727.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@10727.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@10727.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@10727.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@10727.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@10735.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@10735.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@10735.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@10735.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@10735.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@10743.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@10743.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@10743.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@10743.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@10743.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@10751.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@10751.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@10751.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@10751.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@10751.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@10759.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@10759.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@10759.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@10759.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@10759.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@10767.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@10767.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@10767.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@10767.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@10767.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@10807.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@10807.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@10807.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@10807.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@10807.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@10815.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@10815.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@10815.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@10815.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@10815.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@10823.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@10823.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@10823.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@10823.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@10823.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@10831.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@10831.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@10831.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@10831.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@10831.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@10839.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@10839.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@10839.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@10839.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@10839.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@10847.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@10847.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@10847.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@10847.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@10847.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@10855.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@10855.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@10855.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@10855.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@10855.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@10863.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@10863.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@10863.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@10863.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@10863.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@10903.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@10903.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@10903.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@10903.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@10903.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@10911.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@10911.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@10911.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@10911.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@10911.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@10919.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@10919.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@10919.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@10919.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@10919.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@10927.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@10927.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@10927.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@10927.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@10927.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@10935.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@10935.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@10935.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@10935.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@10935.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@10943.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@10943.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@10943.4]
  wire  RetimeWrapper_37_io_in; // @[package.scala 93:22:@10943.4]
  wire  RetimeWrapper_37_io_out; // @[package.scala 93:22:@10943.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@10951.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@10951.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@10951.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@10951.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@10951.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@10959.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@10959.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@10959.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@10959.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@10959.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@10999.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@10999.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@10999.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@10999.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@10999.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@11007.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@11007.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@11007.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@11007.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@11007.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@11015.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@11015.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@11015.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@11015.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@11015.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@11023.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@11023.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@11023.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@11023.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@11023.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@11031.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@11031.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@11031.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@11031.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@11031.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@11039.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@11039.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@11039.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@11039.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@11039.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@11047.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@11047.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@11047.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@11047.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@11047.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@11055.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@11055.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@11055.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@11055.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@11055.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@11095.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@11095.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@11095.4]
  wire  RetimeWrapper_48_io_in; // @[package.scala 93:22:@11095.4]
  wire  RetimeWrapper_48_io_out; // @[package.scala 93:22:@11095.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@11103.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@11103.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@11103.4]
  wire  RetimeWrapper_49_io_in; // @[package.scala 93:22:@11103.4]
  wire  RetimeWrapper_49_io_out; // @[package.scala 93:22:@11103.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@11111.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@11111.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@11111.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@11111.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@11111.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@11119.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@11119.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@11119.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@11119.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@11119.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@11127.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@11127.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@11127.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@11127.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@11127.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@11135.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@11135.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@11135.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@11135.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@11135.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@11143.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@11143.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@11143.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@11143.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@11143.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@11151.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@11151.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@11151.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@11151.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@11151.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@11191.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@11191.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@11191.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@11191.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@11191.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@11199.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@11199.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@11199.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@11199.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@11199.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@11207.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@11207.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@11207.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@11207.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@11207.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@11215.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@11215.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@11215.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@11215.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@11215.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@11223.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@11223.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@11223.4]
  wire  RetimeWrapper_60_io_in; // @[package.scala 93:22:@11223.4]
  wire  RetimeWrapper_60_io_out; // @[package.scala 93:22:@11223.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@11231.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@11231.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@11231.4]
  wire  RetimeWrapper_61_io_in; // @[package.scala 93:22:@11231.4]
  wire  RetimeWrapper_61_io_out; // @[package.scala 93:22:@11231.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@11239.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@11239.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@11239.4]
  wire  RetimeWrapper_62_io_in; // @[package.scala 93:22:@11239.4]
  wire  RetimeWrapper_62_io_out; // @[package.scala 93:22:@11239.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@11247.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@11247.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@11247.4]
  wire  RetimeWrapper_63_io_in; // @[package.scala 93:22:@11247.4]
  wire  RetimeWrapper_63_io_out; // @[package.scala 93:22:@11247.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@11287.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@11287.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@11287.4]
  wire  RetimeWrapper_64_io_in; // @[package.scala 93:22:@11287.4]
  wire  RetimeWrapper_64_io_out; // @[package.scala 93:22:@11287.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@11295.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@11295.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@11295.4]
  wire  RetimeWrapper_65_io_in; // @[package.scala 93:22:@11295.4]
  wire  RetimeWrapper_65_io_out; // @[package.scala 93:22:@11295.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@11303.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@11303.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@11303.4]
  wire  RetimeWrapper_66_io_in; // @[package.scala 93:22:@11303.4]
  wire  RetimeWrapper_66_io_out; // @[package.scala 93:22:@11303.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@11311.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@11311.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@11311.4]
  wire  RetimeWrapper_67_io_in; // @[package.scala 93:22:@11311.4]
  wire  RetimeWrapper_67_io_out; // @[package.scala 93:22:@11311.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@11319.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@11319.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@11319.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@11319.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@11319.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@11327.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@11327.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@11327.4]
  wire  RetimeWrapper_69_io_in; // @[package.scala 93:22:@11327.4]
  wire  RetimeWrapper_69_io_out; // @[package.scala 93:22:@11327.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@11335.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@11335.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@11335.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@11335.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@11335.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@11343.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@11343.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@11343.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@11343.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@11343.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@11383.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@11383.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@11383.4]
  wire  RetimeWrapper_72_io_in; // @[package.scala 93:22:@11383.4]
  wire  RetimeWrapper_72_io_out; // @[package.scala 93:22:@11383.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@11391.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@11391.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@11391.4]
  wire  RetimeWrapper_73_io_in; // @[package.scala 93:22:@11391.4]
  wire  RetimeWrapper_73_io_out; // @[package.scala 93:22:@11391.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@11399.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@11399.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@11399.4]
  wire  RetimeWrapper_74_io_in; // @[package.scala 93:22:@11399.4]
  wire  RetimeWrapper_74_io_out; // @[package.scala 93:22:@11399.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@11407.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@11407.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@11407.4]
  wire  RetimeWrapper_75_io_in; // @[package.scala 93:22:@11407.4]
  wire  RetimeWrapper_75_io_out; // @[package.scala 93:22:@11407.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@11415.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@11415.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@11415.4]
  wire  RetimeWrapper_76_io_in; // @[package.scala 93:22:@11415.4]
  wire  RetimeWrapper_76_io_out; // @[package.scala 93:22:@11415.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@11423.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@11423.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@11423.4]
  wire  RetimeWrapper_77_io_in; // @[package.scala 93:22:@11423.4]
  wire  RetimeWrapper_77_io_out; // @[package.scala 93:22:@11423.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@11431.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@11431.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@11431.4]
  wire  RetimeWrapper_78_io_in; // @[package.scala 93:22:@11431.4]
  wire  RetimeWrapper_78_io_out; // @[package.scala 93:22:@11431.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@11439.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@11439.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@11439.4]
  wire  RetimeWrapper_79_io_in; // @[package.scala 93:22:@11439.4]
  wire  RetimeWrapper_79_io_out; // @[package.scala 93:22:@11439.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@11479.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@11479.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@11479.4]
  wire  RetimeWrapper_80_io_in; // @[package.scala 93:22:@11479.4]
  wire  RetimeWrapper_80_io_out; // @[package.scala 93:22:@11479.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@11487.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@11487.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@11487.4]
  wire  RetimeWrapper_81_io_in; // @[package.scala 93:22:@11487.4]
  wire  RetimeWrapper_81_io_out; // @[package.scala 93:22:@11487.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@11495.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@11495.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@11495.4]
  wire  RetimeWrapper_82_io_in; // @[package.scala 93:22:@11495.4]
  wire  RetimeWrapper_82_io_out; // @[package.scala 93:22:@11495.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@11503.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@11503.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@11503.4]
  wire  RetimeWrapper_83_io_in; // @[package.scala 93:22:@11503.4]
  wire  RetimeWrapper_83_io_out; // @[package.scala 93:22:@11503.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@11511.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@11511.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@11511.4]
  wire  RetimeWrapper_84_io_in; // @[package.scala 93:22:@11511.4]
  wire  RetimeWrapper_84_io_out; // @[package.scala 93:22:@11511.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@11519.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@11519.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@11519.4]
  wire  RetimeWrapper_85_io_in; // @[package.scala 93:22:@11519.4]
  wire  RetimeWrapper_85_io_out; // @[package.scala 93:22:@11519.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@11527.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@11527.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@11527.4]
  wire  RetimeWrapper_86_io_in; // @[package.scala 93:22:@11527.4]
  wire  RetimeWrapper_86_io_out; // @[package.scala 93:22:@11527.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@11535.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@11535.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@11535.4]
  wire  RetimeWrapper_87_io_in; // @[package.scala 93:22:@11535.4]
  wire  RetimeWrapper_87_io_out; // @[package.scala 93:22:@11535.4]
  wire  RetimeWrapper_88_clock; // @[package.scala 93:22:@11575.4]
  wire  RetimeWrapper_88_reset; // @[package.scala 93:22:@11575.4]
  wire  RetimeWrapper_88_io_flow; // @[package.scala 93:22:@11575.4]
  wire  RetimeWrapper_88_io_in; // @[package.scala 93:22:@11575.4]
  wire  RetimeWrapper_88_io_out; // @[package.scala 93:22:@11575.4]
  wire  RetimeWrapper_89_clock; // @[package.scala 93:22:@11583.4]
  wire  RetimeWrapper_89_reset; // @[package.scala 93:22:@11583.4]
  wire  RetimeWrapper_89_io_flow; // @[package.scala 93:22:@11583.4]
  wire  RetimeWrapper_89_io_in; // @[package.scala 93:22:@11583.4]
  wire  RetimeWrapper_89_io_out; // @[package.scala 93:22:@11583.4]
  wire  RetimeWrapper_90_clock; // @[package.scala 93:22:@11591.4]
  wire  RetimeWrapper_90_reset; // @[package.scala 93:22:@11591.4]
  wire  RetimeWrapper_90_io_flow; // @[package.scala 93:22:@11591.4]
  wire  RetimeWrapper_90_io_in; // @[package.scala 93:22:@11591.4]
  wire  RetimeWrapper_90_io_out; // @[package.scala 93:22:@11591.4]
  wire  RetimeWrapper_91_clock; // @[package.scala 93:22:@11599.4]
  wire  RetimeWrapper_91_reset; // @[package.scala 93:22:@11599.4]
  wire  RetimeWrapper_91_io_flow; // @[package.scala 93:22:@11599.4]
  wire  RetimeWrapper_91_io_in; // @[package.scala 93:22:@11599.4]
  wire  RetimeWrapper_91_io_out; // @[package.scala 93:22:@11599.4]
  wire  RetimeWrapper_92_clock; // @[package.scala 93:22:@11607.4]
  wire  RetimeWrapper_92_reset; // @[package.scala 93:22:@11607.4]
  wire  RetimeWrapper_92_io_flow; // @[package.scala 93:22:@11607.4]
  wire  RetimeWrapper_92_io_in; // @[package.scala 93:22:@11607.4]
  wire  RetimeWrapper_92_io_out; // @[package.scala 93:22:@11607.4]
  wire  RetimeWrapper_93_clock; // @[package.scala 93:22:@11615.4]
  wire  RetimeWrapper_93_reset; // @[package.scala 93:22:@11615.4]
  wire  RetimeWrapper_93_io_flow; // @[package.scala 93:22:@11615.4]
  wire  RetimeWrapper_93_io_in; // @[package.scala 93:22:@11615.4]
  wire  RetimeWrapper_93_io_out; // @[package.scala 93:22:@11615.4]
  wire  RetimeWrapper_94_clock; // @[package.scala 93:22:@11623.4]
  wire  RetimeWrapper_94_reset; // @[package.scala 93:22:@11623.4]
  wire  RetimeWrapper_94_io_flow; // @[package.scala 93:22:@11623.4]
  wire  RetimeWrapper_94_io_in; // @[package.scala 93:22:@11623.4]
  wire  RetimeWrapper_94_io_out; // @[package.scala 93:22:@11623.4]
  wire  RetimeWrapper_95_clock; // @[package.scala 93:22:@11631.4]
  wire  RetimeWrapper_95_reset; // @[package.scala 93:22:@11631.4]
  wire  RetimeWrapper_95_io_flow; // @[package.scala 93:22:@11631.4]
  wire  RetimeWrapper_95_io_in; // @[package.scala 93:22:@11631.4]
  wire  RetimeWrapper_95_io_out; // @[package.scala 93:22:@11631.4]
  wire  _T_444; // @[MemPrimitives.scala 82:210:@9310.4]
  wire  _T_446; // @[MemPrimitives.scala 82:210:@9311.4]
  wire  _T_447; // @[MemPrimitives.scala 82:228:@9312.4]
  wire  _T_448; // @[MemPrimitives.scala 83:102:@9313.4]
  wire [9:0] _T_450; // @[Cat.scala 30:58:@9315.4]
  wire  _T_455; // @[MemPrimitives.scala 82:210:@9322.4]
  wire  _T_457; // @[MemPrimitives.scala 82:210:@9323.4]
  wire  _T_458; // @[MemPrimitives.scala 82:228:@9324.4]
  wire  _T_459; // @[MemPrimitives.scala 83:102:@9325.4]
  wire [9:0] _T_461; // @[Cat.scala 30:58:@9327.4]
  wire  _T_468; // @[MemPrimitives.scala 82:210:@9335.4]
  wire  _T_469; // @[MemPrimitives.scala 82:228:@9336.4]
  wire  _T_470; // @[MemPrimitives.scala 83:102:@9337.4]
  wire [9:0] _T_472; // @[Cat.scala 30:58:@9339.4]
  wire  _T_479; // @[MemPrimitives.scala 82:210:@9347.4]
  wire  _T_480; // @[MemPrimitives.scala 82:228:@9348.4]
  wire  _T_481; // @[MemPrimitives.scala 83:102:@9349.4]
  wire [9:0] _T_483; // @[Cat.scala 30:58:@9351.4]
  wire  _T_488; // @[MemPrimitives.scala 82:210:@9358.4]
  wire  _T_491; // @[MemPrimitives.scala 82:228:@9360.4]
  wire  _T_492; // @[MemPrimitives.scala 83:102:@9361.4]
  wire [9:0] _T_494; // @[Cat.scala 30:58:@9363.4]
  wire  _T_499; // @[MemPrimitives.scala 82:210:@9370.4]
  wire  _T_502; // @[MemPrimitives.scala 82:228:@9372.4]
  wire  _T_503; // @[MemPrimitives.scala 83:102:@9373.4]
  wire [9:0] _T_505; // @[Cat.scala 30:58:@9375.4]
  wire  _T_513; // @[MemPrimitives.scala 82:228:@9384.4]
  wire  _T_514; // @[MemPrimitives.scala 83:102:@9385.4]
  wire [9:0] _T_516; // @[Cat.scala 30:58:@9387.4]
  wire  _T_524; // @[MemPrimitives.scala 82:228:@9396.4]
  wire  _T_525; // @[MemPrimitives.scala 83:102:@9397.4]
  wire [9:0] _T_527; // @[Cat.scala 30:58:@9399.4]
  wire  _T_532; // @[MemPrimitives.scala 82:210:@9406.4]
  wire  _T_535; // @[MemPrimitives.scala 82:228:@9408.4]
  wire  _T_536; // @[MemPrimitives.scala 83:102:@9409.4]
  wire [9:0] _T_538; // @[Cat.scala 30:58:@9411.4]
  wire  _T_543; // @[MemPrimitives.scala 82:210:@9418.4]
  wire  _T_546; // @[MemPrimitives.scala 82:228:@9420.4]
  wire  _T_547; // @[MemPrimitives.scala 83:102:@9421.4]
  wire [9:0] _T_549; // @[Cat.scala 30:58:@9423.4]
  wire  _T_557; // @[MemPrimitives.scala 82:228:@9432.4]
  wire  _T_558; // @[MemPrimitives.scala 83:102:@9433.4]
  wire [9:0] _T_560; // @[Cat.scala 30:58:@9435.4]
  wire  _T_568; // @[MemPrimitives.scala 82:228:@9444.4]
  wire  _T_569; // @[MemPrimitives.scala 83:102:@9445.4]
  wire [9:0] _T_571; // @[Cat.scala 30:58:@9447.4]
  wire  _T_576; // @[MemPrimitives.scala 82:210:@9454.4]
  wire  _T_579; // @[MemPrimitives.scala 82:228:@9456.4]
  wire  _T_580; // @[MemPrimitives.scala 83:102:@9457.4]
  wire [9:0] _T_582; // @[Cat.scala 30:58:@9459.4]
  wire  _T_587; // @[MemPrimitives.scala 82:210:@9466.4]
  wire  _T_590; // @[MemPrimitives.scala 82:228:@9468.4]
  wire  _T_591; // @[MemPrimitives.scala 83:102:@9469.4]
  wire [9:0] _T_593; // @[Cat.scala 30:58:@9471.4]
  wire  _T_601; // @[MemPrimitives.scala 82:228:@9480.4]
  wire  _T_602; // @[MemPrimitives.scala 83:102:@9481.4]
  wire [9:0] _T_604; // @[Cat.scala 30:58:@9483.4]
  wire  _T_612; // @[MemPrimitives.scala 82:228:@9492.4]
  wire  _T_613; // @[MemPrimitives.scala 83:102:@9493.4]
  wire [9:0] _T_615; // @[Cat.scala 30:58:@9495.4]
  wire  _T_620; // @[MemPrimitives.scala 110:210:@9502.4]
  wire  _T_622; // @[MemPrimitives.scala 110:210:@9503.4]
  wire  _T_623; // @[MemPrimitives.scala 110:228:@9504.4]
  wire  _T_626; // @[MemPrimitives.scala 110:210:@9506.4]
  wire  _T_628; // @[MemPrimitives.scala 110:210:@9507.4]
  wire  _T_629; // @[MemPrimitives.scala 110:228:@9508.4]
  wire  _T_632; // @[MemPrimitives.scala 110:210:@9510.4]
  wire  _T_634; // @[MemPrimitives.scala 110:210:@9511.4]
  wire  _T_635; // @[MemPrimitives.scala 110:228:@9512.4]
  wire  _T_638; // @[MemPrimitives.scala 110:210:@9514.4]
  wire  _T_640; // @[MemPrimitives.scala 110:210:@9515.4]
  wire  _T_641; // @[MemPrimitives.scala 110:228:@9516.4]
  wire  _T_644; // @[MemPrimitives.scala 110:210:@9518.4]
  wire  _T_646; // @[MemPrimitives.scala 110:210:@9519.4]
  wire  _T_647; // @[MemPrimitives.scala 110:228:@9520.4]
  wire  _T_650; // @[MemPrimitives.scala 110:210:@9522.4]
  wire  _T_652; // @[MemPrimitives.scala 110:210:@9523.4]
  wire  _T_653; // @[MemPrimitives.scala 110:228:@9524.4]
  wire  _T_655; // @[MemPrimitives.scala 123:41:@9535.4]
  wire  _T_656; // @[MemPrimitives.scala 123:41:@9536.4]
  wire  _T_657; // @[MemPrimitives.scala 123:41:@9537.4]
  wire  _T_658; // @[MemPrimitives.scala 123:41:@9538.4]
  wire  _T_659; // @[MemPrimitives.scala 123:41:@9539.4]
  wire  _T_660; // @[MemPrimitives.scala 123:41:@9540.4]
  wire [2:0] _T_662; // @[Cat.scala 30:58:@9542.4]
  wire [2:0] _T_664; // @[Cat.scala 30:58:@9544.4]
  wire [2:0] _T_666; // @[Cat.scala 30:58:@9546.4]
  wire [2:0] _T_668; // @[Cat.scala 30:58:@9548.4]
  wire [2:0] _T_670; // @[Cat.scala 30:58:@9550.4]
  wire [2:0] _T_672; // @[Cat.scala 30:58:@9552.4]
  wire [2:0] _T_673; // @[Mux.scala 31:69:@9553.4]
  wire [2:0] _T_674; // @[Mux.scala 31:69:@9554.4]
  wire [2:0] _T_675; // @[Mux.scala 31:69:@9555.4]
  wire [2:0] _T_676; // @[Mux.scala 31:69:@9556.4]
  wire [2:0] _T_677; // @[Mux.scala 31:69:@9557.4]
  wire  _T_682; // @[MemPrimitives.scala 110:210:@9564.4]
  wire  _T_684; // @[MemPrimitives.scala 110:210:@9565.4]
  wire  _T_685; // @[MemPrimitives.scala 110:228:@9566.4]
  wire  _T_688; // @[MemPrimitives.scala 110:210:@9568.4]
  wire  _T_690; // @[MemPrimitives.scala 110:210:@9569.4]
  wire  _T_691; // @[MemPrimitives.scala 110:228:@9570.4]
  wire  _T_694; // @[MemPrimitives.scala 110:210:@9572.4]
  wire  _T_696; // @[MemPrimitives.scala 110:210:@9573.4]
  wire  _T_697; // @[MemPrimitives.scala 110:228:@9574.4]
  wire  _T_700; // @[MemPrimitives.scala 110:210:@9576.4]
  wire  _T_702; // @[MemPrimitives.scala 110:210:@9577.4]
  wire  _T_703; // @[MemPrimitives.scala 110:228:@9578.4]
  wire  _T_706; // @[MemPrimitives.scala 110:210:@9580.4]
  wire  _T_708; // @[MemPrimitives.scala 110:210:@9581.4]
  wire  _T_709; // @[MemPrimitives.scala 110:228:@9582.4]
  wire  _T_712; // @[MemPrimitives.scala 110:210:@9584.4]
  wire  _T_714; // @[MemPrimitives.scala 110:210:@9585.4]
  wire  _T_715; // @[MemPrimitives.scala 110:228:@9586.4]
  wire  _T_717; // @[MemPrimitives.scala 123:41:@9597.4]
  wire  _T_718; // @[MemPrimitives.scala 123:41:@9598.4]
  wire  _T_719; // @[MemPrimitives.scala 123:41:@9599.4]
  wire  _T_720; // @[MemPrimitives.scala 123:41:@9600.4]
  wire  _T_721; // @[MemPrimitives.scala 123:41:@9601.4]
  wire  _T_722; // @[MemPrimitives.scala 123:41:@9602.4]
  wire [2:0] _T_724; // @[Cat.scala 30:58:@9604.4]
  wire [2:0] _T_726; // @[Cat.scala 30:58:@9606.4]
  wire [2:0] _T_728; // @[Cat.scala 30:58:@9608.4]
  wire [2:0] _T_730; // @[Cat.scala 30:58:@9610.4]
  wire [2:0] _T_732; // @[Cat.scala 30:58:@9612.4]
  wire [2:0] _T_734; // @[Cat.scala 30:58:@9614.4]
  wire [2:0] _T_735; // @[Mux.scala 31:69:@9615.4]
  wire [2:0] _T_736; // @[Mux.scala 31:69:@9616.4]
  wire [2:0] _T_737; // @[Mux.scala 31:69:@9617.4]
  wire [2:0] _T_738; // @[Mux.scala 31:69:@9618.4]
  wire [2:0] _T_739; // @[Mux.scala 31:69:@9619.4]
  wire  _T_746; // @[MemPrimitives.scala 110:210:@9627.4]
  wire  _T_747; // @[MemPrimitives.scala 110:228:@9628.4]
  wire  _T_752; // @[MemPrimitives.scala 110:210:@9631.4]
  wire  _T_753; // @[MemPrimitives.scala 110:228:@9632.4]
  wire  _T_758; // @[MemPrimitives.scala 110:210:@9635.4]
  wire  _T_759; // @[MemPrimitives.scala 110:228:@9636.4]
  wire  _T_764; // @[MemPrimitives.scala 110:210:@9639.4]
  wire  _T_765; // @[MemPrimitives.scala 110:228:@9640.4]
  wire  _T_770; // @[MemPrimitives.scala 110:210:@9643.4]
  wire  _T_771; // @[MemPrimitives.scala 110:228:@9644.4]
  wire  _T_776; // @[MemPrimitives.scala 110:210:@9647.4]
  wire  _T_777; // @[MemPrimitives.scala 110:228:@9648.4]
  wire  _T_779; // @[MemPrimitives.scala 123:41:@9659.4]
  wire  _T_780; // @[MemPrimitives.scala 123:41:@9660.4]
  wire  _T_781; // @[MemPrimitives.scala 123:41:@9661.4]
  wire  _T_782; // @[MemPrimitives.scala 123:41:@9662.4]
  wire  _T_783; // @[MemPrimitives.scala 123:41:@9663.4]
  wire  _T_784; // @[MemPrimitives.scala 123:41:@9664.4]
  wire [2:0] _T_786; // @[Cat.scala 30:58:@9666.4]
  wire [2:0] _T_788; // @[Cat.scala 30:58:@9668.4]
  wire [2:0] _T_790; // @[Cat.scala 30:58:@9670.4]
  wire [2:0] _T_792; // @[Cat.scala 30:58:@9672.4]
  wire [2:0] _T_794; // @[Cat.scala 30:58:@9674.4]
  wire [2:0] _T_796; // @[Cat.scala 30:58:@9676.4]
  wire [2:0] _T_797; // @[Mux.scala 31:69:@9677.4]
  wire [2:0] _T_798; // @[Mux.scala 31:69:@9678.4]
  wire [2:0] _T_799; // @[Mux.scala 31:69:@9679.4]
  wire [2:0] _T_800; // @[Mux.scala 31:69:@9680.4]
  wire [2:0] _T_801; // @[Mux.scala 31:69:@9681.4]
  wire  _T_808; // @[MemPrimitives.scala 110:210:@9689.4]
  wire  _T_809; // @[MemPrimitives.scala 110:228:@9690.4]
  wire  _T_814; // @[MemPrimitives.scala 110:210:@9693.4]
  wire  _T_815; // @[MemPrimitives.scala 110:228:@9694.4]
  wire  _T_820; // @[MemPrimitives.scala 110:210:@9697.4]
  wire  _T_821; // @[MemPrimitives.scala 110:228:@9698.4]
  wire  _T_826; // @[MemPrimitives.scala 110:210:@9701.4]
  wire  _T_827; // @[MemPrimitives.scala 110:228:@9702.4]
  wire  _T_832; // @[MemPrimitives.scala 110:210:@9705.4]
  wire  _T_833; // @[MemPrimitives.scala 110:228:@9706.4]
  wire  _T_838; // @[MemPrimitives.scala 110:210:@9709.4]
  wire  _T_839; // @[MemPrimitives.scala 110:228:@9710.4]
  wire  _T_841; // @[MemPrimitives.scala 123:41:@9721.4]
  wire  _T_842; // @[MemPrimitives.scala 123:41:@9722.4]
  wire  _T_843; // @[MemPrimitives.scala 123:41:@9723.4]
  wire  _T_844; // @[MemPrimitives.scala 123:41:@9724.4]
  wire  _T_845; // @[MemPrimitives.scala 123:41:@9725.4]
  wire  _T_846; // @[MemPrimitives.scala 123:41:@9726.4]
  wire [2:0] _T_848; // @[Cat.scala 30:58:@9728.4]
  wire [2:0] _T_850; // @[Cat.scala 30:58:@9730.4]
  wire [2:0] _T_852; // @[Cat.scala 30:58:@9732.4]
  wire [2:0] _T_854; // @[Cat.scala 30:58:@9734.4]
  wire [2:0] _T_856; // @[Cat.scala 30:58:@9736.4]
  wire [2:0] _T_858; // @[Cat.scala 30:58:@9738.4]
  wire [2:0] _T_859; // @[Mux.scala 31:69:@9739.4]
  wire [2:0] _T_860; // @[Mux.scala 31:69:@9740.4]
  wire [2:0] _T_861; // @[Mux.scala 31:69:@9741.4]
  wire [2:0] _T_862; // @[Mux.scala 31:69:@9742.4]
  wire [2:0] _T_863; // @[Mux.scala 31:69:@9743.4]
  wire  _T_868; // @[MemPrimitives.scala 110:210:@9750.4]
  wire  _T_871; // @[MemPrimitives.scala 110:228:@9752.4]
  wire  _T_874; // @[MemPrimitives.scala 110:210:@9754.4]
  wire  _T_877; // @[MemPrimitives.scala 110:228:@9756.4]
  wire  _T_880; // @[MemPrimitives.scala 110:210:@9758.4]
  wire  _T_883; // @[MemPrimitives.scala 110:228:@9760.4]
  wire  _T_886; // @[MemPrimitives.scala 110:210:@9762.4]
  wire  _T_889; // @[MemPrimitives.scala 110:228:@9764.4]
  wire  _T_892; // @[MemPrimitives.scala 110:210:@9766.4]
  wire  _T_895; // @[MemPrimitives.scala 110:228:@9768.4]
  wire  _T_898; // @[MemPrimitives.scala 110:210:@9770.4]
  wire  _T_901; // @[MemPrimitives.scala 110:228:@9772.4]
  wire  _T_903; // @[MemPrimitives.scala 123:41:@9783.4]
  wire  _T_904; // @[MemPrimitives.scala 123:41:@9784.4]
  wire  _T_905; // @[MemPrimitives.scala 123:41:@9785.4]
  wire  _T_906; // @[MemPrimitives.scala 123:41:@9786.4]
  wire  _T_907; // @[MemPrimitives.scala 123:41:@9787.4]
  wire  _T_908; // @[MemPrimitives.scala 123:41:@9788.4]
  wire [2:0] _T_910; // @[Cat.scala 30:58:@9790.4]
  wire [2:0] _T_912; // @[Cat.scala 30:58:@9792.4]
  wire [2:0] _T_914; // @[Cat.scala 30:58:@9794.4]
  wire [2:0] _T_916; // @[Cat.scala 30:58:@9796.4]
  wire [2:0] _T_918; // @[Cat.scala 30:58:@9798.4]
  wire [2:0] _T_920; // @[Cat.scala 30:58:@9800.4]
  wire [2:0] _T_921; // @[Mux.scala 31:69:@9801.4]
  wire [2:0] _T_922; // @[Mux.scala 31:69:@9802.4]
  wire [2:0] _T_923; // @[Mux.scala 31:69:@9803.4]
  wire [2:0] _T_924; // @[Mux.scala 31:69:@9804.4]
  wire [2:0] _T_925; // @[Mux.scala 31:69:@9805.4]
  wire  _T_930; // @[MemPrimitives.scala 110:210:@9812.4]
  wire  _T_933; // @[MemPrimitives.scala 110:228:@9814.4]
  wire  _T_936; // @[MemPrimitives.scala 110:210:@9816.4]
  wire  _T_939; // @[MemPrimitives.scala 110:228:@9818.4]
  wire  _T_942; // @[MemPrimitives.scala 110:210:@9820.4]
  wire  _T_945; // @[MemPrimitives.scala 110:228:@9822.4]
  wire  _T_948; // @[MemPrimitives.scala 110:210:@9824.4]
  wire  _T_951; // @[MemPrimitives.scala 110:228:@9826.4]
  wire  _T_954; // @[MemPrimitives.scala 110:210:@9828.4]
  wire  _T_957; // @[MemPrimitives.scala 110:228:@9830.4]
  wire  _T_960; // @[MemPrimitives.scala 110:210:@9832.4]
  wire  _T_963; // @[MemPrimitives.scala 110:228:@9834.4]
  wire  _T_965; // @[MemPrimitives.scala 123:41:@9845.4]
  wire  _T_966; // @[MemPrimitives.scala 123:41:@9846.4]
  wire  _T_967; // @[MemPrimitives.scala 123:41:@9847.4]
  wire  _T_968; // @[MemPrimitives.scala 123:41:@9848.4]
  wire  _T_969; // @[MemPrimitives.scala 123:41:@9849.4]
  wire  _T_970; // @[MemPrimitives.scala 123:41:@9850.4]
  wire [2:0] _T_972; // @[Cat.scala 30:58:@9852.4]
  wire [2:0] _T_974; // @[Cat.scala 30:58:@9854.4]
  wire [2:0] _T_976; // @[Cat.scala 30:58:@9856.4]
  wire [2:0] _T_978; // @[Cat.scala 30:58:@9858.4]
  wire [2:0] _T_980; // @[Cat.scala 30:58:@9860.4]
  wire [2:0] _T_982; // @[Cat.scala 30:58:@9862.4]
  wire [2:0] _T_983; // @[Mux.scala 31:69:@9863.4]
  wire [2:0] _T_984; // @[Mux.scala 31:69:@9864.4]
  wire [2:0] _T_985; // @[Mux.scala 31:69:@9865.4]
  wire [2:0] _T_986; // @[Mux.scala 31:69:@9866.4]
  wire [2:0] _T_987; // @[Mux.scala 31:69:@9867.4]
  wire  _T_995; // @[MemPrimitives.scala 110:228:@9876.4]
  wire  _T_1001; // @[MemPrimitives.scala 110:228:@9880.4]
  wire  _T_1007; // @[MemPrimitives.scala 110:228:@9884.4]
  wire  _T_1013; // @[MemPrimitives.scala 110:228:@9888.4]
  wire  _T_1019; // @[MemPrimitives.scala 110:228:@9892.4]
  wire  _T_1025; // @[MemPrimitives.scala 110:228:@9896.4]
  wire  _T_1027; // @[MemPrimitives.scala 123:41:@9907.4]
  wire  _T_1028; // @[MemPrimitives.scala 123:41:@9908.4]
  wire  _T_1029; // @[MemPrimitives.scala 123:41:@9909.4]
  wire  _T_1030; // @[MemPrimitives.scala 123:41:@9910.4]
  wire  _T_1031; // @[MemPrimitives.scala 123:41:@9911.4]
  wire  _T_1032; // @[MemPrimitives.scala 123:41:@9912.4]
  wire [2:0] _T_1034; // @[Cat.scala 30:58:@9914.4]
  wire [2:0] _T_1036; // @[Cat.scala 30:58:@9916.4]
  wire [2:0] _T_1038; // @[Cat.scala 30:58:@9918.4]
  wire [2:0] _T_1040; // @[Cat.scala 30:58:@9920.4]
  wire [2:0] _T_1042; // @[Cat.scala 30:58:@9922.4]
  wire [2:0] _T_1044; // @[Cat.scala 30:58:@9924.4]
  wire [2:0] _T_1045; // @[Mux.scala 31:69:@9925.4]
  wire [2:0] _T_1046; // @[Mux.scala 31:69:@9926.4]
  wire [2:0] _T_1047; // @[Mux.scala 31:69:@9927.4]
  wire [2:0] _T_1048; // @[Mux.scala 31:69:@9928.4]
  wire [2:0] _T_1049; // @[Mux.scala 31:69:@9929.4]
  wire  _T_1057; // @[MemPrimitives.scala 110:228:@9938.4]
  wire  _T_1063; // @[MemPrimitives.scala 110:228:@9942.4]
  wire  _T_1069; // @[MemPrimitives.scala 110:228:@9946.4]
  wire  _T_1075; // @[MemPrimitives.scala 110:228:@9950.4]
  wire  _T_1081; // @[MemPrimitives.scala 110:228:@9954.4]
  wire  _T_1087; // @[MemPrimitives.scala 110:228:@9958.4]
  wire  _T_1089; // @[MemPrimitives.scala 123:41:@9969.4]
  wire  _T_1090; // @[MemPrimitives.scala 123:41:@9970.4]
  wire  _T_1091; // @[MemPrimitives.scala 123:41:@9971.4]
  wire  _T_1092; // @[MemPrimitives.scala 123:41:@9972.4]
  wire  _T_1093; // @[MemPrimitives.scala 123:41:@9973.4]
  wire  _T_1094; // @[MemPrimitives.scala 123:41:@9974.4]
  wire [2:0] _T_1096; // @[Cat.scala 30:58:@9976.4]
  wire [2:0] _T_1098; // @[Cat.scala 30:58:@9978.4]
  wire [2:0] _T_1100; // @[Cat.scala 30:58:@9980.4]
  wire [2:0] _T_1102; // @[Cat.scala 30:58:@9982.4]
  wire [2:0] _T_1104; // @[Cat.scala 30:58:@9984.4]
  wire [2:0] _T_1106; // @[Cat.scala 30:58:@9986.4]
  wire [2:0] _T_1107; // @[Mux.scala 31:69:@9987.4]
  wire [2:0] _T_1108; // @[Mux.scala 31:69:@9988.4]
  wire [2:0] _T_1109; // @[Mux.scala 31:69:@9989.4]
  wire [2:0] _T_1110; // @[Mux.scala 31:69:@9990.4]
  wire [2:0] _T_1111; // @[Mux.scala 31:69:@9991.4]
  wire  _T_1116; // @[MemPrimitives.scala 110:210:@9998.4]
  wire  _T_1119; // @[MemPrimitives.scala 110:228:@10000.4]
  wire  _T_1122; // @[MemPrimitives.scala 110:210:@10002.4]
  wire  _T_1125; // @[MemPrimitives.scala 110:228:@10004.4]
  wire  _T_1128; // @[MemPrimitives.scala 110:210:@10006.4]
  wire  _T_1131; // @[MemPrimitives.scala 110:228:@10008.4]
  wire  _T_1134; // @[MemPrimitives.scala 110:210:@10010.4]
  wire  _T_1137; // @[MemPrimitives.scala 110:228:@10012.4]
  wire  _T_1140; // @[MemPrimitives.scala 110:210:@10014.4]
  wire  _T_1143; // @[MemPrimitives.scala 110:228:@10016.4]
  wire  _T_1146; // @[MemPrimitives.scala 110:210:@10018.4]
  wire  _T_1149; // @[MemPrimitives.scala 110:228:@10020.4]
  wire  _T_1151; // @[MemPrimitives.scala 123:41:@10031.4]
  wire  _T_1152; // @[MemPrimitives.scala 123:41:@10032.4]
  wire  _T_1153; // @[MemPrimitives.scala 123:41:@10033.4]
  wire  _T_1154; // @[MemPrimitives.scala 123:41:@10034.4]
  wire  _T_1155; // @[MemPrimitives.scala 123:41:@10035.4]
  wire  _T_1156; // @[MemPrimitives.scala 123:41:@10036.4]
  wire [2:0] _T_1158; // @[Cat.scala 30:58:@10038.4]
  wire [2:0] _T_1160; // @[Cat.scala 30:58:@10040.4]
  wire [2:0] _T_1162; // @[Cat.scala 30:58:@10042.4]
  wire [2:0] _T_1164; // @[Cat.scala 30:58:@10044.4]
  wire [2:0] _T_1166; // @[Cat.scala 30:58:@10046.4]
  wire [2:0] _T_1168; // @[Cat.scala 30:58:@10048.4]
  wire [2:0] _T_1169; // @[Mux.scala 31:69:@10049.4]
  wire [2:0] _T_1170; // @[Mux.scala 31:69:@10050.4]
  wire [2:0] _T_1171; // @[Mux.scala 31:69:@10051.4]
  wire [2:0] _T_1172; // @[Mux.scala 31:69:@10052.4]
  wire [2:0] _T_1173; // @[Mux.scala 31:69:@10053.4]
  wire  _T_1178; // @[MemPrimitives.scala 110:210:@10060.4]
  wire  _T_1181; // @[MemPrimitives.scala 110:228:@10062.4]
  wire  _T_1184; // @[MemPrimitives.scala 110:210:@10064.4]
  wire  _T_1187; // @[MemPrimitives.scala 110:228:@10066.4]
  wire  _T_1190; // @[MemPrimitives.scala 110:210:@10068.4]
  wire  _T_1193; // @[MemPrimitives.scala 110:228:@10070.4]
  wire  _T_1196; // @[MemPrimitives.scala 110:210:@10072.4]
  wire  _T_1199; // @[MemPrimitives.scala 110:228:@10074.4]
  wire  _T_1202; // @[MemPrimitives.scala 110:210:@10076.4]
  wire  _T_1205; // @[MemPrimitives.scala 110:228:@10078.4]
  wire  _T_1208; // @[MemPrimitives.scala 110:210:@10080.4]
  wire  _T_1211; // @[MemPrimitives.scala 110:228:@10082.4]
  wire  _T_1213; // @[MemPrimitives.scala 123:41:@10093.4]
  wire  _T_1214; // @[MemPrimitives.scala 123:41:@10094.4]
  wire  _T_1215; // @[MemPrimitives.scala 123:41:@10095.4]
  wire  _T_1216; // @[MemPrimitives.scala 123:41:@10096.4]
  wire  _T_1217; // @[MemPrimitives.scala 123:41:@10097.4]
  wire  _T_1218; // @[MemPrimitives.scala 123:41:@10098.4]
  wire [2:0] _T_1220; // @[Cat.scala 30:58:@10100.4]
  wire [2:0] _T_1222; // @[Cat.scala 30:58:@10102.4]
  wire [2:0] _T_1224; // @[Cat.scala 30:58:@10104.4]
  wire [2:0] _T_1226; // @[Cat.scala 30:58:@10106.4]
  wire [2:0] _T_1228; // @[Cat.scala 30:58:@10108.4]
  wire [2:0] _T_1230; // @[Cat.scala 30:58:@10110.4]
  wire [2:0] _T_1231; // @[Mux.scala 31:69:@10111.4]
  wire [2:0] _T_1232; // @[Mux.scala 31:69:@10112.4]
  wire [2:0] _T_1233; // @[Mux.scala 31:69:@10113.4]
  wire [2:0] _T_1234; // @[Mux.scala 31:69:@10114.4]
  wire [2:0] _T_1235; // @[Mux.scala 31:69:@10115.4]
  wire  _T_1243; // @[MemPrimitives.scala 110:228:@10124.4]
  wire  _T_1249; // @[MemPrimitives.scala 110:228:@10128.4]
  wire  _T_1255; // @[MemPrimitives.scala 110:228:@10132.4]
  wire  _T_1261; // @[MemPrimitives.scala 110:228:@10136.4]
  wire  _T_1267; // @[MemPrimitives.scala 110:228:@10140.4]
  wire  _T_1273; // @[MemPrimitives.scala 110:228:@10144.4]
  wire  _T_1275; // @[MemPrimitives.scala 123:41:@10155.4]
  wire  _T_1276; // @[MemPrimitives.scala 123:41:@10156.4]
  wire  _T_1277; // @[MemPrimitives.scala 123:41:@10157.4]
  wire  _T_1278; // @[MemPrimitives.scala 123:41:@10158.4]
  wire  _T_1279; // @[MemPrimitives.scala 123:41:@10159.4]
  wire  _T_1280; // @[MemPrimitives.scala 123:41:@10160.4]
  wire [2:0] _T_1282; // @[Cat.scala 30:58:@10162.4]
  wire [2:0] _T_1284; // @[Cat.scala 30:58:@10164.4]
  wire [2:0] _T_1286; // @[Cat.scala 30:58:@10166.4]
  wire [2:0] _T_1288; // @[Cat.scala 30:58:@10168.4]
  wire [2:0] _T_1290; // @[Cat.scala 30:58:@10170.4]
  wire [2:0] _T_1292; // @[Cat.scala 30:58:@10172.4]
  wire [2:0] _T_1293; // @[Mux.scala 31:69:@10173.4]
  wire [2:0] _T_1294; // @[Mux.scala 31:69:@10174.4]
  wire [2:0] _T_1295; // @[Mux.scala 31:69:@10175.4]
  wire [2:0] _T_1296; // @[Mux.scala 31:69:@10176.4]
  wire [2:0] _T_1297; // @[Mux.scala 31:69:@10177.4]
  wire  _T_1305; // @[MemPrimitives.scala 110:228:@10186.4]
  wire  _T_1311; // @[MemPrimitives.scala 110:228:@10190.4]
  wire  _T_1317; // @[MemPrimitives.scala 110:228:@10194.4]
  wire  _T_1323; // @[MemPrimitives.scala 110:228:@10198.4]
  wire  _T_1329; // @[MemPrimitives.scala 110:228:@10202.4]
  wire  _T_1335; // @[MemPrimitives.scala 110:228:@10206.4]
  wire  _T_1337; // @[MemPrimitives.scala 123:41:@10217.4]
  wire  _T_1338; // @[MemPrimitives.scala 123:41:@10218.4]
  wire  _T_1339; // @[MemPrimitives.scala 123:41:@10219.4]
  wire  _T_1340; // @[MemPrimitives.scala 123:41:@10220.4]
  wire  _T_1341; // @[MemPrimitives.scala 123:41:@10221.4]
  wire  _T_1342; // @[MemPrimitives.scala 123:41:@10222.4]
  wire [2:0] _T_1344; // @[Cat.scala 30:58:@10224.4]
  wire [2:0] _T_1346; // @[Cat.scala 30:58:@10226.4]
  wire [2:0] _T_1348; // @[Cat.scala 30:58:@10228.4]
  wire [2:0] _T_1350; // @[Cat.scala 30:58:@10230.4]
  wire [2:0] _T_1352; // @[Cat.scala 30:58:@10232.4]
  wire [2:0] _T_1354; // @[Cat.scala 30:58:@10234.4]
  wire [2:0] _T_1355; // @[Mux.scala 31:69:@10235.4]
  wire [2:0] _T_1356; // @[Mux.scala 31:69:@10236.4]
  wire [2:0] _T_1357; // @[Mux.scala 31:69:@10237.4]
  wire [2:0] _T_1358; // @[Mux.scala 31:69:@10238.4]
  wire [2:0] _T_1359; // @[Mux.scala 31:69:@10239.4]
  wire  _T_1364; // @[MemPrimitives.scala 110:210:@10246.4]
  wire  _T_1367; // @[MemPrimitives.scala 110:228:@10248.4]
  wire  _T_1370; // @[MemPrimitives.scala 110:210:@10250.4]
  wire  _T_1373; // @[MemPrimitives.scala 110:228:@10252.4]
  wire  _T_1376; // @[MemPrimitives.scala 110:210:@10254.4]
  wire  _T_1379; // @[MemPrimitives.scala 110:228:@10256.4]
  wire  _T_1382; // @[MemPrimitives.scala 110:210:@10258.4]
  wire  _T_1385; // @[MemPrimitives.scala 110:228:@10260.4]
  wire  _T_1388; // @[MemPrimitives.scala 110:210:@10262.4]
  wire  _T_1391; // @[MemPrimitives.scala 110:228:@10264.4]
  wire  _T_1394; // @[MemPrimitives.scala 110:210:@10266.4]
  wire  _T_1397; // @[MemPrimitives.scala 110:228:@10268.4]
  wire  _T_1399; // @[MemPrimitives.scala 123:41:@10279.4]
  wire  _T_1400; // @[MemPrimitives.scala 123:41:@10280.4]
  wire  _T_1401; // @[MemPrimitives.scala 123:41:@10281.4]
  wire  _T_1402; // @[MemPrimitives.scala 123:41:@10282.4]
  wire  _T_1403; // @[MemPrimitives.scala 123:41:@10283.4]
  wire  _T_1404; // @[MemPrimitives.scala 123:41:@10284.4]
  wire [2:0] _T_1406; // @[Cat.scala 30:58:@10286.4]
  wire [2:0] _T_1408; // @[Cat.scala 30:58:@10288.4]
  wire [2:0] _T_1410; // @[Cat.scala 30:58:@10290.4]
  wire [2:0] _T_1412; // @[Cat.scala 30:58:@10292.4]
  wire [2:0] _T_1414; // @[Cat.scala 30:58:@10294.4]
  wire [2:0] _T_1416; // @[Cat.scala 30:58:@10296.4]
  wire [2:0] _T_1417; // @[Mux.scala 31:69:@10297.4]
  wire [2:0] _T_1418; // @[Mux.scala 31:69:@10298.4]
  wire [2:0] _T_1419; // @[Mux.scala 31:69:@10299.4]
  wire [2:0] _T_1420; // @[Mux.scala 31:69:@10300.4]
  wire [2:0] _T_1421; // @[Mux.scala 31:69:@10301.4]
  wire  _T_1426; // @[MemPrimitives.scala 110:210:@10308.4]
  wire  _T_1429; // @[MemPrimitives.scala 110:228:@10310.4]
  wire  _T_1432; // @[MemPrimitives.scala 110:210:@10312.4]
  wire  _T_1435; // @[MemPrimitives.scala 110:228:@10314.4]
  wire  _T_1438; // @[MemPrimitives.scala 110:210:@10316.4]
  wire  _T_1441; // @[MemPrimitives.scala 110:228:@10318.4]
  wire  _T_1444; // @[MemPrimitives.scala 110:210:@10320.4]
  wire  _T_1447; // @[MemPrimitives.scala 110:228:@10322.4]
  wire  _T_1450; // @[MemPrimitives.scala 110:210:@10324.4]
  wire  _T_1453; // @[MemPrimitives.scala 110:228:@10326.4]
  wire  _T_1456; // @[MemPrimitives.scala 110:210:@10328.4]
  wire  _T_1459; // @[MemPrimitives.scala 110:228:@10330.4]
  wire  _T_1461; // @[MemPrimitives.scala 123:41:@10341.4]
  wire  _T_1462; // @[MemPrimitives.scala 123:41:@10342.4]
  wire  _T_1463; // @[MemPrimitives.scala 123:41:@10343.4]
  wire  _T_1464; // @[MemPrimitives.scala 123:41:@10344.4]
  wire  _T_1465; // @[MemPrimitives.scala 123:41:@10345.4]
  wire  _T_1466; // @[MemPrimitives.scala 123:41:@10346.4]
  wire [2:0] _T_1468; // @[Cat.scala 30:58:@10348.4]
  wire [2:0] _T_1470; // @[Cat.scala 30:58:@10350.4]
  wire [2:0] _T_1472; // @[Cat.scala 30:58:@10352.4]
  wire [2:0] _T_1474; // @[Cat.scala 30:58:@10354.4]
  wire [2:0] _T_1476; // @[Cat.scala 30:58:@10356.4]
  wire [2:0] _T_1478; // @[Cat.scala 30:58:@10358.4]
  wire [2:0] _T_1479; // @[Mux.scala 31:69:@10359.4]
  wire [2:0] _T_1480; // @[Mux.scala 31:69:@10360.4]
  wire [2:0] _T_1481; // @[Mux.scala 31:69:@10361.4]
  wire [2:0] _T_1482; // @[Mux.scala 31:69:@10362.4]
  wire [2:0] _T_1483; // @[Mux.scala 31:69:@10363.4]
  wire  _T_1491; // @[MemPrimitives.scala 110:228:@10372.4]
  wire  _T_1497; // @[MemPrimitives.scala 110:228:@10376.4]
  wire  _T_1503; // @[MemPrimitives.scala 110:228:@10380.4]
  wire  _T_1509; // @[MemPrimitives.scala 110:228:@10384.4]
  wire  _T_1515; // @[MemPrimitives.scala 110:228:@10388.4]
  wire  _T_1521; // @[MemPrimitives.scala 110:228:@10392.4]
  wire  _T_1523; // @[MemPrimitives.scala 123:41:@10403.4]
  wire  _T_1524; // @[MemPrimitives.scala 123:41:@10404.4]
  wire  _T_1525; // @[MemPrimitives.scala 123:41:@10405.4]
  wire  _T_1526; // @[MemPrimitives.scala 123:41:@10406.4]
  wire  _T_1527; // @[MemPrimitives.scala 123:41:@10407.4]
  wire  _T_1528; // @[MemPrimitives.scala 123:41:@10408.4]
  wire [2:0] _T_1530; // @[Cat.scala 30:58:@10410.4]
  wire [2:0] _T_1532; // @[Cat.scala 30:58:@10412.4]
  wire [2:0] _T_1534; // @[Cat.scala 30:58:@10414.4]
  wire [2:0] _T_1536; // @[Cat.scala 30:58:@10416.4]
  wire [2:0] _T_1538; // @[Cat.scala 30:58:@10418.4]
  wire [2:0] _T_1540; // @[Cat.scala 30:58:@10420.4]
  wire [2:0] _T_1541; // @[Mux.scala 31:69:@10421.4]
  wire [2:0] _T_1542; // @[Mux.scala 31:69:@10422.4]
  wire [2:0] _T_1543; // @[Mux.scala 31:69:@10423.4]
  wire [2:0] _T_1544; // @[Mux.scala 31:69:@10424.4]
  wire [2:0] _T_1545; // @[Mux.scala 31:69:@10425.4]
  wire  _T_1553; // @[MemPrimitives.scala 110:228:@10434.4]
  wire  _T_1559; // @[MemPrimitives.scala 110:228:@10438.4]
  wire  _T_1565; // @[MemPrimitives.scala 110:228:@10442.4]
  wire  _T_1571; // @[MemPrimitives.scala 110:228:@10446.4]
  wire  _T_1577; // @[MemPrimitives.scala 110:228:@10450.4]
  wire  _T_1583; // @[MemPrimitives.scala 110:228:@10454.4]
  wire  _T_1585; // @[MemPrimitives.scala 123:41:@10465.4]
  wire  _T_1586; // @[MemPrimitives.scala 123:41:@10466.4]
  wire  _T_1587; // @[MemPrimitives.scala 123:41:@10467.4]
  wire  _T_1588; // @[MemPrimitives.scala 123:41:@10468.4]
  wire  _T_1589; // @[MemPrimitives.scala 123:41:@10469.4]
  wire  _T_1590; // @[MemPrimitives.scala 123:41:@10470.4]
  wire [2:0] _T_1592; // @[Cat.scala 30:58:@10472.4]
  wire [2:0] _T_1594; // @[Cat.scala 30:58:@10474.4]
  wire [2:0] _T_1596; // @[Cat.scala 30:58:@10476.4]
  wire [2:0] _T_1598; // @[Cat.scala 30:58:@10478.4]
  wire [2:0] _T_1600; // @[Cat.scala 30:58:@10480.4]
  wire [2:0] _T_1602; // @[Cat.scala 30:58:@10482.4]
  wire [2:0] _T_1603; // @[Mux.scala 31:69:@10483.4]
  wire [2:0] _T_1604; // @[Mux.scala 31:69:@10484.4]
  wire [2:0] _T_1605; // @[Mux.scala 31:69:@10485.4]
  wire [2:0] _T_1606; // @[Mux.scala 31:69:@10486.4]
  wire [2:0] _T_1607; // @[Mux.scala 31:69:@10487.4]
  wire  _T_1671; // @[package.scala 96:25:@10572.4 package.scala 96:25:@10573.4]
  wire [7:0] _T_1675; // @[Mux.scala 31:69:@10582.4]
  wire  _T_1668; // @[package.scala 96:25:@10564.4 package.scala 96:25:@10565.4]
  wire [7:0] _T_1676; // @[Mux.scala 31:69:@10583.4]
  wire  _T_1665; // @[package.scala 96:25:@10556.4 package.scala 96:25:@10557.4]
  wire [7:0] _T_1677; // @[Mux.scala 31:69:@10584.4]
  wire  _T_1662; // @[package.scala 96:25:@10548.4 package.scala 96:25:@10549.4]
  wire [7:0] _T_1678; // @[Mux.scala 31:69:@10585.4]
  wire  _T_1659; // @[package.scala 96:25:@10540.4 package.scala 96:25:@10541.4]
  wire [7:0] _T_1679; // @[Mux.scala 31:69:@10586.4]
  wire  _T_1656; // @[package.scala 96:25:@10532.4 package.scala 96:25:@10533.4]
  wire [7:0] _T_1680; // @[Mux.scala 31:69:@10587.4]
  wire  _T_1653; // @[package.scala 96:25:@10524.4 package.scala 96:25:@10525.4]
  wire  _T_1742; // @[package.scala 96:25:@10668.4 package.scala 96:25:@10669.4]
  wire [7:0] _T_1746; // @[Mux.scala 31:69:@10678.4]
  wire  _T_1739; // @[package.scala 96:25:@10660.4 package.scala 96:25:@10661.4]
  wire [7:0] _T_1747; // @[Mux.scala 31:69:@10679.4]
  wire  _T_1736; // @[package.scala 96:25:@10652.4 package.scala 96:25:@10653.4]
  wire [7:0] _T_1748; // @[Mux.scala 31:69:@10680.4]
  wire  _T_1733; // @[package.scala 96:25:@10644.4 package.scala 96:25:@10645.4]
  wire [7:0] _T_1749; // @[Mux.scala 31:69:@10681.4]
  wire  _T_1730; // @[package.scala 96:25:@10636.4 package.scala 96:25:@10637.4]
  wire [7:0] _T_1750; // @[Mux.scala 31:69:@10682.4]
  wire  _T_1727; // @[package.scala 96:25:@10628.4 package.scala 96:25:@10629.4]
  wire [7:0] _T_1751; // @[Mux.scala 31:69:@10683.4]
  wire  _T_1724; // @[package.scala 96:25:@10620.4 package.scala 96:25:@10621.4]
  wire  _T_1813; // @[package.scala 96:25:@10764.4 package.scala 96:25:@10765.4]
  wire [7:0] _T_1817; // @[Mux.scala 31:69:@10774.4]
  wire  _T_1810; // @[package.scala 96:25:@10756.4 package.scala 96:25:@10757.4]
  wire [7:0] _T_1818; // @[Mux.scala 31:69:@10775.4]
  wire  _T_1807; // @[package.scala 96:25:@10748.4 package.scala 96:25:@10749.4]
  wire [7:0] _T_1819; // @[Mux.scala 31:69:@10776.4]
  wire  _T_1804; // @[package.scala 96:25:@10740.4 package.scala 96:25:@10741.4]
  wire [7:0] _T_1820; // @[Mux.scala 31:69:@10777.4]
  wire  _T_1801; // @[package.scala 96:25:@10732.4 package.scala 96:25:@10733.4]
  wire [7:0] _T_1821; // @[Mux.scala 31:69:@10778.4]
  wire  _T_1798; // @[package.scala 96:25:@10724.4 package.scala 96:25:@10725.4]
  wire [7:0] _T_1822; // @[Mux.scala 31:69:@10779.4]
  wire  _T_1795; // @[package.scala 96:25:@10716.4 package.scala 96:25:@10717.4]
  wire  _T_1884; // @[package.scala 96:25:@10860.4 package.scala 96:25:@10861.4]
  wire [7:0] _T_1888; // @[Mux.scala 31:69:@10870.4]
  wire  _T_1881; // @[package.scala 96:25:@10852.4 package.scala 96:25:@10853.4]
  wire [7:0] _T_1889; // @[Mux.scala 31:69:@10871.4]
  wire  _T_1878; // @[package.scala 96:25:@10844.4 package.scala 96:25:@10845.4]
  wire [7:0] _T_1890; // @[Mux.scala 31:69:@10872.4]
  wire  _T_1875; // @[package.scala 96:25:@10836.4 package.scala 96:25:@10837.4]
  wire [7:0] _T_1891; // @[Mux.scala 31:69:@10873.4]
  wire  _T_1872; // @[package.scala 96:25:@10828.4 package.scala 96:25:@10829.4]
  wire [7:0] _T_1892; // @[Mux.scala 31:69:@10874.4]
  wire  _T_1869; // @[package.scala 96:25:@10820.4 package.scala 96:25:@10821.4]
  wire [7:0] _T_1893; // @[Mux.scala 31:69:@10875.4]
  wire  _T_1866; // @[package.scala 96:25:@10812.4 package.scala 96:25:@10813.4]
  wire  _T_1955; // @[package.scala 96:25:@10956.4 package.scala 96:25:@10957.4]
  wire [7:0] _T_1959; // @[Mux.scala 31:69:@10966.4]
  wire  _T_1952; // @[package.scala 96:25:@10948.4 package.scala 96:25:@10949.4]
  wire [7:0] _T_1960; // @[Mux.scala 31:69:@10967.4]
  wire  _T_1949; // @[package.scala 96:25:@10940.4 package.scala 96:25:@10941.4]
  wire [7:0] _T_1961; // @[Mux.scala 31:69:@10968.4]
  wire  _T_1946; // @[package.scala 96:25:@10932.4 package.scala 96:25:@10933.4]
  wire [7:0] _T_1962; // @[Mux.scala 31:69:@10969.4]
  wire  _T_1943; // @[package.scala 96:25:@10924.4 package.scala 96:25:@10925.4]
  wire [7:0] _T_1963; // @[Mux.scala 31:69:@10970.4]
  wire  _T_1940; // @[package.scala 96:25:@10916.4 package.scala 96:25:@10917.4]
  wire [7:0] _T_1964; // @[Mux.scala 31:69:@10971.4]
  wire  _T_1937; // @[package.scala 96:25:@10908.4 package.scala 96:25:@10909.4]
  wire  _T_2026; // @[package.scala 96:25:@11052.4 package.scala 96:25:@11053.4]
  wire [7:0] _T_2030; // @[Mux.scala 31:69:@11062.4]
  wire  _T_2023; // @[package.scala 96:25:@11044.4 package.scala 96:25:@11045.4]
  wire [7:0] _T_2031; // @[Mux.scala 31:69:@11063.4]
  wire  _T_2020; // @[package.scala 96:25:@11036.4 package.scala 96:25:@11037.4]
  wire [7:0] _T_2032; // @[Mux.scala 31:69:@11064.4]
  wire  _T_2017; // @[package.scala 96:25:@11028.4 package.scala 96:25:@11029.4]
  wire [7:0] _T_2033; // @[Mux.scala 31:69:@11065.4]
  wire  _T_2014; // @[package.scala 96:25:@11020.4 package.scala 96:25:@11021.4]
  wire [7:0] _T_2034; // @[Mux.scala 31:69:@11066.4]
  wire  _T_2011; // @[package.scala 96:25:@11012.4 package.scala 96:25:@11013.4]
  wire [7:0] _T_2035; // @[Mux.scala 31:69:@11067.4]
  wire  _T_2008; // @[package.scala 96:25:@11004.4 package.scala 96:25:@11005.4]
  wire  _T_2097; // @[package.scala 96:25:@11148.4 package.scala 96:25:@11149.4]
  wire [7:0] _T_2101; // @[Mux.scala 31:69:@11158.4]
  wire  _T_2094; // @[package.scala 96:25:@11140.4 package.scala 96:25:@11141.4]
  wire [7:0] _T_2102; // @[Mux.scala 31:69:@11159.4]
  wire  _T_2091; // @[package.scala 96:25:@11132.4 package.scala 96:25:@11133.4]
  wire [7:0] _T_2103; // @[Mux.scala 31:69:@11160.4]
  wire  _T_2088; // @[package.scala 96:25:@11124.4 package.scala 96:25:@11125.4]
  wire [7:0] _T_2104; // @[Mux.scala 31:69:@11161.4]
  wire  _T_2085; // @[package.scala 96:25:@11116.4 package.scala 96:25:@11117.4]
  wire [7:0] _T_2105; // @[Mux.scala 31:69:@11162.4]
  wire  _T_2082; // @[package.scala 96:25:@11108.4 package.scala 96:25:@11109.4]
  wire [7:0] _T_2106; // @[Mux.scala 31:69:@11163.4]
  wire  _T_2079; // @[package.scala 96:25:@11100.4 package.scala 96:25:@11101.4]
  wire  _T_2168; // @[package.scala 96:25:@11244.4 package.scala 96:25:@11245.4]
  wire [7:0] _T_2172; // @[Mux.scala 31:69:@11254.4]
  wire  _T_2165; // @[package.scala 96:25:@11236.4 package.scala 96:25:@11237.4]
  wire [7:0] _T_2173; // @[Mux.scala 31:69:@11255.4]
  wire  _T_2162; // @[package.scala 96:25:@11228.4 package.scala 96:25:@11229.4]
  wire [7:0] _T_2174; // @[Mux.scala 31:69:@11256.4]
  wire  _T_2159; // @[package.scala 96:25:@11220.4 package.scala 96:25:@11221.4]
  wire [7:0] _T_2175; // @[Mux.scala 31:69:@11257.4]
  wire  _T_2156; // @[package.scala 96:25:@11212.4 package.scala 96:25:@11213.4]
  wire [7:0] _T_2176; // @[Mux.scala 31:69:@11258.4]
  wire  _T_2153; // @[package.scala 96:25:@11204.4 package.scala 96:25:@11205.4]
  wire [7:0] _T_2177; // @[Mux.scala 31:69:@11259.4]
  wire  _T_2150; // @[package.scala 96:25:@11196.4 package.scala 96:25:@11197.4]
  wire  _T_2239; // @[package.scala 96:25:@11340.4 package.scala 96:25:@11341.4]
  wire [7:0] _T_2243; // @[Mux.scala 31:69:@11350.4]
  wire  _T_2236; // @[package.scala 96:25:@11332.4 package.scala 96:25:@11333.4]
  wire [7:0] _T_2244; // @[Mux.scala 31:69:@11351.4]
  wire  _T_2233; // @[package.scala 96:25:@11324.4 package.scala 96:25:@11325.4]
  wire [7:0] _T_2245; // @[Mux.scala 31:69:@11352.4]
  wire  _T_2230; // @[package.scala 96:25:@11316.4 package.scala 96:25:@11317.4]
  wire [7:0] _T_2246; // @[Mux.scala 31:69:@11353.4]
  wire  _T_2227; // @[package.scala 96:25:@11308.4 package.scala 96:25:@11309.4]
  wire [7:0] _T_2247; // @[Mux.scala 31:69:@11354.4]
  wire  _T_2224; // @[package.scala 96:25:@11300.4 package.scala 96:25:@11301.4]
  wire [7:0] _T_2248; // @[Mux.scala 31:69:@11355.4]
  wire  _T_2221; // @[package.scala 96:25:@11292.4 package.scala 96:25:@11293.4]
  wire  _T_2310; // @[package.scala 96:25:@11436.4 package.scala 96:25:@11437.4]
  wire [7:0] _T_2314; // @[Mux.scala 31:69:@11446.4]
  wire  _T_2307; // @[package.scala 96:25:@11428.4 package.scala 96:25:@11429.4]
  wire [7:0] _T_2315; // @[Mux.scala 31:69:@11447.4]
  wire  _T_2304; // @[package.scala 96:25:@11420.4 package.scala 96:25:@11421.4]
  wire [7:0] _T_2316; // @[Mux.scala 31:69:@11448.4]
  wire  _T_2301; // @[package.scala 96:25:@11412.4 package.scala 96:25:@11413.4]
  wire [7:0] _T_2317; // @[Mux.scala 31:69:@11449.4]
  wire  _T_2298; // @[package.scala 96:25:@11404.4 package.scala 96:25:@11405.4]
  wire [7:0] _T_2318; // @[Mux.scala 31:69:@11450.4]
  wire  _T_2295; // @[package.scala 96:25:@11396.4 package.scala 96:25:@11397.4]
  wire [7:0] _T_2319; // @[Mux.scala 31:69:@11451.4]
  wire  _T_2292; // @[package.scala 96:25:@11388.4 package.scala 96:25:@11389.4]
  wire  _T_2381; // @[package.scala 96:25:@11532.4 package.scala 96:25:@11533.4]
  wire [7:0] _T_2385; // @[Mux.scala 31:69:@11542.4]
  wire  _T_2378; // @[package.scala 96:25:@11524.4 package.scala 96:25:@11525.4]
  wire [7:0] _T_2386; // @[Mux.scala 31:69:@11543.4]
  wire  _T_2375; // @[package.scala 96:25:@11516.4 package.scala 96:25:@11517.4]
  wire [7:0] _T_2387; // @[Mux.scala 31:69:@11544.4]
  wire  _T_2372; // @[package.scala 96:25:@11508.4 package.scala 96:25:@11509.4]
  wire [7:0] _T_2388; // @[Mux.scala 31:69:@11545.4]
  wire  _T_2369; // @[package.scala 96:25:@11500.4 package.scala 96:25:@11501.4]
  wire [7:0] _T_2389; // @[Mux.scala 31:69:@11546.4]
  wire  _T_2366; // @[package.scala 96:25:@11492.4 package.scala 96:25:@11493.4]
  wire [7:0] _T_2390; // @[Mux.scala 31:69:@11547.4]
  wire  _T_2363; // @[package.scala 96:25:@11484.4 package.scala 96:25:@11485.4]
  wire  _T_2452; // @[package.scala 96:25:@11628.4 package.scala 96:25:@11629.4]
  wire [7:0] _T_2456; // @[Mux.scala 31:69:@11638.4]
  wire  _T_2449; // @[package.scala 96:25:@11620.4 package.scala 96:25:@11621.4]
  wire [7:0] _T_2457; // @[Mux.scala 31:69:@11639.4]
  wire  _T_2446; // @[package.scala 96:25:@11612.4 package.scala 96:25:@11613.4]
  wire [7:0] _T_2458; // @[Mux.scala 31:69:@11640.4]
  wire  _T_2443; // @[package.scala 96:25:@11604.4 package.scala 96:25:@11605.4]
  wire [7:0] _T_2459; // @[Mux.scala 31:69:@11641.4]
  wire  _T_2440; // @[package.scala 96:25:@11596.4 package.scala 96:25:@11597.4]
  wire [7:0] _T_2460; // @[Mux.scala 31:69:@11642.4]
  wire  _T_2437; // @[package.scala 96:25:@11588.4 package.scala 96:25:@11589.4]
  wire [7:0] _T_2461; // @[Mux.scala 31:69:@11643.4]
  wire  _T_2434; // @[package.scala 96:25:@11580.4 package.scala 96:25:@11581.4]
  Mem1D_4 Mem1D ( // @[MemPrimitives.scala 64:21:@9054.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  Mem1D_4 Mem1D_1 ( // @[MemPrimitives.scala 64:21:@9070.4]
    .clock(Mem1D_1_clock),
    .reset(Mem1D_1_reset),
    .io_r_ofs_0(Mem1D_1_io_r_ofs_0),
    .io_r_backpressure(Mem1D_1_io_r_backpressure),
    .io_w_ofs_0(Mem1D_1_io_w_ofs_0),
    .io_w_data_0(Mem1D_1_io_w_data_0),
    .io_w_en_0(Mem1D_1_io_w_en_0),
    .io_output(Mem1D_1_io_output)
  );
  Mem1D_4 Mem1D_2 ( // @[MemPrimitives.scala 64:21:@9086.4]
    .clock(Mem1D_2_clock),
    .reset(Mem1D_2_reset),
    .io_r_ofs_0(Mem1D_2_io_r_ofs_0),
    .io_r_backpressure(Mem1D_2_io_r_backpressure),
    .io_w_ofs_0(Mem1D_2_io_w_ofs_0),
    .io_w_data_0(Mem1D_2_io_w_data_0),
    .io_w_en_0(Mem1D_2_io_w_en_0),
    .io_output(Mem1D_2_io_output)
  );
  Mem1D_4 Mem1D_3 ( // @[MemPrimitives.scala 64:21:@9102.4]
    .clock(Mem1D_3_clock),
    .reset(Mem1D_3_reset),
    .io_r_ofs_0(Mem1D_3_io_r_ofs_0),
    .io_r_backpressure(Mem1D_3_io_r_backpressure),
    .io_w_ofs_0(Mem1D_3_io_w_ofs_0),
    .io_w_data_0(Mem1D_3_io_w_data_0),
    .io_w_en_0(Mem1D_3_io_w_en_0),
    .io_output(Mem1D_3_io_output)
  );
  Mem1D_4 Mem1D_4 ( // @[MemPrimitives.scala 64:21:@9118.4]
    .clock(Mem1D_4_clock),
    .reset(Mem1D_4_reset),
    .io_r_ofs_0(Mem1D_4_io_r_ofs_0),
    .io_r_backpressure(Mem1D_4_io_r_backpressure),
    .io_w_ofs_0(Mem1D_4_io_w_ofs_0),
    .io_w_data_0(Mem1D_4_io_w_data_0),
    .io_w_en_0(Mem1D_4_io_w_en_0),
    .io_output(Mem1D_4_io_output)
  );
  Mem1D_4 Mem1D_5 ( // @[MemPrimitives.scala 64:21:@9134.4]
    .clock(Mem1D_5_clock),
    .reset(Mem1D_5_reset),
    .io_r_ofs_0(Mem1D_5_io_r_ofs_0),
    .io_r_backpressure(Mem1D_5_io_r_backpressure),
    .io_w_ofs_0(Mem1D_5_io_w_ofs_0),
    .io_w_data_0(Mem1D_5_io_w_data_0),
    .io_w_en_0(Mem1D_5_io_w_en_0),
    .io_output(Mem1D_5_io_output)
  );
  Mem1D_4 Mem1D_6 ( // @[MemPrimitives.scala 64:21:@9150.4]
    .clock(Mem1D_6_clock),
    .reset(Mem1D_6_reset),
    .io_r_ofs_0(Mem1D_6_io_r_ofs_0),
    .io_r_backpressure(Mem1D_6_io_r_backpressure),
    .io_w_ofs_0(Mem1D_6_io_w_ofs_0),
    .io_w_data_0(Mem1D_6_io_w_data_0),
    .io_w_en_0(Mem1D_6_io_w_en_0),
    .io_output(Mem1D_6_io_output)
  );
  Mem1D_4 Mem1D_7 ( // @[MemPrimitives.scala 64:21:@9166.4]
    .clock(Mem1D_7_clock),
    .reset(Mem1D_7_reset),
    .io_r_ofs_0(Mem1D_7_io_r_ofs_0),
    .io_r_backpressure(Mem1D_7_io_r_backpressure),
    .io_w_ofs_0(Mem1D_7_io_w_ofs_0),
    .io_w_data_0(Mem1D_7_io_w_data_0),
    .io_w_en_0(Mem1D_7_io_w_en_0),
    .io_output(Mem1D_7_io_output)
  );
  Mem1D_4 Mem1D_8 ( // @[MemPrimitives.scala 64:21:@9182.4]
    .clock(Mem1D_8_clock),
    .reset(Mem1D_8_reset),
    .io_r_ofs_0(Mem1D_8_io_r_ofs_0),
    .io_r_backpressure(Mem1D_8_io_r_backpressure),
    .io_w_ofs_0(Mem1D_8_io_w_ofs_0),
    .io_w_data_0(Mem1D_8_io_w_data_0),
    .io_w_en_0(Mem1D_8_io_w_en_0),
    .io_output(Mem1D_8_io_output)
  );
  Mem1D_4 Mem1D_9 ( // @[MemPrimitives.scala 64:21:@9198.4]
    .clock(Mem1D_9_clock),
    .reset(Mem1D_9_reset),
    .io_r_ofs_0(Mem1D_9_io_r_ofs_0),
    .io_r_backpressure(Mem1D_9_io_r_backpressure),
    .io_w_ofs_0(Mem1D_9_io_w_ofs_0),
    .io_w_data_0(Mem1D_9_io_w_data_0),
    .io_w_en_0(Mem1D_9_io_w_en_0),
    .io_output(Mem1D_9_io_output)
  );
  Mem1D_4 Mem1D_10 ( // @[MemPrimitives.scala 64:21:@9214.4]
    .clock(Mem1D_10_clock),
    .reset(Mem1D_10_reset),
    .io_r_ofs_0(Mem1D_10_io_r_ofs_0),
    .io_r_backpressure(Mem1D_10_io_r_backpressure),
    .io_w_ofs_0(Mem1D_10_io_w_ofs_0),
    .io_w_data_0(Mem1D_10_io_w_data_0),
    .io_w_en_0(Mem1D_10_io_w_en_0),
    .io_output(Mem1D_10_io_output)
  );
  Mem1D_4 Mem1D_11 ( // @[MemPrimitives.scala 64:21:@9230.4]
    .clock(Mem1D_11_clock),
    .reset(Mem1D_11_reset),
    .io_r_ofs_0(Mem1D_11_io_r_ofs_0),
    .io_r_backpressure(Mem1D_11_io_r_backpressure),
    .io_w_ofs_0(Mem1D_11_io_w_ofs_0),
    .io_w_data_0(Mem1D_11_io_w_data_0),
    .io_w_en_0(Mem1D_11_io_w_en_0),
    .io_output(Mem1D_11_io_output)
  );
  Mem1D_4 Mem1D_12 ( // @[MemPrimitives.scala 64:21:@9246.4]
    .clock(Mem1D_12_clock),
    .reset(Mem1D_12_reset),
    .io_r_ofs_0(Mem1D_12_io_r_ofs_0),
    .io_r_backpressure(Mem1D_12_io_r_backpressure),
    .io_w_ofs_0(Mem1D_12_io_w_ofs_0),
    .io_w_data_0(Mem1D_12_io_w_data_0),
    .io_w_en_0(Mem1D_12_io_w_en_0),
    .io_output(Mem1D_12_io_output)
  );
  Mem1D_4 Mem1D_13 ( // @[MemPrimitives.scala 64:21:@9262.4]
    .clock(Mem1D_13_clock),
    .reset(Mem1D_13_reset),
    .io_r_ofs_0(Mem1D_13_io_r_ofs_0),
    .io_r_backpressure(Mem1D_13_io_r_backpressure),
    .io_w_ofs_0(Mem1D_13_io_w_ofs_0),
    .io_w_data_0(Mem1D_13_io_w_data_0),
    .io_w_en_0(Mem1D_13_io_w_en_0),
    .io_output(Mem1D_13_io_output)
  );
  Mem1D_4 Mem1D_14 ( // @[MemPrimitives.scala 64:21:@9278.4]
    .clock(Mem1D_14_clock),
    .reset(Mem1D_14_reset),
    .io_r_ofs_0(Mem1D_14_io_r_ofs_0),
    .io_r_backpressure(Mem1D_14_io_r_backpressure),
    .io_w_ofs_0(Mem1D_14_io_w_ofs_0),
    .io_w_data_0(Mem1D_14_io_w_data_0),
    .io_w_en_0(Mem1D_14_io_w_en_0),
    .io_output(Mem1D_14_io_output)
  );
  Mem1D_4 Mem1D_15 ( // @[MemPrimitives.scala 64:21:@9294.4]
    .clock(Mem1D_15_clock),
    .reset(Mem1D_15_reset),
    .io_r_ofs_0(Mem1D_15_io_r_ofs_0),
    .io_r_backpressure(Mem1D_15_io_r_backpressure),
    .io_w_ofs_0(Mem1D_15_io_w_ofs_0),
    .io_w_data_0(Mem1D_15_io_w_data_0),
    .io_w_en_0(Mem1D_15_io_w_en_0),
    .io_output(Mem1D_15_io_output)
  );
  StickySelects StickySelects ( // @[MemPrimitives.scala 121:29:@9526.4]
    .clock(StickySelects_clock),
    .reset(StickySelects_reset),
    .io_ins_0(StickySelects_io_ins_0),
    .io_ins_1(StickySelects_io_ins_1),
    .io_ins_2(StickySelects_io_ins_2),
    .io_ins_3(StickySelects_io_ins_3),
    .io_ins_4(StickySelects_io_ins_4),
    .io_ins_5(StickySelects_io_ins_5),
    .io_outs_0(StickySelects_io_outs_0),
    .io_outs_1(StickySelects_io_outs_1),
    .io_outs_2(StickySelects_io_outs_2),
    .io_outs_3(StickySelects_io_outs_3),
    .io_outs_4(StickySelects_io_outs_4),
    .io_outs_5(StickySelects_io_outs_5)
  );
  StickySelects StickySelects_1 ( // @[MemPrimitives.scala 121:29:@9588.4]
    .clock(StickySelects_1_clock),
    .reset(StickySelects_1_reset),
    .io_ins_0(StickySelects_1_io_ins_0),
    .io_ins_1(StickySelects_1_io_ins_1),
    .io_ins_2(StickySelects_1_io_ins_2),
    .io_ins_3(StickySelects_1_io_ins_3),
    .io_ins_4(StickySelects_1_io_ins_4),
    .io_ins_5(StickySelects_1_io_ins_5),
    .io_outs_0(StickySelects_1_io_outs_0),
    .io_outs_1(StickySelects_1_io_outs_1),
    .io_outs_2(StickySelects_1_io_outs_2),
    .io_outs_3(StickySelects_1_io_outs_3),
    .io_outs_4(StickySelects_1_io_outs_4),
    .io_outs_5(StickySelects_1_io_outs_5)
  );
  StickySelects StickySelects_2 ( // @[MemPrimitives.scala 121:29:@9650.4]
    .clock(StickySelects_2_clock),
    .reset(StickySelects_2_reset),
    .io_ins_0(StickySelects_2_io_ins_0),
    .io_ins_1(StickySelects_2_io_ins_1),
    .io_ins_2(StickySelects_2_io_ins_2),
    .io_ins_3(StickySelects_2_io_ins_3),
    .io_ins_4(StickySelects_2_io_ins_4),
    .io_ins_5(StickySelects_2_io_ins_5),
    .io_outs_0(StickySelects_2_io_outs_0),
    .io_outs_1(StickySelects_2_io_outs_1),
    .io_outs_2(StickySelects_2_io_outs_2),
    .io_outs_3(StickySelects_2_io_outs_3),
    .io_outs_4(StickySelects_2_io_outs_4),
    .io_outs_5(StickySelects_2_io_outs_5)
  );
  StickySelects StickySelects_3 ( // @[MemPrimitives.scala 121:29:@9712.4]
    .clock(StickySelects_3_clock),
    .reset(StickySelects_3_reset),
    .io_ins_0(StickySelects_3_io_ins_0),
    .io_ins_1(StickySelects_3_io_ins_1),
    .io_ins_2(StickySelects_3_io_ins_2),
    .io_ins_3(StickySelects_3_io_ins_3),
    .io_ins_4(StickySelects_3_io_ins_4),
    .io_ins_5(StickySelects_3_io_ins_5),
    .io_outs_0(StickySelects_3_io_outs_0),
    .io_outs_1(StickySelects_3_io_outs_1),
    .io_outs_2(StickySelects_3_io_outs_2),
    .io_outs_3(StickySelects_3_io_outs_3),
    .io_outs_4(StickySelects_3_io_outs_4),
    .io_outs_5(StickySelects_3_io_outs_5)
  );
  StickySelects StickySelects_4 ( // @[MemPrimitives.scala 121:29:@9774.4]
    .clock(StickySelects_4_clock),
    .reset(StickySelects_4_reset),
    .io_ins_0(StickySelects_4_io_ins_0),
    .io_ins_1(StickySelects_4_io_ins_1),
    .io_ins_2(StickySelects_4_io_ins_2),
    .io_ins_3(StickySelects_4_io_ins_3),
    .io_ins_4(StickySelects_4_io_ins_4),
    .io_ins_5(StickySelects_4_io_ins_5),
    .io_outs_0(StickySelects_4_io_outs_0),
    .io_outs_1(StickySelects_4_io_outs_1),
    .io_outs_2(StickySelects_4_io_outs_2),
    .io_outs_3(StickySelects_4_io_outs_3),
    .io_outs_4(StickySelects_4_io_outs_4),
    .io_outs_5(StickySelects_4_io_outs_5)
  );
  StickySelects StickySelects_5 ( // @[MemPrimitives.scala 121:29:@9836.4]
    .clock(StickySelects_5_clock),
    .reset(StickySelects_5_reset),
    .io_ins_0(StickySelects_5_io_ins_0),
    .io_ins_1(StickySelects_5_io_ins_1),
    .io_ins_2(StickySelects_5_io_ins_2),
    .io_ins_3(StickySelects_5_io_ins_3),
    .io_ins_4(StickySelects_5_io_ins_4),
    .io_ins_5(StickySelects_5_io_ins_5),
    .io_outs_0(StickySelects_5_io_outs_0),
    .io_outs_1(StickySelects_5_io_outs_1),
    .io_outs_2(StickySelects_5_io_outs_2),
    .io_outs_3(StickySelects_5_io_outs_3),
    .io_outs_4(StickySelects_5_io_outs_4),
    .io_outs_5(StickySelects_5_io_outs_5)
  );
  StickySelects StickySelects_6 ( // @[MemPrimitives.scala 121:29:@9898.4]
    .clock(StickySelects_6_clock),
    .reset(StickySelects_6_reset),
    .io_ins_0(StickySelects_6_io_ins_0),
    .io_ins_1(StickySelects_6_io_ins_1),
    .io_ins_2(StickySelects_6_io_ins_2),
    .io_ins_3(StickySelects_6_io_ins_3),
    .io_ins_4(StickySelects_6_io_ins_4),
    .io_ins_5(StickySelects_6_io_ins_5),
    .io_outs_0(StickySelects_6_io_outs_0),
    .io_outs_1(StickySelects_6_io_outs_1),
    .io_outs_2(StickySelects_6_io_outs_2),
    .io_outs_3(StickySelects_6_io_outs_3),
    .io_outs_4(StickySelects_6_io_outs_4),
    .io_outs_5(StickySelects_6_io_outs_5)
  );
  StickySelects StickySelects_7 ( // @[MemPrimitives.scala 121:29:@9960.4]
    .clock(StickySelects_7_clock),
    .reset(StickySelects_7_reset),
    .io_ins_0(StickySelects_7_io_ins_0),
    .io_ins_1(StickySelects_7_io_ins_1),
    .io_ins_2(StickySelects_7_io_ins_2),
    .io_ins_3(StickySelects_7_io_ins_3),
    .io_ins_4(StickySelects_7_io_ins_4),
    .io_ins_5(StickySelects_7_io_ins_5),
    .io_outs_0(StickySelects_7_io_outs_0),
    .io_outs_1(StickySelects_7_io_outs_1),
    .io_outs_2(StickySelects_7_io_outs_2),
    .io_outs_3(StickySelects_7_io_outs_3),
    .io_outs_4(StickySelects_7_io_outs_4),
    .io_outs_5(StickySelects_7_io_outs_5)
  );
  StickySelects StickySelects_8 ( // @[MemPrimitives.scala 121:29:@10022.4]
    .clock(StickySelects_8_clock),
    .reset(StickySelects_8_reset),
    .io_ins_0(StickySelects_8_io_ins_0),
    .io_ins_1(StickySelects_8_io_ins_1),
    .io_ins_2(StickySelects_8_io_ins_2),
    .io_ins_3(StickySelects_8_io_ins_3),
    .io_ins_4(StickySelects_8_io_ins_4),
    .io_ins_5(StickySelects_8_io_ins_5),
    .io_outs_0(StickySelects_8_io_outs_0),
    .io_outs_1(StickySelects_8_io_outs_1),
    .io_outs_2(StickySelects_8_io_outs_2),
    .io_outs_3(StickySelects_8_io_outs_3),
    .io_outs_4(StickySelects_8_io_outs_4),
    .io_outs_5(StickySelects_8_io_outs_5)
  );
  StickySelects StickySelects_9 ( // @[MemPrimitives.scala 121:29:@10084.4]
    .clock(StickySelects_9_clock),
    .reset(StickySelects_9_reset),
    .io_ins_0(StickySelects_9_io_ins_0),
    .io_ins_1(StickySelects_9_io_ins_1),
    .io_ins_2(StickySelects_9_io_ins_2),
    .io_ins_3(StickySelects_9_io_ins_3),
    .io_ins_4(StickySelects_9_io_ins_4),
    .io_ins_5(StickySelects_9_io_ins_5),
    .io_outs_0(StickySelects_9_io_outs_0),
    .io_outs_1(StickySelects_9_io_outs_1),
    .io_outs_2(StickySelects_9_io_outs_2),
    .io_outs_3(StickySelects_9_io_outs_3),
    .io_outs_4(StickySelects_9_io_outs_4),
    .io_outs_5(StickySelects_9_io_outs_5)
  );
  StickySelects StickySelects_10 ( // @[MemPrimitives.scala 121:29:@10146.4]
    .clock(StickySelects_10_clock),
    .reset(StickySelects_10_reset),
    .io_ins_0(StickySelects_10_io_ins_0),
    .io_ins_1(StickySelects_10_io_ins_1),
    .io_ins_2(StickySelects_10_io_ins_2),
    .io_ins_3(StickySelects_10_io_ins_3),
    .io_ins_4(StickySelects_10_io_ins_4),
    .io_ins_5(StickySelects_10_io_ins_5),
    .io_outs_0(StickySelects_10_io_outs_0),
    .io_outs_1(StickySelects_10_io_outs_1),
    .io_outs_2(StickySelects_10_io_outs_2),
    .io_outs_3(StickySelects_10_io_outs_3),
    .io_outs_4(StickySelects_10_io_outs_4),
    .io_outs_5(StickySelects_10_io_outs_5)
  );
  StickySelects StickySelects_11 ( // @[MemPrimitives.scala 121:29:@10208.4]
    .clock(StickySelects_11_clock),
    .reset(StickySelects_11_reset),
    .io_ins_0(StickySelects_11_io_ins_0),
    .io_ins_1(StickySelects_11_io_ins_1),
    .io_ins_2(StickySelects_11_io_ins_2),
    .io_ins_3(StickySelects_11_io_ins_3),
    .io_ins_4(StickySelects_11_io_ins_4),
    .io_ins_5(StickySelects_11_io_ins_5),
    .io_outs_0(StickySelects_11_io_outs_0),
    .io_outs_1(StickySelects_11_io_outs_1),
    .io_outs_2(StickySelects_11_io_outs_2),
    .io_outs_3(StickySelects_11_io_outs_3),
    .io_outs_4(StickySelects_11_io_outs_4),
    .io_outs_5(StickySelects_11_io_outs_5)
  );
  StickySelects StickySelects_12 ( // @[MemPrimitives.scala 121:29:@10270.4]
    .clock(StickySelects_12_clock),
    .reset(StickySelects_12_reset),
    .io_ins_0(StickySelects_12_io_ins_0),
    .io_ins_1(StickySelects_12_io_ins_1),
    .io_ins_2(StickySelects_12_io_ins_2),
    .io_ins_3(StickySelects_12_io_ins_3),
    .io_ins_4(StickySelects_12_io_ins_4),
    .io_ins_5(StickySelects_12_io_ins_5),
    .io_outs_0(StickySelects_12_io_outs_0),
    .io_outs_1(StickySelects_12_io_outs_1),
    .io_outs_2(StickySelects_12_io_outs_2),
    .io_outs_3(StickySelects_12_io_outs_3),
    .io_outs_4(StickySelects_12_io_outs_4),
    .io_outs_5(StickySelects_12_io_outs_5)
  );
  StickySelects StickySelects_13 ( // @[MemPrimitives.scala 121:29:@10332.4]
    .clock(StickySelects_13_clock),
    .reset(StickySelects_13_reset),
    .io_ins_0(StickySelects_13_io_ins_0),
    .io_ins_1(StickySelects_13_io_ins_1),
    .io_ins_2(StickySelects_13_io_ins_2),
    .io_ins_3(StickySelects_13_io_ins_3),
    .io_ins_4(StickySelects_13_io_ins_4),
    .io_ins_5(StickySelects_13_io_ins_5),
    .io_outs_0(StickySelects_13_io_outs_0),
    .io_outs_1(StickySelects_13_io_outs_1),
    .io_outs_2(StickySelects_13_io_outs_2),
    .io_outs_3(StickySelects_13_io_outs_3),
    .io_outs_4(StickySelects_13_io_outs_4),
    .io_outs_5(StickySelects_13_io_outs_5)
  );
  StickySelects StickySelects_14 ( // @[MemPrimitives.scala 121:29:@10394.4]
    .clock(StickySelects_14_clock),
    .reset(StickySelects_14_reset),
    .io_ins_0(StickySelects_14_io_ins_0),
    .io_ins_1(StickySelects_14_io_ins_1),
    .io_ins_2(StickySelects_14_io_ins_2),
    .io_ins_3(StickySelects_14_io_ins_3),
    .io_ins_4(StickySelects_14_io_ins_4),
    .io_ins_5(StickySelects_14_io_ins_5),
    .io_outs_0(StickySelects_14_io_outs_0),
    .io_outs_1(StickySelects_14_io_outs_1),
    .io_outs_2(StickySelects_14_io_outs_2),
    .io_outs_3(StickySelects_14_io_outs_3),
    .io_outs_4(StickySelects_14_io_outs_4),
    .io_outs_5(StickySelects_14_io_outs_5)
  );
  StickySelects StickySelects_15 ( // @[MemPrimitives.scala 121:29:@10456.4]
    .clock(StickySelects_15_clock),
    .reset(StickySelects_15_reset),
    .io_ins_0(StickySelects_15_io_ins_0),
    .io_ins_1(StickySelects_15_io_ins_1),
    .io_ins_2(StickySelects_15_io_ins_2),
    .io_ins_3(StickySelects_15_io_ins_3),
    .io_ins_4(StickySelects_15_io_ins_4),
    .io_ins_5(StickySelects_15_io_ins_5),
    .io_outs_0(StickySelects_15_io_outs_0),
    .io_outs_1(StickySelects_15_io_outs_1),
    .io_outs_2(StickySelects_15_io_outs_2),
    .io_outs_3(StickySelects_15_io_outs_3),
    .io_outs_4(StickySelects_15_io_outs_4),
    .io_outs_5(StickySelects_15_io_outs_5)
  );
  RetimeWrapper_52 RetimeWrapper ( // @[package.scala 93:22:@10519.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_1 ( // @[package.scala 93:22:@10527.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_2 ( // @[package.scala 93:22:@10535.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_3 ( // @[package.scala 93:22:@10543.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_4 ( // @[package.scala 93:22:@10551.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_5 ( // @[package.scala 93:22:@10559.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_6 ( // @[package.scala 93:22:@10567.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_7 ( // @[package.scala 93:22:@10575.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_8 ( // @[package.scala 93:22:@10615.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_9 ( // @[package.scala 93:22:@10623.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_10 ( // @[package.scala 93:22:@10631.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_11 ( // @[package.scala 93:22:@10639.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_12 ( // @[package.scala 93:22:@10647.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_13 ( // @[package.scala 93:22:@10655.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_14 ( // @[package.scala 93:22:@10663.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_15 ( // @[package.scala 93:22:@10671.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_16 ( // @[package.scala 93:22:@10711.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_17 ( // @[package.scala 93:22:@10719.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_18 ( // @[package.scala 93:22:@10727.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_19 ( // @[package.scala 93:22:@10735.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_20 ( // @[package.scala 93:22:@10743.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_21 ( // @[package.scala 93:22:@10751.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_22 ( // @[package.scala 93:22:@10759.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_23 ( // @[package.scala 93:22:@10767.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_24 ( // @[package.scala 93:22:@10807.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_25 ( // @[package.scala 93:22:@10815.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_26 ( // @[package.scala 93:22:@10823.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_27 ( // @[package.scala 93:22:@10831.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_28 ( // @[package.scala 93:22:@10839.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_29 ( // @[package.scala 93:22:@10847.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_30 ( // @[package.scala 93:22:@10855.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_31 ( // @[package.scala 93:22:@10863.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_32 ( // @[package.scala 93:22:@10903.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_33 ( // @[package.scala 93:22:@10911.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_34 ( // @[package.scala 93:22:@10919.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_35 ( // @[package.scala 93:22:@10927.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_36 ( // @[package.scala 93:22:@10935.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_37 ( // @[package.scala 93:22:@10943.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_38 ( // @[package.scala 93:22:@10951.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_39 ( // @[package.scala 93:22:@10959.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_40 ( // @[package.scala 93:22:@10999.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_41 ( // @[package.scala 93:22:@11007.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_42 ( // @[package.scala 93:22:@11015.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_43 ( // @[package.scala 93:22:@11023.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_44 ( // @[package.scala 93:22:@11031.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_45 ( // @[package.scala 93:22:@11039.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_46 ( // @[package.scala 93:22:@11047.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_47 ( // @[package.scala 93:22:@11055.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_48 ( // @[package.scala 93:22:@11095.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_49 ( // @[package.scala 93:22:@11103.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_50 ( // @[package.scala 93:22:@11111.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_51 ( // @[package.scala 93:22:@11119.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_52 ( // @[package.scala 93:22:@11127.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_53 ( // @[package.scala 93:22:@11135.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_54 ( // @[package.scala 93:22:@11143.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_55 ( // @[package.scala 93:22:@11151.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_56 ( // @[package.scala 93:22:@11191.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_57 ( // @[package.scala 93:22:@11199.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_58 ( // @[package.scala 93:22:@11207.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_59 ( // @[package.scala 93:22:@11215.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_60 ( // @[package.scala 93:22:@11223.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_61 ( // @[package.scala 93:22:@11231.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_62 ( // @[package.scala 93:22:@11239.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_63 ( // @[package.scala 93:22:@11247.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_64 ( // @[package.scala 93:22:@11287.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_65 ( // @[package.scala 93:22:@11295.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_66 ( // @[package.scala 93:22:@11303.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_67 ( // @[package.scala 93:22:@11311.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_68 ( // @[package.scala 93:22:@11319.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_69 ( // @[package.scala 93:22:@11327.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_70 ( // @[package.scala 93:22:@11335.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_71 ( // @[package.scala 93:22:@11343.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_72 ( // @[package.scala 93:22:@11383.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_73 ( // @[package.scala 93:22:@11391.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_74 ( // @[package.scala 93:22:@11399.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_75 ( // @[package.scala 93:22:@11407.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_76 ( // @[package.scala 93:22:@11415.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_77 ( // @[package.scala 93:22:@11423.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_78 ( // @[package.scala 93:22:@11431.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_79 ( // @[package.scala 93:22:@11439.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_80 ( // @[package.scala 93:22:@11479.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_81 ( // @[package.scala 93:22:@11487.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_82 ( // @[package.scala 93:22:@11495.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_83 ( // @[package.scala 93:22:@11503.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_84 ( // @[package.scala 93:22:@11511.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_85 ( // @[package.scala 93:22:@11519.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_86 ( // @[package.scala 93:22:@11527.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_87 ( // @[package.scala 93:22:@11535.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_88 ( // @[package.scala 93:22:@11575.4]
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_89 ( // @[package.scala 93:22:@11583.4]
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_90 ( // @[package.scala 93:22:@11591.4]
    .clock(RetimeWrapper_90_clock),
    .reset(RetimeWrapper_90_reset),
    .io_flow(RetimeWrapper_90_io_flow),
    .io_in(RetimeWrapper_90_io_in),
    .io_out(RetimeWrapper_90_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_91 ( // @[package.scala 93:22:@11599.4]
    .clock(RetimeWrapper_91_clock),
    .reset(RetimeWrapper_91_reset),
    .io_flow(RetimeWrapper_91_io_flow),
    .io_in(RetimeWrapper_91_io_in),
    .io_out(RetimeWrapper_91_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_92 ( // @[package.scala 93:22:@11607.4]
    .clock(RetimeWrapper_92_clock),
    .reset(RetimeWrapper_92_reset),
    .io_flow(RetimeWrapper_92_io_flow),
    .io_in(RetimeWrapper_92_io_in),
    .io_out(RetimeWrapper_92_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_93 ( // @[package.scala 93:22:@11615.4]
    .clock(RetimeWrapper_93_clock),
    .reset(RetimeWrapper_93_reset),
    .io_flow(RetimeWrapper_93_io_flow),
    .io_in(RetimeWrapper_93_io_in),
    .io_out(RetimeWrapper_93_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_94 ( // @[package.scala 93:22:@11623.4]
    .clock(RetimeWrapper_94_clock),
    .reset(RetimeWrapper_94_reset),
    .io_flow(RetimeWrapper_94_io_flow),
    .io_in(RetimeWrapper_94_io_in),
    .io_out(RetimeWrapper_94_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_95 ( // @[package.scala 93:22:@11631.4]
    .clock(RetimeWrapper_95_clock),
    .reset(RetimeWrapper_95_reset),
    .io_flow(RetimeWrapper_95_io_flow),
    .io_in(RetimeWrapper_95_io_in),
    .io_out(RetimeWrapper_95_io_out)
  );
  assign _T_444 = io_wPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@9310.4]
  assign _T_446 = io_wPort_0_banks_1 == 3'h0; // @[MemPrimitives.scala 82:210:@9311.4]
  assign _T_447 = _T_444 & _T_446; // @[MemPrimitives.scala 82:228:@9312.4]
  assign _T_448 = io_wPort_0_en_0 & _T_447; // @[MemPrimitives.scala 83:102:@9313.4]
  assign _T_450 = {_T_448,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9315.4]
  assign _T_455 = io_wPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@9322.4]
  assign _T_457 = io_wPort_1_banks_1 == 3'h1; // @[MemPrimitives.scala 82:210:@9323.4]
  assign _T_458 = _T_455 & _T_457; // @[MemPrimitives.scala 82:228:@9324.4]
  assign _T_459 = io_wPort_1_en_0 & _T_458; // @[MemPrimitives.scala 83:102:@9325.4]
  assign _T_461 = {_T_459,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@9327.4]
  assign _T_468 = io_wPort_0_banks_1 == 3'h2; // @[MemPrimitives.scala 82:210:@9335.4]
  assign _T_469 = _T_444 & _T_468; // @[MemPrimitives.scala 82:228:@9336.4]
  assign _T_470 = io_wPort_0_en_0 & _T_469; // @[MemPrimitives.scala 83:102:@9337.4]
  assign _T_472 = {_T_470,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9339.4]
  assign _T_479 = io_wPort_1_banks_1 == 3'h3; // @[MemPrimitives.scala 82:210:@9347.4]
  assign _T_480 = _T_455 & _T_479; // @[MemPrimitives.scala 82:228:@9348.4]
  assign _T_481 = io_wPort_1_en_0 & _T_480; // @[MemPrimitives.scala 83:102:@9349.4]
  assign _T_483 = {_T_481,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@9351.4]
  assign _T_488 = io_wPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@9358.4]
  assign _T_491 = _T_488 & _T_446; // @[MemPrimitives.scala 82:228:@9360.4]
  assign _T_492 = io_wPort_0_en_0 & _T_491; // @[MemPrimitives.scala 83:102:@9361.4]
  assign _T_494 = {_T_492,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9363.4]
  assign _T_499 = io_wPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@9370.4]
  assign _T_502 = _T_499 & _T_457; // @[MemPrimitives.scala 82:228:@9372.4]
  assign _T_503 = io_wPort_1_en_0 & _T_502; // @[MemPrimitives.scala 83:102:@9373.4]
  assign _T_505 = {_T_503,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@9375.4]
  assign _T_513 = _T_488 & _T_468; // @[MemPrimitives.scala 82:228:@9384.4]
  assign _T_514 = io_wPort_0_en_0 & _T_513; // @[MemPrimitives.scala 83:102:@9385.4]
  assign _T_516 = {_T_514,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9387.4]
  assign _T_524 = _T_499 & _T_479; // @[MemPrimitives.scala 82:228:@9396.4]
  assign _T_525 = io_wPort_1_en_0 & _T_524; // @[MemPrimitives.scala 83:102:@9397.4]
  assign _T_527 = {_T_525,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@9399.4]
  assign _T_532 = io_wPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@9406.4]
  assign _T_535 = _T_532 & _T_446; // @[MemPrimitives.scala 82:228:@9408.4]
  assign _T_536 = io_wPort_0_en_0 & _T_535; // @[MemPrimitives.scala 83:102:@9409.4]
  assign _T_538 = {_T_536,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9411.4]
  assign _T_543 = io_wPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@9418.4]
  assign _T_546 = _T_543 & _T_457; // @[MemPrimitives.scala 82:228:@9420.4]
  assign _T_547 = io_wPort_1_en_0 & _T_546; // @[MemPrimitives.scala 83:102:@9421.4]
  assign _T_549 = {_T_547,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@9423.4]
  assign _T_557 = _T_532 & _T_468; // @[MemPrimitives.scala 82:228:@9432.4]
  assign _T_558 = io_wPort_0_en_0 & _T_557; // @[MemPrimitives.scala 83:102:@9433.4]
  assign _T_560 = {_T_558,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9435.4]
  assign _T_568 = _T_543 & _T_479; // @[MemPrimitives.scala 82:228:@9444.4]
  assign _T_569 = io_wPort_1_en_0 & _T_568; // @[MemPrimitives.scala 83:102:@9445.4]
  assign _T_571 = {_T_569,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@9447.4]
  assign _T_576 = io_wPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@9454.4]
  assign _T_579 = _T_576 & _T_446; // @[MemPrimitives.scala 82:228:@9456.4]
  assign _T_580 = io_wPort_0_en_0 & _T_579; // @[MemPrimitives.scala 83:102:@9457.4]
  assign _T_582 = {_T_580,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9459.4]
  assign _T_587 = io_wPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@9466.4]
  assign _T_590 = _T_587 & _T_457; // @[MemPrimitives.scala 82:228:@9468.4]
  assign _T_591 = io_wPort_1_en_0 & _T_590; // @[MemPrimitives.scala 83:102:@9469.4]
  assign _T_593 = {_T_591,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@9471.4]
  assign _T_601 = _T_576 & _T_468; // @[MemPrimitives.scala 82:228:@9480.4]
  assign _T_602 = io_wPort_0_en_0 & _T_601; // @[MemPrimitives.scala 83:102:@9481.4]
  assign _T_604 = {_T_602,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9483.4]
  assign _T_612 = _T_587 & _T_479; // @[MemPrimitives.scala 82:228:@9492.4]
  assign _T_613 = io_wPort_1_en_0 & _T_612; // @[MemPrimitives.scala 83:102:@9493.4]
  assign _T_615 = {_T_613,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@9495.4]
  assign _T_620 = io_rPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9502.4]
  assign _T_622 = io_rPort_2_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@9503.4]
  assign _T_623 = _T_620 & _T_622; // @[MemPrimitives.scala 110:228:@9504.4]
  assign _T_626 = io_rPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9506.4]
  assign _T_628 = io_rPort_3_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@9507.4]
  assign _T_629 = _T_626 & _T_628; // @[MemPrimitives.scala 110:228:@9508.4]
  assign _T_632 = io_rPort_6_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9510.4]
  assign _T_634 = io_rPort_6_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@9511.4]
  assign _T_635 = _T_632 & _T_634; // @[MemPrimitives.scala 110:228:@9512.4]
  assign _T_638 = io_rPort_7_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9514.4]
  assign _T_640 = io_rPort_7_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@9515.4]
  assign _T_641 = _T_638 & _T_640; // @[MemPrimitives.scala 110:228:@9516.4]
  assign _T_644 = io_rPort_9_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9518.4]
  assign _T_646 = io_rPort_9_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@9519.4]
  assign _T_647 = _T_644 & _T_646; // @[MemPrimitives.scala 110:228:@9520.4]
  assign _T_650 = io_rPort_10_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9522.4]
  assign _T_652 = io_rPort_10_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@9523.4]
  assign _T_653 = _T_650 & _T_652; // @[MemPrimitives.scala 110:228:@9524.4]
  assign _T_655 = StickySelects_io_outs_0; // @[MemPrimitives.scala 123:41:@9535.4]
  assign _T_656 = StickySelects_io_outs_1; // @[MemPrimitives.scala 123:41:@9536.4]
  assign _T_657 = StickySelects_io_outs_2; // @[MemPrimitives.scala 123:41:@9537.4]
  assign _T_658 = StickySelects_io_outs_3; // @[MemPrimitives.scala 123:41:@9538.4]
  assign _T_659 = StickySelects_io_outs_4; // @[MemPrimitives.scala 123:41:@9539.4]
  assign _T_660 = StickySelects_io_outs_5; // @[MemPrimitives.scala 123:41:@9540.4]
  assign _T_662 = {_T_655,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@9542.4]
  assign _T_664 = {_T_656,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@9544.4]
  assign _T_666 = {_T_657,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@9546.4]
  assign _T_668 = {_T_658,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@9548.4]
  assign _T_670 = {_T_659,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@9550.4]
  assign _T_672 = {_T_660,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@9552.4]
  assign _T_673 = _T_659 ? _T_670 : _T_672; // @[Mux.scala 31:69:@9553.4]
  assign _T_674 = _T_658 ? _T_668 : _T_673; // @[Mux.scala 31:69:@9554.4]
  assign _T_675 = _T_657 ? _T_666 : _T_674; // @[Mux.scala 31:69:@9555.4]
  assign _T_676 = _T_656 ? _T_664 : _T_675; // @[Mux.scala 31:69:@9556.4]
  assign _T_677 = _T_655 ? _T_662 : _T_676; // @[Mux.scala 31:69:@9557.4]
  assign _T_682 = io_rPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9564.4]
  assign _T_684 = io_rPort_0_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@9565.4]
  assign _T_685 = _T_682 & _T_684; // @[MemPrimitives.scala 110:228:@9566.4]
  assign _T_688 = io_rPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9568.4]
  assign _T_690 = io_rPort_1_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@9569.4]
  assign _T_691 = _T_688 & _T_690; // @[MemPrimitives.scala 110:228:@9570.4]
  assign _T_694 = io_rPort_4_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9572.4]
  assign _T_696 = io_rPort_4_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@9573.4]
  assign _T_697 = _T_694 & _T_696; // @[MemPrimitives.scala 110:228:@9574.4]
  assign _T_700 = io_rPort_5_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9576.4]
  assign _T_702 = io_rPort_5_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@9577.4]
  assign _T_703 = _T_700 & _T_702; // @[MemPrimitives.scala 110:228:@9578.4]
  assign _T_706 = io_rPort_8_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9580.4]
  assign _T_708 = io_rPort_8_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@9581.4]
  assign _T_709 = _T_706 & _T_708; // @[MemPrimitives.scala 110:228:@9582.4]
  assign _T_712 = io_rPort_11_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9584.4]
  assign _T_714 = io_rPort_11_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@9585.4]
  assign _T_715 = _T_712 & _T_714; // @[MemPrimitives.scala 110:228:@9586.4]
  assign _T_717 = StickySelects_1_io_outs_0; // @[MemPrimitives.scala 123:41:@9597.4]
  assign _T_718 = StickySelects_1_io_outs_1; // @[MemPrimitives.scala 123:41:@9598.4]
  assign _T_719 = StickySelects_1_io_outs_2; // @[MemPrimitives.scala 123:41:@9599.4]
  assign _T_720 = StickySelects_1_io_outs_3; // @[MemPrimitives.scala 123:41:@9600.4]
  assign _T_721 = StickySelects_1_io_outs_4; // @[MemPrimitives.scala 123:41:@9601.4]
  assign _T_722 = StickySelects_1_io_outs_5; // @[MemPrimitives.scala 123:41:@9602.4]
  assign _T_724 = {_T_717,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@9604.4]
  assign _T_726 = {_T_718,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@9606.4]
  assign _T_728 = {_T_719,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@9608.4]
  assign _T_730 = {_T_720,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@9610.4]
  assign _T_732 = {_T_721,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@9612.4]
  assign _T_734 = {_T_722,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@9614.4]
  assign _T_735 = _T_721 ? _T_732 : _T_734; // @[Mux.scala 31:69:@9615.4]
  assign _T_736 = _T_720 ? _T_730 : _T_735; // @[Mux.scala 31:69:@9616.4]
  assign _T_737 = _T_719 ? _T_728 : _T_736; // @[Mux.scala 31:69:@9617.4]
  assign _T_738 = _T_718 ? _T_726 : _T_737; // @[Mux.scala 31:69:@9618.4]
  assign _T_739 = _T_717 ? _T_724 : _T_738; // @[Mux.scala 31:69:@9619.4]
  assign _T_746 = io_rPort_2_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@9627.4]
  assign _T_747 = _T_620 & _T_746; // @[MemPrimitives.scala 110:228:@9628.4]
  assign _T_752 = io_rPort_3_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@9631.4]
  assign _T_753 = _T_626 & _T_752; // @[MemPrimitives.scala 110:228:@9632.4]
  assign _T_758 = io_rPort_6_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@9635.4]
  assign _T_759 = _T_632 & _T_758; // @[MemPrimitives.scala 110:228:@9636.4]
  assign _T_764 = io_rPort_7_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@9639.4]
  assign _T_765 = _T_638 & _T_764; // @[MemPrimitives.scala 110:228:@9640.4]
  assign _T_770 = io_rPort_9_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@9643.4]
  assign _T_771 = _T_644 & _T_770; // @[MemPrimitives.scala 110:228:@9644.4]
  assign _T_776 = io_rPort_10_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@9647.4]
  assign _T_777 = _T_650 & _T_776; // @[MemPrimitives.scala 110:228:@9648.4]
  assign _T_779 = StickySelects_2_io_outs_0; // @[MemPrimitives.scala 123:41:@9659.4]
  assign _T_780 = StickySelects_2_io_outs_1; // @[MemPrimitives.scala 123:41:@9660.4]
  assign _T_781 = StickySelects_2_io_outs_2; // @[MemPrimitives.scala 123:41:@9661.4]
  assign _T_782 = StickySelects_2_io_outs_3; // @[MemPrimitives.scala 123:41:@9662.4]
  assign _T_783 = StickySelects_2_io_outs_4; // @[MemPrimitives.scala 123:41:@9663.4]
  assign _T_784 = StickySelects_2_io_outs_5; // @[MemPrimitives.scala 123:41:@9664.4]
  assign _T_786 = {_T_779,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@9666.4]
  assign _T_788 = {_T_780,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@9668.4]
  assign _T_790 = {_T_781,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@9670.4]
  assign _T_792 = {_T_782,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@9672.4]
  assign _T_794 = {_T_783,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@9674.4]
  assign _T_796 = {_T_784,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@9676.4]
  assign _T_797 = _T_783 ? _T_794 : _T_796; // @[Mux.scala 31:69:@9677.4]
  assign _T_798 = _T_782 ? _T_792 : _T_797; // @[Mux.scala 31:69:@9678.4]
  assign _T_799 = _T_781 ? _T_790 : _T_798; // @[Mux.scala 31:69:@9679.4]
  assign _T_800 = _T_780 ? _T_788 : _T_799; // @[Mux.scala 31:69:@9680.4]
  assign _T_801 = _T_779 ? _T_786 : _T_800; // @[Mux.scala 31:69:@9681.4]
  assign _T_808 = io_rPort_0_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@9689.4]
  assign _T_809 = _T_682 & _T_808; // @[MemPrimitives.scala 110:228:@9690.4]
  assign _T_814 = io_rPort_1_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@9693.4]
  assign _T_815 = _T_688 & _T_814; // @[MemPrimitives.scala 110:228:@9694.4]
  assign _T_820 = io_rPort_4_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@9697.4]
  assign _T_821 = _T_694 & _T_820; // @[MemPrimitives.scala 110:228:@9698.4]
  assign _T_826 = io_rPort_5_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@9701.4]
  assign _T_827 = _T_700 & _T_826; // @[MemPrimitives.scala 110:228:@9702.4]
  assign _T_832 = io_rPort_8_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@9705.4]
  assign _T_833 = _T_706 & _T_832; // @[MemPrimitives.scala 110:228:@9706.4]
  assign _T_838 = io_rPort_11_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@9709.4]
  assign _T_839 = _T_712 & _T_838; // @[MemPrimitives.scala 110:228:@9710.4]
  assign _T_841 = StickySelects_3_io_outs_0; // @[MemPrimitives.scala 123:41:@9721.4]
  assign _T_842 = StickySelects_3_io_outs_1; // @[MemPrimitives.scala 123:41:@9722.4]
  assign _T_843 = StickySelects_3_io_outs_2; // @[MemPrimitives.scala 123:41:@9723.4]
  assign _T_844 = StickySelects_3_io_outs_3; // @[MemPrimitives.scala 123:41:@9724.4]
  assign _T_845 = StickySelects_3_io_outs_4; // @[MemPrimitives.scala 123:41:@9725.4]
  assign _T_846 = StickySelects_3_io_outs_5; // @[MemPrimitives.scala 123:41:@9726.4]
  assign _T_848 = {_T_841,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@9728.4]
  assign _T_850 = {_T_842,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@9730.4]
  assign _T_852 = {_T_843,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@9732.4]
  assign _T_854 = {_T_844,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@9734.4]
  assign _T_856 = {_T_845,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@9736.4]
  assign _T_858 = {_T_846,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@9738.4]
  assign _T_859 = _T_845 ? _T_856 : _T_858; // @[Mux.scala 31:69:@9739.4]
  assign _T_860 = _T_844 ? _T_854 : _T_859; // @[Mux.scala 31:69:@9740.4]
  assign _T_861 = _T_843 ? _T_852 : _T_860; // @[Mux.scala 31:69:@9741.4]
  assign _T_862 = _T_842 ? _T_850 : _T_861; // @[Mux.scala 31:69:@9742.4]
  assign _T_863 = _T_841 ? _T_848 : _T_862; // @[Mux.scala 31:69:@9743.4]
  assign _T_868 = io_rPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9750.4]
  assign _T_871 = _T_868 & _T_622; // @[MemPrimitives.scala 110:228:@9752.4]
  assign _T_874 = io_rPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9754.4]
  assign _T_877 = _T_874 & _T_628; // @[MemPrimitives.scala 110:228:@9756.4]
  assign _T_880 = io_rPort_6_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9758.4]
  assign _T_883 = _T_880 & _T_634; // @[MemPrimitives.scala 110:228:@9760.4]
  assign _T_886 = io_rPort_7_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9762.4]
  assign _T_889 = _T_886 & _T_640; // @[MemPrimitives.scala 110:228:@9764.4]
  assign _T_892 = io_rPort_9_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9766.4]
  assign _T_895 = _T_892 & _T_646; // @[MemPrimitives.scala 110:228:@9768.4]
  assign _T_898 = io_rPort_10_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9770.4]
  assign _T_901 = _T_898 & _T_652; // @[MemPrimitives.scala 110:228:@9772.4]
  assign _T_903 = StickySelects_4_io_outs_0; // @[MemPrimitives.scala 123:41:@9783.4]
  assign _T_904 = StickySelects_4_io_outs_1; // @[MemPrimitives.scala 123:41:@9784.4]
  assign _T_905 = StickySelects_4_io_outs_2; // @[MemPrimitives.scala 123:41:@9785.4]
  assign _T_906 = StickySelects_4_io_outs_3; // @[MemPrimitives.scala 123:41:@9786.4]
  assign _T_907 = StickySelects_4_io_outs_4; // @[MemPrimitives.scala 123:41:@9787.4]
  assign _T_908 = StickySelects_4_io_outs_5; // @[MemPrimitives.scala 123:41:@9788.4]
  assign _T_910 = {_T_903,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@9790.4]
  assign _T_912 = {_T_904,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@9792.4]
  assign _T_914 = {_T_905,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@9794.4]
  assign _T_916 = {_T_906,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@9796.4]
  assign _T_918 = {_T_907,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@9798.4]
  assign _T_920 = {_T_908,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@9800.4]
  assign _T_921 = _T_907 ? _T_918 : _T_920; // @[Mux.scala 31:69:@9801.4]
  assign _T_922 = _T_906 ? _T_916 : _T_921; // @[Mux.scala 31:69:@9802.4]
  assign _T_923 = _T_905 ? _T_914 : _T_922; // @[Mux.scala 31:69:@9803.4]
  assign _T_924 = _T_904 ? _T_912 : _T_923; // @[Mux.scala 31:69:@9804.4]
  assign _T_925 = _T_903 ? _T_910 : _T_924; // @[Mux.scala 31:69:@9805.4]
  assign _T_930 = io_rPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9812.4]
  assign _T_933 = _T_930 & _T_684; // @[MemPrimitives.scala 110:228:@9814.4]
  assign _T_936 = io_rPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9816.4]
  assign _T_939 = _T_936 & _T_690; // @[MemPrimitives.scala 110:228:@9818.4]
  assign _T_942 = io_rPort_4_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9820.4]
  assign _T_945 = _T_942 & _T_696; // @[MemPrimitives.scala 110:228:@9822.4]
  assign _T_948 = io_rPort_5_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9824.4]
  assign _T_951 = _T_948 & _T_702; // @[MemPrimitives.scala 110:228:@9826.4]
  assign _T_954 = io_rPort_8_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9828.4]
  assign _T_957 = _T_954 & _T_708; // @[MemPrimitives.scala 110:228:@9830.4]
  assign _T_960 = io_rPort_11_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9832.4]
  assign _T_963 = _T_960 & _T_714; // @[MemPrimitives.scala 110:228:@9834.4]
  assign _T_965 = StickySelects_5_io_outs_0; // @[MemPrimitives.scala 123:41:@9845.4]
  assign _T_966 = StickySelects_5_io_outs_1; // @[MemPrimitives.scala 123:41:@9846.4]
  assign _T_967 = StickySelects_5_io_outs_2; // @[MemPrimitives.scala 123:41:@9847.4]
  assign _T_968 = StickySelects_5_io_outs_3; // @[MemPrimitives.scala 123:41:@9848.4]
  assign _T_969 = StickySelects_5_io_outs_4; // @[MemPrimitives.scala 123:41:@9849.4]
  assign _T_970 = StickySelects_5_io_outs_5; // @[MemPrimitives.scala 123:41:@9850.4]
  assign _T_972 = {_T_965,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@9852.4]
  assign _T_974 = {_T_966,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@9854.4]
  assign _T_976 = {_T_967,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@9856.4]
  assign _T_978 = {_T_968,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@9858.4]
  assign _T_980 = {_T_969,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@9860.4]
  assign _T_982 = {_T_970,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@9862.4]
  assign _T_983 = _T_969 ? _T_980 : _T_982; // @[Mux.scala 31:69:@9863.4]
  assign _T_984 = _T_968 ? _T_978 : _T_983; // @[Mux.scala 31:69:@9864.4]
  assign _T_985 = _T_967 ? _T_976 : _T_984; // @[Mux.scala 31:69:@9865.4]
  assign _T_986 = _T_966 ? _T_974 : _T_985; // @[Mux.scala 31:69:@9866.4]
  assign _T_987 = _T_965 ? _T_972 : _T_986; // @[Mux.scala 31:69:@9867.4]
  assign _T_995 = _T_868 & _T_746; // @[MemPrimitives.scala 110:228:@9876.4]
  assign _T_1001 = _T_874 & _T_752; // @[MemPrimitives.scala 110:228:@9880.4]
  assign _T_1007 = _T_880 & _T_758; // @[MemPrimitives.scala 110:228:@9884.4]
  assign _T_1013 = _T_886 & _T_764; // @[MemPrimitives.scala 110:228:@9888.4]
  assign _T_1019 = _T_892 & _T_770; // @[MemPrimitives.scala 110:228:@9892.4]
  assign _T_1025 = _T_898 & _T_776; // @[MemPrimitives.scala 110:228:@9896.4]
  assign _T_1027 = StickySelects_6_io_outs_0; // @[MemPrimitives.scala 123:41:@9907.4]
  assign _T_1028 = StickySelects_6_io_outs_1; // @[MemPrimitives.scala 123:41:@9908.4]
  assign _T_1029 = StickySelects_6_io_outs_2; // @[MemPrimitives.scala 123:41:@9909.4]
  assign _T_1030 = StickySelects_6_io_outs_3; // @[MemPrimitives.scala 123:41:@9910.4]
  assign _T_1031 = StickySelects_6_io_outs_4; // @[MemPrimitives.scala 123:41:@9911.4]
  assign _T_1032 = StickySelects_6_io_outs_5; // @[MemPrimitives.scala 123:41:@9912.4]
  assign _T_1034 = {_T_1027,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@9914.4]
  assign _T_1036 = {_T_1028,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@9916.4]
  assign _T_1038 = {_T_1029,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@9918.4]
  assign _T_1040 = {_T_1030,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@9920.4]
  assign _T_1042 = {_T_1031,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@9922.4]
  assign _T_1044 = {_T_1032,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@9924.4]
  assign _T_1045 = _T_1031 ? _T_1042 : _T_1044; // @[Mux.scala 31:69:@9925.4]
  assign _T_1046 = _T_1030 ? _T_1040 : _T_1045; // @[Mux.scala 31:69:@9926.4]
  assign _T_1047 = _T_1029 ? _T_1038 : _T_1046; // @[Mux.scala 31:69:@9927.4]
  assign _T_1048 = _T_1028 ? _T_1036 : _T_1047; // @[Mux.scala 31:69:@9928.4]
  assign _T_1049 = _T_1027 ? _T_1034 : _T_1048; // @[Mux.scala 31:69:@9929.4]
  assign _T_1057 = _T_930 & _T_808; // @[MemPrimitives.scala 110:228:@9938.4]
  assign _T_1063 = _T_936 & _T_814; // @[MemPrimitives.scala 110:228:@9942.4]
  assign _T_1069 = _T_942 & _T_820; // @[MemPrimitives.scala 110:228:@9946.4]
  assign _T_1075 = _T_948 & _T_826; // @[MemPrimitives.scala 110:228:@9950.4]
  assign _T_1081 = _T_954 & _T_832; // @[MemPrimitives.scala 110:228:@9954.4]
  assign _T_1087 = _T_960 & _T_838; // @[MemPrimitives.scala 110:228:@9958.4]
  assign _T_1089 = StickySelects_7_io_outs_0; // @[MemPrimitives.scala 123:41:@9969.4]
  assign _T_1090 = StickySelects_7_io_outs_1; // @[MemPrimitives.scala 123:41:@9970.4]
  assign _T_1091 = StickySelects_7_io_outs_2; // @[MemPrimitives.scala 123:41:@9971.4]
  assign _T_1092 = StickySelects_7_io_outs_3; // @[MemPrimitives.scala 123:41:@9972.4]
  assign _T_1093 = StickySelects_7_io_outs_4; // @[MemPrimitives.scala 123:41:@9973.4]
  assign _T_1094 = StickySelects_7_io_outs_5; // @[MemPrimitives.scala 123:41:@9974.4]
  assign _T_1096 = {_T_1089,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@9976.4]
  assign _T_1098 = {_T_1090,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@9978.4]
  assign _T_1100 = {_T_1091,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@9980.4]
  assign _T_1102 = {_T_1092,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@9982.4]
  assign _T_1104 = {_T_1093,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@9984.4]
  assign _T_1106 = {_T_1094,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@9986.4]
  assign _T_1107 = _T_1093 ? _T_1104 : _T_1106; // @[Mux.scala 31:69:@9987.4]
  assign _T_1108 = _T_1092 ? _T_1102 : _T_1107; // @[Mux.scala 31:69:@9988.4]
  assign _T_1109 = _T_1091 ? _T_1100 : _T_1108; // @[Mux.scala 31:69:@9989.4]
  assign _T_1110 = _T_1090 ? _T_1098 : _T_1109; // @[Mux.scala 31:69:@9990.4]
  assign _T_1111 = _T_1089 ? _T_1096 : _T_1110; // @[Mux.scala 31:69:@9991.4]
  assign _T_1116 = io_rPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@9998.4]
  assign _T_1119 = _T_1116 & _T_622; // @[MemPrimitives.scala 110:228:@10000.4]
  assign _T_1122 = io_rPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10002.4]
  assign _T_1125 = _T_1122 & _T_628; // @[MemPrimitives.scala 110:228:@10004.4]
  assign _T_1128 = io_rPort_6_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10006.4]
  assign _T_1131 = _T_1128 & _T_634; // @[MemPrimitives.scala 110:228:@10008.4]
  assign _T_1134 = io_rPort_7_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10010.4]
  assign _T_1137 = _T_1134 & _T_640; // @[MemPrimitives.scala 110:228:@10012.4]
  assign _T_1140 = io_rPort_9_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10014.4]
  assign _T_1143 = _T_1140 & _T_646; // @[MemPrimitives.scala 110:228:@10016.4]
  assign _T_1146 = io_rPort_10_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10018.4]
  assign _T_1149 = _T_1146 & _T_652; // @[MemPrimitives.scala 110:228:@10020.4]
  assign _T_1151 = StickySelects_8_io_outs_0; // @[MemPrimitives.scala 123:41:@10031.4]
  assign _T_1152 = StickySelects_8_io_outs_1; // @[MemPrimitives.scala 123:41:@10032.4]
  assign _T_1153 = StickySelects_8_io_outs_2; // @[MemPrimitives.scala 123:41:@10033.4]
  assign _T_1154 = StickySelects_8_io_outs_3; // @[MemPrimitives.scala 123:41:@10034.4]
  assign _T_1155 = StickySelects_8_io_outs_4; // @[MemPrimitives.scala 123:41:@10035.4]
  assign _T_1156 = StickySelects_8_io_outs_5; // @[MemPrimitives.scala 123:41:@10036.4]
  assign _T_1158 = {_T_1151,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@10038.4]
  assign _T_1160 = {_T_1152,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@10040.4]
  assign _T_1162 = {_T_1153,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@10042.4]
  assign _T_1164 = {_T_1154,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@10044.4]
  assign _T_1166 = {_T_1155,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@10046.4]
  assign _T_1168 = {_T_1156,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@10048.4]
  assign _T_1169 = _T_1155 ? _T_1166 : _T_1168; // @[Mux.scala 31:69:@10049.4]
  assign _T_1170 = _T_1154 ? _T_1164 : _T_1169; // @[Mux.scala 31:69:@10050.4]
  assign _T_1171 = _T_1153 ? _T_1162 : _T_1170; // @[Mux.scala 31:69:@10051.4]
  assign _T_1172 = _T_1152 ? _T_1160 : _T_1171; // @[Mux.scala 31:69:@10052.4]
  assign _T_1173 = _T_1151 ? _T_1158 : _T_1172; // @[Mux.scala 31:69:@10053.4]
  assign _T_1178 = io_rPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10060.4]
  assign _T_1181 = _T_1178 & _T_684; // @[MemPrimitives.scala 110:228:@10062.4]
  assign _T_1184 = io_rPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10064.4]
  assign _T_1187 = _T_1184 & _T_690; // @[MemPrimitives.scala 110:228:@10066.4]
  assign _T_1190 = io_rPort_4_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10068.4]
  assign _T_1193 = _T_1190 & _T_696; // @[MemPrimitives.scala 110:228:@10070.4]
  assign _T_1196 = io_rPort_5_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10072.4]
  assign _T_1199 = _T_1196 & _T_702; // @[MemPrimitives.scala 110:228:@10074.4]
  assign _T_1202 = io_rPort_8_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10076.4]
  assign _T_1205 = _T_1202 & _T_708; // @[MemPrimitives.scala 110:228:@10078.4]
  assign _T_1208 = io_rPort_11_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10080.4]
  assign _T_1211 = _T_1208 & _T_714; // @[MemPrimitives.scala 110:228:@10082.4]
  assign _T_1213 = StickySelects_9_io_outs_0; // @[MemPrimitives.scala 123:41:@10093.4]
  assign _T_1214 = StickySelects_9_io_outs_1; // @[MemPrimitives.scala 123:41:@10094.4]
  assign _T_1215 = StickySelects_9_io_outs_2; // @[MemPrimitives.scala 123:41:@10095.4]
  assign _T_1216 = StickySelects_9_io_outs_3; // @[MemPrimitives.scala 123:41:@10096.4]
  assign _T_1217 = StickySelects_9_io_outs_4; // @[MemPrimitives.scala 123:41:@10097.4]
  assign _T_1218 = StickySelects_9_io_outs_5; // @[MemPrimitives.scala 123:41:@10098.4]
  assign _T_1220 = {_T_1213,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@10100.4]
  assign _T_1222 = {_T_1214,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@10102.4]
  assign _T_1224 = {_T_1215,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@10104.4]
  assign _T_1226 = {_T_1216,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@10106.4]
  assign _T_1228 = {_T_1217,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@10108.4]
  assign _T_1230 = {_T_1218,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@10110.4]
  assign _T_1231 = _T_1217 ? _T_1228 : _T_1230; // @[Mux.scala 31:69:@10111.4]
  assign _T_1232 = _T_1216 ? _T_1226 : _T_1231; // @[Mux.scala 31:69:@10112.4]
  assign _T_1233 = _T_1215 ? _T_1224 : _T_1232; // @[Mux.scala 31:69:@10113.4]
  assign _T_1234 = _T_1214 ? _T_1222 : _T_1233; // @[Mux.scala 31:69:@10114.4]
  assign _T_1235 = _T_1213 ? _T_1220 : _T_1234; // @[Mux.scala 31:69:@10115.4]
  assign _T_1243 = _T_1116 & _T_746; // @[MemPrimitives.scala 110:228:@10124.4]
  assign _T_1249 = _T_1122 & _T_752; // @[MemPrimitives.scala 110:228:@10128.4]
  assign _T_1255 = _T_1128 & _T_758; // @[MemPrimitives.scala 110:228:@10132.4]
  assign _T_1261 = _T_1134 & _T_764; // @[MemPrimitives.scala 110:228:@10136.4]
  assign _T_1267 = _T_1140 & _T_770; // @[MemPrimitives.scala 110:228:@10140.4]
  assign _T_1273 = _T_1146 & _T_776; // @[MemPrimitives.scala 110:228:@10144.4]
  assign _T_1275 = StickySelects_10_io_outs_0; // @[MemPrimitives.scala 123:41:@10155.4]
  assign _T_1276 = StickySelects_10_io_outs_1; // @[MemPrimitives.scala 123:41:@10156.4]
  assign _T_1277 = StickySelects_10_io_outs_2; // @[MemPrimitives.scala 123:41:@10157.4]
  assign _T_1278 = StickySelects_10_io_outs_3; // @[MemPrimitives.scala 123:41:@10158.4]
  assign _T_1279 = StickySelects_10_io_outs_4; // @[MemPrimitives.scala 123:41:@10159.4]
  assign _T_1280 = StickySelects_10_io_outs_5; // @[MemPrimitives.scala 123:41:@10160.4]
  assign _T_1282 = {_T_1275,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@10162.4]
  assign _T_1284 = {_T_1276,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@10164.4]
  assign _T_1286 = {_T_1277,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@10166.4]
  assign _T_1288 = {_T_1278,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@10168.4]
  assign _T_1290 = {_T_1279,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@10170.4]
  assign _T_1292 = {_T_1280,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@10172.4]
  assign _T_1293 = _T_1279 ? _T_1290 : _T_1292; // @[Mux.scala 31:69:@10173.4]
  assign _T_1294 = _T_1278 ? _T_1288 : _T_1293; // @[Mux.scala 31:69:@10174.4]
  assign _T_1295 = _T_1277 ? _T_1286 : _T_1294; // @[Mux.scala 31:69:@10175.4]
  assign _T_1296 = _T_1276 ? _T_1284 : _T_1295; // @[Mux.scala 31:69:@10176.4]
  assign _T_1297 = _T_1275 ? _T_1282 : _T_1296; // @[Mux.scala 31:69:@10177.4]
  assign _T_1305 = _T_1178 & _T_808; // @[MemPrimitives.scala 110:228:@10186.4]
  assign _T_1311 = _T_1184 & _T_814; // @[MemPrimitives.scala 110:228:@10190.4]
  assign _T_1317 = _T_1190 & _T_820; // @[MemPrimitives.scala 110:228:@10194.4]
  assign _T_1323 = _T_1196 & _T_826; // @[MemPrimitives.scala 110:228:@10198.4]
  assign _T_1329 = _T_1202 & _T_832; // @[MemPrimitives.scala 110:228:@10202.4]
  assign _T_1335 = _T_1208 & _T_838; // @[MemPrimitives.scala 110:228:@10206.4]
  assign _T_1337 = StickySelects_11_io_outs_0; // @[MemPrimitives.scala 123:41:@10217.4]
  assign _T_1338 = StickySelects_11_io_outs_1; // @[MemPrimitives.scala 123:41:@10218.4]
  assign _T_1339 = StickySelects_11_io_outs_2; // @[MemPrimitives.scala 123:41:@10219.4]
  assign _T_1340 = StickySelects_11_io_outs_3; // @[MemPrimitives.scala 123:41:@10220.4]
  assign _T_1341 = StickySelects_11_io_outs_4; // @[MemPrimitives.scala 123:41:@10221.4]
  assign _T_1342 = StickySelects_11_io_outs_5; // @[MemPrimitives.scala 123:41:@10222.4]
  assign _T_1344 = {_T_1337,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@10224.4]
  assign _T_1346 = {_T_1338,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@10226.4]
  assign _T_1348 = {_T_1339,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@10228.4]
  assign _T_1350 = {_T_1340,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@10230.4]
  assign _T_1352 = {_T_1341,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@10232.4]
  assign _T_1354 = {_T_1342,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@10234.4]
  assign _T_1355 = _T_1341 ? _T_1352 : _T_1354; // @[Mux.scala 31:69:@10235.4]
  assign _T_1356 = _T_1340 ? _T_1350 : _T_1355; // @[Mux.scala 31:69:@10236.4]
  assign _T_1357 = _T_1339 ? _T_1348 : _T_1356; // @[Mux.scala 31:69:@10237.4]
  assign _T_1358 = _T_1338 ? _T_1346 : _T_1357; // @[Mux.scala 31:69:@10238.4]
  assign _T_1359 = _T_1337 ? _T_1344 : _T_1358; // @[Mux.scala 31:69:@10239.4]
  assign _T_1364 = io_rPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10246.4]
  assign _T_1367 = _T_1364 & _T_622; // @[MemPrimitives.scala 110:228:@10248.4]
  assign _T_1370 = io_rPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10250.4]
  assign _T_1373 = _T_1370 & _T_628; // @[MemPrimitives.scala 110:228:@10252.4]
  assign _T_1376 = io_rPort_6_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10254.4]
  assign _T_1379 = _T_1376 & _T_634; // @[MemPrimitives.scala 110:228:@10256.4]
  assign _T_1382 = io_rPort_7_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10258.4]
  assign _T_1385 = _T_1382 & _T_640; // @[MemPrimitives.scala 110:228:@10260.4]
  assign _T_1388 = io_rPort_9_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10262.4]
  assign _T_1391 = _T_1388 & _T_646; // @[MemPrimitives.scala 110:228:@10264.4]
  assign _T_1394 = io_rPort_10_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10266.4]
  assign _T_1397 = _T_1394 & _T_652; // @[MemPrimitives.scala 110:228:@10268.4]
  assign _T_1399 = StickySelects_12_io_outs_0; // @[MemPrimitives.scala 123:41:@10279.4]
  assign _T_1400 = StickySelects_12_io_outs_1; // @[MemPrimitives.scala 123:41:@10280.4]
  assign _T_1401 = StickySelects_12_io_outs_2; // @[MemPrimitives.scala 123:41:@10281.4]
  assign _T_1402 = StickySelects_12_io_outs_3; // @[MemPrimitives.scala 123:41:@10282.4]
  assign _T_1403 = StickySelects_12_io_outs_4; // @[MemPrimitives.scala 123:41:@10283.4]
  assign _T_1404 = StickySelects_12_io_outs_5; // @[MemPrimitives.scala 123:41:@10284.4]
  assign _T_1406 = {_T_1399,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@10286.4]
  assign _T_1408 = {_T_1400,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@10288.4]
  assign _T_1410 = {_T_1401,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@10290.4]
  assign _T_1412 = {_T_1402,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@10292.4]
  assign _T_1414 = {_T_1403,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@10294.4]
  assign _T_1416 = {_T_1404,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@10296.4]
  assign _T_1417 = _T_1403 ? _T_1414 : _T_1416; // @[Mux.scala 31:69:@10297.4]
  assign _T_1418 = _T_1402 ? _T_1412 : _T_1417; // @[Mux.scala 31:69:@10298.4]
  assign _T_1419 = _T_1401 ? _T_1410 : _T_1418; // @[Mux.scala 31:69:@10299.4]
  assign _T_1420 = _T_1400 ? _T_1408 : _T_1419; // @[Mux.scala 31:69:@10300.4]
  assign _T_1421 = _T_1399 ? _T_1406 : _T_1420; // @[Mux.scala 31:69:@10301.4]
  assign _T_1426 = io_rPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10308.4]
  assign _T_1429 = _T_1426 & _T_684; // @[MemPrimitives.scala 110:228:@10310.4]
  assign _T_1432 = io_rPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10312.4]
  assign _T_1435 = _T_1432 & _T_690; // @[MemPrimitives.scala 110:228:@10314.4]
  assign _T_1438 = io_rPort_4_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10316.4]
  assign _T_1441 = _T_1438 & _T_696; // @[MemPrimitives.scala 110:228:@10318.4]
  assign _T_1444 = io_rPort_5_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10320.4]
  assign _T_1447 = _T_1444 & _T_702; // @[MemPrimitives.scala 110:228:@10322.4]
  assign _T_1450 = io_rPort_8_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10324.4]
  assign _T_1453 = _T_1450 & _T_708; // @[MemPrimitives.scala 110:228:@10326.4]
  assign _T_1456 = io_rPort_11_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10328.4]
  assign _T_1459 = _T_1456 & _T_714; // @[MemPrimitives.scala 110:228:@10330.4]
  assign _T_1461 = StickySelects_13_io_outs_0; // @[MemPrimitives.scala 123:41:@10341.4]
  assign _T_1462 = StickySelects_13_io_outs_1; // @[MemPrimitives.scala 123:41:@10342.4]
  assign _T_1463 = StickySelects_13_io_outs_2; // @[MemPrimitives.scala 123:41:@10343.4]
  assign _T_1464 = StickySelects_13_io_outs_3; // @[MemPrimitives.scala 123:41:@10344.4]
  assign _T_1465 = StickySelects_13_io_outs_4; // @[MemPrimitives.scala 123:41:@10345.4]
  assign _T_1466 = StickySelects_13_io_outs_5; // @[MemPrimitives.scala 123:41:@10346.4]
  assign _T_1468 = {_T_1461,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@10348.4]
  assign _T_1470 = {_T_1462,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@10350.4]
  assign _T_1472 = {_T_1463,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@10352.4]
  assign _T_1474 = {_T_1464,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@10354.4]
  assign _T_1476 = {_T_1465,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@10356.4]
  assign _T_1478 = {_T_1466,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@10358.4]
  assign _T_1479 = _T_1465 ? _T_1476 : _T_1478; // @[Mux.scala 31:69:@10359.4]
  assign _T_1480 = _T_1464 ? _T_1474 : _T_1479; // @[Mux.scala 31:69:@10360.4]
  assign _T_1481 = _T_1463 ? _T_1472 : _T_1480; // @[Mux.scala 31:69:@10361.4]
  assign _T_1482 = _T_1462 ? _T_1470 : _T_1481; // @[Mux.scala 31:69:@10362.4]
  assign _T_1483 = _T_1461 ? _T_1468 : _T_1482; // @[Mux.scala 31:69:@10363.4]
  assign _T_1491 = _T_1364 & _T_746; // @[MemPrimitives.scala 110:228:@10372.4]
  assign _T_1497 = _T_1370 & _T_752; // @[MemPrimitives.scala 110:228:@10376.4]
  assign _T_1503 = _T_1376 & _T_758; // @[MemPrimitives.scala 110:228:@10380.4]
  assign _T_1509 = _T_1382 & _T_764; // @[MemPrimitives.scala 110:228:@10384.4]
  assign _T_1515 = _T_1388 & _T_770; // @[MemPrimitives.scala 110:228:@10388.4]
  assign _T_1521 = _T_1394 & _T_776; // @[MemPrimitives.scala 110:228:@10392.4]
  assign _T_1523 = StickySelects_14_io_outs_0; // @[MemPrimitives.scala 123:41:@10403.4]
  assign _T_1524 = StickySelects_14_io_outs_1; // @[MemPrimitives.scala 123:41:@10404.4]
  assign _T_1525 = StickySelects_14_io_outs_2; // @[MemPrimitives.scala 123:41:@10405.4]
  assign _T_1526 = StickySelects_14_io_outs_3; // @[MemPrimitives.scala 123:41:@10406.4]
  assign _T_1527 = StickySelects_14_io_outs_4; // @[MemPrimitives.scala 123:41:@10407.4]
  assign _T_1528 = StickySelects_14_io_outs_5; // @[MemPrimitives.scala 123:41:@10408.4]
  assign _T_1530 = {_T_1523,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@10410.4]
  assign _T_1532 = {_T_1524,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@10412.4]
  assign _T_1534 = {_T_1525,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@10414.4]
  assign _T_1536 = {_T_1526,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@10416.4]
  assign _T_1538 = {_T_1527,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@10418.4]
  assign _T_1540 = {_T_1528,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@10420.4]
  assign _T_1541 = _T_1527 ? _T_1538 : _T_1540; // @[Mux.scala 31:69:@10421.4]
  assign _T_1542 = _T_1526 ? _T_1536 : _T_1541; // @[Mux.scala 31:69:@10422.4]
  assign _T_1543 = _T_1525 ? _T_1534 : _T_1542; // @[Mux.scala 31:69:@10423.4]
  assign _T_1544 = _T_1524 ? _T_1532 : _T_1543; // @[Mux.scala 31:69:@10424.4]
  assign _T_1545 = _T_1523 ? _T_1530 : _T_1544; // @[Mux.scala 31:69:@10425.4]
  assign _T_1553 = _T_1426 & _T_808; // @[MemPrimitives.scala 110:228:@10434.4]
  assign _T_1559 = _T_1432 & _T_814; // @[MemPrimitives.scala 110:228:@10438.4]
  assign _T_1565 = _T_1438 & _T_820; // @[MemPrimitives.scala 110:228:@10442.4]
  assign _T_1571 = _T_1444 & _T_826; // @[MemPrimitives.scala 110:228:@10446.4]
  assign _T_1577 = _T_1450 & _T_832; // @[MemPrimitives.scala 110:228:@10450.4]
  assign _T_1583 = _T_1456 & _T_838; // @[MemPrimitives.scala 110:228:@10454.4]
  assign _T_1585 = StickySelects_15_io_outs_0; // @[MemPrimitives.scala 123:41:@10465.4]
  assign _T_1586 = StickySelects_15_io_outs_1; // @[MemPrimitives.scala 123:41:@10466.4]
  assign _T_1587 = StickySelects_15_io_outs_2; // @[MemPrimitives.scala 123:41:@10467.4]
  assign _T_1588 = StickySelects_15_io_outs_3; // @[MemPrimitives.scala 123:41:@10468.4]
  assign _T_1589 = StickySelects_15_io_outs_4; // @[MemPrimitives.scala 123:41:@10469.4]
  assign _T_1590 = StickySelects_15_io_outs_5; // @[MemPrimitives.scala 123:41:@10470.4]
  assign _T_1592 = {_T_1585,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@10472.4]
  assign _T_1594 = {_T_1586,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@10474.4]
  assign _T_1596 = {_T_1587,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@10476.4]
  assign _T_1598 = {_T_1588,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@10478.4]
  assign _T_1600 = {_T_1589,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@10480.4]
  assign _T_1602 = {_T_1590,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@10482.4]
  assign _T_1603 = _T_1589 ? _T_1600 : _T_1602; // @[Mux.scala 31:69:@10483.4]
  assign _T_1604 = _T_1588 ? _T_1598 : _T_1603; // @[Mux.scala 31:69:@10484.4]
  assign _T_1605 = _T_1587 ? _T_1596 : _T_1604; // @[Mux.scala 31:69:@10485.4]
  assign _T_1606 = _T_1586 ? _T_1594 : _T_1605; // @[Mux.scala 31:69:@10486.4]
  assign _T_1607 = _T_1585 ? _T_1592 : _T_1606; // @[Mux.scala 31:69:@10487.4]
  assign _T_1671 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@10572.4 package.scala 96:25:@10573.4]
  assign _T_1675 = _T_1671 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@10582.4]
  assign _T_1668 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@10564.4 package.scala 96:25:@10565.4]
  assign _T_1676 = _T_1668 ? Mem1D_11_io_output : _T_1675; // @[Mux.scala 31:69:@10583.4]
  assign _T_1665 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@10556.4 package.scala 96:25:@10557.4]
  assign _T_1677 = _T_1665 ? Mem1D_9_io_output : _T_1676; // @[Mux.scala 31:69:@10584.4]
  assign _T_1662 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@10548.4 package.scala 96:25:@10549.4]
  assign _T_1678 = _T_1662 ? Mem1D_7_io_output : _T_1677; // @[Mux.scala 31:69:@10585.4]
  assign _T_1659 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@10540.4 package.scala 96:25:@10541.4]
  assign _T_1679 = _T_1659 ? Mem1D_5_io_output : _T_1678; // @[Mux.scala 31:69:@10586.4]
  assign _T_1656 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@10532.4 package.scala 96:25:@10533.4]
  assign _T_1680 = _T_1656 ? Mem1D_3_io_output : _T_1679; // @[Mux.scala 31:69:@10587.4]
  assign _T_1653 = RetimeWrapper_io_out; // @[package.scala 96:25:@10524.4 package.scala 96:25:@10525.4]
  assign _T_1742 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@10668.4 package.scala 96:25:@10669.4]
  assign _T_1746 = _T_1742 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@10678.4]
  assign _T_1739 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@10660.4 package.scala 96:25:@10661.4]
  assign _T_1747 = _T_1739 ? Mem1D_11_io_output : _T_1746; // @[Mux.scala 31:69:@10679.4]
  assign _T_1736 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@10652.4 package.scala 96:25:@10653.4]
  assign _T_1748 = _T_1736 ? Mem1D_9_io_output : _T_1747; // @[Mux.scala 31:69:@10680.4]
  assign _T_1733 = RetimeWrapper_11_io_out; // @[package.scala 96:25:@10644.4 package.scala 96:25:@10645.4]
  assign _T_1749 = _T_1733 ? Mem1D_7_io_output : _T_1748; // @[Mux.scala 31:69:@10681.4]
  assign _T_1730 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@10636.4 package.scala 96:25:@10637.4]
  assign _T_1750 = _T_1730 ? Mem1D_5_io_output : _T_1749; // @[Mux.scala 31:69:@10682.4]
  assign _T_1727 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@10628.4 package.scala 96:25:@10629.4]
  assign _T_1751 = _T_1727 ? Mem1D_3_io_output : _T_1750; // @[Mux.scala 31:69:@10683.4]
  assign _T_1724 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@10620.4 package.scala 96:25:@10621.4]
  assign _T_1813 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@10764.4 package.scala 96:25:@10765.4]
  assign _T_1817 = _T_1813 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@10774.4]
  assign _T_1810 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@10756.4 package.scala 96:25:@10757.4]
  assign _T_1818 = _T_1810 ? Mem1D_10_io_output : _T_1817; // @[Mux.scala 31:69:@10775.4]
  assign _T_1807 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@10748.4 package.scala 96:25:@10749.4]
  assign _T_1819 = _T_1807 ? Mem1D_8_io_output : _T_1818; // @[Mux.scala 31:69:@10776.4]
  assign _T_1804 = RetimeWrapper_19_io_out; // @[package.scala 96:25:@10740.4 package.scala 96:25:@10741.4]
  assign _T_1820 = _T_1804 ? Mem1D_6_io_output : _T_1819; // @[Mux.scala 31:69:@10777.4]
  assign _T_1801 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@10732.4 package.scala 96:25:@10733.4]
  assign _T_1821 = _T_1801 ? Mem1D_4_io_output : _T_1820; // @[Mux.scala 31:69:@10778.4]
  assign _T_1798 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@10724.4 package.scala 96:25:@10725.4]
  assign _T_1822 = _T_1798 ? Mem1D_2_io_output : _T_1821; // @[Mux.scala 31:69:@10779.4]
  assign _T_1795 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@10716.4 package.scala 96:25:@10717.4]
  assign _T_1884 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@10860.4 package.scala 96:25:@10861.4]
  assign _T_1888 = _T_1884 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@10870.4]
  assign _T_1881 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@10852.4 package.scala 96:25:@10853.4]
  assign _T_1889 = _T_1881 ? Mem1D_10_io_output : _T_1888; // @[Mux.scala 31:69:@10871.4]
  assign _T_1878 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@10844.4 package.scala 96:25:@10845.4]
  assign _T_1890 = _T_1878 ? Mem1D_8_io_output : _T_1889; // @[Mux.scala 31:69:@10872.4]
  assign _T_1875 = RetimeWrapper_27_io_out; // @[package.scala 96:25:@10836.4 package.scala 96:25:@10837.4]
  assign _T_1891 = _T_1875 ? Mem1D_6_io_output : _T_1890; // @[Mux.scala 31:69:@10873.4]
  assign _T_1872 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@10828.4 package.scala 96:25:@10829.4]
  assign _T_1892 = _T_1872 ? Mem1D_4_io_output : _T_1891; // @[Mux.scala 31:69:@10874.4]
  assign _T_1869 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@10820.4 package.scala 96:25:@10821.4]
  assign _T_1893 = _T_1869 ? Mem1D_2_io_output : _T_1892; // @[Mux.scala 31:69:@10875.4]
  assign _T_1866 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@10812.4 package.scala 96:25:@10813.4]
  assign _T_1955 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@10956.4 package.scala 96:25:@10957.4]
  assign _T_1959 = _T_1955 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@10966.4]
  assign _T_1952 = RetimeWrapper_37_io_out; // @[package.scala 96:25:@10948.4 package.scala 96:25:@10949.4]
  assign _T_1960 = _T_1952 ? Mem1D_11_io_output : _T_1959; // @[Mux.scala 31:69:@10967.4]
  assign _T_1949 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@10940.4 package.scala 96:25:@10941.4]
  assign _T_1961 = _T_1949 ? Mem1D_9_io_output : _T_1960; // @[Mux.scala 31:69:@10968.4]
  assign _T_1946 = RetimeWrapper_35_io_out; // @[package.scala 96:25:@10932.4 package.scala 96:25:@10933.4]
  assign _T_1962 = _T_1946 ? Mem1D_7_io_output : _T_1961; // @[Mux.scala 31:69:@10969.4]
  assign _T_1943 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@10924.4 package.scala 96:25:@10925.4]
  assign _T_1963 = _T_1943 ? Mem1D_5_io_output : _T_1962; // @[Mux.scala 31:69:@10970.4]
  assign _T_1940 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@10916.4 package.scala 96:25:@10917.4]
  assign _T_1964 = _T_1940 ? Mem1D_3_io_output : _T_1963; // @[Mux.scala 31:69:@10971.4]
  assign _T_1937 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@10908.4 package.scala 96:25:@10909.4]
  assign _T_2026 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@11052.4 package.scala 96:25:@11053.4]
  assign _T_2030 = _T_2026 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@11062.4]
  assign _T_2023 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@11044.4 package.scala 96:25:@11045.4]
  assign _T_2031 = _T_2023 ? Mem1D_11_io_output : _T_2030; // @[Mux.scala 31:69:@11063.4]
  assign _T_2020 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@11036.4 package.scala 96:25:@11037.4]
  assign _T_2032 = _T_2020 ? Mem1D_9_io_output : _T_2031; // @[Mux.scala 31:69:@11064.4]
  assign _T_2017 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@11028.4 package.scala 96:25:@11029.4]
  assign _T_2033 = _T_2017 ? Mem1D_7_io_output : _T_2032; // @[Mux.scala 31:69:@11065.4]
  assign _T_2014 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@11020.4 package.scala 96:25:@11021.4]
  assign _T_2034 = _T_2014 ? Mem1D_5_io_output : _T_2033; // @[Mux.scala 31:69:@11066.4]
  assign _T_2011 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@11012.4 package.scala 96:25:@11013.4]
  assign _T_2035 = _T_2011 ? Mem1D_3_io_output : _T_2034; // @[Mux.scala 31:69:@11067.4]
  assign _T_2008 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@11004.4 package.scala 96:25:@11005.4]
  assign _T_2097 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@11148.4 package.scala 96:25:@11149.4]
  assign _T_2101 = _T_2097 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@11158.4]
  assign _T_2094 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@11140.4 package.scala 96:25:@11141.4]
  assign _T_2102 = _T_2094 ? Mem1D_10_io_output : _T_2101; // @[Mux.scala 31:69:@11159.4]
  assign _T_2091 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@11132.4 package.scala 96:25:@11133.4]
  assign _T_2103 = _T_2091 ? Mem1D_8_io_output : _T_2102; // @[Mux.scala 31:69:@11160.4]
  assign _T_2088 = RetimeWrapper_51_io_out; // @[package.scala 96:25:@11124.4 package.scala 96:25:@11125.4]
  assign _T_2104 = _T_2088 ? Mem1D_6_io_output : _T_2103; // @[Mux.scala 31:69:@11161.4]
  assign _T_2085 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@11116.4 package.scala 96:25:@11117.4]
  assign _T_2105 = _T_2085 ? Mem1D_4_io_output : _T_2104; // @[Mux.scala 31:69:@11162.4]
  assign _T_2082 = RetimeWrapper_49_io_out; // @[package.scala 96:25:@11108.4 package.scala 96:25:@11109.4]
  assign _T_2106 = _T_2082 ? Mem1D_2_io_output : _T_2105; // @[Mux.scala 31:69:@11163.4]
  assign _T_2079 = RetimeWrapper_48_io_out; // @[package.scala 96:25:@11100.4 package.scala 96:25:@11101.4]
  assign _T_2168 = RetimeWrapper_62_io_out; // @[package.scala 96:25:@11244.4 package.scala 96:25:@11245.4]
  assign _T_2172 = _T_2168 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@11254.4]
  assign _T_2165 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@11236.4 package.scala 96:25:@11237.4]
  assign _T_2173 = _T_2165 ? Mem1D_10_io_output : _T_2172; // @[Mux.scala 31:69:@11255.4]
  assign _T_2162 = RetimeWrapper_60_io_out; // @[package.scala 96:25:@11228.4 package.scala 96:25:@11229.4]
  assign _T_2174 = _T_2162 ? Mem1D_8_io_output : _T_2173; // @[Mux.scala 31:69:@11256.4]
  assign _T_2159 = RetimeWrapper_59_io_out; // @[package.scala 96:25:@11220.4 package.scala 96:25:@11221.4]
  assign _T_2175 = _T_2159 ? Mem1D_6_io_output : _T_2174; // @[Mux.scala 31:69:@11257.4]
  assign _T_2156 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@11212.4 package.scala 96:25:@11213.4]
  assign _T_2176 = _T_2156 ? Mem1D_4_io_output : _T_2175; // @[Mux.scala 31:69:@11258.4]
  assign _T_2153 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@11204.4 package.scala 96:25:@11205.4]
  assign _T_2177 = _T_2153 ? Mem1D_2_io_output : _T_2176; // @[Mux.scala 31:69:@11259.4]
  assign _T_2150 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@11196.4 package.scala 96:25:@11197.4]
  assign _T_2239 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@11340.4 package.scala 96:25:@11341.4]
  assign _T_2243 = _T_2239 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@11350.4]
  assign _T_2236 = RetimeWrapper_69_io_out; // @[package.scala 96:25:@11332.4 package.scala 96:25:@11333.4]
  assign _T_2244 = _T_2236 ? Mem1D_11_io_output : _T_2243; // @[Mux.scala 31:69:@11351.4]
  assign _T_2233 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@11324.4 package.scala 96:25:@11325.4]
  assign _T_2245 = _T_2233 ? Mem1D_9_io_output : _T_2244; // @[Mux.scala 31:69:@11352.4]
  assign _T_2230 = RetimeWrapper_67_io_out; // @[package.scala 96:25:@11316.4 package.scala 96:25:@11317.4]
  assign _T_2246 = _T_2230 ? Mem1D_7_io_output : _T_2245; // @[Mux.scala 31:69:@11353.4]
  assign _T_2227 = RetimeWrapper_66_io_out; // @[package.scala 96:25:@11308.4 package.scala 96:25:@11309.4]
  assign _T_2247 = _T_2227 ? Mem1D_5_io_output : _T_2246; // @[Mux.scala 31:69:@11354.4]
  assign _T_2224 = RetimeWrapper_65_io_out; // @[package.scala 96:25:@11300.4 package.scala 96:25:@11301.4]
  assign _T_2248 = _T_2224 ? Mem1D_3_io_output : _T_2247; // @[Mux.scala 31:69:@11355.4]
  assign _T_2221 = RetimeWrapper_64_io_out; // @[package.scala 96:25:@11292.4 package.scala 96:25:@11293.4]
  assign _T_2310 = RetimeWrapper_78_io_out; // @[package.scala 96:25:@11436.4 package.scala 96:25:@11437.4]
  assign _T_2314 = _T_2310 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@11446.4]
  assign _T_2307 = RetimeWrapper_77_io_out; // @[package.scala 96:25:@11428.4 package.scala 96:25:@11429.4]
  assign _T_2315 = _T_2307 ? Mem1D_10_io_output : _T_2314; // @[Mux.scala 31:69:@11447.4]
  assign _T_2304 = RetimeWrapper_76_io_out; // @[package.scala 96:25:@11420.4 package.scala 96:25:@11421.4]
  assign _T_2316 = _T_2304 ? Mem1D_8_io_output : _T_2315; // @[Mux.scala 31:69:@11448.4]
  assign _T_2301 = RetimeWrapper_75_io_out; // @[package.scala 96:25:@11412.4 package.scala 96:25:@11413.4]
  assign _T_2317 = _T_2301 ? Mem1D_6_io_output : _T_2316; // @[Mux.scala 31:69:@11449.4]
  assign _T_2298 = RetimeWrapper_74_io_out; // @[package.scala 96:25:@11404.4 package.scala 96:25:@11405.4]
  assign _T_2318 = _T_2298 ? Mem1D_4_io_output : _T_2317; // @[Mux.scala 31:69:@11450.4]
  assign _T_2295 = RetimeWrapper_73_io_out; // @[package.scala 96:25:@11396.4 package.scala 96:25:@11397.4]
  assign _T_2319 = _T_2295 ? Mem1D_2_io_output : _T_2318; // @[Mux.scala 31:69:@11451.4]
  assign _T_2292 = RetimeWrapper_72_io_out; // @[package.scala 96:25:@11388.4 package.scala 96:25:@11389.4]
  assign _T_2381 = RetimeWrapper_86_io_out; // @[package.scala 96:25:@11532.4 package.scala 96:25:@11533.4]
  assign _T_2385 = _T_2381 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@11542.4]
  assign _T_2378 = RetimeWrapper_85_io_out; // @[package.scala 96:25:@11524.4 package.scala 96:25:@11525.4]
  assign _T_2386 = _T_2378 ? Mem1D_10_io_output : _T_2385; // @[Mux.scala 31:69:@11543.4]
  assign _T_2375 = RetimeWrapper_84_io_out; // @[package.scala 96:25:@11516.4 package.scala 96:25:@11517.4]
  assign _T_2387 = _T_2375 ? Mem1D_8_io_output : _T_2386; // @[Mux.scala 31:69:@11544.4]
  assign _T_2372 = RetimeWrapper_83_io_out; // @[package.scala 96:25:@11508.4 package.scala 96:25:@11509.4]
  assign _T_2388 = _T_2372 ? Mem1D_6_io_output : _T_2387; // @[Mux.scala 31:69:@11545.4]
  assign _T_2369 = RetimeWrapper_82_io_out; // @[package.scala 96:25:@11500.4 package.scala 96:25:@11501.4]
  assign _T_2389 = _T_2369 ? Mem1D_4_io_output : _T_2388; // @[Mux.scala 31:69:@11546.4]
  assign _T_2366 = RetimeWrapper_81_io_out; // @[package.scala 96:25:@11492.4 package.scala 96:25:@11493.4]
  assign _T_2390 = _T_2366 ? Mem1D_2_io_output : _T_2389; // @[Mux.scala 31:69:@11547.4]
  assign _T_2363 = RetimeWrapper_80_io_out; // @[package.scala 96:25:@11484.4 package.scala 96:25:@11485.4]
  assign _T_2452 = RetimeWrapper_94_io_out; // @[package.scala 96:25:@11628.4 package.scala 96:25:@11629.4]
  assign _T_2456 = _T_2452 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@11638.4]
  assign _T_2449 = RetimeWrapper_93_io_out; // @[package.scala 96:25:@11620.4 package.scala 96:25:@11621.4]
  assign _T_2457 = _T_2449 ? Mem1D_11_io_output : _T_2456; // @[Mux.scala 31:69:@11639.4]
  assign _T_2446 = RetimeWrapper_92_io_out; // @[package.scala 96:25:@11612.4 package.scala 96:25:@11613.4]
  assign _T_2458 = _T_2446 ? Mem1D_9_io_output : _T_2457; // @[Mux.scala 31:69:@11640.4]
  assign _T_2443 = RetimeWrapper_91_io_out; // @[package.scala 96:25:@11604.4 package.scala 96:25:@11605.4]
  assign _T_2459 = _T_2443 ? Mem1D_7_io_output : _T_2458; // @[Mux.scala 31:69:@11641.4]
  assign _T_2440 = RetimeWrapper_90_io_out; // @[package.scala 96:25:@11596.4 package.scala 96:25:@11597.4]
  assign _T_2460 = _T_2440 ? Mem1D_5_io_output : _T_2459; // @[Mux.scala 31:69:@11642.4]
  assign _T_2437 = RetimeWrapper_89_io_out; // @[package.scala 96:25:@11588.4 package.scala 96:25:@11589.4]
  assign _T_2461 = _T_2437 ? Mem1D_3_io_output : _T_2460; // @[Mux.scala 31:69:@11643.4]
  assign _T_2434 = RetimeWrapper_88_io_out; // @[package.scala 96:25:@11580.4 package.scala 96:25:@11581.4]
  assign io_rPort_11_output_0 = _T_2434 ? Mem1D_1_io_output : _T_2461; // @[MemPrimitives.scala 148:13:@11645.4]
  assign io_rPort_10_output_0 = _T_2363 ? Mem1D_io_output : _T_2390; // @[MemPrimitives.scala 148:13:@11549.4]
  assign io_rPort_9_output_0 = _T_2292 ? Mem1D_io_output : _T_2319; // @[MemPrimitives.scala 148:13:@11453.4]
  assign io_rPort_8_output_0 = _T_2221 ? Mem1D_1_io_output : _T_2248; // @[MemPrimitives.scala 148:13:@11357.4]
  assign io_rPort_7_output_0 = _T_2150 ? Mem1D_io_output : _T_2177; // @[MemPrimitives.scala 148:13:@11261.4]
  assign io_rPort_6_output_0 = _T_2079 ? Mem1D_io_output : _T_2106; // @[MemPrimitives.scala 148:13:@11165.4]
  assign io_rPort_5_output_0 = _T_2008 ? Mem1D_1_io_output : _T_2035; // @[MemPrimitives.scala 148:13:@11069.4]
  assign io_rPort_4_output_0 = _T_1937 ? Mem1D_1_io_output : _T_1964; // @[MemPrimitives.scala 148:13:@10973.4]
  assign io_rPort_3_output_0 = _T_1866 ? Mem1D_io_output : _T_1893; // @[MemPrimitives.scala 148:13:@10877.4]
  assign io_rPort_2_output_0 = _T_1795 ? Mem1D_io_output : _T_1822; // @[MemPrimitives.scala 148:13:@10781.4]
  assign io_rPort_1_output_0 = _T_1724 ? Mem1D_1_io_output : _T_1751; // @[MemPrimitives.scala 148:13:@10685.4]
  assign io_rPort_0_output_0 = _T_1653 ? Mem1D_1_io_output : _T_1680; // @[MemPrimitives.scala 148:13:@10589.4]
  assign Mem1D_clock = clock; // @[:@9055.4]
  assign Mem1D_reset = reset; // @[:@9056.4]
  assign Mem1D_io_r_ofs_0 = _T_677[0]; // @[MemPrimitives.scala 127:28:@9561.4]
  assign Mem1D_io_r_backpressure = _T_677[1]; // @[MemPrimitives.scala 128:32:@9562.4]
  assign Mem1D_io_w_ofs_0 = _T_450[0]; // @[MemPrimitives.scala 94:28:@9319.4]
  assign Mem1D_io_w_data_0 = _T_450[8:1]; // @[MemPrimitives.scala 95:29:@9320.4]
  assign Mem1D_io_w_en_0 = _T_450[9]; // @[MemPrimitives.scala 96:27:@9321.4]
  assign Mem1D_1_clock = clock; // @[:@9071.4]
  assign Mem1D_1_reset = reset; // @[:@9072.4]
  assign Mem1D_1_io_r_ofs_0 = _T_739[0]; // @[MemPrimitives.scala 127:28:@9623.4]
  assign Mem1D_1_io_r_backpressure = _T_739[1]; // @[MemPrimitives.scala 128:32:@9624.4]
  assign Mem1D_1_io_w_ofs_0 = _T_461[0]; // @[MemPrimitives.scala 94:28:@9331.4]
  assign Mem1D_1_io_w_data_0 = _T_461[8:1]; // @[MemPrimitives.scala 95:29:@9332.4]
  assign Mem1D_1_io_w_en_0 = _T_461[9]; // @[MemPrimitives.scala 96:27:@9333.4]
  assign Mem1D_2_clock = clock; // @[:@9087.4]
  assign Mem1D_2_reset = reset; // @[:@9088.4]
  assign Mem1D_2_io_r_ofs_0 = _T_801[0]; // @[MemPrimitives.scala 127:28:@9685.4]
  assign Mem1D_2_io_r_backpressure = _T_801[1]; // @[MemPrimitives.scala 128:32:@9686.4]
  assign Mem1D_2_io_w_ofs_0 = _T_472[0]; // @[MemPrimitives.scala 94:28:@9343.4]
  assign Mem1D_2_io_w_data_0 = _T_472[8:1]; // @[MemPrimitives.scala 95:29:@9344.4]
  assign Mem1D_2_io_w_en_0 = _T_472[9]; // @[MemPrimitives.scala 96:27:@9345.4]
  assign Mem1D_3_clock = clock; // @[:@9103.4]
  assign Mem1D_3_reset = reset; // @[:@9104.4]
  assign Mem1D_3_io_r_ofs_0 = _T_863[0]; // @[MemPrimitives.scala 127:28:@9747.4]
  assign Mem1D_3_io_r_backpressure = _T_863[1]; // @[MemPrimitives.scala 128:32:@9748.4]
  assign Mem1D_3_io_w_ofs_0 = _T_483[0]; // @[MemPrimitives.scala 94:28:@9355.4]
  assign Mem1D_3_io_w_data_0 = _T_483[8:1]; // @[MemPrimitives.scala 95:29:@9356.4]
  assign Mem1D_3_io_w_en_0 = _T_483[9]; // @[MemPrimitives.scala 96:27:@9357.4]
  assign Mem1D_4_clock = clock; // @[:@9119.4]
  assign Mem1D_4_reset = reset; // @[:@9120.4]
  assign Mem1D_4_io_r_ofs_0 = _T_925[0]; // @[MemPrimitives.scala 127:28:@9809.4]
  assign Mem1D_4_io_r_backpressure = _T_925[1]; // @[MemPrimitives.scala 128:32:@9810.4]
  assign Mem1D_4_io_w_ofs_0 = _T_494[0]; // @[MemPrimitives.scala 94:28:@9367.4]
  assign Mem1D_4_io_w_data_0 = _T_494[8:1]; // @[MemPrimitives.scala 95:29:@9368.4]
  assign Mem1D_4_io_w_en_0 = _T_494[9]; // @[MemPrimitives.scala 96:27:@9369.4]
  assign Mem1D_5_clock = clock; // @[:@9135.4]
  assign Mem1D_5_reset = reset; // @[:@9136.4]
  assign Mem1D_5_io_r_ofs_0 = _T_987[0]; // @[MemPrimitives.scala 127:28:@9871.4]
  assign Mem1D_5_io_r_backpressure = _T_987[1]; // @[MemPrimitives.scala 128:32:@9872.4]
  assign Mem1D_5_io_w_ofs_0 = _T_505[0]; // @[MemPrimitives.scala 94:28:@9379.4]
  assign Mem1D_5_io_w_data_0 = _T_505[8:1]; // @[MemPrimitives.scala 95:29:@9380.4]
  assign Mem1D_5_io_w_en_0 = _T_505[9]; // @[MemPrimitives.scala 96:27:@9381.4]
  assign Mem1D_6_clock = clock; // @[:@9151.4]
  assign Mem1D_6_reset = reset; // @[:@9152.4]
  assign Mem1D_6_io_r_ofs_0 = _T_1049[0]; // @[MemPrimitives.scala 127:28:@9933.4]
  assign Mem1D_6_io_r_backpressure = _T_1049[1]; // @[MemPrimitives.scala 128:32:@9934.4]
  assign Mem1D_6_io_w_ofs_0 = _T_516[0]; // @[MemPrimitives.scala 94:28:@9391.4]
  assign Mem1D_6_io_w_data_0 = _T_516[8:1]; // @[MemPrimitives.scala 95:29:@9392.4]
  assign Mem1D_6_io_w_en_0 = _T_516[9]; // @[MemPrimitives.scala 96:27:@9393.4]
  assign Mem1D_7_clock = clock; // @[:@9167.4]
  assign Mem1D_7_reset = reset; // @[:@9168.4]
  assign Mem1D_7_io_r_ofs_0 = _T_1111[0]; // @[MemPrimitives.scala 127:28:@9995.4]
  assign Mem1D_7_io_r_backpressure = _T_1111[1]; // @[MemPrimitives.scala 128:32:@9996.4]
  assign Mem1D_7_io_w_ofs_0 = _T_527[0]; // @[MemPrimitives.scala 94:28:@9403.4]
  assign Mem1D_7_io_w_data_0 = _T_527[8:1]; // @[MemPrimitives.scala 95:29:@9404.4]
  assign Mem1D_7_io_w_en_0 = _T_527[9]; // @[MemPrimitives.scala 96:27:@9405.4]
  assign Mem1D_8_clock = clock; // @[:@9183.4]
  assign Mem1D_8_reset = reset; // @[:@9184.4]
  assign Mem1D_8_io_r_ofs_0 = _T_1173[0]; // @[MemPrimitives.scala 127:28:@10057.4]
  assign Mem1D_8_io_r_backpressure = _T_1173[1]; // @[MemPrimitives.scala 128:32:@10058.4]
  assign Mem1D_8_io_w_ofs_0 = _T_538[0]; // @[MemPrimitives.scala 94:28:@9415.4]
  assign Mem1D_8_io_w_data_0 = _T_538[8:1]; // @[MemPrimitives.scala 95:29:@9416.4]
  assign Mem1D_8_io_w_en_0 = _T_538[9]; // @[MemPrimitives.scala 96:27:@9417.4]
  assign Mem1D_9_clock = clock; // @[:@9199.4]
  assign Mem1D_9_reset = reset; // @[:@9200.4]
  assign Mem1D_9_io_r_ofs_0 = _T_1235[0]; // @[MemPrimitives.scala 127:28:@10119.4]
  assign Mem1D_9_io_r_backpressure = _T_1235[1]; // @[MemPrimitives.scala 128:32:@10120.4]
  assign Mem1D_9_io_w_ofs_0 = _T_549[0]; // @[MemPrimitives.scala 94:28:@9427.4]
  assign Mem1D_9_io_w_data_0 = _T_549[8:1]; // @[MemPrimitives.scala 95:29:@9428.4]
  assign Mem1D_9_io_w_en_0 = _T_549[9]; // @[MemPrimitives.scala 96:27:@9429.4]
  assign Mem1D_10_clock = clock; // @[:@9215.4]
  assign Mem1D_10_reset = reset; // @[:@9216.4]
  assign Mem1D_10_io_r_ofs_0 = _T_1297[0]; // @[MemPrimitives.scala 127:28:@10181.4]
  assign Mem1D_10_io_r_backpressure = _T_1297[1]; // @[MemPrimitives.scala 128:32:@10182.4]
  assign Mem1D_10_io_w_ofs_0 = _T_560[0]; // @[MemPrimitives.scala 94:28:@9439.4]
  assign Mem1D_10_io_w_data_0 = _T_560[8:1]; // @[MemPrimitives.scala 95:29:@9440.4]
  assign Mem1D_10_io_w_en_0 = _T_560[9]; // @[MemPrimitives.scala 96:27:@9441.4]
  assign Mem1D_11_clock = clock; // @[:@9231.4]
  assign Mem1D_11_reset = reset; // @[:@9232.4]
  assign Mem1D_11_io_r_ofs_0 = _T_1359[0]; // @[MemPrimitives.scala 127:28:@10243.4]
  assign Mem1D_11_io_r_backpressure = _T_1359[1]; // @[MemPrimitives.scala 128:32:@10244.4]
  assign Mem1D_11_io_w_ofs_0 = _T_571[0]; // @[MemPrimitives.scala 94:28:@9451.4]
  assign Mem1D_11_io_w_data_0 = _T_571[8:1]; // @[MemPrimitives.scala 95:29:@9452.4]
  assign Mem1D_11_io_w_en_0 = _T_571[9]; // @[MemPrimitives.scala 96:27:@9453.4]
  assign Mem1D_12_clock = clock; // @[:@9247.4]
  assign Mem1D_12_reset = reset; // @[:@9248.4]
  assign Mem1D_12_io_r_ofs_0 = _T_1421[0]; // @[MemPrimitives.scala 127:28:@10305.4]
  assign Mem1D_12_io_r_backpressure = _T_1421[1]; // @[MemPrimitives.scala 128:32:@10306.4]
  assign Mem1D_12_io_w_ofs_0 = _T_582[0]; // @[MemPrimitives.scala 94:28:@9463.4]
  assign Mem1D_12_io_w_data_0 = _T_582[8:1]; // @[MemPrimitives.scala 95:29:@9464.4]
  assign Mem1D_12_io_w_en_0 = _T_582[9]; // @[MemPrimitives.scala 96:27:@9465.4]
  assign Mem1D_13_clock = clock; // @[:@9263.4]
  assign Mem1D_13_reset = reset; // @[:@9264.4]
  assign Mem1D_13_io_r_ofs_0 = _T_1483[0]; // @[MemPrimitives.scala 127:28:@10367.4]
  assign Mem1D_13_io_r_backpressure = _T_1483[1]; // @[MemPrimitives.scala 128:32:@10368.4]
  assign Mem1D_13_io_w_ofs_0 = _T_593[0]; // @[MemPrimitives.scala 94:28:@9475.4]
  assign Mem1D_13_io_w_data_0 = _T_593[8:1]; // @[MemPrimitives.scala 95:29:@9476.4]
  assign Mem1D_13_io_w_en_0 = _T_593[9]; // @[MemPrimitives.scala 96:27:@9477.4]
  assign Mem1D_14_clock = clock; // @[:@9279.4]
  assign Mem1D_14_reset = reset; // @[:@9280.4]
  assign Mem1D_14_io_r_ofs_0 = _T_1545[0]; // @[MemPrimitives.scala 127:28:@10429.4]
  assign Mem1D_14_io_r_backpressure = _T_1545[1]; // @[MemPrimitives.scala 128:32:@10430.4]
  assign Mem1D_14_io_w_ofs_0 = _T_604[0]; // @[MemPrimitives.scala 94:28:@9487.4]
  assign Mem1D_14_io_w_data_0 = _T_604[8:1]; // @[MemPrimitives.scala 95:29:@9488.4]
  assign Mem1D_14_io_w_en_0 = _T_604[9]; // @[MemPrimitives.scala 96:27:@9489.4]
  assign Mem1D_15_clock = clock; // @[:@9295.4]
  assign Mem1D_15_reset = reset; // @[:@9296.4]
  assign Mem1D_15_io_r_ofs_0 = _T_1607[0]; // @[MemPrimitives.scala 127:28:@10491.4]
  assign Mem1D_15_io_r_backpressure = _T_1607[1]; // @[MemPrimitives.scala 128:32:@10492.4]
  assign Mem1D_15_io_w_ofs_0 = _T_615[0]; // @[MemPrimitives.scala 94:28:@9499.4]
  assign Mem1D_15_io_w_data_0 = _T_615[8:1]; // @[MemPrimitives.scala 95:29:@9500.4]
  assign Mem1D_15_io_w_en_0 = _T_615[9]; // @[MemPrimitives.scala 96:27:@9501.4]
  assign StickySelects_clock = clock; // @[:@9527.4]
  assign StickySelects_reset = reset; // @[:@9528.4]
  assign StickySelects_io_ins_0 = io_rPort_2_en_0 & _T_623; // @[MemPrimitives.scala 122:60:@9529.4]
  assign StickySelects_io_ins_1 = io_rPort_3_en_0 & _T_629; // @[MemPrimitives.scala 122:60:@9530.4]
  assign StickySelects_io_ins_2 = io_rPort_6_en_0 & _T_635; // @[MemPrimitives.scala 122:60:@9531.4]
  assign StickySelects_io_ins_3 = io_rPort_7_en_0 & _T_641; // @[MemPrimitives.scala 122:60:@9532.4]
  assign StickySelects_io_ins_4 = io_rPort_9_en_0 & _T_647; // @[MemPrimitives.scala 122:60:@9533.4]
  assign StickySelects_io_ins_5 = io_rPort_10_en_0 & _T_653; // @[MemPrimitives.scala 122:60:@9534.4]
  assign StickySelects_1_clock = clock; // @[:@9589.4]
  assign StickySelects_1_reset = reset; // @[:@9590.4]
  assign StickySelects_1_io_ins_0 = io_rPort_0_en_0 & _T_685; // @[MemPrimitives.scala 122:60:@9591.4]
  assign StickySelects_1_io_ins_1 = io_rPort_1_en_0 & _T_691; // @[MemPrimitives.scala 122:60:@9592.4]
  assign StickySelects_1_io_ins_2 = io_rPort_4_en_0 & _T_697; // @[MemPrimitives.scala 122:60:@9593.4]
  assign StickySelects_1_io_ins_3 = io_rPort_5_en_0 & _T_703; // @[MemPrimitives.scala 122:60:@9594.4]
  assign StickySelects_1_io_ins_4 = io_rPort_8_en_0 & _T_709; // @[MemPrimitives.scala 122:60:@9595.4]
  assign StickySelects_1_io_ins_5 = io_rPort_11_en_0 & _T_715; // @[MemPrimitives.scala 122:60:@9596.4]
  assign StickySelects_2_clock = clock; // @[:@9651.4]
  assign StickySelects_2_reset = reset; // @[:@9652.4]
  assign StickySelects_2_io_ins_0 = io_rPort_2_en_0 & _T_747; // @[MemPrimitives.scala 122:60:@9653.4]
  assign StickySelects_2_io_ins_1 = io_rPort_3_en_0 & _T_753; // @[MemPrimitives.scala 122:60:@9654.4]
  assign StickySelects_2_io_ins_2 = io_rPort_6_en_0 & _T_759; // @[MemPrimitives.scala 122:60:@9655.4]
  assign StickySelects_2_io_ins_3 = io_rPort_7_en_0 & _T_765; // @[MemPrimitives.scala 122:60:@9656.4]
  assign StickySelects_2_io_ins_4 = io_rPort_9_en_0 & _T_771; // @[MemPrimitives.scala 122:60:@9657.4]
  assign StickySelects_2_io_ins_5 = io_rPort_10_en_0 & _T_777; // @[MemPrimitives.scala 122:60:@9658.4]
  assign StickySelects_3_clock = clock; // @[:@9713.4]
  assign StickySelects_3_reset = reset; // @[:@9714.4]
  assign StickySelects_3_io_ins_0 = io_rPort_0_en_0 & _T_809; // @[MemPrimitives.scala 122:60:@9715.4]
  assign StickySelects_3_io_ins_1 = io_rPort_1_en_0 & _T_815; // @[MemPrimitives.scala 122:60:@9716.4]
  assign StickySelects_3_io_ins_2 = io_rPort_4_en_0 & _T_821; // @[MemPrimitives.scala 122:60:@9717.4]
  assign StickySelects_3_io_ins_3 = io_rPort_5_en_0 & _T_827; // @[MemPrimitives.scala 122:60:@9718.4]
  assign StickySelects_3_io_ins_4 = io_rPort_8_en_0 & _T_833; // @[MemPrimitives.scala 122:60:@9719.4]
  assign StickySelects_3_io_ins_5 = io_rPort_11_en_0 & _T_839; // @[MemPrimitives.scala 122:60:@9720.4]
  assign StickySelects_4_clock = clock; // @[:@9775.4]
  assign StickySelects_4_reset = reset; // @[:@9776.4]
  assign StickySelects_4_io_ins_0 = io_rPort_2_en_0 & _T_871; // @[MemPrimitives.scala 122:60:@9777.4]
  assign StickySelects_4_io_ins_1 = io_rPort_3_en_0 & _T_877; // @[MemPrimitives.scala 122:60:@9778.4]
  assign StickySelects_4_io_ins_2 = io_rPort_6_en_0 & _T_883; // @[MemPrimitives.scala 122:60:@9779.4]
  assign StickySelects_4_io_ins_3 = io_rPort_7_en_0 & _T_889; // @[MemPrimitives.scala 122:60:@9780.4]
  assign StickySelects_4_io_ins_4 = io_rPort_9_en_0 & _T_895; // @[MemPrimitives.scala 122:60:@9781.4]
  assign StickySelects_4_io_ins_5 = io_rPort_10_en_0 & _T_901; // @[MemPrimitives.scala 122:60:@9782.4]
  assign StickySelects_5_clock = clock; // @[:@9837.4]
  assign StickySelects_5_reset = reset; // @[:@9838.4]
  assign StickySelects_5_io_ins_0 = io_rPort_0_en_0 & _T_933; // @[MemPrimitives.scala 122:60:@9839.4]
  assign StickySelects_5_io_ins_1 = io_rPort_1_en_0 & _T_939; // @[MemPrimitives.scala 122:60:@9840.4]
  assign StickySelects_5_io_ins_2 = io_rPort_4_en_0 & _T_945; // @[MemPrimitives.scala 122:60:@9841.4]
  assign StickySelects_5_io_ins_3 = io_rPort_5_en_0 & _T_951; // @[MemPrimitives.scala 122:60:@9842.4]
  assign StickySelects_5_io_ins_4 = io_rPort_8_en_0 & _T_957; // @[MemPrimitives.scala 122:60:@9843.4]
  assign StickySelects_5_io_ins_5 = io_rPort_11_en_0 & _T_963; // @[MemPrimitives.scala 122:60:@9844.4]
  assign StickySelects_6_clock = clock; // @[:@9899.4]
  assign StickySelects_6_reset = reset; // @[:@9900.4]
  assign StickySelects_6_io_ins_0 = io_rPort_2_en_0 & _T_995; // @[MemPrimitives.scala 122:60:@9901.4]
  assign StickySelects_6_io_ins_1 = io_rPort_3_en_0 & _T_1001; // @[MemPrimitives.scala 122:60:@9902.4]
  assign StickySelects_6_io_ins_2 = io_rPort_6_en_0 & _T_1007; // @[MemPrimitives.scala 122:60:@9903.4]
  assign StickySelects_6_io_ins_3 = io_rPort_7_en_0 & _T_1013; // @[MemPrimitives.scala 122:60:@9904.4]
  assign StickySelects_6_io_ins_4 = io_rPort_9_en_0 & _T_1019; // @[MemPrimitives.scala 122:60:@9905.4]
  assign StickySelects_6_io_ins_5 = io_rPort_10_en_0 & _T_1025; // @[MemPrimitives.scala 122:60:@9906.4]
  assign StickySelects_7_clock = clock; // @[:@9961.4]
  assign StickySelects_7_reset = reset; // @[:@9962.4]
  assign StickySelects_7_io_ins_0 = io_rPort_0_en_0 & _T_1057; // @[MemPrimitives.scala 122:60:@9963.4]
  assign StickySelects_7_io_ins_1 = io_rPort_1_en_0 & _T_1063; // @[MemPrimitives.scala 122:60:@9964.4]
  assign StickySelects_7_io_ins_2 = io_rPort_4_en_0 & _T_1069; // @[MemPrimitives.scala 122:60:@9965.4]
  assign StickySelects_7_io_ins_3 = io_rPort_5_en_0 & _T_1075; // @[MemPrimitives.scala 122:60:@9966.4]
  assign StickySelects_7_io_ins_4 = io_rPort_8_en_0 & _T_1081; // @[MemPrimitives.scala 122:60:@9967.4]
  assign StickySelects_7_io_ins_5 = io_rPort_11_en_0 & _T_1087; // @[MemPrimitives.scala 122:60:@9968.4]
  assign StickySelects_8_clock = clock; // @[:@10023.4]
  assign StickySelects_8_reset = reset; // @[:@10024.4]
  assign StickySelects_8_io_ins_0 = io_rPort_2_en_0 & _T_1119; // @[MemPrimitives.scala 122:60:@10025.4]
  assign StickySelects_8_io_ins_1 = io_rPort_3_en_0 & _T_1125; // @[MemPrimitives.scala 122:60:@10026.4]
  assign StickySelects_8_io_ins_2 = io_rPort_6_en_0 & _T_1131; // @[MemPrimitives.scala 122:60:@10027.4]
  assign StickySelects_8_io_ins_3 = io_rPort_7_en_0 & _T_1137; // @[MemPrimitives.scala 122:60:@10028.4]
  assign StickySelects_8_io_ins_4 = io_rPort_9_en_0 & _T_1143; // @[MemPrimitives.scala 122:60:@10029.4]
  assign StickySelects_8_io_ins_5 = io_rPort_10_en_0 & _T_1149; // @[MemPrimitives.scala 122:60:@10030.4]
  assign StickySelects_9_clock = clock; // @[:@10085.4]
  assign StickySelects_9_reset = reset; // @[:@10086.4]
  assign StickySelects_9_io_ins_0 = io_rPort_0_en_0 & _T_1181; // @[MemPrimitives.scala 122:60:@10087.4]
  assign StickySelects_9_io_ins_1 = io_rPort_1_en_0 & _T_1187; // @[MemPrimitives.scala 122:60:@10088.4]
  assign StickySelects_9_io_ins_2 = io_rPort_4_en_0 & _T_1193; // @[MemPrimitives.scala 122:60:@10089.4]
  assign StickySelects_9_io_ins_3 = io_rPort_5_en_0 & _T_1199; // @[MemPrimitives.scala 122:60:@10090.4]
  assign StickySelects_9_io_ins_4 = io_rPort_8_en_0 & _T_1205; // @[MemPrimitives.scala 122:60:@10091.4]
  assign StickySelects_9_io_ins_5 = io_rPort_11_en_0 & _T_1211; // @[MemPrimitives.scala 122:60:@10092.4]
  assign StickySelects_10_clock = clock; // @[:@10147.4]
  assign StickySelects_10_reset = reset; // @[:@10148.4]
  assign StickySelects_10_io_ins_0 = io_rPort_2_en_0 & _T_1243; // @[MemPrimitives.scala 122:60:@10149.4]
  assign StickySelects_10_io_ins_1 = io_rPort_3_en_0 & _T_1249; // @[MemPrimitives.scala 122:60:@10150.4]
  assign StickySelects_10_io_ins_2 = io_rPort_6_en_0 & _T_1255; // @[MemPrimitives.scala 122:60:@10151.4]
  assign StickySelects_10_io_ins_3 = io_rPort_7_en_0 & _T_1261; // @[MemPrimitives.scala 122:60:@10152.4]
  assign StickySelects_10_io_ins_4 = io_rPort_9_en_0 & _T_1267; // @[MemPrimitives.scala 122:60:@10153.4]
  assign StickySelects_10_io_ins_5 = io_rPort_10_en_0 & _T_1273; // @[MemPrimitives.scala 122:60:@10154.4]
  assign StickySelects_11_clock = clock; // @[:@10209.4]
  assign StickySelects_11_reset = reset; // @[:@10210.4]
  assign StickySelects_11_io_ins_0 = io_rPort_0_en_0 & _T_1305; // @[MemPrimitives.scala 122:60:@10211.4]
  assign StickySelects_11_io_ins_1 = io_rPort_1_en_0 & _T_1311; // @[MemPrimitives.scala 122:60:@10212.4]
  assign StickySelects_11_io_ins_2 = io_rPort_4_en_0 & _T_1317; // @[MemPrimitives.scala 122:60:@10213.4]
  assign StickySelects_11_io_ins_3 = io_rPort_5_en_0 & _T_1323; // @[MemPrimitives.scala 122:60:@10214.4]
  assign StickySelects_11_io_ins_4 = io_rPort_8_en_0 & _T_1329; // @[MemPrimitives.scala 122:60:@10215.4]
  assign StickySelects_11_io_ins_5 = io_rPort_11_en_0 & _T_1335; // @[MemPrimitives.scala 122:60:@10216.4]
  assign StickySelects_12_clock = clock; // @[:@10271.4]
  assign StickySelects_12_reset = reset; // @[:@10272.4]
  assign StickySelects_12_io_ins_0 = io_rPort_2_en_0 & _T_1367; // @[MemPrimitives.scala 122:60:@10273.4]
  assign StickySelects_12_io_ins_1 = io_rPort_3_en_0 & _T_1373; // @[MemPrimitives.scala 122:60:@10274.4]
  assign StickySelects_12_io_ins_2 = io_rPort_6_en_0 & _T_1379; // @[MemPrimitives.scala 122:60:@10275.4]
  assign StickySelects_12_io_ins_3 = io_rPort_7_en_0 & _T_1385; // @[MemPrimitives.scala 122:60:@10276.4]
  assign StickySelects_12_io_ins_4 = io_rPort_9_en_0 & _T_1391; // @[MemPrimitives.scala 122:60:@10277.4]
  assign StickySelects_12_io_ins_5 = io_rPort_10_en_0 & _T_1397; // @[MemPrimitives.scala 122:60:@10278.4]
  assign StickySelects_13_clock = clock; // @[:@10333.4]
  assign StickySelects_13_reset = reset; // @[:@10334.4]
  assign StickySelects_13_io_ins_0 = io_rPort_0_en_0 & _T_1429; // @[MemPrimitives.scala 122:60:@10335.4]
  assign StickySelects_13_io_ins_1 = io_rPort_1_en_0 & _T_1435; // @[MemPrimitives.scala 122:60:@10336.4]
  assign StickySelects_13_io_ins_2 = io_rPort_4_en_0 & _T_1441; // @[MemPrimitives.scala 122:60:@10337.4]
  assign StickySelects_13_io_ins_3 = io_rPort_5_en_0 & _T_1447; // @[MemPrimitives.scala 122:60:@10338.4]
  assign StickySelects_13_io_ins_4 = io_rPort_8_en_0 & _T_1453; // @[MemPrimitives.scala 122:60:@10339.4]
  assign StickySelects_13_io_ins_5 = io_rPort_11_en_0 & _T_1459; // @[MemPrimitives.scala 122:60:@10340.4]
  assign StickySelects_14_clock = clock; // @[:@10395.4]
  assign StickySelects_14_reset = reset; // @[:@10396.4]
  assign StickySelects_14_io_ins_0 = io_rPort_2_en_0 & _T_1491; // @[MemPrimitives.scala 122:60:@10397.4]
  assign StickySelects_14_io_ins_1 = io_rPort_3_en_0 & _T_1497; // @[MemPrimitives.scala 122:60:@10398.4]
  assign StickySelects_14_io_ins_2 = io_rPort_6_en_0 & _T_1503; // @[MemPrimitives.scala 122:60:@10399.4]
  assign StickySelects_14_io_ins_3 = io_rPort_7_en_0 & _T_1509; // @[MemPrimitives.scala 122:60:@10400.4]
  assign StickySelects_14_io_ins_4 = io_rPort_9_en_0 & _T_1515; // @[MemPrimitives.scala 122:60:@10401.4]
  assign StickySelects_14_io_ins_5 = io_rPort_10_en_0 & _T_1521; // @[MemPrimitives.scala 122:60:@10402.4]
  assign StickySelects_15_clock = clock; // @[:@10457.4]
  assign StickySelects_15_reset = reset; // @[:@10458.4]
  assign StickySelects_15_io_ins_0 = io_rPort_0_en_0 & _T_1553; // @[MemPrimitives.scala 122:60:@10459.4]
  assign StickySelects_15_io_ins_1 = io_rPort_1_en_0 & _T_1559; // @[MemPrimitives.scala 122:60:@10460.4]
  assign StickySelects_15_io_ins_2 = io_rPort_4_en_0 & _T_1565; // @[MemPrimitives.scala 122:60:@10461.4]
  assign StickySelects_15_io_ins_3 = io_rPort_5_en_0 & _T_1571; // @[MemPrimitives.scala 122:60:@10462.4]
  assign StickySelects_15_io_ins_4 = io_rPort_8_en_0 & _T_1577; // @[MemPrimitives.scala 122:60:@10463.4]
  assign StickySelects_15_io_ins_5 = io_rPort_11_en_0 & _T_1583; // @[MemPrimitives.scala 122:60:@10464.4]
  assign RetimeWrapper_clock = clock; // @[:@10520.4]
  assign RetimeWrapper_reset = reset; // @[:@10521.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@10523.4]
  assign RetimeWrapper_io_in = _T_685 & io_rPort_0_en_0; // @[package.scala 94:16:@10522.4]
  assign RetimeWrapper_1_clock = clock; // @[:@10528.4]
  assign RetimeWrapper_1_reset = reset; // @[:@10529.4]
  assign RetimeWrapper_1_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@10531.4]
  assign RetimeWrapper_1_io_in = _T_809 & io_rPort_0_en_0; // @[package.scala 94:16:@10530.4]
  assign RetimeWrapper_2_clock = clock; // @[:@10536.4]
  assign RetimeWrapper_2_reset = reset; // @[:@10537.4]
  assign RetimeWrapper_2_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@10539.4]
  assign RetimeWrapper_2_io_in = _T_933 & io_rPort_0_en_0; // @[package.scala 94:16:@10538.4]
  assign RetimeWrapper_3_clock = clock; // @[:@10544.4]
  assign RetimeWrapper_3_reset = reset; // @[:@10545.4]
  assign RetimeWrapper_3_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@10547.4]
  assign RetimeWrapper_3_io_in = _T_1057 & io_rPort_0_en_0; // @[package.scala 94:16:@10546.4]
  assign RetimeWrapper_4_clock = clock; // @[:@10552.4]
  assign RetimeWrapper_4_reset = reset; // @[:@10553.4]
  assign RetimeWrapper_4_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@10555.4]
  assign RetimeWrapper_4_io_in = _T_1181 & io_rPort_0_en_0; // @[package.scala 94:16:@10554.4]
  assign RetimeWrapper_5_clock = clock; // @[:@10560.4]
  assign RetimeWrapper_5_reset = reset; // @[:@10561.4]
  assign RetimeWrapper_5_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@10563.4]
  assign RetimeWrapper_5_io_in = _T_1305 & io_rPort_0_en_0; // @[package.scala 94:16:@10562.4]
  assign RetimeWrapper_6_clock = clock; // @[:@10568.4]
  assign RetimeWrapper_6_reset = reset; // @[:@10569.4]
  assign RetimeWrapper_6_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@10571.4]
  assign RetimeWrapper_6_io_in = _T_1429 & io_rPort_0_en_0; // @[package.scala 94:16:@10570.4]
  assign RetimeWrapper_7_clock = clock; // @[:@10576.4]
  assign RetimeWrapper_7_reset = reset; // @[:@10577.4]
  assign RetimeWrapper_7_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@10579.4]
  assign RetimeWrapper_7_io_in = _T_1553 & io_rPort_0_en_0; // @[package.scala 94:16:@10578.4]
  assign RetimeWrapper_8_clock = clock; // @[:@10616.4]
  assign RetimeWrapper_8_reset = reset; // @[:@10617.4]
  assign RetimeWrapper_8_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@10619.4]
  assign RetimeWrapper_8_io_in = _T_691 & io_rPort_1_en_0; // @[package.scala 94:16:@10618.4]
  assign RetimeWrapper_9_clock = clock; // @[:@10624.4]
  assign RetimeWrapper_9_reset = reset; // @[:@10625.4]
  assign RetimeWrapper_9_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@10627.4]
  assign RetimeWrapper_9_io_in = _T_815 & io_rPort_1_en_0; // @[package.scala 94:16:@10626.4]
  assign RetimeWrapper_10_clock = clock; // @[:@10632.4]
  assign RetimeWrapper_10_reset = reset; // @[:@10633.4]
  assign RetimeWrapper_10_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@10635.4]
  assign RetimeWrapper_10_io_in = _T_939 & io_rPort_1_en_0; // @[package.scala 94:16:@10634.4]
  assign RetimeWrapper_11_clock = clock; // @[:@10640.4]
  assign RetimeWrapper_11_reset = reset; // @[:@10641.4]
  assign RetimeWrapper_11_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@10643.4]
  assign RetimeWrapper_11_io_in = _T_1063 & io_rPort_1_en_0; // @[package.scala 94:16:@10642.4]
  assign RetimeWrapper_12_clock = clock; // @[:@10648.4]
  assign RetimeWrapper_12_reset = reset; // @[:@10649.4]
  assign RetimeWrapper_12_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@10651.4]
  assign RetimeWrapper_12_io_in = _T_1187 & io_rPort_1_en_0; // @[package.scala 94:16:@10650.4]
  assign RetimeWrapper_13_clock = clock; // @[:@10656.4]
  assign RetimeWrapper_13_reset = reset; // @[:@10657.4]
  assign RetimeWrapper_13_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@10659.4]
  assign RetimeWrapper_13_io_in = _T_1311 & io_rPort_1_en_0; // @[package.scala 94:16:@10658.4]
  assign RetimeWrapper_14_clock = clock; // @[:@10664.4]
  assign RetimeWrapper_14_reset = reset; // @[:@10665.4]
  assign RetimeWrapper_14_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@10667.4]
  assign RetimeWrapper_14_io_in = _T_1435 & io_rPort_1_en_0; // @[package.scala 94:16:@10666.4]
  assign RetimeWrapper_15_clock = clock; // @[:@10672.4]
  assign RetimeWrapper_15_reset = reset; // @[:@10673.4]
  assign RetimeWrapper_15_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@10675.4]
  assign RetimeWrapper_15_io_in = _T_1559 & io_rPort_1_en_0; // @[package.scala 94:16:@10674.4]
  assign RetimeWrapper_16_clock = clock; // @[:@10712.4]
  assign RetimeWrapper_16_reset = reset; // @[:@10713.4]
  assign RetimeWrapper_16_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@10715.4]
  assign RetimeWrapper_16_io_in = _T_623 & io_rPort_2_en_0; // @[package.scala 94:16:@10714.4]
  assign RetimeWrapper_17_clock = clock; // @[:@10720.4]
  assign RetimeWrapper_17_reset = reset; // @[:@10721.4]
  assign RetimeWrapper_17_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@10723.4]
  assign RetimeWrapper_17_io_in = _T_747 & io_rPort_2_en_0; // @[package.scala 94:16:@10722.4]
  assign RetimeWrapper_18_clock = clock; // @[:@10728.4]
  assign RetimeWrapper_18_reset = reset; // @[:@10729.4]
  assign RetimeWrapper_18_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@10731.4]
  assign RetimeWrapper_18_io_in = _T_871 & io_rPort_2_en_0; // @[package.scala 94:16:@10730.4]
  assign RetimeWrapper_19_clock = clock; // @[:@10736.4]
  assign RetimeWrapper_19_reset = reset; // @[:@10737.4]
  assign RetimeWrapper_19_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@10739.4]
  assign RetimeWrapper_19_io_in = _T_995 & io_rPort_2_en_0; // @[package.scala 94:16:@10738.4]
  assign RetimeWrapper_20_clock = clock; // @[:@10744.4]
  assign RetimeWrapper_20_reset = reset; // @[:@10745.4]
  assign RetimeWrapper_20_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@10747.4]
  assign RetimeWrapper_20_io_in = _T_1119 & io_rPort_2_en_0; // @[package.scala 94:16:@10746.4]
  assign RetimeWrapper_21_clock = clock; // @[:@10752.4]
  assign RetimeWrapper_21_reset = reset; // @[:@10753.4]
  assign RetimeWrapper_21_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@10755.4]
  assign RetimeWrapper_21_io_in = _T_1243 & io_rPort_2_en_0; // @[package.scala 94:16:@10754.4]
  assign RetimeWrapper_22_clock = clock; // @[:@10760.4]
  assign RetimeWrapper_22_reset = reset; // @[:@10761.4]
  assign RetimeWrapper_22_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@10763.4]
  assign RetimeWrapper_22_io_in = _T_1367 & io_rPort_2_en_0; // @[package.scala 94:16:@10762.4]
  assign RetimeWrapper_23_clock = clock; // @[:@10768.4]
  assign RetimeWrapper_23_reset = reset; // @[:@10769.4]
  assign RetimeWrapper_23_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@10771.4]
  assign RetimeWrapper_23_io_in = _T_1491 & io_rPort_2_en_0; // @[package.scala 94:16:@10770.4]
  assign RetimeWrapper_24_clock = clock; // @[:@10808.4]
  assign RetimeWrapper_24_reset = reset; // @[:@10809.4]
  assign RetimeWrapper_24_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@10811.4]
  assign RetimeWrapper_24_io_in = _T_629 & io_rPort_3_en_0; // @[package.scala 94:16:@10810.4]
  assign RetimeWrapper_25_clock = clock; // @[:@10816.4]
  assign RetimeWrapper_25_reset = reset; // @[:@10817.4]
  assign RetimeWrapper_25_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@10819.4]
  assign RetimeWrapper_25_io_in = _T_753 & io_rPort_3_en_0; // @[package.scala 94:16:@10818.4]
  assign RetimeWrapper_26_clock = clock; // @[:@10824.4]
  assign RetimeWrapper_26_reset = reset; // @[:@10825.4]
  assign RetimeWrapper_26_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@10827.4]
  assign RetimeWrapper_26_io_in = _T_877 & io_rPort_3_en_0; // @[package.scala 94:16:@10826.4]
  assign RetimeWrapper_27_clock = clock; // @[:@10832.4]
  assign RetimeWrapper_27_reset = reset; // @[:@10833.4]
  assign RetimeWrapper_27_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@10835.4]
  assign RetimeWrapper_27_io_in = _T_1001 & io_rPort_3_en_0; // @[package.scala 94:16:@10834.4]
  assign RetimeWrapper_28_clock = clock; // @[:@10840.4]
  assign RetimeWrapper_28_reset = reset; // @[:@10841.4]
  assign RetimeWrapper_28_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@10843.4]
  assign RetimeWrapper_28_io_in = _T_1125 & io_rPort_3_en_0; // @[package.scala 94:16:@10842.4]
  assign RetimeWrapper_29_clock = clock; // @[:@10848.4]
  assign RetimeWrapper_29_reset = reset; // @[:@10849.4]
  assign RetimeWrapper_29_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@10851.4]
  assign RetimeWrapper_29_io_in = _T_1249 & io_rPort_3_en_0; // @[package.scala 94:16:@10850.4]
  assign RetimeWrapper_30_clock = clock; // @[:@10856.4]
  assign RetimeWrapper_30_reset = reset; // @[:@10857.4]
  assign RetimeWrapper_30_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@10859.4]
  assign RetimeWrapper_30_io_in = _T_1373 & io_rPort_3_en_0; // @[package.scala 94:16:@10858.4]
  assign RetimeWrapper_31_clock = clock; // @[:@10864.4]
  assign RetimeWrapper_31_reset = reset; // @[:@10865.4]
  assign RetimeWrapper_31_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@10867.4]
  assign RetimeWrapper_31_io_in = _T_1497 & io_rPort_3_en_0; // @[package.scala 94:16:@10866.4]
  assign RetimeWrapper_32_clock = clock; // @[:@10904.4]
  assign RetimeWrapper_32_reset = reset; // @[:@10905.4]
  assign RetimeWrapper_32_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@10907.4]
  assign RetimeWrapper_32_io_in = _T_697 & io_rPort_4_en_0; // @[package.scala 94:16:@10906.4]
  assign RetimeWrapper_33_clock = clock; // @[:@10912.4]
  assign RetimeWrapper_33_reset = reset; // @[:@10913.4]
  assign RetimeWrapper_33_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@10915.4]
  assign RetimeWrapper_33_io_in = _T_821 & io_rPort_4_en_0; // @[package.scala 94:16:@10914.4]
  assign RetimeWrapper_34_clock = clock; // @[:@10920.4]
  assign RetimeWrapper_34_reset = reset; // @[:@10921.4]
  assign RetimeWrapper_34_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@10923.4]
  assign RetimeWrapper_34_io_in = _T_945 & io_rPort_4_en_0; // @[package.scala 94:16:@10922.4]
  assign RetimeWrapper_35_clock = clock; // @[:@10928.4]
  assign RetimeWrapper_35_reset = reset; // @[:@10929.4]
  assign RetimeWrapper_35_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@10931.4]
  assign RetimeWrapper_35_io_in = _T_1069 & io_rPort_4_en_0; // @[package.scala 94:16:@10930.4]
  assign RetimeWrapper_36_clock = clock; // @[:@10936.4]
  assign RetimeWrapper_36_reset = reset; // @[:@10937.4]
  assign RetimeWrapper_36_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@10939.4]
  assign RetimeWrapper_36_io_in = _T_1193 & io_rPort_4_en_0; // @[package.scala 94:16:@10938.4]
  assign RetimeWrapper_37_clock = clock; // @[:@10944.4]
  assign RetimeWrapper_37_reset = reset; // @[:@10945.4]
  assign RetimeWrapper_37_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@10947.4]
  assign RetimeWrapper_37_io_in = _T_1317 & io_rPort_4_en_0; // @[package.scala 94:16:@10946.4]
  assign RetimeWrapper_38_clock = clock; // @[:@10952.4]
  assign RetimeWrapper_38_reset = reset; // @[:@10953.4]
  assign RetimeWrapper_38_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@10955.4]
  assign RetimeWrapper_38_io_in = _T_1441 & io_rPort_4_en_0; // @[package.scala 94:16:@10954.4]
  assign RetimeWrapper_39_clock = clock; // @[:@10960.4]
  assign RetimeWrapper_39_reset = reset; // @[:@10961.4]
  assign RetimeWrapper_39_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@10963.4]
  assign RetimeWrapper_39_io_in = _T_1565 & io_rPort_4_en_0; // @[package.scala 94:16:@10962.4]
  assign RetimeWrapper_40_clock = clock; // @[:@11000.4]
  assign RetimeWrapper_40_reset = reset; // @[:@11001.4]
  assign RetimeWrapper_40_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@11003.4]
  assign RetimeWrapper_40_io_in = _T_703 & io_rPort_5_en_0; // @[package.scala 94:16:@11002.4]
  assign RetimeWrapper_41_clock = clock; // @[:@11008.4]
  assign RetimeWrapper_41_reset = reset; // @[:@11009.4]
  assign RetimeWrapper_41_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@11011.4]
  assign RetimeWrapper_41_io_in = _T_827 & io_rPort_5_en_0; // @[package.scala 94:16:@11010.4]
  assign RetimeWrapper_42_clock = clock; // @[:@11016.4]
  assign RetimeWrapper_42_reset = reset; // @[:@11017.4]
  assign RetimeWrapper_42_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@11019.4]
  assign RetimeWrapper_42_io_in = _T_951 & io_rPort_5_en_0; // @[package.scala 94:16:@11018.4]
  assign RetimeWrapper_43_clock = clock; // @[:@11024.4]
  assign RetimeWrapper_43_reset = reset; // @[:@11025.4]
  assign RetimeWrapper_43_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@11027.4]
  assign RetimeWrapper_43_io_in = _T_1075 & io_rPort_5_en_0; // @[package.scala 94:16:@11026.4]
  assign RetimeWrapper_44_clock = clock; // @[:@11032.4]
  assign RetimeWrapper_44_reset = reset; // @[:@11033.4]
  assign RetimeWrapper_44_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@11035.4]
  assign RetimeWrapper_44_io_in = _T_1199 & io_rPort_5_en_0; // @[package.scala 94:16:@11034.4]
  assign RetimeWrapper_45_clock = clock; // @[:@11040.4]
  assign RetimeWrapper_45_reset = reset; // @[:@11041.4]
  assign RetimeWrapper_45_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@11043.4]
  assign RetimeWrapper_45_io_in = _T_1323 & io_rPort_5_en_0; // @[package.scala 94:16:@11042.4]
  assign RetimeWrapper_46_clock = clock; // @[:@11048.4]
  assign RetimeWrapper_46_reset = reset; // @[:@11049.4]
  assign RetimeWrapper_46_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@11051.4]
  assign RetimeWrapper_46_io_in = _T_1447 & io_rPort_5_en_0; // @[package.scala 94:16:@11050.4]
  assign RetimeWrapper_47_clock = clock; // @[:@11056.4]
  assign RetimeWrapper_47_reset = reset; // @[:@11057.4]
  assign RetimeWrapper_47_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@11059.4]
  assign RetimeWrapper_47_io_in = _T_1571 & io_rPort_5_en_0; // @[package.scala 94:16:@11058.4]
  assign RetimeWrapper_48_clock = clock; // @[:@11096.4]
  assign RetimeWrapper_48_reset = reset; // @[:@11097.4]
  assign RetimeWrapper_48_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@11099.4]
  assign RetimeWrapper_48_io_in = _T_635 & io_rPort_6_en_0; // @[package.scala 94:16:@11098.4]
  assign RetimeWrapper_49_clock = clock; // @[:@11104.4]
  assign RetimeWrapper_49_reset = reset; // @[:@11105.4]
  assign RetimeWrapper_49_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@11107.4]
  assign RetimeWrapper_49_io_in = _T_759 & io_rPort_6_en_0; // @[package.scala 94:16:@11106.4]
  assign RetimeWrapper_50_clock = clock; // @[:@11112.4]
  assign RetimeWrapper_50_reset = reset; // @[:@11113.4]
  assign RetimeWrapper_50_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@11115.4]
  assign RetimeWrapper_50_io_in = _T_883 & io_rPort_6_en_0; // @[package.scala 94:16:@11114.4]
  assign RetimeWrapper_51_clock = clock; // @[:@11120.4]
  assign RetimeWrapper_51_reset = reset; // @[:@11121.4]
  assign RetimeWrapper_51_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@11123.4]
  assign RetimeWrapper_51_io_in = _T_1007 & io_rPort_6_en_0; // @[package.scala 94:16:@11122.4]
  assign RetimeWrapper_52_clock = clock; // @[:@11128.4]
  assign RetimeWrapper_52_reset = reset; // @[:@11129.4]
  assign RetimeWrapper_52_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@11131.4]
  assign RetimeWrapper_52_io_in = _T_1131 & io_rPort_6_en_0; // @[package.scala 94:16:@11130.4]
  assign RetimeWrapper_53_clock = clock; // @[:@11136.4]
  assign RetimeWrapper_53_reset = reset; // @[:@11137.4]
  assign RetimeWrapper_53_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@11139.4]
  assign RetimeWrapper_53_io_in = _T_1255 & io_rPort_6_en_0; // @[package.scala 94:16:@11138.4]
  assign RetimeWrapper_54_clock = clock; // @[:@11144.4]
  assign RetimeWrapper_54_reset = reset; // @[:@11145.4]
  assign RetimeWrapper_54_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@11147.4]
  assign RetimeWrapper_54_io_in = _T_1379 & io_rPort_6_en_0; // @[package.scala 94:16:@11146.4]
  assign RetimeWrapper_55_clock = clock; // @[:@11152.4]
  assign RetimeWrapper_55_reset = reset; // @[:@11153.4]
  assign RetimeWrapper_55_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@11155.4]
  assign RetimeWrapper_55_io_in = _T_1503 & io_rPort_6_en_0; // @[package.scala 94:16:@11154.4]
  assign RetimeWrapper_56_clock = clock; // @[:@11192.4]
  assign RetimeWrapper_56_reset = reset; // @[:@11193.4]
  assign RetimeWrapper_56_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@11195.4]
  assign RetimeWrapper_56_io_in = _T_641 & io_rPort_7_en_0; // @[package.scala 94:16:@11194.4]
  assign RetimeWrapper_57_clock = clock; // @[:@11200.4]
  assign RetimeWrapper_57_reset = reset; // @[:@11201.4]
  assign RetimeWrapper_57_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@11203.4]
  assign RetimeWrapper_57_io_in = _T_765 & io_rPort_7_en_0; // @[package.scala 94:16:@11202.4]
  assign RetimeWrapper_58_clock = clock; // @[:@11208.4]
  assign RetimeWrapper_58_reset = reset; // @[:@11209.4]
  assign RetimeWrapper_58_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@11211.4]
  assign RetimeWrapper_58_io_in = _T_889 & io_rPort_7_en_0; // @[package.scala 94:16:@11210.4]
  assign RetimeWrapper_59_clock = clock; // @[:@11216.4]
  assign RetimeWrapper_59_reset = reset; // @[:@11217.4]
  assign RetimeWrapper_59_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@11219.4]
  assign RetimeWrapper_59_io_in = _T_1013 & io_rPort_7_en_0; // @[package.scala 94:16:@11218.4]
  assign RetimeWrapper_60_clock = clock; // @[:@11224.4]
  assign RetimeWrapper_60_reset = reset; // @[:@11225.4]
  assign RetimeWrapper_60_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@11227.4]
  assign RetimeWrapper_60_io_in = _T_1137 & io_rPort_7_en_0; // @[package.scala 94:16:@11226.4]
  assign RetimeWrapper_61_clock = clock; // @[:@11232.4]
  assign RetimeWrapper_61_reset = reset; // @[:@11233.4]
  assign RetimeWrapper_61_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@11235.4]
  assign RetimeWrapper_61_io_in = _T_1261 & io_rPort_7_en_0; // @[package.scala 94:16:@11234.4]
  assign RetimeWrapper_62_clock = clock; // @[:@11240.4]
  assign RetimeWrapper_62_reset = reset; // @[:@11241.4]
  assign RetimeWrapper_62_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@11243.4]
  assign RetimeWrapper_62_io_in = _T_1385 & io_rPort_7_en_0; // @[package.scala 94:16:@11242.4]
  assign RetimeWrapper_63_clock = clock; // @[:@11248.4]
  assign RetimeWrapper_63_reset = reset; // @[:@11249.4]
  assign RetimeWrapper_63_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@11251.4]
  assign RetimeWrapper_63_io_in = _T_1509 & io_rPort_7_en_0; // @[package.scala 94:16:@11250.4]
  assign RetimeWrapper_64_clock = clock; // @[:@11288.4]
  assign RetimeWrapper_64_reset = reset; // @[:@11289.4]
  assign RetimeWrapper_64_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@11291.4]
  assign RetimeWrapper_64_io_in = _T_709 & io_rPort_8_en_0; // @[package.scala 94:16:@11290.4]
  assign RetimeWrapper_65_clock = clock; // @[:@11296.4]
  assign RetimeWrapper_65_reset = reset; // @[:@11297.4]
  assign RetimeWrapper_65_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@11299.4]
  assign RetimeWrapper_65_io_in = _T_833 & io_rPort_8_en_0; // @[package.scala 94:16:@11298.4]
  assign RetimeWrapper_66_clock = clock; // @[:@11304.4]
  assign RetimeWrapper_66_reset = reset; // @[:@11305.4]
  assign RetimeWrapper_66_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@11307.4]
  assign RetimeWrapper_66_io_in = _T_957 & io_rPort_8_en_0; // @[package.scala 94:16:@11306.4]
  assign RetimeWrapper_67_clock = clock; // @[:@11312.4]
  assign RetimeWrapper_67_reset = reset; // @[:@11313.4]
  assign RetimeWrapper_67_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@11315.4]
  assign RetimeWrapper_67_io_in = _T_1081 & io_rPort_8_en_0; // @[package.scala 94:16:@11314.4]
  assign RetimeWrapper_68_clock = clock; // @[:@11320.4]
  assign RetimeWrapper_68_reset = reset; // @[:@11321.4]
  assign RetimeWrapper_68_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@11323.4]
  assign RetimeWrapper_68_io_in = _T_1205 & io_rPort_8_en_0; // @[package.scala 94:16:@11322.4]
  assign RetimeWrapper_69_clock = clock; // @[:@11328.4]
  assign RetimeWrapper_69_reset = reset; // @[:@11329.4]
  assign RetimeWrapper_69_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@11331.4]
  assign RetimeWrapper_69_io_in = _T_1329 & io_rPort_8_en_0; // @[package.scala 94:16:@11330.4]
  assign RetimeWrapper_70_clock = clock; // @[:@11336.4]
  assign RetimeWrapper_70_reset = reset; // @[:@11337.4]
  assign RetimeWrapper_70_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@11339.4]
  assign RetimeWrapper_70_io_in = _T_1453 & io_rPort_8_en_0; // @[package.scala 94:16:@11338.4]
  assign RetimeWrapper_71_clock = clock; // @[:@11344.4]
  assign RetimeWrapper_71_reset = reset; // @[:@11345.4]
  assign RetimeWrapper_71_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@11347.4]
  assign RetimeWrapper_71_io_in = _T_1577 & io_rPort_8_en_0; // @[package.scala 94:16:@11346.4]
  assign RetimeWrapper_72_clock = clock; // @[:@11384.4]
  assign RetimeWrapper_72_reset = reset; // @[:@11385.4]
  assign RetimeWrapper_72_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@11387.4]
  assign RetimeWrapper_72_io_in = _T_647 & io_rPort_9_en_0; // @[package.scala 94:16:@11386.4]
  assign RetimeWrapper_73_clock = clock; // @[:@11392.4]
  assign RetimeWrapper_73_reset = reset; // @[:@11393.4]
  assign RetimeWrapper_73_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@11395.4]
  assign RetimeWrapper_73_io_in = _T_771 & io_rPort_9_en_0; // @[package.scala 94:16:@11394.4]
  assign RetimeWrapper_74_clock = clock; // @[:@11400.4]
  assign RetimeWrapper_74_reset = reset; // @[:@11401.4]
  assign RetimeWrapper_74_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@11403.4]
  assign RetimeWrapper_74_io_in = _T_895 & io_rPort_9_en_0; // @[package.scala 94:16:@11402.4]
  assign RetimeWrapper_75_clock = clock; // @[:@11408.4]
  assign RetimeWrapper_75_reset = reset; // @[:@11409.4]
  assign RetimeWrapper_75_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@11411.4]
  assign RetimeWrapper_75_io_in = _T_1019 & io_rPort_9_en_0; // @[package.scala 94:16:@11410.4]
  assign RetimeWrapper_76_clock = clock; // @[:@11416.4]
  assign RetimeWrapper_76_reset = reset; // @[:@11417.4]
  assign RetimeWrapper_76_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@11419.4]
  assign RetimeWrapper_76_io_in = _T_1143 & io_rPort_9_en_0; // @[package.scala 94:16:@11418.4]
  assign RetimeWrapper_77_clock = clock; // @[:@11424.4]
  assign RetimeWrapper_77_reset = reset; // @[:@11425.4]
  assign RetimeWrapper_77_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@11427.4]
  assign RetimeWrapper_77_io_in = _T_1267 & io_rPort_9_en_0; // @[package.scala 94:16:@11426.4]
  assign RetimeWrapper_78_clock = clock; // @[:@11432.4]
  assign RetimeWrapper_78_reset = reset; // @[:@11433.4]
  assign RetimeWrapper_78_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@11435.4]
  assign RetimeWrapper_78_io_in = _T_1391 & io_rPort_9_en_0; // @[package.scala 94:16:@11434.4]
  assign RetimeWrapper_79_clock = clock; // @[:@11440.4]
  assign RetimeWrapper_79_reset = reset; // @[:@11441.4]
  assign RetimeWrapper_79_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@11443.4]
  assign RetimeWrapper_79_io_in = _T_1515 & io_rPort_9_en_0; // @[package.scala 94:16:@11442.4]
  assign RetimeWrapper_80_clock = clock; // @[:@11480.4]
  assign RetimeWrapper_80_reset = reset; // @[:@11481.4]
  assign RetimeWrapper_80_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@11483.4]
  assign RetimeWrapper_80_io_in = _T_653 & io_rPort_10_en_0; // @[package.scala 94:16:@11482.4]
  assign RetimeWrapper_81_clock = clock; // @[:@11488.4]
  assign RetimeWrapper_81_reset = reset; // @[:@11489.4]
  assign RetimeWrapper_81_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@11491.4]
  assign RetimeWrapper_81_io_in = _T_777 & io_rPort_10_en_0; // @[package.scala 94:16:@11490.4]
  assign RetimeWrapper_82_clock = clock; // @[:@11496.4]
  assign RetimeWrapper_82_reset = reset; // @[:@11497.4]
  assign RetimeWrapper_82_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@11499.4]
  assign RetimeWrapper_82_io_in = _T_901 & io_rPort_10_en_0; // @[package.scala 94:16:@11498.4]
  assign RetimeWrapper_83_clock = clock; // @[:@11504.4]
  assign RetimeWrapper_83_reset = reset; // @[:@11505.4]
  assign RetimeWrapper_83_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@11507.4]
  assign RetimeWrapper_83_io_in = _T_1025 & io_rPort_10_en_0; // @[package.scala 94:16:@11506.4]
  assign RetimeWrapper_84_clock = clock; // @[:@11512.4]
  assign RetimeWrapper_84_reset = reset; // @[:@11513.4]
  assign RetimeWrapper_84_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@11515.4]
  assign RetimeWrapper_84_io_in = _T_1149 & io_rPort_10_en_0; // @[package.scala 94:16:@11514.4]
  assign RetimeWrapper_85_clock = clock; // @[:@11520.4]
  assign RetimeWrapper_85_reset = reset; // @[:@11521.4]
  assign RetimeWrapper_85_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@11523.4]
  assign RetimeWrapper_85_io_in = _T_1273 & io_rPort_10_en_0; // @[package.scala 94:16:@11522.4]
  assign RetimeWrapper_86_clock = clock; // @[:@11528.4]
  assign RetimeWrapper_86_reset = reset; // @[:@11529.4]
  assign RetimeWrapper_86_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@11531.4]
  assign RetimeWrapper_86_io_in = _T_1397 & io_rPort_10_en_0; // @[package.scala 94:16:@11530.4]
  assign RetimeWrapper_87_clock = clock; // @[:@11536.4]
  assign RetimeWrapper_87_reset = reset; // @[:@11537.4]
  assign RetimeWrapper_87_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@11539.4]
  assign RetimeWrapper_87_io_in = _T_1521 & io_rPort_10_en_0; // @[package.scala 94:16:@11538.4]
  assign RetimeWrapper_88_clock = clock; // @[:@11576.4]
  assign RetimeWrapper_88_reset = reset; // @[:@11577.4]
  assign RetimeWrapper_88_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@11579.4]
  assign RetimeWrapper_88_io_in = _T_715 & io_rPort_11_en_0; // @[package.scala 94:16:@11578.4]
  assign RetimeWrapper_89_clock = clock; // @[:@11584.4]
  assign RetimeWrapper_89_reset = reset; // @[:@11585.4]
  assign RetimeWrapper_89_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@11587.4]
  assign RetimeWrapper_89_io_in = _T_839 & io_rPort_11_en_0; // @[package.scala 94:16:@11586.4]
  assign RetimeWrapper_90_clock = clock; // @[:@11592.4]
  assign RetimeWrapper_90_reset = reset; // @[:@11593.4]
  assign RetimeWrapper_90_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@11595.4]
  assign RetimeWrapper_90_io_in = _T_963 & io_rPort_11_en_0; // @[package.scala 94:16:@11594.4]
  assign RetimeWrapper_91_clock = clock; // @[:@11600.4]
  assign RetimeWrapper_91_reset = reset; // @[:@11601.4]
  assign RetimeWrapper_91_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@11603.4]
  assign RetimeWrapper_91_io_in = _T_1087 & io_rPort_11_en_0; // @[package.scala 94:16:@11602.4]
  assign RetimeWrapper_92_clock = clock; // @[:@11608.4]
  assign RetimeWrapper_92_reset = reset; // @[:@11609.4]
  assign RetimeWrapper_92_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@11611.4]
  assign RetimeWrapper_92_io_in = _T_1211 & io_rPort_11_en_0; // @[package.scala 94:16:@11610.4]
  assign RetimeWrapper_93_clock = clock; // @[:@11616.4]
  assign RetimeWrapper_93_reset = reset; // @[:@11617.4]
  assign RetimeWrapper_93_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@11619.4]
  assign RetimeWrapper_93_io_in = _T_1335 & io_rPort_11_en_0; // @[package.scala 94:16:@11618.4]
  assign RetimeWrapper_94_clock = clock; // @[:@11624.4]
  assign RetimeWrapper_94_reset = reset; // @[:@11625.4]
  assign RetimeWrapper_94_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@11627.4]
  assign RetimeWrapper_94_io_in = _T_1459 & io_rPort_11_en_0; // @[package.scala 94:16:@11626.4]
  assign RetimeWrapper_95_clock = clock; // @[:@11632.4]
  assign RetimeWrapper_95_reset = reset; // @[:@11633.4]
  assign RetimeWrapper_95_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@11635.4]
  assign RetimeWrapper_95_io_in = _T_1583 & io_rPort_11_en_0; // @[package.scala 94:16:@11634.4]
endmodule
module RetimeWrapper_148( // @[:@11659.2]
  input         clock, // @[:@11660.4]
  input         reset, // @[:@11661.4]
  input         io_flow, // @[:@11662.4]
  input  [15:0] io_in, // @[:@11662.4]
  output [15:0] io_out // @[:@11662.4]
);
  wire [15:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@11664.4]
  wire [15:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@11664.4]
  wire [15:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@11664.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@11664.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@11664.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@11664.4]
  RetimeShiftRegister #(.WIDTH(16), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@11664.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@11677.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@11676.4]
  assign sr_init = 16'h0; // @[RetimeShiftRegister.scala 19:16:@11675.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@11674.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@11673.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@11671.4]
endmodule
module SimBlackBoxesfix2fixBox_2( // @[:@11679.2]
  input  [31:0] io_a, // @[:@11682.4]
  output [32:0] io_b // @[:@11682.4]
);
  wire  _T_20; // @[implicits.scala 69:16:@11689.4]
  assign _T_20 = io_a[31]; // @[implicits.scala 69:16:@11689.4]
  assign io_b = {_T_20,io_a}; // @[SimBlackBoxes.scala 99:40:@11694.4]
endmodule
module __2( // @[:@11696.2]
  input  [31:0] io_b, // @[:@11699.4]
  output [32:0] io_result // @[:@11699.4]
);
  wire [31:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@11704.4]
  wire [32:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@11704.4]
  SimBlackBoxesfix2fixBox_2 SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@11704.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@11717.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@11712.4]
endmodule
module RetimeWrapper_149( // @[:@11771.2]
  input         clock, // @[:@11772.4]
  input         reset, // @[:@11773.4]
  input         io_flow, // @[:@11774.4]
  input  [31:0] io_in, // @[:@11774.4]
  output [31:0] io_out // @[:@11774.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@11776.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@11776.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@11776.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@11776.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@11776.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@11776.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@11776.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@11789.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@11788.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@11787.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@11786.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@11785.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@11783.4]
endmodule
module fix2fixBox( // @[:@11791.2]
  input         clock, // @[:@11792.4]
  input         reset, // @[:@11793.4]
  input  [32:0] io_a, // @[:@11794.4]
  input         io_flow, // @[:@11794.4]
  output [31:0] io_b // @[:@11794.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@11804.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@11804.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@11804.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@11804.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@11804.4]
  RetimeWrapper_149 RetimeWrapper ( // @[package.scala 93:22:@11804.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@11811.4]
  assign RetimeWrapper_clock = clock; // @[:@11805.4]
  assign RetimeWrapper_reset = reset; // @[:@11806.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@11808.4]
  assign RetimeWrapper_io_in = io_a[31:0]; // @[package.scala 94:16:@11807.4]
endmodule
module x297_sum( // @[:@11813.2]
  input         clock, // @[:@11814.4]
  input         reset, // @[:@11815.4]
  input  [31:0] io_a, // @[:@11816.4]
  input  [31:0] io_b, // @[:@11816.4]
  input         io_flow, // @[:@11816.4]
  output [31:0] io_result // @[:@11816.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@11824.4]
  wire [32:0] __io_result; // @[Math.scala 709:24:@11824.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@11831.4]
  wire [32:0] __1_io_result; // @[Math.scala 709:24:@11831.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@11849.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@11849.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@11849.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@11849.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@11849.4]
  wire [32:0] a_upcast_number; // @[Math.scala 712:22:@11829.4 Math.scala 713:14:@11830.4]
  wire [32:0] b_upcast_number; // @[Math.scala 712:22:@11836.4 Math.scala 713:14:@11837.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@11838.4]
  __2 _ ( // @[Math.scala 709:24:@11824.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 709:24:@11831.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox fix2fixBox ( // @[Math.scala 141:30:@11849.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@11829.4 Math.scala 713:14:@11830.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@11836.4 Math.scala 713:14:@11837.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@11838.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@11857.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@11827.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@11834.4]
  assign fix2fixBox_clock = clock; // @[:@11850.4]
  assign fix2fixBox_reset = reset; // @[:@11851.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@11852.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@11855.4]
endmodule
module RetimeWrapper_152( // @[:@11935.2]
  input         clock, // @[:@11936.4]
  input         reset, // @[:@11937.4]
  input         io_flow, // @[:@11938.4]
  input  [31:0] io_in, // @[:@11938.4]
  output [31:0] io_out // @[:@11938.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@11940.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@11940.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@11940.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@11940.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@11940.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@11940.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@11940.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@11953.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@11952.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@11951.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@11950.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@11949.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@11947.4]
endmodule
module RetimeWrapper_163( // @[:@12583.2]
  input         clock, // @[:@12584.4]
  input         reset, // @[:@12585.4]
  input         io_flow, // @[:@12586.4]
  input  [31:0] io_in, // @[:@12586.4]
  output [31:0] io_out // @[:@12586.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@12588.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@12588.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@12588.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@12588.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@12588.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@12588.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(4)) sr ( // @[RetimeShiftRegister.scala 15:20:@12588.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@12601.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@12600.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@12599.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@12598.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@12597.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@12595.4]
endmodule
module RetimeWrapper_169( // @[:@12923.2]
  input         clock, // @[:@12924.4]
  input         reset, // @[:@12925.4]
  input         io_flow, // @[:@12926.4]
  input  [31:0] io_in, // @[:@12926.4]
  output [31:0] io_out // @[:@12926.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@12928.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@12928.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@12928.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@12928.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@12928.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@12928.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(5)) sr ( // @[RetimeShiftRegister.scala 15:20:@12928.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@12941.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@12940.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@12939.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@12938.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@12937.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@12935.4]
endmodule
module RetimeWrapper_171( // @[:@12987.2]
  input   clock, // @[:@12988.4]
  input   reset, // @[:@12989.4]
  input   io_flow, // @[:@12990.4]
  input   io_in, // @[:@12990.4]
  output  io_out // @[:@12990.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@12992.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@12992.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@12992.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@12992.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@12992.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@12992.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(6)) sr ( // @[RetimeShiftRegister.scala 15:20:@12992.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@13005.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@13004.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@13003.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@13002.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@13001.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@12999.4]
endmodule
module RetimeWrapper_180( // @[:@13423.2]
  input         clock, // @[:@13424.4]
  input         reset, // @[:@13425.4]
  input         io_flow, // @[:@13426.4]
  input  [31:0] io_in, // @[:@13426.4]
  output [31:0] io_out // @[:@13426.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@13428.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@13428.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@13428.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@13428.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@13428.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@13428.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(6)) sr ( // @[RetimeShiftRegister.scala 15:20:@13428.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@13441.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@13440.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@13439.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@13438.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@13437.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@13435.4]
endmodule
module x358_rdrow( // @[:@14521.2]
  input         clock, // @[:@14522.4]
  input         reset, // @[:@14523.4]
  input  [31:0] io_a, // @[:@14524.4]
  input  [31:0] io_b, // @[:@14524.4]
  input         io_flow, // @[:@14524.4]
  output [31:0] io_result // @[:@14524.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@14532.4]
  wire [32:0] __io_result; // @[Math.scala 709:24:@14532.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@14539.4]
  wire [32:0] __1_io_result; // @[Math.scala 709:24:@14539.4]
  wire  fix2fixBox_clock; // @[Math.scala 182:30:@14558.4]
  wire  fix2fixBox_reset; // @[Math.scala 182:30:@14558.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 182:30:@14558.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 182:30:@14558.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 182:30:@14558.4]
  wire [32:0] a_upcast_number; // @[Math.scala 712:22:@14537.4 Math.scala 713:14:@14538.4]
  wire [32:0] b_upcast_number; // @[Math.scala 712:22:@14544.4 Math.scala 713:14:@14545.4]
  wire [33:0] _T_21; // @[Math.scala 177:37:@14546.4]
  wire [33:0] _T_22; // @[Math.scala 177:37:@14547.4]
  __2 _ ( // @[Math.scala 709:24:@14532.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 709:24:@14539.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox fix2fixBox ( // @[Math.scala 182:30:@14558.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@14537.4 Math.scala 713:14:@14538.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@14544.4 Math.scala 713:14:@14545.4]
  assign _T_21 = a_upcast_number - b_upcast_number; // @[Math.scala 177:37:@14546.4]
  assign _T_22 = $unsigned(_T_21); // @[Math.scala 177:37:@14547.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 188:17:@14566.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@14535.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@14542.4]
  assign fix2fixBox_clock = clock; // @[:@14559.4]
  assign fix2fixBox_reset = reset; // @[:@14560.4]
  assign fix2fixBox_io_a = _T_22[32:0]; // @[Math.scala 183:23:@14561.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 186:26:@14564.4]
endmodule
module SimBlackBoxesfix2fixBox_40( // @[:@16829.2]
  input  [7:0] io_a, // @[:@16832.4]
  output [8:0] io_b // @[:@16832.4]
);
  assign io_b = {1'h0,io_a}; // @[SimBlackBoxes.scala 99:40:@16843.4]
endmodule
module __40( // @[:@16845.2]
  input  [7:0] io_b, // @[:@16848.4]
  output [8:0] io_result // @[:@16848.4]
);
  wire [7:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@16853.4]
  wire [8:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@16853.4]
  SimBlackBoxesfix2fixBox_40 SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@16853.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@16866.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@16861.4]
endmodule
module fix2fixBox_19( // @[:@16939.2]
  input        clock, // @[:@16940.4]
  input        reset, // @[:@16941.4]
  input  [8:0] io_a, // @[:@16942.4]
  input        io_flow, // @[:@16942.4]
  output [7:0] io_b // @[:@16942.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@16952.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@16952.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@16952.4]
  wire [7:0] RetimeWrapper_io_in; // @[package.scala 93:22:@16952.4]
  wire [7:0] RetimeWrapper_io_out; // @[package.scala 93:22:@16952.4]
  RetimeWrapper_21 RetimeWrapper ( // @[package.scala 93:22:@16952.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@16959.4]
  assign RetimeWrapper_clock = clock; // @[:@16953.4]
  assign RetimeWrapper_reset = reset; // @[:@16954.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@16956.4]
  assign RetimeWrapper_io_in = io_a[7:0]; // @[package.scala 94:16:@16955.4]
endmodule
module x431_x17( // @[:@16961.2]
  input        clock, // @[:@16962.4]
  input        reset, // @[:@16963.4]
  input  [7:0] io_a, // @[:@16964.4]
  input  [7:0] io_b, // @[:@16964.4]
  input        io_flow, // @[:@16964.4]
  output [7:0] io_result // @[:@16964.4]
);
  wire [7:0] __io_b; // @[Math.scala 709:24:@16972.4]
  wire [8:0] __io_result; // @[Math.scala 709:24:@16972.4]
  wire [7:0] __1_io_b; // @[Math.scala 709:24:@16979.4]
  wire [8:0] __1_io_result; // @[Math.scala 709:24:@16979.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@16989.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@16989.4]
  wire [8:0] fix2fixBox_io_a; // @[Math.scala 141:30:@16989.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@16989.4]
  wire [7:0] fix2fixBox_io_b; // @[Math.scala 141:30:@16989.4]
  wire [8:0] a_upcast_number; // @[Math.scala 712:22:@16977.4 Math.scala 713:14:@16978.4]
  wire [8:0] b_upcast_number; // @[Math.scala 712:22:@16984.4 Math.scala 713:14:@16985.4]
  wire [9:0] _T_21; // @[Math.scala 136:37:@16986.4]
  __40 _ ( // @[Math.scala 709:24:@16972.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __40 __1 ( // @[Math.scala 709:24:@16979.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_19 fix2fixBox ( // @[Math.scala 141:30:@16989.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@16977.4 Math.scala 713:14:@16978.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@16984.4 Math.scala 713:14:@16985.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@16986.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@16997.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@16975.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@16982.4]
  assign fix2fixBox_clock = clock; // @[:@16990.4]
  assign fix2fixBox_reset = reset; // @[:@16991.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@16992.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@16995.4]
endmodule
module fix2fixBox_23( // @[:@17587.2]
  input  [8:0] io_a, // @[:@17590.4]
  output [7:0] io_b // @[:@17590.4]
);
  assign io_b = io_a[7:0]; // @[Converter.scala 95:38:@17600.4]
endmodule
module x435_x17( // @[:@17602.2]
  input  [7:0] io_a, // @[:@17605.4]
  input  [7:0] io_b, // @[:@17605.4]
  output [7:0] io_result // @[:@17605.4]
);
  wire [7:0] __io_b; // @[Math.scala 709:24:@17613.4]
  wire [8:0] __io_result; // @[Math.scala 709:24:@17613.4]
  wire [7:0] __1_io_b; // @[Math.scala 709:24:@17620.4]
  wire [8:0] __1_io_result; // @[Math.scala 709:24:@17620.4]
  wire [8:0] fix2fixBox_io_a; // @[Math.scala 141:30:@17630.4]
  wire [7:0] fix2fixBox_io_b; // @[Math.scala 141:30:@17630.4]
  wire [8:0] a_upcast_number; // @[Math.scala 712:22:@17618.4 Math.scala 713:14:@17619.4]
  wire [8:0] b_upcast_number; // @[Math.scala 712:22:@17625.4 Math.scala 713:14:@17626.4]
  wire [9:0] _T_21; // @[Math.scala 136:37:@17627.4]
  __40 _ ( // @[Math.scala 709:24:@17613.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __40 __1 ( // @[Math.scala 709:24:@17620.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_23 fix2fixBox ( // @[Math.scala 141:30:@17630.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@17618.4 Math.scala 713:14:@17619.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@17625.4 Math.scala 713:14:@17626.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@17627.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@17638.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@17616.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@17623.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@17633.4]
endmodule
module RetimeWrapper_228( // @[:@18109.2]
  input        clock, // @[:@18110.4]
  input        reset, // @[:@18111.4]
  input        io_flow, // @[:@18112.4]
  input  [7:0] io_in, // @[:@18112.4]
  output [7:0] io_out // @[:@18112.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@18114.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@18114.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@18114.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@18114.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@18114.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@18114.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@18114.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@18127.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@18126.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@18125.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@18124.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@18123.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@18121.4]
endmodule
module x440_sub( // @[:@18222.2]
  input  [7:0] io_a, // @[:@18225.4]
  input  [7:0] io_b, // @[:@18225.4]
  output [7:0] io_result // @[:@18225.4]
);
  wire [7:0] __io_b; // @[Math.scala 709:24:@18233.4]
  wire [8:0] __io_result; // @[Math.scala 709:24:@18233.4]
  wire [7:0] __1_io_b; // @[Math.scala 709:24:@18240.4]
  wire [8:0] __1_io_result; // @[Math.scala 709:24:@18240.4]
  wire [8:0] fix2fixBox_io_a; // @[Math.scala 182:30:@18251.4]
  wire [7:0] fix2fixBox_io_b; // @[Math.scala 182:30:@18251.4]
  wire [8:0] a_upcast_number; // @[Math.scala 712:22:@18238.4 Math.scala 713:14:@18239.4]
  wire [8:0] b_upcast_number; // @[Math.scala 712:22:@18245.4 Math.scala 713:14:@18246.4]
  wire [9:0] _T_21; // @[Math.scala 177:37:@18247.4]
  wire [9:0] _T_22; // @[Math.scala 177:37:@18248.4]
  __40 _ ( // @[Math.scala 709:24:@18233.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __40 __1 ( // @[Math.scala 709:24:@18240.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_23 fix2fixBox ( // @[Math.scala 182:30:@18251.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@18238.4 Math.scala 713:14:@18239.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@18245.4 Math.scala 713:14:@18246.4]
  assign _T_21 = a_upcast_number - b_upcast_number; // @[Math.scala 177:37:@18247.4]
  assign _T_22 = $unsigned(_T_21); // @[Math.scala 177:37:@18248.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 188:17:@18259.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@18236.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@18243.4]
  assign fix2fixBox_io_a = _T_22[8:0]; // @[Math.scala 183:23:@18254.4]
endmodule
module RetimeWrapper_230( // @[:@18305.2]
  input        clock, // @[:@18306.4]
  input        reset, // @[:@18307.4]
  input        io_flow, // @[:@18308.4]
  input  [7:0] io_in, // @[:@18308.4]
  output [7:0] io_out // @[:@18308.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@18310.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@18310.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@18310.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@18310.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@18310.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@18310.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(5)) sr ( // @[RetimeShiftRegister.scala 15:20:@18310.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@18323.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@18322.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@18321.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@18320.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@18319.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@18317.4]
endmodule
module SimBlackBoxesfix2fixBox_58( // @[:@18325.2]
  input  [7:0] io_a, // @[:@18328.4]
  output [7:0] io_b // @[:@18328.4]
);
  assign io_b = io_a; // @[SimBlackBoxes.scala 99:40:@18338.4]
endmodule
module __58( // @[:@18340.2]
  input  [7:0] io_b, // @[:@18343.4]
  output [7:0] io_result // @[:@18343.4]
);
  wire [7:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@18348.4]
  wire [7:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@18348.4]
  SimBlackBoxesfix2fixBox_58 SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@18348.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@18361.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@18356.4]
endmodule
module x444_div( // @[:@18363.2]
  input        clock, // @[:@18364.4]
  input        reset, // @[:@18365.4]
  input  [7:0] io_a, // @[:@18366.4]
  input        io_flow, // @[:@18366.4]
  output [7:0] io_result // @[:@18366.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@18373.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@18373.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@18373.4]
  wire [7:0] RetimeWrapper_io_in; // @[package.scala 93:22:@18373.4]
  wire [7:0] RetimeWrapper_io_out; // @[package.scala 93:22:@18373.4]
  wire [7:0] __io_b; // @[Math.scala 709:24:@18383.4]
  wire [7:0] __io_result; // @[Math.scala 709:24:@18383.4]
  RetimeWrapper_230 RetimeWrapper ( // @[package.scala 93:22:@18373.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  __58 _ ( // @[Math.scala 709:24:@18383.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  assign io_result = __io_result; // @[Math.scala 291:34:@18391.4]
  assign RetimeWrapper_clock = clock; // @[:@18374.4]
  assign RetimeWrapper_reset = reset; // @[:@18375.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@18377.4]
  assign RetimeWrapper_io_in = io_a / 8'h5; // @[package.scala 94:16:@18376.4]
  assign __io_b = RetimeWrapper_io_out; // @[Math.scala 710:17:@18386.4]
endmodule
module RetimeWrapper_231( // @[:@18405.2]
  input        clock, // @[:@18406.4]
  input        reset, // @[:@18407.4]
  input        io_flow, // @[:@18408.4]
  input  [7:0] io_in, // @[:@18408.4]
  output [7:0] io_out // @[:@18408.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@18410.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@18410.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@18410.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@18410.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@18410.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@18410.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(8)) sr ( // @[RetimeShiftRegister.scala 15:20:@18410.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@18423.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@18422.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@18421.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@18420.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@18419.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@18417.4]
endmodule
module RetimeWrapper_232( // @[:@18568.2]
  input        clock, // @[:@18569.4]
  input        reset, // @[:@18570.4]
  input        io_flow, // @[:@18571.4]
  input  [7:0] io_in, // @[:@18571.4]
  output [7:0] io_out // @[:@18571.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@18573.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@18573.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@18573.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@18573.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@18573.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@18573.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(6)) sr ( // @[RetimeShiftRegister.scala 15:20:@18573.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@18586.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@18585.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@18584.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@18583.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@18582.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@18580.4]
endmodule
module RetimeWrapper_246( // @[:@20423.2]
  input         clock, // @[:@20424.4]
  input         reset, // @[:@20425.4]
  input         io_flow, // @[:@20426.4]
  input  [15:0] io_in, // @[:@20426.4]
  output [15:0] io_out // @[:@20426.4]
);
  wire [15:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@20428.4]
  wire [15:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@20428.4]
  wire [15:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@20428.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@20428.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@20428.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@20428.4]
  RetimeShiftRegister #(.WIDTH(16), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@20428.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@20441.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@20440.4]
  assign sr_init = 16'h0; // @[RetimeShiftRegister.scala 19:16:@20439.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@20438.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@20437.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@20435.4]
endmodule
module x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1( // @[:@20539.2]
  input          clock, // @[:@20540.4]
  input          reset, // @[:@20541.4]
  output         io_in_x270_TREADY, // @[:@20542.4]
  input  [255:0] io_in_x270_TDATA, // @[:@20542.4]
  input  [7:0]   io_in_x270_TID, // @[:@20542.4]
  input  [7:0]   io_in_x270_TDEST, // @[:@20542.4]
  output         io_in_x271_TVALID, // @[:@20542.4]
  input          io_in_x271_TREADY, // @[:@20542.4]
  output [255:0] io_in_x271_TDATA, // @[:@20542.4]
  input          io_sigsIn_backpressure, // @[:@20542.4]
  input          io_sigsIn_datapathEn, // @[:@20542.4]
  input          io_sigsIn_break, // @[:@20542.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_1, // @[:@20542.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_0, // @[:@20542.4]
  input          io_sigsIn_cchainOutputs_0_oobs_0, // @[:@20542.4]
  input          io_sigsIn_cchainOutputs_0_oobs_1, // @[:@20542.4]
  input          io_rr // @[:@20542.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@20556.4]
  wire [31:0] __io_result; // @[Math.scala 709:24:@20556.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@20568.4]
  wire [31:0] __1_io_result; // @[Math.scala 709:24:@20568.4]
  wire  x283_lb_0_clock; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire  x283_lb_0_reset; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire [2:0] x283_lb_0_io_rPort_11_banks_1; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire [2:0] x283_lb_0_io_rPort_11_banks_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire  x283_lb_0_io_rPort_11_ofs_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire  x283_lb_0_io_rPort_11_en_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire  x283_lb_0_io_rPort_11_backpressure; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire [7:0] x283_lb_0_io_rPort_11_output_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire [2:0] x283_lb_0_io_rPort_10_banks_1; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire [2:0] x283_lb_0_io_rPort_10_banks_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire  x283_lb_0_io_rPort_10_ofs_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire  x283_lb_0_io_rPort_10_en_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire  x283_lb_0_io_rPort_10_backpressure; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire [7:0] x283_lb_0_io_rPort_10_output_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire [2:0] x283_lb_0_io_rPort_9_banks_1; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire [2:0] x283_lb_0_io_rPort_9_banks_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire  x283_lb_0_io_rPort_9_ofs_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire  x283_lb_0_io_rPort_9_en_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire  x283_lb_0_io_rPort_9_backpressure; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire [7:0] x283_lb_0_io_rPort_9_output_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire [2:0] x283_lb_0_io_rPort_8_banks_1; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire [2:0] x283_lb_0_io_rPort_8_banks_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire  x283_lb_0_io_rPort_8_ofs_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire  x283_lb_0_io_rPort_8_en_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire  x283_lb_0_io_rPort_8_backpressure; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire [7:0] x283_lb_0_io_rPort_8_output_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire [2:0] x283_lb_0_io_rPort_7_banks_1; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire [2:0] x283_lb_0_io_rPort_7_banks_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire  x283_lb_0_io_rPort_7_ofs_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire  x283_lb_0_io_rPort_7_en_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire  x283_lb_0_io_rPort_7_backpressure; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire [7:0] x283_lb_0_io_rPort_7_output_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire [2:0] x283_lb_0_io_rPort_6_banks_1; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire [2:0] x283_lb_0_io_rPort_6_banks_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire  x283_lb_0_io_rPort_6_ofs_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire  x283_lb_0_io_rPort_6_en_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire  x283_lb_0_io_rPort_6_backpressure; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire [7:0] x283_lb_0_io_rPort_6_output_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire [2:0] x283_lb_0_io_rPort_5_banks_1; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire [2:0] x283_lb_0_io_rPort_5_banks_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire  x283_lb_0_io_rPort_5_ofs_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire  x283_lb_0_io_rPort_5_en_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire  x283_lb_0_io_rPort_5_backpressure; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire [7:0] x283_lb_0_io_rPort_5_output_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire [2:0] x283_lb_0_io_rPort_4_banks_1; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire [2:0] x283_lb_0_io_rPort_4_banks_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire  x283_lb_0_io_rPort_4_ofs_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire  x283_lb_0_io_rPort_4_en_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire  x283_lb_0_io_rPort_4_backpressure; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire [7:0] x283_lb_0_io_rPort_4_output_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire [2:0] x283_lb_0_io_rPort_3_banks_1; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire [2:0] x283_lb_0_io_rPort_3_banks_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire  x283_lb_0_io_rPort_3_ofs_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire  x283_lb_0_io_rPort_3_en_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire  x283_lb_0_io_rPort_3_backpressure; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire [7:0] x283_lb_0_io_rPort_3_output_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire [2:0] x283_lb_0_io_rPort_2_banks_1; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire [2:0] x283_lb_0_io_rPort_2_banks_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire  x283_lb_0_io_rPort_2_ofs_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire  x283_lb_0_io_rPort_2_en_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire  x283_lb_0_io_rPort_2_backpressure; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire [7:0] x283_lb_0_io_rPort_2_output_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire [2:0] x283_lb_0_io_rPort_1_banks_1; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire [2:0] x283_lb_0_io_rPort_1_banks_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire  x283_lb_0_io_rPort_1_ofs_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire  x283_lb_0_io_rPort_1_en_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire  x283_lb_0_io_rPort_1_backpressure; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire [7:0] x283_lb_0_io_rPort_1_output_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire [2:0] x283_lb_0_io_rPort_0_banks_1; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire [2:0] x283_lb_0_io_rPort_0_banks_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire  x283_lb_0_io_rPort_0_ofs_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire  x283_lb_0_io_rPort_0_en_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire  x283_lb_0_io_rPort_0_backpressure; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire [7:0] x283_lb_0_io_rPort_0_output_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire [2:0] x283_lb_0_io_wPort_1_banks_1; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire [2:0] x283_lb_0_io_wPort_1_banks_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire  x283_lb_0_io_wPort_1_ofs_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire [7:0] x283_lb_0_io_wPort_1_data_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire  x283_lb_0_io_wPort_1_en_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire [2:0] x283_lb_0_io_wPort_0_banks_1; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire [2:0] x283_lb_0_io_wPort_0_banks_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire  x283_lb_0_io_wPort_0_ofs_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire [7:0] x283_lb_0_io_wPort_0_data_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire  x283_lb_0_io_wPort_0_en_0; // @[m_x283_lb_0.scala 39:17:@20578.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@20684.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@20684.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@20684.4]
  wire [15:0] RetimeWrapper_io_in; // @[package.scala 93:22:@20684.4]
  wire [15:0] RetimeWrapper_io_out; // @[package.scala 93:22:@20684.4]
  wire  x297_sum_1_clock; // @[Math.scala 150:24:@20791.4]
  wire  x297_sum_1_reset; // @[Math.scala 150:24:@20791.4]
  wire [31:0] x297_sum_1_io_a; // @[Math.scala 150:24:@20791.4]
  wire [31:0] x297_sum_1_io_b; // @[Math.scala 150:24:@20791.4]
  wire  x297_sum_1_io_flow; // @[Math.scala 150:24:@20791.4]
  wire [31:0] x297_sum_1_io_result; // @[Math.scala 150:24:@20791.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@20801.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@20801.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@20801.4]
  wire [7:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@20801.4]
  wire [7:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@20801.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@20810.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@20810.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@20810.4]
  wire [31:0] RetimeWrapper_2_io_in; // @[package.scala 93:22:@20810.4]
  wire [31:0] RetimeWrapper_2_io_out; // @[package.scala 93:22:@20810.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@20819.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@20819.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@20819.4]
  wire [31:0] RetimeWrapper_3_io_in; // @[package.scala 93:22:@20819.4]
  wire [31:0] RetimeWrapper_3_io_out; // @[package.scala 93:22:@20819.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@20828.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@20828.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@20828.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@20828.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@20828.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@20837.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@20837.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@20837.4]
  wire [31:0] RetimeWrapper_5_io_in; // @[package.scala 93:22:@20837.4]
  wire [31:0] RetimeWrapper_5_io_out; // @[package.scala 93:22:@20837.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@20846.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@20846.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@20846.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@20846.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@20846.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@20857.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@20857.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@20857.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@20857.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@20857.4]
  wire  x303_rdcol_1_clock; // @[Math.scala 150:24:@20880.4]
  wire  x303_rdcol_1_reset; // @[Math.scala 150:24:@20880.4]
  wire [31:0] x303_rdcol_1_io_a; // @[Math.scala 150:24:@20880.4]
  wire [31:0] x303_rdcol_1_io_b; // @[Math.scala 150:24:@20880.4]
  wire  x303_rdcol_1_io_flow; // @[Math.scala 150:24:@20880.4]
  wire [31:0] x303_rdcol_1_io_result; // @[Math.scala 150:24:@20880.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@20912.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@20912.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@20912.4]
  wire [31:0] RetimeWrapper_8_io_in; // @[package.scala 93:22:@20912.4]
  wire [31:0] RetimeWrapper_8_io_out; // @[package.scala 93:22:@20912.4]
  wire  x307_sum_1_clock; // @[Math.scala 150:24:@20921.4]
  wire  x307_sum_1_reset; // @[Math.scala 150:24:@20921.4]
  wire [31:0] x307_sum_1_io_a; // @[Math.scala 150:24:@20921.4]
  wire [31:0] x307_sum_1_io_b; // @[Math.scala 150:24:@20921.4]
  wire  x307_sum_1_io_flow; // @[Math.scala 150:24:@20921.4]
  wire [31:0] x307_sum_1_io_result; // @[Math.scala 150:24:@20921.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@20931.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@20931.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@20931.4]
  wire [31:0] RetimeWrapper_9_io_in; // @[package.scala 93:22:@20931.4]
  wire [31:0] RetimeWrapper_9_io_out; // @[package.scala 93:22:@20931.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@20940.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@20940.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@20940.4]
  wire [7:0] RetimeWrapper_10_io_in; // @[package.scala 93:22:@20940.4]
  wire [7:0] RetimeWrapper_10_io_out; // @[package.scala 93:22:@20940.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@20951.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@20951.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@20951.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@20951.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@20951.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@20972.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@20972.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@20972.4]
  wire [31:0] RetimeWrapper_12_io_in; // @[package.scala 93:22:@20972.4]
  wire [31:0] RetimeWrapper_12_io_out; // @[package.scala 93:22:@20972.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@20999.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@20999.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@20999.4]
  wire [31:0] RetimeWrapper_13_io_in; // @[package.scala 93:22:@20999.4]
  wire [31:0] RetimeWrapper_13_io_out; // @[package.scala 93:22:@20999.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@21015.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@21015.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@21015.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@21015.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@21015.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@21050.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@21050.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@21050.4]
  wire [31:0] RetimeWrapper_15_io_in; // @[package.scala 93:22:@21050.4]
  wire [31:0] RetimeWrapper_15_io_out; // @[package.scala 93:22:@21050.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@21059.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@21059.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@21059.4]
  wire [31:0] RetimeWrapper_16_io_in; // @[package.scala 93:22:@21059.4]
  wire [31:0] RetimeWrapper_16_io_out; // @[package.scala 93:22:@21059.4]
  wire  x320_sum_1_clock; // @[Math.scala 150:24:@21068.4]
  wire  x320_sum_1_reset; // @[Math.scala 150:24:@21068.4]
  wire [31:0] x320_sum_1_io_a; // @[Math.scala 150:24:@21068.4]
  wire [31:0] x320_sum_1_io_b; // @[Math.scala 150:24:@21068.4]
  wire  x320_sum_1_io_flow; // @[Math.scala 150:24:@21068.4]
  wire [31:0] x320_sum_1_io_result; // @[Math.scala 150:24:@21068.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@21078.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@21078.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@21078.4]
  wire [31:0] RetimeWrapper_17_io_in; // @[package.scala 93:22:@21078.4]
  wire [31:0] RetimeWrapper_17_io_out; // @[package.scala 93:22:@21078.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@21087.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@21087.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@21087.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@21087.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@21087.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@21096.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@21096.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@21096.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@21096.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@21096.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@21105.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@21105.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@21105.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@21105.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@21105.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@21114.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@21114.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@21114.4]
  wire [31:0] RetimeWrapper_21_io_in; // @[package.scala 93:22:@21114.4]
  wire [31:0] RetimeWrapper_21_io_out; // @[package.scala 93:22:@21114.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@21126.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@21126.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@21126.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@21126.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@21126.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@21147.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@21147.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@21147.4]
  wire [31:0] RetimeWrapper_23_io_in; // @[package.scala 93:22:@21147.4]
  wire [31:0] RetimeWrapper_23_io_out; // @[package.scala 93:22:@21147.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@21171.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@21171.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@21171.4]
  wire [31:0] RetimeWrapper_24_io_in; // @[package.scala 93:22:@21171.4]
  wire [31:0] RetimeWrapper_24_io_out; // @[package.scala 93:22:@21171.4]
  wire  x329_sum_1_clock; // @[Math.scala 150:24:@21180.4]
  wire  x329_sum_1_reset; // @[Math.scala 150:24:@21180.4]
  wire [31:0] x329_sum_1_io_a; // @[Math.scala 150:24:@21180.4]
  wire [31:0] x329_sum_1_io_b; // @[Math.scala 150:24:@21180.4]
  wire  x329_sum_1_io_flow; // @[Math.scala 150:24:@21180.4]
  wire [31:0] x329_sum_1_io_result; // @[Math.scala 150:24:@21180.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@21190.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@21190.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@21190.4]
  wire [31:0] RetimeWrapper_25_io_in; // @[package.scala 93:22:@21190.4]
  wire [31:0] RetimeWrapper_25_io_out; // @[package.scala 93:22:@21190.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@21199.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@21199.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@21199.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@21199.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@21199.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@21208.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@21208.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@21208.4]
  wire [31:0] RetimeWrapper_27_io_in; // @[package.scala 93:22:@21208.4]
  wire [31:0] RetimeWrapper_27_io_out; // @[package.scala 93:22:@21208.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@21220.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@21220.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@21220.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@21220.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@21220.4]
  wire  x334_rdcol_1_clock; // @[Math.scala 150:24:@21243.4]
  wire  x334_rdcol_1_reset; // @[Math.scala 150:24:@21243.4]
  wire [31:0] x334_rdcol_1_io_a; // @[Math.scala 150:24:@21243.4]
  wire [31:0] x334_rdcol_1_io_b; // @[Math.scala 150:24:@21243.4]
  wire  x334_rdcol_1_io_flow; // @[Math.scala 150:24:@21243.4]
  wire [31:0] x334_rdcol_1_io_result; // @[Math.scala 150:24:@21243.4]
  wire  x340_sum_1_clock; // @[Math.scala 150:24:@21286.4]
  wire  x340_sum_1_reset; // @[Math.scala 150:24:@21286.4]
  wire [31:0] x340_sum_1_io_a; // @[Math.scala 150:24:@21286.4]
  wire [31:0] x340_sum_1_io_b; // @[Math.scala 150:24:@21286.4]
  wire  x340_sum_1_io_flow; // @[Math.scala 150:24:@21286.4]
  wire [31:0] x340_sum_1_io_result; // @[Math.scala 150:24:@21286.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@21296.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@21296.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@21296.4]
  wire [31:0] RetimeWrapper_29_io_in; // @[package.scala 93:22:@21296.4]
  wire [31:0] RetimeWrapper_29_io_out; // @[package.scala 93:22:@21296.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@21305.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@21305.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@21305.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@21305.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@21305.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@21317.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@21317.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@21317.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@21317.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@21317.4]
  wire  x346_rdcol_1_clock; // @[Math.scala 150:24:@21340.4]
  wire  x346_rdcol_1_reset; // @[Math.scala 150:24:@21340.4]
  wire [31:0] x346_rdcol_1_io_a; // @[Math.scala 150:24:@21340.4]
  wire [31:0] x346_rdcol_1_io_b; // @[Math.scala 150:24:@21340.4]
  wire  x346_rdcol_1_io_flow; // @[Math.scala 150:24:@21340.4]
  wire [31:0] x346_rdcol_1_io_result; // @[Math.scala 150:24:@21340.4]
  wire  x352_sum_1_clock; // @[Math.scala 150:24:@21383.4]
  wire  x352_sum_1_reset; // @[Math.scala 150:24:@21383.4]
  wire [31:0] x352_sum_1_io_a; // @[Math.scala 150:24:@21383.4]
  wire [31:0] x352_sum_1_io_b; // @[Math.scala 150:24:@21383.4]
  wire  x352_sum_1_io_flow; // @[Math.scala 150:24:@21383.4]
  wire [31:0] x352_sum_1_io_result; // @[Math.scala 150:24:@21383.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@21393.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@21393.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@21393.4]
  wire [31:0] RetimeWrapper_32_io_in; // @[package.scala 93:22:@21393.4]
  wire [31:0] RetimeWrapper_32_io_out; // @[package.scala 93:22:@21393.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@21402.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@21402.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@21402.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@21402.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@21402.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@21414.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@21414.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@21414.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@21414.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@21414.4]
  wire  x358_rdrow_1_clock; // @[Math.scala 191:24:@21437.4]
  wire  x358_rdrow_1_reset; // @[Math.scala 191:24:@21437.4]
  wire [31:0] x358_rdrow_1_io_a; // @[Math.scala 191:24:@21437.4]
  wire [31:0] x358_rdrow_1_io_b; // @[Math.scala 191:24:@21437.4]
  wire  x358_rdrow_1_io_flow; // @[Math.scala 191:24:@21437.4]
  wire [31:0] x358_rdrow_1_io_result; // @[Math.scala 191:24:@21437.4]
  wire  x365_sum_1_clock; // @[Math.scala 150:24:@21491.4]
  wire  x365_sum_1_reset; // @[Math.scala 150:24:@21491.4]
  wire [31:0] x365_sum_1_io_a; // @[Math.scala 150:24:@21491.4]
  wire [31:0] x365_sum_1_io_b; // @[Math.scala 150:24:@21491.4]
  wire  x365_sum_1_io_flow; // @[Math.scala 150:24:@21491.4]
  wire [31:0] x365_sum_1_io_result; // @[Math.scala 150:24:@21491.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@21501.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@21501.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@21501.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@21501.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@21501.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@21510.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@21510.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@21510.4]
  wire [31:0] RetimeWrapper_36_io_in; // @[package.scala 93:22:@21510.4]
  wire [31:0] RetimeWrapper_36_io_out; // @[package.scala 93:22:@21510.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@21522.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@21522.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@21522.4]
  wire  RetimeWrapper_37_io_in; // @[package.scala 93:22:@21522.4]
  wire  RetimeWrapper_37_io_out; // @[package.scala 93:22:@21522.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@21543.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@21543.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@21543.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@21543.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@21543.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@21558.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@21558.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@21558.4]
  wire [31:0] RetimeWrapper_39_io_in; // @[package.scala 93:22:@21558.4]
  wire [31:0] RetimeWrapper_39_io_out; // @[package.scala 93:22:@21558.4]
  wire  x373_sum_1_clock; // @[Math.scala 150:24:@21569.4]
  wire  x373_sum_1_reset; // @[Math.scala 150:24:@21569.4]
  wire [31:0] x373_sum_1_io_a; // @[Math.scala 150:24:@21569.4]
  wire [31:0] x373_sum_1_io_b; // @[Math.scala 150:24:@21569.4]
  wire  x373_sum_1_io_flow; // @[Math.scala 150:24:@21569.4]
  wire [31:0] x373_sum_1_io_result; // @[Math.scala 150:24:@21569.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@21579.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@21579.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@21579.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@21579.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@21579.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@21591.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@21591.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@21591.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@21591.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@21591.4]
  wire  x380_sum_1_clock; // @[Math.scala 150:24:@21618.4]
  wire  x380_sum_1_reset; // @[Math.scala 150:24:@21618.4]
  wire [31:0] x380_sum_1_io_a; // @[Math.scala 150:24:@21618.4]
  wire [31:0] x380_sum_1_io_b; // @[Math.scala 150:24:@21618.4]
  wire  x380_sum_1_io_flow; // @[Math.scala 150:24:@21618.4]
  wire [31:0] x380_sum_1_io_result; // @[Math.scala 150:24:@21618.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@21628.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@21628.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@21628.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@21628.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@21628.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@21640.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@21640.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@21640.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@21640.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@21640.4]
  wire  x387_sum_1_clock; // @[Math.scala 150:24:@21667.4]
  wire  x387_sum_1_reset; // @[Math.scala 150:24:@21667.4]
  wire [31:0] x387_sum_1_io_a; // @[Math.scala 150:24:@21667.4]
  wire [31:0] x387_sum_1_io_b; // @[Math.scala 150:24:@21667.4]
  wire  x387_sum_1_io_flow; // @[Math.scala 150:24:@21667.4]
  wire [31:0] x387_sum_1_io_result; // @[Math.scala 150:24:@21667.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@21677.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@21677.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@21677.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@21677.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@21677.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@21689.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@21689.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@21689.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@21689.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@21689.4]
  wire  x392_rdrow_1_clock; // @[Math.scala 191:24:@21712.4]
  wire  x392_rdrow_1_reset; // @[Math.scala 191:24:@21712.4]
  wire [31:0] x392_rdrow_1_io_a; // @[Math.scala 191:24:@21712.4]
  wire [31:0] x392_rdrow_1_io_b; // @[Math.scala 191:24:@21712.4]
  wire  x392_rdrow_1_io_flow; // @[Math.scala 191:24:@21712.4]
  wire [31:0] x392_rdrow_1_io_result; // @[Math.scala 191:24:@21712.4]
  wire  x399_sum_1_clock; // @[Math.scala 150:24:@21766.4]
  wire  x399_sum_1_reset; // @[Math.scala 150:24:@21766.4]
  wire [31:0] x399_sum_1_io_a; // @[Math.scala 150:24:@21766.4]
  wire [31:0] x399_sum_1_io_b; // @[Math.scala 150:24:@21766.4]
  wire  x399_sum_1_io_flow; // @[Math.scala 150:24:@21766.4]
  wire [31:0] x399_sum_1_io_result; // @[Math.scala 150:24:@21766.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@21776.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@21776.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@21776.4]
  wire [31:0] RetimeWrapper_46_io_in; // @[package.scala 93:22:@21776.4]
  wire [31:0] RetimeWrapper_46_io_out; // @[package.scala 93:22:@21776.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@21785.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@21785.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@21785.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@21785.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@21785.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@21797.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@21797.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@21797.4]
  wire  RetimeWrapper_48_io_in; // @[package.scala 93:22:@21797.4]
  wire  RetimeWrapper_48_io_out; // @[package.scala 93:22:@21797.4]
  wire  x407_sum_1_clock; // @[Math.scala 150:24:@21824.4]
  wire  x407_sum_1_reset; // @[Math.scala 150:24:@21824.4]
  wire [31:0] x407_sum_1_io_a; // @[Math.scala 150:24:@21824.4]
  wire [31:0] x407_sum_1_io_b; // @[Math.scala 150:24:@21824.4]
  wire  x407_sum_1_io_flow; // @[Math.scala 150:24:@21824.4]
  wire [31:0] x407_sum_1_io_result; // @[Math.scala 150:24:@21824.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@21834.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@21834.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@21834.4]
  wire  RetimeWrapper_49_io_in; // @[package.scala 93:22:@21834.4]
  wire  RetimeWrapper_49_io_out; // @[package.scala 93:22:@21834.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@21846.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@21846.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@21846.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@21846.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@21846.4]
  wire  x414_sum_1_clock; // @[Math.scala 150:24:@21873.4]
  wire  x414_sum_1_reset; // @[Math.scala 150:24:@21873.4]
  wire [31:0] x414_sum_1_io_a; // @[Math.scala 150:24:@21873.4]
  wire [31:0] x414_sum_1_io_b; // @[Math.scala 150:24:@21873.4]
  wire  x414_sum_1_io_flow; // @[Math.scala 150:24:@21873.4]
  wire [31:0] x414_sum_1_io_result; // @[Math.scala 150:24:@21873.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@21883.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@21883.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@21883.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@21883.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@21883.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@21895.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@21895.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@21895.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@21895.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@21895.4]
  wire  x421_sum_1_clock; // @[Math.scala 150:24:@21922.4]
  wire  x421_sum_1_reset; // @[Math.scala 150:24:@21922.4]
  wire [31:0] x421_sum_1_io_a; // @[Math.scala 150:24:@21922.4]
  wire [31:0] x421_sum_1_io_b; // @[Math.scala 150:24:@21922.4]
  wire  x421_sum_1_io_flow; // @[Math.scala 150:24:@21922.4]
  wire [31:0] x421_sum_1_io_result; // @[Math.scala 150:24:@21922.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@21932.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@21932.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@21932.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@21932.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@21932.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@21944.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@21944.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@21944.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@21944.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@21944.4]
  wire  x431_x17_1_clock; // @[Math.scala 150:24:@21992.4]
  wire  x431_x17_1_reset; // @[Math.scala 150:24:@21992.4]
  wire [7:0] x431_x17_1_io_a; // @[Math.scala 150:24:@21992.4]
  wire [7:0] x431_x17_1_io_b; // @[Math.scala 150:24:@21992.4]
  wire  x431_x17_1_io_flow; // @[Math.scala 150:24:@21992.4]
  wire [7:0] x431_x17_1_io_result; // @[Math.scala 150:24:@21992.4]
  wire  x432_x18_1_clock; // @[Math.scala 150:24:@22002.4]
  wire  x432_x18_1_reset; // @[Math.scala 150:24:@22002.4]
  wire [7:0] x432_x18_1_io_a; // @[Math.scala 150:24:@22002.4]
  wire [7:0] x432_x18_1_io_b; // @[Math.scala 150:24:@22002.4]
  wire  x432_x18_1_io_flow; // @[Math.scala 150:24:@22002.4]
  wire [7:0] x432_x18_1_io_result; // @[Math.scala 150:24:@22002.4]
  wire  x433_x17_1_clock; // @[Math.scala 150:24:@22012.4]
  wire  x433_x17_1_reset; // @[Math.scala 150:24:@22012.4]
  wire [7:0] x433_x17_1_io_a; // @[Math.scala 150:24:@22012.4]
  wire [7:0] x433_x17_1_io_b; // @[Math.scala 150:24:@22012.4]
  wire  x433_x17_1_io_flow; // @[Math.scala 150:24:@22012.4]
  wire [7:0] x433_x17_1_io_result; // @[Math.scala 150:24:@22012.4]
  wire  x434_x18_1_clock; // @[Math.scala 150:24:@22022.4]
  wire  x434_x18_1_reset; // @[Math.scala 150:24:@22022.4]
  wire [7:0] x434_x18_1_io_a; // @[Math.scala 150:24:@22022.4]
  wire [7:0] x434_x18_1_io_b; // @[Math.scala 150:24:@22022.4]
  wire  x434_x18_1_io_flow; // @[Math.scala 150:24:@22022.4]
  wire [7:0] x434_x18_1_io_result; // @[Math.scala 150:24:@22022.4]
  wire [7:0] x435_x17_1_io_a; // @[Math.scala 150:24:@22032.4]
  wire [7:0] x435_x17_1_io_b; // @[Math.scala 150:24:@22032.4]
  wire [7:0] x435_x17_1_io_result; // @[Math.scala 150:24:@22032.4]
  wire [7:0] x436_x18_1_io_a; // @[Math.scala 150:24:@22042.4]
  wire [7:0] x436_x18_1_io_b; // @[Math.scala 150:24:@22042.4]
  wire [7:0] x436_x18_1_io_result; // @[Math.scala 150:24:@22042.4]
  wire [7:0] x437_x17_1_io_a; // @[Math.scala 150:24:@22052.4]
  wire [7:0] x437_x17_1_io_b; // @[Math.scala 150:24:@22052.4]
  wire [7:0] x437_x17_1_io_result; // @[Math.scala 150:24:@22052.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@22062.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@22062.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@22062.4]
  wire [7:0] RetimeWrapper_55_io_in; // @[package.scala 93:22:@22062.4]
  wire [7:0] RetimeWrapper_55_io_out; // @[package.scala 93:22:@22062.4]
  wire [7:0] x438_sum_1_io_a; // @[Math.scala 150:24:@22071.4]
  wire [7:0] x438_sum_1_io_b; // @[Math.scala 150:24:@22071.4]
  wire [7:0] x438_sum_1_io_result; // @[Math.scala 150:24:@22071.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@22085.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@22085.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@22085.4]
  wire [7:0] RetimeWrapper_56_io_in; // @[package.scala 93:22:@22085.4]
  wire [7:0] RetimeWrapper_56_io_out; // @[package.scala 93:22:@22085.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@22095.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@22095.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@22095.4]
  wire [7:0] RetimeWrapper_57_io_in; // @[package.scala 93:22:@22095.4]
  wire [7:0] RetimeWrapper_57_io_out; // @[package.scala 93:22:@22095.4]
  wire [7:0] x440_sub_1_io_a; // @[Math.scala 191:24:@22104.4]
  wire [7:0] x440_sub_1_io_b; // @[Math.scala 191:24:@22104.4]
  wire [7:0] x440_sub_1_io_result; // @[Math.scala 191:24:@22104.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@22129.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@22129.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@22129.4]
  wire [7:0] RetimeWrapper_58_io_in; // @[package.scala 93:22:@22129.4]
  wire [7:0] RetimeWrapper_58_io_out; // @[package.scala 93:22:@22129.4]
  wire  x444_div_1_clock; // @[Math.scala 327:24:@22140.4]
  wire  x444_div_1_reset; // @[Math.scala 327:24:@22140.4]
  wire [7:0] x444_div_1_io_a; // @[Math.scala 327:24:@22140.4]
  wire  x444_div_1_io_flow; // @[Math.scala 327:24:@22140.4]
  wire [7:0] x444_div_1_io_result; // @[Math.scala 327:24:@22140.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@22150.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@22150.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@22150.4]
  wire [7:0] RetimeWrapper_59_io_in; // @[package.scala 93:22:@22150.4]
  wire [7:0] RetimeWrapper_59_io_out; // @[package.scala 93:22:@22150.4]
  wire [7:0] x445_sum_1_io_a; // @[Math.scala 150:24:@22159.4]
  wire [7:0] x445_sum_1_io_b; // @[Math.scala 150:24:@22159.4]
  wire [7:0] x445_sum_1_io_result; // @[Math.scala 150:24:@22159.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@22169.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@22169.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@22169.4]
  wire [7:0] RetimeWrapper_60_io_in; // @[package.scala 93:22:@22169.4]
  wire [7:0] RetimeWrapper_60_io_out; // @[package.scala 93:22:@22169.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@22178.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@22178.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@22178.4]
  wire  RetimeWrapper_61_io_in; // @[package.scala 93:22:@22178.4]
  wire  RetimeWrapper_61_io_out; // @[package.scala 93:22:@22178.4]
  wire  x452_x17_1_clock; // @[Math.scala 150:24:@22215.4]
  wire  x452_x17_1_reset; // @[Math.scala 150:24:@22215.4]
  wire [7:0] x452_x17_1_io_a; // @[Math.scala 150:24:@22215.4]
  wire [7:0] x452_x17_1_io_b; // @[Math.scala 150:24:@22215.4]
  wire  x452_x17_1_io_flow; // @[Math.scala 150:24:@22215.4]
  wire [7:0] x452_x17_1_io_result; // @[Math.scala 150:24:@22215.4]
  wire  x453_x18_1_clock; // @[Math.scala 150:24:@22225.4]
  wire  x453_x18_1_reset; // @[Math.scala 150:24:@22225.4]
  wire [7:0] x453_x18_1_io_a; // @[Math.scala 150:24:@22225.4]
  wire [7:0] x453_x18_1_io_b; // @[Math.scala 150:24:@22225.4]
  wire  x453_x18_1_io_flow; // @[Math.scala 150:24:@22225.4]
  wire [7:0] x453_x18_1_io_result; // @[Math.scala 150:24:@22225.4]
  wire  x454_x17_1_clock; // @[Math.scala 150:24:@22235.4]
  wire  x454_x17_1_reset; // @[Math.scala 150:24:@22235.4]
  wire [7:0] x454_x17_1_io_a; // @[Math.scala 150:24:@22235.4]
  wire [7:0] x454_x17_1_io_b; // @[Math.scala 150:24:@22235.4]
  wire  x454_x17_1_io_flow; // @[Math.scala 150:24:@22235.4]
  wire [7:0] x454_x17_1_io_result; // @[Math.scala 150:24:@22235.4]
  wire  x455_x18_1_clock; // @[Math.scala 150:24:@22245.4]
  wire  x455_x18_1_reset; // @[Math.scala 150:24:@22245.4]
  wire [7:0] x455_x18_1_io_a; // @[Math.scala 150:24:@22245.4]
  wire [7:0] x455_x18_1_io_b; // @[Math.scala 150:24:@22245.4]
  wire  x455_x18_1_io_flow; // @[Math.scala 150:24:@22245.4]
  wire [7:0] x455_x18_1_io_result; // @[Math.scala 150:24:@22245.4]
  wire [7:0] x456_x17_1_io_a; // @[Math.scala 150:24:@22255.4]
  wire [7:0] x456_x17_1_io_b; // @[Math.scala 150:24:@22255.4]
  wire [7:0] x456_x17_1_io_result; // @[Math.scala 150:24:@22255.4]
  wire [7:0] x457_x18_1_io_a; // @[Math.scala 150:24:@22265.4]
  wire [7:0] x457_x18_1_io_b; // @[Math.scala 150:24:@22265.4]
  wire [7:0] x457_x18_1_io_result; // @[Math.scala 150:24:@22265.4]
  wire [7:0] x458_x17_1_io_a; // @[Math.scala 150:24:@22275.4]
  wire [7:0] x458_x17_1_io_b; // @[Math.scala 150:24:@22275.4]
  wire [7:0] x458_x17_1_io_result; // @[Math.scala 150:24:@22275.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@22285.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@22285.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@22285.4]
  wire [7:0] RetimeWrapper_62_io_in; // @[package.scala 93:22:@22285.4]
  wire [7:0] RetimeWrapper_62_io_out; // @[package.scala 93:22:@22285.4]
  wire [7:0] x459_sum_1_io_a; // @[Math.scala 150:24:@22294.4]
  wire [7:0] x459_sum_1_io_b; // @[Math.scala 150:24:@22294.4]
  wire [7:0] x459_sum_1_io_result; // @[Math.scala 150:24:@22294.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@22308.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@22308.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@22308.4]
  wire [7:0] RetimeWrapper_63_io_in; // @[package.scala 93:22:@22308.4]
  wire [7:0] RetimeWrapper_63_io_out; // @[package.scala 93:22:@22308.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@22318.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@22318.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@22318.4]
  wire [7:0] RetimeWrapper_64_io_in; // @[package.scala 93:22:@22318.4]
  wire [7:0] RetimeWrapper_64_io_out; // @[package.scala 93:22:@22318.4]
  wire [7:0] x461_sub_1_io_a; // @[Math.scala 191:24:@22327.4]
  wire [7:0] x461_sub_1_io_b; // @[Math.scala 191:24:@22327.4]
  wire [7:0] x461_sub_1_io_result; // @[Math.scala 191:24:@22327.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@22352.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@22352.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@22352.4]
  wire [7:0] RetimeWrapper_65_io_in; // @[package.scala 93:22:@22352.4]
  wire [7:0] RetimeWrapper_65_io_out; // @[package.scala 93:22:@22352.4]
  wire  x465_div_1_clock; // @[Math.scala 327:24:@22365.4]
  wire  x465_div_1_reset; // @[Math.scala 327:24:@22365.4]
  wire [7:0] x465_div_1_io_a; // @[Math.scala 327:24:@22365.4]
  wire  x465_div_1_io_flow; // @[Math.scala 327:24:@22365.4]
  wire [7:0] x465_div_1_io_result; // @[Math.scala 327:24:@22365.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@22375.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@22375.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@22375.4]
  wire [7:0] RetimeWrapper_66_io_in; // @[package.scala 93:22:@22375.4]
  wire [7:0] RetimeWrapper_66_io_out; // @[package.scala 93:22:@22375.4]
  wire [7:0] x466_sum_1_io_a; // @[Math.scala 150:24:@22384.4]
  wire [7:0] x466_sum_1_io_b; // @[Math.scala 150:24:@22384.4]
  wire [7:0] x466_sum_1_io_result; // @[Math.scala 150:24:@22384.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@22394.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@22394.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@22394.4]
  wire  RetimeWrapper_67_io_in; // @[package.scala 93:22:@22394.4]
  wire  RetimeWrapper_67_io_out; // @[package.scala 93:22:@22394.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@22403.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@22403.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@22403.4]
  wire [7:0] RetimeWrapper_68_io_in; // @[package.scala 93:22:@22403.4]
  wire [7:0] RetimeWrapper_68_io_out; // @[package.scala 93:22:@22403.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@22421.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@22421.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@22421.4]
  wire [15:0] RetimeWrapper_69_io_in; // @[package.scala 93:22:@22421.4]
  wire [15:0] RetimeWrapper_69_io_out; // @[package.scala 93:22:@22421.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@22430.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@22430.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@22430.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@22430.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@22430.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@22439.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@22439.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@22439.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@22439.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@22439.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@22448.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@22448.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@22448.4]
  wire  RetimeWrapper_72_io_in; // @[package.scala 93:22:@22448.4]
  wire  RetimeWrapper_72_io_out; // @[package.scala 93:22:@22448.4]
  wire  b281; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 62:18:@20576.4]
  wire  b282; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 63:18:@20577.4]
  wire  _T_206; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 68:30:@20672.4]
  wire  _T_207; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 68:37:@20673.4]
  wire  _T_211; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 70:76:@20678.4]
  wire  _T_212; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 70:62:@20679.4]
  wire  _T_214; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 70:101:@20680.4]
  wire [15:0] x551_x284_D1_0_number; // @[package.scala 96:25:@20689.4 package.scala 96:25:@20690.4]
  wire [31:0] b279_number; // @[Math.scala 712:22:@20561.4 Math.scala 713:14:@20562.4]
  wire [31:0] _T_242; // @[Math.scala 499:52:@20705.4]
  wire  x288; // @[Math.scala 499:44:@20713.4]
  wire  x289; // @[Math.scala 499:44:@20720.4]
  wire  x290; // @[Math.scala 499:44:@20727.4]
  wire [31:0] _T_289; // @[Mux.scala 19:72:@20739.4]
  wire [31:0] _T_291; // @[Mux.scala 19:72:@20740.4]
  wire [31:0] _T_293; // @[Mux.scala 19:72:@20741.4]
  wire [31:0] _T_295; // @[Mux.scala 19:72:@20743.4]
  wire [31:0] x291_number; // @[Mux.scala 19:72:@20744.4]
  wire [31:0] _T_307; // @[Math.scala 406:49:@20754.4]
  wire [31:0] _T_309; // @[Math.scala 406:56:@20756.4]
  wire [31:0] _T_310; // @[Math.scala 406:56:@20757.4]
  wire [31:0] b280_number; // @[Math.scala 712:22:@20573.4 Math.scala 713:14:@20574.4]
  wire [31:0] _T_319; // @[Math.scala 406:49:@20765.4]
  wire [31:0] _T_321; // @[Math.scala 406:56:@20767.4]
  wire [31:0] _T_322; // @[Math.scala 406:56:@20768.4]
  wire  _T_327; // @[FixedPoint.scala 50:25:@20774.4]
  wire [1:0] _T_331; // @[Bitwise.scala 72:12:@20776.4]
  wire [29:0] _T_332; // @[FixedPoint.scala 18:52:@20777.4]
  wire  _T_337; // @[FixedPoint.scala 50:25:@20783.4]
  wire [1:0] _T_341; // @[Bitwise.scala 72:12:@20785.4]
  wire [29:0] _T_342; // @[FixedPoint.scala 18:52:@20786.4]
  wire  _T_366; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 117:101:@20854.4]
  wire  _T_370; // @[package.scala 96:25:@20862.4 package.scala 96:25:@20863.4]
  wire  _T_372; // @[implicits.scala 55:10:@20864.4]
  wire  _T_373; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 117:118:@20865.4]
  wire  _T_375; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 117:205:@20867.4]
  wire  _T_376; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 117:224:@20868.4]
  wire  x555_b281_D2; // @[package.scala 96:25:@20833.4 package.scala 96:25:@20834.4]
  wire  _T_377; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 117:250:@20869.4]
  wire  x557_b282_D2; // @[package.scala 96:25:@20851.4 package.scala 96:25:@20852.4]
  wire [31:0] x303_rdcol_number; // @[Math.scala 154:22:@20886.4 Math.scala 155:14:@20887.4]
  wire [31:0] _T_394; // @[Math.scala 406:49:@20895.4]
  wire [31:0] _T_396; // @[Math.scala 406:56:@20897.4]
  wire [31:0] _T_397; // @[Math.scala 406:56:@20898.4]
  wire  _T_402; // @[FixedPoint.scala 50:25:@20904.4]
  wire [1:0] _T_406; // @[Bitwise.scala 72:12:@20906.4]
  wire [29:0] _T_407; // @[FixedPoint.scala 18:52:@20907.4]
  wire  _T_426; // @[package.scala 96:25:@20956.4 package.scala 96:25:@20957.4]
  wire  _T_428; // @[implicits.scala 55:10:@20958.4]
  wire  _T_429; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 138:118:@20959.4]
  wire  _T_431; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 138:205:@20961.4]
  wire  _T_432; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 138:224:@20962.4]
  wire  _T_433; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 138:250:@20963.4]
  wire [31:0] x561_b279_D4_number; // @[package.scala 96:25:@20977.4 package.scala 96:25:@20978.4]
  wire [31:0] _T_445; // @[Math.scala 406:49:@20984.4]
  wire [31:0] _T_447; // @[Math.scala 406:56:@20986.4]
  wire [31:0] _T_448; // @[Math.scala 406:56:@20987.4]
  wire [31:0] x543_number; // @[implicits.scala 133:21:@20988.4]
  wire  x314; // @[Math.scala 465:44:@20996.4]
  wire [31:0] x562_x303_rdcol_D4_number; // @[package.scala 96:25:@21004.4 package.scala 96:25:@21005.4]
  wire [31:0] _T_466; // @[Math.scala 465:37:@21010.4]
  wire  x315; // @[Math.scala 465:44:@21012.4]
  wire  x563_x314_D1; // @[package.scala 96:25:@21020.4 package.scala 96:25:@21021.4]
  wire  x316; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 153:24:@21024.4]
  wire [31:0] _T_483; // @[Math.scala 406:49:@21033.4]
  wire [31:0] _T_485; // @[Math.scala 406:56:@21035.4]
  wire [31:0] _T_486; // @[Math.scala 406:56:@21036.4]
  wire  _T_491; // @[FixedPoint.scala 50:25:@21042.4]
  wire [1:0] _T_495; // @[Bitwise.scala 72:12:@21044.4]
  wire [29:0] _T_496; // @[FixedPoint.scala 18:52:@21045.4]
  wire  _T_533; // @[package.scala 96:25:@21131.4 package.scala 96:25:@21132.4]
  wire  _T_535; // @[implicits.scala 55:10:@21133.4]
  wire  _T_536; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 186:194:@21134.4]
  wire  x567_x317_D1; // @[package.scala 96:25:@21092.4 package.scala 96:25:@21093.4]
  wire  _T_537; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 186:281:@21135.4]
  wire  x568_b281_D6; // @[package.scala 96:25:@21101.4 package.scala 96:25:@21102.4]
  wire  _T_538; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 186:324:@21136.4]
  wire  x569_b282_D6; // @[package.scala 96:25:@21110.4 package.scala 96:25:@21111.4]
  wire [31:0] x571_b280_D4_number; // @[package.scala 96:25:@21152.4 package.scala 96:25:@21153.4]
  wire [31:0] _T_551; // @[Math.scala 465:37:@21160.4]
  wire  x326; // @[Math.scala 465:44:@21162.4]
  wire  x327; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 196:59:@21165.4]
  wire  _T_584; // @[package.scala 96:25:@21225.4 package.scala 96:25:@21226.4]
  wire  _T_586; // @[implicits.scala 55:10:@21227.4]
  wire  _T_587; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 213:194:@21228.4]
  wire  x574_x328_D2; // @[package.scala 96:25:@21204.4 package.scala 96:25:@21205.4]
  wire  _T_588; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 213:281:@21229.4]
  wire  _T_589; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 213:289:@21230.4]
  wire [31:0] x334_rdcol_number; // @[Math.scala 154:22:@21249.4 Math.scala 155:14:@21250.4]
  wire [31:0] _T_604; // @[Math.scala 465:37:@21255.4]
  wire  x335; // @[Math.scala 465:44:@21257.4]
  wire  x336; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 221:59:@21260.4]
  wire [31:0] _T_620; // @[Math.scala 406:56:@21271.4]
  wire [31:0] _T_621; // @[Math.scala 406:56:@21272.4]
  wire  _T_626; // @[FixedPoint.scala 50:25:@21278.4]
  wire [1:0] _T_630; // @[Bitwise.scala 72:12:@21280.4]
  wire [29:0] _T_631; // @[FixedPoint.scala 18:52:@21281.4]
  wire  _T_653; // @[package.scala 96:25:@21322.4 package.scala 96:25:@21323.4]
  wire  _T_655; // @[implicits.scala 55:10:@21324.4]
  wire  _T_656; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 238:194:@21325.4]
  wire  x577_x337_D1; // @[package.scala 96:25:@21310.4 package.scala 96:25:@21311.4]
  wire  _T_657; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 238:281:@21326.4]
  wire  _T_658; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 238:289:@21327.4]
  wire [31:0] x346_rdcol_number; // @[Math.scala 154:22:@21346.4 Math.scala 155:14:@21347.4]
  wire [31:0] _T_673; // @[Math.scala 465:37:@21352.4]
  wire  x347; // @[Math.scala 465:44:@21354.4]
  wire  x348; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 246:59:@21357.4]
  wire [31:0] _T_689; // @[Math.scala 406:56:@21368.4]
  wire [31:0] _T_690; // @[Math.scala 406:56:@21369.4]
  wire  _T_695; // @[FixedPoint.scala 50:25:@21375.4]
  wire [1:0] _T_699; // @[Bitwise.scala 72:12:@21377.4]
  wire [29:0] _T_700; // @[FixedPoint.scala 18:52:@21378.4]
  wire  _T_722; // @[package.scala 96:25:@21419.4 package.scala 96:25:@21420.4]
  wire  _T_724; // @[implicits.scala 55:10:@21421.4]
  wire  _T_725; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 263:194:@21422.4]
  wire  x579_x349_D1; // @[package.scala 96:25:@21407.4 package.scala 96:25:@21408.4]
  wire  _T_726; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 263:281:@21423.4]
  wire  _T_727; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 263:289:@21424.4]
  wire [31:0] x358_rdrow_number; // @[Math.scala 195:22:@21443.4 Math.scala 196:14:@21444.4]
  wire [31:0] _T_744; // @[Math.scala 406:49:@21450.4]
  wire [31:0] _T_746; // @[Math.scala 406:56:@21452.4]
  wire [31:0] _T_747; // @[Math.scala 406:56:@21453.4]
  wire [31:0] x547_number; // @[implicits.scala 133:21:@21454.4]
  wire  x360; // @[Math.scala 465:44:@21462.4]
  wire  x361; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 273:24:@21465.4]
  wire [31:0] _T_768; // @[Math.scala 406:49:@21474.4]
  wire [31:0] _T_770; // @[Math.scala 406:56:@21476.4]
  wire [31:0] _T_771; // @[Math.scala 406:56:@21477.4]
  wire  _T_776; // @[FixedPoint.scala 50:25:@21483.4]
  wire [1:0] _T_780; // @[Bitwise.scala 72:12:@21485.4]
  wire [29:0] _T_781; // @[FixedPoint.scala 18:52:@21486.4]
  wire  _T_803; // @[package.scala 96:25:@21527.4 package.scala 96:25:@21528.4]
  wire  _T_805; // @[implicits.scala 55:10:@21529.4]
  wire  _T_806; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 290:194:@21530.4]
  wire  x580_x362_D1; // @[package.scala 96:25:@21506.4 package.scala 96:25:@21507.4]
  wire  _T_807; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 290:281:@21531.4]
  wire  _T_808; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 290:289:@21532.4]
  wire  x582_x326_D1; // @[package.scala 96:25:@21548.4 package.scala 96:25:@21549.4]
  wire  x371; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 302:59:@21552.4]
  wire  _T_840; // @[package.scala 96:25:@21596.4 package.scala 96:25:@21597.4]
  wire  _T_842; // @[implicits.scala 55:10:@21598.4]
  wire  _T_843; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 317:194:@21599.4]
  wire  x584_x372_D1; // @[package.scala 96:25:@21584.4 package.scala 96:25:@21585.4]
  wire  _T_844; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 317:281:@21600.4]
  wire  _T_845; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 317:289:@21601.4]
  wire  x378; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 321:59:@21612.4]
  wire  _T_869; // @[package.scala 96:25:@21645.4 package.scala 96:25:@21646.4]
  wire  _T_871; // @[implicits.scala 55:10:@21647.4]
  wire  _T_872; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 332:194:@21648.4]
  wire  x585_x379_D1; // @[package.scala 96:25:@21633.4 package.scala 96:25:@21634.4]
  wire  _T_873; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 332:281:@21649.4]
  wire  _T_874; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 332:289:@21650.4]
  wire  x385; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 336:59:@21661.4]
  wire  _T_898; // @[package.scala 96:25:@21694.4 package.scala 96:25:@21695.4]
  wire  _T_900; // @[implicits.scala 55:10:@21696.4]
  wire  _T_901; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 347:194:@21697.4]
  wire  x586_x386_D1; // @[package.scala 96:25:@21682.4 package.scala 96:25:@21683.4]
  wire  _T_902; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 347:281:@21698.4]
  wire  _T_903; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 347:289:@21699.4]
  wire [31:0] x392_rdrow_number; // @[Math.scala 195:22:@21718.4 Math.scala 196:14:@21719.4]
  wire [31:0] _T_920; // @[Math.scala 406:49:@21725.4]
  wire [31:0] _T_922; // @[Math.scala 406:56:@21727.4]
  wire [31:0] _T_923; // @[Math.scala 406:56:@21728.4]
  wire [31:0] x549_number; // @[implicits.scala 133:21:@21729.4]
  wire  x394; // @[Math.scala 465:44:@21737.4]
  wire  x395; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 357:24:@21740.4]
  wire [31:0] _T_944; // @[Math.scala 406:49:@21749.4]
  wire [31:0] _T_946; // @[Math.scala 406:56:@21751.4]
  wire [31:0] _T_947; // @[Math.scala 406:56:@21752.4]
  wire  _T_952; // @[FixedPoint.scala 50:25:@21758.4]
  wire [1:0] _T_956; // @[Bitwise.scala 72:12:@21760.4]
  wire [29:0] _T_957; // @[FixedPoint.scala 18:52:@21761.4]
  wire  _T_979; // @[package.scala 96:25:@21802.4 package.scala 96:25:@21803.4]
  wire  _T_981; // @[implicits.scala 55:10:@21804.4]
  wire  _T_982; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 374:194:@21805.4]
  wire  x588_x396_D1; // @[package.scala 96:25:@21790.4 package.scala 96:25:@21791.4]
  wire  _T_983; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 374:281:@21806.4]
  wire  _T_984; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 374:289:@21807.4]
  wire  x405; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 378:24:@21818.4]
  wire  _T_1008; // @[package.scala 96:25:@21851.4 package.scala 96:25:@21852.4]
  wire  _T_1010; // @[implicits.scala 55:10:@21853.4]
  wire  _T_1011; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 389:194:@21854.4]
  wire  x589_x406_D1; // @[package.scala 96:25:@21839.4 package.scala 96:25:@21840.4]
  wire  _T_1012; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 389:281:@21855.4]
  wire  _T_1013; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 389:289:@21856.4]
  wire  x412; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 393:24:@21867.4]
  wire  _T_1037; // @[package.scala 96:25:@21900.4 package.scala 96:25:@21901.4]
  wire  _T_1039; // @[implicits.scala 55:10:@21902.4]
  wire  _T_1040; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 404:194:@21903.4]
  wire  x590_x413_D1; // @[package.scala 96:25:@21888.4 package.scala 96:25:@21889.4]
  wire  _T_1041; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 404:281:@21904.4]
  wire  _T_1042; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 404:289:@21905.4]
  wire  x419; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 408:24:@21916.4]
  wire  _T_1066; // @[package.scala 96:25:@21949.4 package.scala 96:25:@21950.4]
  wire  _T_1068; // @[implicits.scala 55:10:@21951.4]
  wire  _T_1069; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 419:194:@21952.4]
  wire  x591_x420_D1; // @[package.scala 96:25:@21937.4 package.scala 96:25:@21938.4]
  wire  _T_1070; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 419:281:@21953.4]
  wire  _T_1071; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 419:289:@21954.4]
  wire [7:0] x332_rd_0_number; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 209:29:@21216.4 sm_x472_inr_Foreach_SAMPLER_BOX.scala 213:371:@21237.4]
  wire [8:0] _GEN_0; // @[Math.scala 450:32:@21968.4]
  wire [8:0] _T_1079; // @[Math.scala 450:32:@21968.4]
  wire [7:0] x369_rd_0_number; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 286:29:@21518.4 sm_x472_inr_Foreach_SAMPLER_BOX.scala 290:371:@21539.4]
  wire [8:0] _GEN_1; // @[Math.scala 450:32:@21973.4]
  wire [8:0] _T_1083; // @[Math.scala 450:32:@21973.4]
  wire [7:0] x376_rd_0_number; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 313:29:@21587.4 sm_x472_inr_Foreach_SAMPLER_BOX.scala 317:406:@21608.4]
  wire [9:0] _GEN_2; // @[Math.scala 450:32:@21978.4]
  wire [9:0] _T_1087; // @[Math.scala 450:32:@21978.4]
  wire [7:0] x383_rd_0_number; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 328:29:@21636.4 sm_x472_inr_Foreach_SAMPLER_BOX.scala 332:406:@21657.4]
  wire [8:0] _GEN_3; // @[Math.scala 450:32:@21983.4]
  wire [8:0] _T_1091; // @[Math.scala 450:32:@21983.4]
  wire [7:0] x410_rd_0_number; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 385:29:@21842.4 sm_x472_inr_Foreach_SAMPLER_BOX.scala 389:406:@21863.4]
  wire [8:0] _GEN_4; // @[Math.scala 450:32:@21988.4]
  wire [8:0] _T_1095; // @[Math.scala 450:32:@21988.4]
  wire [7:0] x438_sum_number; // @[Math.scala 154:22:@22077.4 Math.scala 155:14:@22078.4]
  wire [3:0] _T_1131; // @[FixedPoint.scala 18:52:@22083.4]
  wire [7:0] x440_sub_number; // @[Math.scala 195:22:@22110.4 Math.scala 196:14:@22111.4]
  wire  x441; // @[Math.scala 466:37:@22116.4]
  wire [7:0] x439_number; // @[package.scala 96:25:@22090.4 package.scala 96:25:@22091.4]
  wire  x597_x443_D6; // @[package.scala 96:25:@22183.4 package.scala 96:25:@22184.4]
  wire [7:0] x596_x439_D6_number; // @[package.scala 96:25:@22174.4 package.scala 96:25:@22175.4]
  wire [7:0] x445_sum_number; // @[Math.scala 154:22:@22165.4 Math.scala 155:14:@22166.4]
  wire [7:0] x446_number; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 483:24:@22187.4]
  wire [7:0] x344_rd_0_number; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 234:29:@21313.4 sm_x472_inr_Foreach_SAMPLER_BOX.scala 238:371:@21334.4]
  wire [8:0] _GEN_5; // @[Math.scala 450:32:@22191.4]
  wire [8:0] _T_1186; // @[Math.scala 450:32:@22191.4]
  wire [8:0] _GEN_6; // @[Math.scala 450:32:@22196.4]
  wire [8:0] _T_1190; // @[Math.scala 450:32:@22196.4]
  wire [9:0] _GEN_7; // @[Math.scala 450:32:@22201.4]
  wire [9:0] _T_1194; // @[Math.scala 450:32:@22201.4]
  wire [7:0] x390_rd_0_number; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 343:29:@21685.4 sm_x472_inr_Foreach_SAMPLER_BOX.scala 347:406:@21706.4]
  wire [8:0] _GEN_8; // @[Math.scala 450:32:@22206.4]
  wire [8:0] _T_1198; // @[Math.scala 450:32:@22206.4]
  wire [7:0] x417_rd_0_number; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 400:29:@21891.4 sm_x472_inr_Foreach_SAMPLER_BOX.scala 404:406:@21912.4]
  wire [8:0] _GEN_9; // @[Math.scala 450:32:@22211.4]
  wire [8:0] _T_1202; // @[Math.scala 450:32:@22211.4]
  wire [7:0] x459_sum_number; // @[Math.scala 154:22:@22300.4 Math.scala 155:14:@22301.4]
  wire [3:0] _T_1238; // @[FixedPoint.scala 18:52:@22306.4]
  wire [7:0] x461_sub_number; // @[Math.scala 195:22:@22333.4 Math.scala 196:14:@22334.4]
  wire  x462; // @[Math.scala 466:37:@22339.4]
  wire [7:0] x460_number; // @[package.scala 96:25:@22313.4 package.scala 96:25:@22314.4]
  wire  x602_x464_D6; // @[package.scala 96:25:@22399.4 package.scala 96:25:@22400.4]
  wire [7:0] x603_x460_D6_number; // @[package.scala 96:25:@22408.4 package.scala 96:25:@22409.4]
  wire [7:0] x466_sum_number; // @[Math.scala 154:22:@22390.4 Math.scala 155:14:@22391.4]
  wire [7:0] x467_number; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 545:24:@22412.4]
  wire  _T_1313; // @[package.scala 96:25:@22453.4 package.scala 96:25:@22454.4]
  wire  _T_1315; // @[implicits.scala 55:10:@22455.4]
  wire  x605_b281_D19; // @[package.scala 96:25:@22444.4 package.scala 96:25:@22445.4]
  wire  _T_1316; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 555:116:@22456.4]
  wire  x604_b282_D19; // @[package.scala 96:25:@22435.4 package.scala 96:25:@22436.4]
  wire  _T_1317; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 555:122:@22457.4]
  wire [31:0] x553_x297_sum_D1_number; // @[package.scala 96:25:@20815.4 package.scala 96:25:@20816.4]
  wire [31:0] x554_x541_D2_number; // @[package.scala 96:25:@20824.4 package.scala 96:25:@20825.4]
  wire [31:0] x556_x540_D2_number; // @[package.scala 96:25:@20842.4 package.scala 96:25:@20843.4]
  wire [31:0] x307_sum_number; // @[Math.scala 154:22:@20927.4 Math.scala 155:14:@20928.4]
  wire [31:0] x559_x542_D1_number; // @[package.scala 96:25:@20936.4 package.scala 96:25:@20937.4]
  wire [31:0] x320_sum_number; // @[Math.scala 154:22:@21074.4 Math.scala 155:14:@21075.4]
  wire [31:0] x566_x542_D5_number; // @[package.scala 96:25:@21083.4 package.scala 96:25:@21084.4]
  wire [31:0] x570_x544_D2_number; // @[package.scala 96:25:@21119.4 package.scala 96:25:@21120.4]
  wire [31:0] x573_x329_sum_D1_number; // @[package.scala 96:25:@21195.4 package.scala 96:25:@21196.4]
  wire [31:0] x575_x541_D6_number; // @[package.scala 96:25:@21213.4 package.scala 96:25:@21214.4]
  wire [31:0] x340_sum_number; // @[Math.scala 154:22:@21292.4 Math.scala 155:14:@21293.4]
  wire [31:0] x576_x545_D1_number; // @[package.scala 96:25:@21301.4 package.scala 96:25:@21302.4]
  wire [31:0] x352_sum_number; // @[Math.scala 154:22:@21389.4 Math.scala 155:14:@21390.4]
  wire [31:0] x578_x546_D1_number; // @[package.scala 96:25:@21398.4 package.scala 96:25:@21399.4]
  wire [31:0] x365_sum_number; // @[Math.scala 154:22:@21497.4 Math.scala 155:14:@21498.4]
  wire [31:0] x581_x548_D1_number; // @[package.scala 96:25:@21515.4 package.scala 96:25:@21516.4]
  wire [31:0] x373_sum_number; // @[Math.scala 154:22:@21575.4 Math.scala 155:14:@21576.4]
  wire [31:0] x380_sum_number; // @[Math.scala 154:22:@21624.4 Math.scala 155:14:@21625.4]
  wire [31:0] x387_sum_number; // @[Math.scala 154:22:@21673.4 Math.scala 155:14:@21674.4]
  wire [31:0] x399_sum_number; // @[Math.scala 154:22:@21772.4 Math.scala 155:14:@21773.4]
  wire [31:0] x587_x550_D1_number; // @[package.scala 96:25:@21781.4 package.scala 96:25:@21782.4]
  wire [31:0] x407_sum_number; // @[Math.scala 154:22:@21830.4 Math.scala 155:14:@21831.4]
  wire [31:0] x414_sum_number; // @[Math.scala 154:22:@21879.4 Math.scala 155:14:@21880.4]
  wire [31:0] x421_sum_number; // @[Math.scala 154:22:@21928.4 Math.scala 155:14:@21929.4]
  _ _ ( // @[Math.scala 709:24:@20556.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 709:24:@20568.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  x283_lb_0 x283_lb_0 ( // @[m_x283_lb_0.scala 39:17:@20578.4]
    .clock(x283_lb_0_clock),
    .reset(x283_lb_0_reset),
    .io_rPort_11_banks_1(x283_lb_0_io_rPort_11_banks_1),
    .io_rPort_11_banks_0(x283_lb_0_io_rPort_11_banks_0),
    .io_rPort_11_ofs_0(x283_lb_0_io_rPort_11_ofs_0),
    .io_rPort_11_en_0(x283_lb_0_io_rPort_11_en_0),
    .io_rPort_11_backpressure(x283_lb_0_io_rPort_11_backpressure),
    .io_rPort_11_output_0(x283_lb_0_io_rPort_11_output_0),
    .io_rPort_10_banks_1(x283_lb_0_io_rPort_10_banks_1),
    .io_rPort_10_banks_0(x283_lb_0_io_rPort_10_banks_0),
    .io_rPort_10_ofs_0(x283_lb_0_io_rPort_10_ofs_0),
    .io_rPort_10_en_0(x283_lb_0_io_rPort_10_en_0),
    .io_rPort_10_backpressure(x283_lb_0_io_rPort_10_backpressure),
    .io_rPort_10_output_0(x283_lb_0_io_rPort_10_output_0),
    .io_rPort_9_banks_1(x283_lb_0_io_rPort_9_banks_1),
    .io_rPort_9_banks_0(x283_lb_0_io_rPort_9_banks_0),
    .io_rPort_9_ofs_0(x283_lb_0_io_rPort_9_ofs_0),
    .io_rPort_9_en_0(x283_lb_0_io_rPort_9_en_0),
    .io_rPort_9_backpressure(x283_lb_0_io_rPort_9_backpressure),
    .io_rPort_9_output_0(x283_lb_0_io_rPort_9_output_0),
    .io_rPort_8_banks_1(x283_lb_0_io_rPort_8_banks_1),
    .io_rPort_8_banks_0(x283_lb_0_io_rPort_8_banks_0),
    .io_rPort_8_ofs_0(x283_lb_0_io_rPort_8_ofs_0),
    .io_rPort_8_en_0(x283_lb_0_io_rPort_8_en_0),
    .io_rPort_8_backpressure(x283_lb_0_io_rPort_8_backpressure),
    .io_rPort_8_output_0(x283_lb_0_io_rPort_8_output_0),
    .io_rPort_7_banks_1(x283_lb_0_io_rPort_7_banks_1),
    .io_rPort_7_banks_0(x283_lb_0_io_rPort_7_banks_0),
    .io_rPort_7_ofs_0(x283_lb_0_io_rPort_7_ofs_0),
    .io_rPort_7_en_0(x283_lb_0_io_rPort_7_en_0),
    .io_rPort_7_backpressure(x283_lb_0_io_rPort_7_backpressure),
    .io_rPort_7_output_0(x283_lb_0_io_rPort_7_output_0),
    .io_rPort_6_banks_1(x283_lb_0_io_rPort_6_banks_1),
    .io_rPort_6_banks_0(x283_lb_0_io_rPort_6_banks_0),
    .io_rPort_6_ofs_0(x283_lb_0_io_rPort_6_ofs_0),
    .io_rPort_6_en_0(x283_lb_0_io_rPort_6_en_0),
    .io_rPort_6_backpressure(x283_lb_0_io_rPort_6_backpressure),
    .io_rPort_6_output_0(x283_lb_0_io_rPort_6_output_0),
    .io_rPort_5_banks_1(x283_lb_0_io_rPort_5_banks_1),
    .io_rPort_5_banks_0(x283_lb_0_io_rPort_5_banks_0),
    .io_rPort_5_ofs_0(x283_lb_0_io_rPort_5_ofs_0),
    .io_rPort_5_en_0(x283_lb_0_io_rPort_5_en_0),
    .io_rPort_5_backpressure(x283_lb_0_io_rPort_5_backpressure),
    .io_rPort_5_output_0(x283_lb_0_io_rPort_5_output_0),
    .io_rPort_4_banks_1(x283_lb_0_io_rPort_4_banks_1),
    .io_rPort_4_banks_0(x283_lb_0_io_rPort_4_banks_0),
    .io_rPort_4_ofs_0(x283_lb_0_io_rPort_4_ofs_0),
    .io_rPort_4_en_0(x283_lb_0_io_rPort_4_en_0),
    .io_rPort_4_backpressure(x283_lb_0_io_rPort_4_backpressure),
    .io_rPort_4_output_0(x283_lb_0_io_rPort_4_output_0),
    .io_rPort_3_banks_1(x283_lb_0_io_rPort_3_banks_1),
    .io_rPort_3_banks_0(x283_lb_0_io_rPort_3_banks_0),
    .io_rPort_3_ofs_0(x283_lb_0_io_rPort_3_ofs_0),
    .io_rPort_3_en_0(x283_lb_0_io_rPort_3_en_0),
    .io_rPort_3_backpressure(x283_lb_0_io_rPort_3_backpressure),
    .io_rPort_3_output_0(x283_lb_0_io_rPort_3_output_0),
    .io_rPort_2_banks_1(x283_lb_0_io_rPort_2_banks_1),
    .io_rPort_2_banks_0(x283_lb_0_io_rPort_2_banks_0),
    .io_rPort_2_ofs_0(x283_lb_0_io_rPort_2_ofs_0),
    .io_rPort_2_en_0(x283_lb_0_io_rPort_2_en_0),
    .io_rPort_2_backpressure(x283_lb_0_io_rPort_2_backpressure),
    .io_rPort_2_output_0(x283_lb_0_io_rPort_2_output_0),
    .io_rPort_1_banks_1(x283_lb_0_io_rPort_1_banks_1),
    .io_rPort_1_banks_0(x283_lb_0_io_rPort_1_banks_0),
    .io_rPort_1_ofs_0(x283_lb_0_io_rPort_1_ofs_0),
    .io_rPort_1_en_0(x283_lb_0_io_rPort_1_en_0),
    .io_rPort_1_backpressure(x283_lb_0_io_rPort_1_backpressure),
    .io_rPort_1_output_0(x283_lb_0_io_rPort_1_output_0),
    .io_rPort_0_banks_1(x283_lb_0_io_rPort_0_banks_1),
    .io_rPort_0_banks_0(x283_lb_0_io_rPort_0_banks_0),
    .io_rPort_0_ofs_0(x283_lb_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x283_lb_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x283_lb_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x283_lb_0_io_rPort_0_output_0),
    .io_wPort_1_banks_1(x283_lb_0_io_wPort_1_banks_1),
    .io_wPort_1_banks_0(x283_lb_0_io_wPort_1_banks_0),
    .io_wPort_1_ofs_0(x283_lb_0_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(x283_lb_0_io_wPort_1_data_0),
    .io_wPort_1_en_0(x283_lb_0_io_wPort_1_en_0),
    .io_wPort_0_banks_1(x283_lb_0_io_wPort_0_banks_1),
    .io_wPort_0_banks_0(x283_lb_0_io_wPort_0_banks_0),
    .io_wPort_0_ofs_0(x283_lb_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x283_lb_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x283_lb_0_io_wPort_0_en_0)
  );
  RetimeWrapper_148 RetimeWrapper ( // @[package.scala 93:22:@20684.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x297_sum x297_sum_1 ( // @[Math.scala 150:24:@20791.4]
    .clock(x297_sum_1_clock),
    .reset(x297_sum_1_reset),
    .io_a(x297_sum_1_io_a),
    .io_b(x297_sum_1_io_b),
    .io_flow(x297_sum_1_io_flow),
    .io_result(x297_sum_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_1 ( // @[package.scala 93:22:@20801.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_149 RetimeWrapper_2 ( // @[package.scala 93:22:@20810.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_152 RetimeWrapper_3 ( // @[package.scala 93:22:@20819.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_4 ( // @[package.scala 93:22:@20828.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_152 RetimeWrapper_5 ( // @[package.scala 93:22:@20837.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_6 ( // @[package.scala 93:22:@20846.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_7 ( // @[package.scala 93:22:@20857.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  x297_sum x303_rdcol_1 ( // @[Math.scala 150:24:@20880.4]
    .clock(x303_rdcol_1_clock),
    .reset(x303_rdcol_1_reset),
    .io_a(x303_rdcol_1_io_a),
    .io_b(x303_rdcol_1_io_b),
    .io_flow(x303_rdcol_1_io_flow),
    .io_result(x303_rdcol_1_io_result)
  );
  RetimeWrapper_149 RetimeWrapper_8 ( // @[package.scala 93:22:@20912.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  x297_sum x307_sum_1 ( // @[Math.scala 150:24:@20921.4]
    .clock(x307_sum_1_clock),
    .reset(x307_sum_1_reset),
    .io_a(x307_sum_1_io_a),
    .io_b(x307_sum_1_io_b),
    .io_flow(x307_sum_1_io_flow),
    .io_result(x307_sum_1_io_result)
  );
  RetimeWrapper_149 RetimeWrapper_9 ( // @[package.scala 93:22:@20931.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_10 ( // @[package.scala 93:22:@20940.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_11 ( // @[package.scala 93:22:@20951.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_163 RetimeWrapper_12 ( // @[package.scala 93:22:@20972.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_163 RetimeWrapper_13 ( // @[package.scala 93:22:@20999.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper RetimeWrapper_14 ( // @[package.scala 93:22:@21015.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_149 RetimeWrapper_15 ( // @[package.scala 93:22:@21050.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_163 RetimeWrapper_16 ( // @[package.scala 93:22:@21059.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  x297_sum x320_sum_1 ( // @[Math.scala 150:24:@21068.4]
    .clock(x320_sum_1_clock),
    .reset(x320_sum_1_reset),
    .io_a(x320_sum_1_io_a),
    .io_b(x320_sum_1_io_b),
    .io_flow(x320_sum_1_io_flow),
    .io_result(x320_sum_1_io_result)
  );
  RetimeWrapper_169 RetimeWrapper_17 ( // @[package.scala 93:22:@21078.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper RetimeWrapper_18 ( // @[package.scala 93:22:@21087.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_171 RetimeWrapper_19 ( // @[package.scala 93:22:@21096.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_171 RetimeWrapper_20 ( // @[package.scala 93:22:@21105.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_152 RetimeWrapper_21 ( // @[package.scala 93:22:@21114.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_171 RetimeWrapper_22 ( // @[package.scala 93:22:@21126.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_163 RetimeWrapper_23 ( // @[package.scala 93:22:@21147.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_163 RetimeWrapper_24 ( // @[package.scala 93:22:@21171.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  x297_sum x329_sum_1 ( // @[Math.scala 150:24:@21180.4]
    .clock(x329_sum_1_clock),
    .reset(x329_sum_1_reset),
    .io_a(x329_sum_1_io_a),
    .io_b(x329_sum_1_io_b),
    .io_flow(x329_sum_1_io_flow),
    .io_result(x329_sum_1_io_result)
  );
  RetimeWrapper_149 RetimeWrapper_25 ( // @[package.scala 93:22:@21190.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_26 ( // @[package.scala 93:22:@21199.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_180 RetimeWrapper_27 ( // @[package.scala 93:22:@21208.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_171 RetimeWrapper_28 ( // @[package.scala 93:22:@21220.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  x297_sum x334_rdcol_1 ( // @[Math.scala 150:24:@21243.4]
    .clock(x334_rdcol_1_clock),
    .reset(x334_rdcol_1_reset),
    .io_a(x334_rdcol_1_io_a),
    .io_b(x334_rdcol_1_io_b),
    .io_flow(x334_rdcol_1_io_flow),
    .io_result(x334_rdcol_1_io_result)
  );
  x297_sum x340_sum_1 ( // @[Math.scala 150:24:@21286.4]
    .clock(x340_sum_1_clock),
    .reset(x340_sum_1_reset),
    .io_a(x340_sum_1_io_a),
    .io_b(x340_sum_1_io_b),
    .io_flow(x340_sum_1_io_flow),
    .io_result(x340_sum_1_io_result)
  );
  RetimeWrapper_149 RetimeWrapper_29 ( // @[package.scala 93:22:@21296.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper RetimeWrapper_30 ( // @[package.scala 93:22:@21305.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_171 RetimeWrapper_31 ( // @[package.scala 93:22:@21317.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  x297_sum x346_rdcol_1 ( // @[Math.scala 150:24:@21340.4]
    .clock(x346_rdcol_1_clock),
    .reset(x346_rdcol_1_reset),
    .io_a(x346_rdcol_1_io_a),
    .io_b(x346_rdcol_1_io_b),
    .io_flow(x346_rdcol_1_io_flow),
    .io_result(x346_rdcol_1_io_result)
  );
  x297_sum x352_sum_1 ( // @[Math.scala 150:24:@21383.4]
    .clock(x352_sum_1_clock),
    .reset(x352_sum_1_reset),
    .io_a(x352_sum_1_io_a),
    .io_b(x352_sum_1_io_b),
    .io_flow(x352_sum_1_io_flow),
    .io_result(x352_sum_1_io_result)
  );
  RetimeWrapper_149 RetimeWrapper_32 ( // @[package.scala 93:22:@21393.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper RetimeWrapper_33 ( // @[package.scala 93:22:@21402.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_171 RetimeWrapper_34 ( // @[package.scala 93:22:@21414.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  x358_rdrow x358_rdrow_1 ( // @[Math.scala 191:24:@21437.4]
    .clock(x358_rdrow_1_clock),
    .reset(x358_rdrow_1_reset),
    .io_a(x358_rdrow_1_io_a),
    .io_b(x358_rdrow_1_io_b),
    .io_flow(x358_rdrow_1_io_flow),
    .io_result(x358_rdrow_1_io_result)
  );
  x297_sum x365_sum_1 ( // @[Math.scala 150:24:@21491.4]
    .clock(x365_sum_1_clock),
    .reset(x365_sum_1_reset),
    .io_a(x365_sum_1_io_a),
    .io_b(x365_sum_1_io_b),
    .io_flow(x365_sum_1_io_flow),
    .io_result(x365_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_35 ( // @[package.scala 93:22:@21501.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_149 RetimeWrapper_36 ( // @[package.scala 93:22:@21510.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_171 RetimeWrapper_37 ( // @[package.scala 93:22:@21522.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper RetimeWrapper_38 ( // @[package.scala 93:22:@21543.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_169 RetimeWrapper_39 ( // @[package.scala 93:22:@21558.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  x297_sum x373_sum_1 ( // @[Math.scala 150:24:@21569.4]
    .clock(x373_sum_1_clock),
    .reset(x373_sum_1_reset),
    .io_a(x373_sum_1_io_a),
    .io_b(x373_sum_1_io_b),
    .io_flow(x373_sum_1_io_flow),
    .io_result(x373_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_40 ( // @[package.scala 93:22:@21579.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper_171 RetimeWrapper_41 ( // @[package.scala 93:22:@21591.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  x297_sum x380_sum_1 ( // @[Math.scala 150:24:@21618.4]
    .clock(x380_sum_1_clock),
    .reset(x380_sum_1_reset),
    .io_a(x380_sum_1_io_a),
    .io_b(x380_sum_1_io_b),
    .io_flow(x380_sum_1_io_flow),
    .io_result(x380_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_42 ( // @[package.scala 93:22:@21628.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_171 RetimeWrapper_43 ( // @[package.scala 93:22:@21640.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  x297_sum x387_sum_1 ( // @[Math.scala 150:24:@21667.4]
    .clock(x387_sum_1_clock),
    .reset(x387_sum_1_reset),
    .io_a(x387_sum_1_io_a),
    .io_b(x387_sum_1_io_b),
    .io_flow(x387_sum_1_io_flow),
    .io_result(x387_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_44 ( // @[package.scala 93:22:@21677.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_171 RetimeWrapper_45 ( // @[package.scala 93:22:@21689.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  x358_rdrow x392_rdrow_1 ( // @[Math.scala 191:24:@21712.4]
    .clock(x392_rdrow_1_clock),
    .reset(x392_rdrow_1_reset),
    .io_a(x392_rdrow_1_io_a),
    .io_b(x392_rdrow_1_io_b),
    .io_flow(x392_rdrow_1_io_flow),
    .io_result(x392_rdrow_1_io_result)
  );
  x297_sum x399_sum_1 ( // @[Math.scala 150:24:@21766.4]
    .clock(x399_sum_1_clock),
    .reset(x399_sum_1_reset),
    .io_a(x399_sum_1_io_a),
    .io_b(x399_sum_1_io_b),
    .io_flow(x399_sum_1_io_flow),
    .io_result(x399_sum_1_io_result)
  );
  RetimeWrapper_149 RetimeWrapper_46 ( // @[package.scala 93:22:@21776.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper RetimeWrapper_47 ( // @[package.scala 93:22:@21785.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_171 RetimeWrapper_48 ( // @[package.scala 93:22:@21797.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  x297_sum x407_sum_1 ( // @[Math.scala 150:24:@21824.4]
    .clock(x407_sum_1_clock),
    .reset(x407_sum_1_reset),
    .io_a(x407_sum_1_io_a),
    .io_b(x407_sum_1_io_b),
    .io_flow(x407_sum_1_io_flow),
    .io_result(x407_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_49 ( // @[package.scala 93:22:@21834.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_171 RetimeWrapper_50 ( // @[package.scala 93:22:@21846.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  x297_sum x414_sum_1 ( // @[Math.scala 150:24:@21873.4]
    .clock(x414_sum_1_clock),
    .reset(x414_sum_1_reset),
    .io_a(x414_sum_1_io_a),
    .io_b(x414_sum_1_io_b),
    .io_flow(x414_sum_1_io_flow),
    .io_result(x414_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_51 ( // @[package.scala 93:22:@21883.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_171 RetimeWrapper_52 ( // @[package.scala 93:22:@21895.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  x297_sum x421_sum_1 ( // @[Math.scala 150:24:@21922.4]
    .clock(x421_sum_1_clock),
    .reset(x421_sum_1_reset),
    .io_a(x421_sum_1_io_a),
    .io_b(x421_sum_1_io_b),
    .io_flow(x421_sum_1_io_flow),
    .io_result(x421_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_53 ( // @[package.scala 93:22:@21932.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper_171 RetimeWrapper_54 ( // @[package.scala 93:22:@21944.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  x431_x17 x431_x17_1 ( // @[Math.scala 150:24:@21992.4]
    .clock(x431_x17_1_clock),
    .reset(x431_x17_1_reset),
    .io_a(x431_x17_1_io_a),
    .io_b(x431_x17_1_io_b),
    .io_flow(x431_x17_1_io_flow),
    .io_result(x431_x17_1_io_result)
  );
  x431_x17 x432_x18_1 ( // @[Math.scala 150:24:@22002.4]
    .clock(x432_x18_1_clock),
    .reset(x432_x18_1_reset),
    .io_a(x432_x18_1_io_a),
    .io_b(x432_x18_1_io_b),
    .io_flow(x432_x18_1_io_flow),
    .io_result(x432_x18_1_io_result)
  );
  x431_x17 x433_x17_1 ( // @[Math.scala 150:24:@22012.4]
    .clock(x433_x17_1_clock),
    .reset(x433_x17_1_reset),
    .io_a(x433_x17_1_io_a),
    .io_b(x433_x17_1_io_b),
    .io_flow(x433_x17_1_io_flow),
    .io_result(x433_x17_1_io_result)
  );
  x431_x17 x434_x18_1 ( // @[Math.scala 150:24:@22022.4]
    .clock(x434_x18_1_clock),
    .reset(x434_x18_1_reset),
    .io_a(x434_x18_1_io_a),
    .io_b(x434_x18_1_io_b),
    .io_flow(x434_x18_1_io_flow),
    .io_result(x434_x18_1_io_result)
  );
  x435_x17 x435_x17_1 ( // @[Math.scala 150:24:@22032.4]
    .io_a(x435_x17_1_io_a),
    .io_b(x435_x17_1_io_b),
    .io_result(x435_x17_1_io_result)
  );
  x435_x17 x436_x18_1 ( // @[Math.scala 150:24:@22042.4]
    .io_a(x436_x18_1_io_a),
    .io_b(x436_x18_1_io_b),
    .io_result(x436_x18_1_io_result)
  );
  x435_x17 x437_x17_1 ( // @[Math.scala 150:24:@22052.4]
    .io_a(x437_x17_1_io_a),
    .io_b(x437_x17_1_io_b),
    .io_result(x437_x17_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_55 ( // @[package.scala 93:22:@22062.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  x435_x17 x438_sum_1 ( // @[Math.scala 150:24:@22071.4]
    .io_a(x438_sum_1_io_a),
    .io_b(x438_sum_1_io_b),
    .io_result(x438_sum_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_56 ( // @[package.scala 93:22:@22085.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper_228 RetimeWrapper_57 ( // @[package.scala 93:22:@22095.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  x440_sub x440_sub_1 ( // @[Math.scala 191:24:@22104.4]
    .io_a(x440_sub_1_io_a),
    .io_b(x440_sub_1_io_b),
    .io_result(x440_sub_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_58 ( // @[package.scala 93:22:@22129.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  x444_div x444_div_1 ( // @[Math.scala 327:24:@22140.4]
    .clock(x444_div_1_clock),
    .reset(x444_div_1_reset),
    .io_a(x444_div_1_io_a),
    .io_flow(x444_div_1_io_flow),
    .io_result(x444_div_1_io_result)
  );
  RetimeWrapper_231 RetimeWrapper_59 ( // @[package.scala 93:22:@22150.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  x435_x17 x445_sum_1 ( // @[Math.scala 150:24:@22159.4]
    .io_a(x445_sum_1_io_a),
    .io_b(x445_sum_1_io_b),
    .io_result(x445_sum_1_io_result)
  );
  RetimeWrapper_232 RetimeWrapper_60 ( // @[package.scala 93:22:@22169.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_171 RetimeWrapper_61 ( // @[package.scala 93:22:@22178.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  x431_x17 x452_x17_1 ( // @[Math.scala 150:24:@22215.4]
    .clock(x452_x17_1_clock),
    .reset(x452_x17_1_reset),
    .io_a(x452_x17_1_io_a),
    .io_b(x452_x17_1_io_b),
    .io_flow(x452_x17_1_io_flow),
    .io_result(x452_x17_1_io_result)
  );
  x431_x17 x453_x18_1 ( // @[Math.scala 150:24:@22225.4]
    .clock(x453_x18_1_clock),
    .reset(x453_x18_1_reset),
    .io_a(x453_x18_1_io_a),
    .io_b(x453_x18_1_io_b),
    .io_flow(x453_x18_1_io_flow),
    .io_result(x453_x18_1_io_result)
  );
  x431_x17 x454_x17_1 ( // @[Math.scala 150:24:@22235.4]
    .clock(x454_x17_1_clock),
    .reset(x454_x17_1_reset),
    .io_a(x454_x17_1_io_a),
    .io_b(x454_x17_1_io_b),
    .io_flow(x454_x17_1_io_flow),
    .io_result(x454_x17_1_io_result)
  );
  x431_x17 x455_x18_1 ( // @[Math.scala 150:24:@22245.4]
    .clock(x455_x18_1_clock),
    .reset(x455_x18_1_reset),
    .io_a(x455_x18_1_io_a),
    .io_b(x455_x18_1_io_b),
    .io_flow(x455_x18_1_io_flow),
    .io_result(x455_x18_1_io_result)
  );
  x435_x17 x456_x17_1 ( // @[Math.scala 150:24:@22255.4]
    .io_a(x456_x17_1_io_a),
    .io_b(x456_x17_1_io_b),
    .io_result(x456_x17_1_io_result)
  );
  x435_x17 x457_x18_1 ( // @[Math.scala 150:24:@22265.4]
    .io_a(x457_x18_1_io_a),
    .io_b(x457_x18_1_io_b),
    .io_result(x457_x18_1_io_result)
  );
  x435_x17 x458_x17_1 ( // @[Math.scala 150:24:@22275.4]
    .io_a(x458_x17_1_io_a),
    .io_b(x458_x17_1_io_b),
    .io_result(x458_x17_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_62 ( // @[package.scala 93:22:@22285.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  x435_x17 x459_sum_1 ( // @[Math.scala 150:24:@22294.4]
    .io_a(x459_sum_1_io_a),
    .io_b(x459_sum_1_io_b),
    .io_result(x459_sum_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_63 ( // @[package.scala 93:22:@22308.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  RetimeWrapper_228 RetimeWrapper_64 ( // @[package.scala 93:22:@22318.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  x440_sub x461_sub_1 ( // @[Math.scala 191:24:@22327.4]
    .io_a(x461_sub_1_io_a),
    .io_b(x461_sub_1_io_b),
    .io_result(x461_sub_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_65 ( // @[package.scala 93:22:@22352.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  x444_div x465_div_1 ( // @[Math.scala 327:24:@22365.4]
    .clock(x465_div_1_clock),
    .reset(x465_div_1_reset),
    .io_a(x465_div_1_io_a),
    .io_flow(x465_div_1_io_flow),
    .io_result(x465_div_1_io_result)
  );
  RetimeWrapper_231 RetimeWrapper_66 ( // @[package.scala 93:22:@22375.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  x435_x17 x466_sum_1 ( // @[Math.scala 150:24:@22384.4]
    .io_a(x466_sum_1_io_a),
    .io_b(x466_sum_1_io_b),
    .io_result(x466_sum_1_io_result)
  );
  RetimeWrapper_171 RetimeWrapper_67 ( // @[package.scala 93:22:@22394.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  RetimeWrapper_232 RetimeWrapper_68 ( // @[package.scala 93:22:@22403.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_246 RetimeWrapper_69 ( // @[package.scala 93:22:@22421.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  RetimeWrapper_16 RetimeWrapper_70 ( // @[package.scala 93:22:@22430.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_16 RetimeWrapper_71 ( // @[package.scala 93:22:@22439.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  RetimeWrapper_16 RetimeWrapper_72 ( // @[package.scala 93:22:@22448.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  assign b281 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 62:18:@20576.4]
  assign b282 = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 63:18:@20577.4]
  assign _T_206 = b281 & b282; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 68:30:@20672.4]
  assign _T_207 = _T_206 & io_sigsIn_datapathEn; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 68:37:@20673.4]
  assign _T_211 = io_in_x270_TID == 8'h0; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 70:76:@20678.4]
  assign _T_212 = _T_207 & _T_211; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 70:62:@20679.4]
  assign _T_214 = io_in_x270_TDEST == 8'h0; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 70:101:@20680.4]
  assign x551_x284_D1_0_number = RetimeWrapper_io_out; // @[package.scala 96:25:@20689.4 package.scala 96:25:@20690.4]
  assign b279_number = __io_result; // @[Math.scala 712:22:@20561.4 Math.scala 713:14:@20562.4]
  assign _T_242 = $signed(b279_number); // @[Math.scala 499:52:@20705.4]
  assign x288 = $signed(32'sh1) == $signed(_T_242); // @[Math.scala 499:44:@20713.4]
  assign x289 = $signed(32'sh2) == $signed(_T_242); // @[Math.scala 499:44:@20720.4]
  assign x290 = $signed(32'sh3) == $signed(_T_242); // @[Math.scala 499:44:@20727.4]
  assign _T_289 = x288 ? 32'h1 : 32'h0; // @[Mux.scala 19:72:@20739.4]
  assign _T_291 = x289 ? 32'h2 : 32'h0; // @[Mux.scala 19:72:@20740.4]
  assign _T_293 = x290 ? 32'h3 : 32'h0; // @[Mux.scala 19:72:@20741.4]
  assign _T_295 = _T_289 | _T_291; // @[Mux.scala 19:72:@20743.4]
  assign x291_number = _T_295 | _T_293; // @[Mux.scala 19:72:@20744.4]
  assign _T_307 = $signed(x291_number); // @[Math.scala 406:49:@20754.4]
  assign _T_309 = $signed(_T_307) & $signed(32'sh3); // @[Math.scala 406:56:@20756.4]
  assign _T_310 = $signed(_T_309); // @[Math.scala 406:56:@20757.4]
  assign b280_number = __1_io_result; // @[Math.scala 712:22:@20573.4 Math.scala 713:14:@20574.4]
  assign _T_319 = $signed(b280_number); // @[Math.scala 406:49:@20765.4]
  assign _T_321 = $signed(_T_319) & $signed(32'sh3); // @[Math.scala 406:56:@20767.4]
  assign _T_322 = $signed(_T_321); // @[Math.scala 406:56:@20768.4]
  assign _T_327 = x291_number[31]; // @[FixedPoint.scala 50:25:@20774.4]
  assign _T_331 = _T_327 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@20776.4]
  assign _T_332 = x291_number[31:2]; // @[FixedPoint.scala 18:52:@20777.4]
  assign _T_337 = b280_number[31]; // @[FixedPoint.scala 50:25:@20783.4]
  assign _T_341 = _T_337 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@20785.4]
  assign _T_342 = b280_number[31:2]; // @[FixedPoint.scala 18:52:@20786.4]
  assign _T_366 = ~ io_sigsIn_break; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 117:101:@20854.4]
  assign _T_370 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@20862.4 package.scala 96:25:@20863.4]
  assign _T_372 = io_rr ? _T_370 : 1'h0; // @[implicits.scala 55:10:@20864.4]
  assign _T_373 = _T_366 & _T_372; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 117:118:@20865.4]
  assign _T_375 = _T_373 & _T_366; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 117:205:@20867.4]
  assign _T_376 = _T_375 & io_sigsIn_backpressure; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 117:224:@20868.4]
  assign x555_b281_D2 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@20833.4 package.scala 96:25:@20834.4]
  assign _T_377 = _T_376 & x555_b281_D2; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 117:250:@20869.4]
  assign x557_b282_D2 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@20851.4 package.scala 96:25:@20852.4]
  assign x303_rdcol_number = x303_rdcol_1_io_result; // @[Math.scala 154:22:@20886.4 Math.scala 155:14:@20887.4]
  assign _T_394 = $signed(x303_rdcol_number); // @[Math.scala 406:49:@20895.4]
  assign _T_396 = $signed(_T_394) & $signed(32'sh3); // @[Math.scala 406:56:@20897.4]
  assign _T_397 = $signed(_T_396); // @[Math.scala 406:56:@20898.4]
  assign _T_402 = x303_rdcol_number[31]; // @[FixedPoint.scala 50:25:@20904.4]
  assign _T_406 = _T_402 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@20906.4]
  assign _T_407 = x303_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@20907.4]
  assign _T_426 = RetimeWrapper_11_io_out; // @[package.scala 96:25:@20956.4 package.scala 96:25:@20957.4]
  assign _T_428 = io_rr ? _T_426 : 1'h0; // @[implicits.scala 55:10:@20958.4]
  assign _T_429 = _T_366 & _T_428; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 138:118:@20959.4]
  assign _T_431 = _T_429 & _T_366; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 138:205:@20961.4]
  assign _T_432 = _T_431 & io_sigsIn_backpressure; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 138:224:@20962.4]
  assign _T_433 = _T_432 & x555_b281_D2; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 138:250:@20963.4]
  assign x561_b279_D4_number = RetimeWrapper_12_io_out; // @[package.scala 96:25:@20977.4 package.scala 96:25:@20978.4]
  assign _T_445 = $signed(x561_b279_D4_number); // @[Math.scala 406:49:@20984.4]
  assign _T_447 = $signed(_T_445) & $signed(32'sh3); // @[Math.scala 406:56:@20986.4]
  assign _T_448 = $signed(_T_447); // @[Math.scala 406:56:@20987.4]
  assign x543_number = $unsigned(_T_448); // @[implicits.scala 133:21:@20988.4]
  assign x314 = $signed(_T_445) < $signed(32'sh0); // @[Math.scala 465:44:@20996.4]
  assign x562_x303_rdcol_D4_number = RetimeWrapper_13_io_out; // @[package.scala 96:25:@21004.4 package.scala 96:25:@21005.4]
  assign _T_466 = $signed(x562_x303_rdcol_D4_number); // @[Math.scala 465:37:@21010.4]
  assign x315 = $signed(_T_466) < $signed(32'sh0); // @[Math.scala 465:44:@21012.4]
  assign x563_x314_D1 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@21020.4 package.scala 96:25:@21021.4]
  assign x316 = x563_x314_D1 | x315; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 153:24:@21024.4]
  assign _T_483 = $signed(x543_number); // @[Math.scala 406:49:@21033.4]
  assign _T_485 = $signed(_T_483) & $signed(32'sh3); // @[Math.scala 406:56:@21035.4]
  assign _T_486 = $signed(_T_485); // @[Math.scala 406:56:@21036.4]
  assign _T_491 = x543_number[31]; // @[FixedPoint.scala 50:25:@21042.4]
  assign _T_495 = _T_491 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@21044.4]
  assign _T_496 = x543_number[31:2]; // @[FixedPoint.scala 18:52:@21045.4]
  assign _T_533 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@21131.4 package.scala 96:25:@21132.4]
  assign _T_535 = io_rr ? _T_533 : 1'h0; // @[implicits.scala 55:10:@21133.4]
  assign _T_536 = _T_366 & _T_535; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 186:194:@21134.4]
  assign x567_x317_D1 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@21092.4 package.scala 96:25:@21093.4]
  assign _T_537 = _T_536 & x567_x317_D1; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 186:281:@21135.4]
  assign x568_b281_D6 = RetimeWrapper_19_io_out; // @[package.scala 96:25:@21101.4 package.scala 96:25:@21102.4]
  assign _T_538 = _T_537 & x568_b281_D6; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 186:324:@21136.4]
  assign x569_b282_D6 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@21110.4 package.scala 96:25:@21111.4]
  assign x571_b280_D4_number = RetimeWrapper_23_io_out; // @[package.scala 96:25:@21152.4 package.scala 96:25:@21153.4]
  assign _T_551 = $signed(x571_b280_D4_number); // @[Math.scala 465:37:@21160.4]
  assign x326 = $signed(_T_551) < $signed(32'sh0); // @[Math.scala 465:44:@21162.4]
  assign x327 = x314 | x326; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 196:59:@21165.4]
  assign _T_584 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@21225.4 package.scala 96:25:@21226.4]
  assign _T_586 = io_rr ? _T_584 : 1'h0; // @[implicits.scala 55:10:@21227.4]
  assign _T_587 = _T_366 & _T_586; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 213:194:@21228.4]
  assign x574_x328_D2 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@21204.4 package.scala 96:25:@21205.4]
  assign _T_588 = _T_587 & x574_x328_D2; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 213:281:@21229.4]
  assign _T_589 = _T_588 & x568_b281_D6; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 213:289:@21230.4]
  assign x334_rdcol_number = x334_rdcol_1_io_result; // @[Math.scala 154:22:@21249.4 Math.scala 155:14:@21250.4]
  assign _T_604 = $signed(x334_rdcol_number); // @[Math.scala 465:37:@21255.4]
  assign x335 = $signed(_T_604) < $signed(32'sh0); // @[Math.scala 465:44:@21257.4]
  assign x336 = x563_x314_D1 | x335; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 221:59:@21260.4]
  assign _T_620 = $signed(_T_604) & $signed(32'sh3); // @[Math.scala 406:56:@21271.4]
  assign _T_621 = $signed(_T_620); // @[Math.scala 406:56:@21272.4]
  assign _T_626 = x334_rdcol_number[31]; // @[FixedPoint.scala 50:25:@21278.4]
  assign _T_630 = _T_626 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@21280.4]
  assign _T_631 = x334_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@21281.4]
  assign _T_653 = RetimeWrapper_31_io_out; // @[package.scala 96:25:@21322.4 package.scala 96:25:@21323.4]
  assign _T_655 = io_rr ? _T_653 : 1'h0; // @[implicits.scala 55:10:@21324.4]
  assign _T_656 = _T_366 & _T_655; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 238:194:@21325.4]
  assign x577_x337_D1 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@21310.4 package.scala 96:25:@21311.4]
  assign _T_657 = _T_656 & x577_x337_D1; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 238:281:@21326.4]
  assign _T_658 = _T_657 & x568_b281_D6; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 238:289:@21327.4]
  assign x346_rdcol_number = x346_rdcol_1_io_result; // @[Math.scala 154:22:@21346.4 Math.scala 155:14:@21347.4]
  assign _T_673 = $signed(x346_rdcol_number); // @[Math.scala 465:37:@21352.4]
  assign x347 = $signed(_T_673) < $signed(32'sh0); // @[Math.scala 465:44:@21354.4]
  assign x348 = x563_x314_D1 | x347; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 246:59:@21357.4]
  assign _T_689 = $signed(_T_673) & $signed(32'sh3); // @[Math.scala 406:56:@21368.4]
  assign _T_690 = $signed(_T_689); // @[Math.scala 406:56:@21369.4]
  assign _T_695 = x346_rdcol_number[31]; // @[FixedPoint.scala 50:25:@21375.4]
  assign _T_699 = _T_695 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@21377.4]
  assign _T_700 = x346_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@21378.4]
  assign _T_722 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@21419.4 package.scala 96:25:@21420.4]
  assign _T_724 = io_rr ? _T_722 : 1'h0; // @[implicits.scala 55:10:@21421.4]
  assign _T_725 = _T_366 & _T_724; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 263:194:@21422.4]
  assign x579_x349_D1 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@21407.4 package.scala 96:25:@21408.4]
  assign _T_726 = _T_725 & x579_x349_D1; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 263:281:@21423.4]
  assign _T_727 = _T_726 & x568_b281_D6; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 263:289:@21424.4]
  assign x358_rdrow_number = x358_rdrow_1_io_result; // @[Math.scala 195:22:@21443.4 Math.scala 196:14:@21444.4]
  assign _T_744 = $signed(x358_rdrow_number); // @[Math.scala 406:49:@21450.4]
  assign _T_746 = $signed(_T_744) & $signed(32'sh3); // @[Math.scala 406:56:@21452.4]
  assign _T_747 = $signed(_T_746); // @[Math.scala 406:56:@21453.4]
  assign x547_number = $unsigned(_T_747); // @[implicits.scala 133:21:@21454.4]
  assign x360 = $signed(_T_744) < $signed(32'sh0); // @[Math.scala 465:44:@21462.4]
  assign x361 = x360 | x315; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 273:24:@21465.4]
  assign _T_768 = $signed(x547_number); // @[Math.scala 406:49:@21474.4]
  assign _T_770 = $signed(_T_768) & $signed(32'sh3); // @[Math.scala 406:56:@21476.4]
  assign _T_771 = $signed(_T_770); // @[Math.scala 406:56:@21477.4]
  assign _T_776 = x547_number[31]; // @[FixedPoint.scala 50:25:@21483.4]
  assign _T_780 = _T_776 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@21485.4]
  assign _T_781 = x547_number[31:2]; // @[FixedPoint.scala 18:52:@21486.4]
  assign _T_803 = RetimeWrapper_37_io_out; // @[package.scala 96:25:@21527.4 package.scala 96:25:@21528.4]
  assign _T_805 = io_rr ? _T_803 : 1'h0; // @[implicits.scala 55:10:@21529.4]
  assign _T_806 = _T_366 & _T_805; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 290:194:@21530.4]
  assign x580_x362_D1 = RetimeWrapper_35_io_out; // @[package.scala 96:25:@21506.4 package.scala 96:25:@21507.4]
  assign _T_807 = _T_806 & x580_x362_D1; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 290:281:@21531.4]
  assign _T_808 = _T_807 & x568_b281_D6; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 290:289:@21532.4]
  assign x582_x326_D1 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@21548.4 package.scala 96:25:@21549.4]
  assign x371 = x360 | x582_x326_D1; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 302:59:@21552.4]
  assign _T_840 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@21596.4 package.scala 96:25:@21597.4]
  assign _T_842 = io_rr ? _T_840 : 1'h0; // @[implicits.scala 55:10:@21598.4]
  assign _T_843 = _T_366 & _T_842; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 317:194:@21599.4]
  assign x584_x372_D1 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@21584.4 package.scala 96:25:@21585.4]
  assign _T_844 = _T_843 & x584_x372_D1; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 317:281:@21600.4]
  assign _T_845 = _T_844 & x568_b281_D6; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 317:289:@21601.4]
  assign x378 = x360 | x335; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 321:59:@21612.4]
  assign _T_869 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@21645.4 package.scala 96:25:@21646.4]
  assign _T_871 = io_rr ? _T_869 : 1'h0; // @[implicits.scala 55:10:@21647.4]
  assign _T_872 = _T_366 & _T_871; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 332:194:@21648.4]
  assign x585_x379_D1 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@21633.4 package.scala 96:25:@21634.4]
  assign _T_873 = _T_872 & x585_x379_D1; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 332:281:@21649.4]
  assign _T_874 = _T_873 & x568_b281_D6; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 332:289:@21650.4]
  assign x385 = x360 | x347; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 336:59:@21661.4]
  assign _T_898 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@21694.4 package.scala 96:25:@21695.4]
  assign _T_900 = io_rr ? _T_898 : 1'h0; // @[implicits.scala 55:10:@21696.4]
  assign _T_901 = _T_366 & _T_900; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 347:194:@21697.4]
  assign x586_x386_D1 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@21682.4 package.scala 96:25:@21683.4]
  assign _T_902 = _T_901 & x586_x386_D1; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 347:281:@21698.4]
  assign _T_903 = _T_902 & x568_b281_D6; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 347:289:@21699.4]
  assign x392_rdrow_number = x392_rdrow_1_io_result; // @[Math.scala 195:22:@21718.4 Math.scala 196:14:@21719.4]
  assign _T_920 = $signed(x392_rdrow_number); // @[Math.scala 406:49:@21725.4]
  assign _T_922 = $signed(_T_920) & $signed(32'sh3); // @[Math.scala 406:56:@21727.4]
  assign _T_923 = $signed(_T_922); // @[Math.scala 406:56:@21728.4]
  assign x549_number = $unsigned(_T_923); // @[implicits.scala 133:21:@21729.4]
  assign x394 = $signed(_T_920) < $signed(32'sh0); // @[Math.scala 465:44:@21737.4]
  assign x395 = x394 | x315; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 357:24:@21740.4]
  assign _T_944 = $signed(x549_number); // @[Math.scala 406:49:@21749.4]
  assign _T_946 = $signed(_T_944) & $signed(32'sh3); // @[Math.scala 406:56:@21751.4]
  assign _T_947 = $signed(_T_946); // @[Math.scala 406:56:@21752.4]
  assign _T_952 = x549_number[31]; // @[FixedPoint.scala 50:25:@21758.4]
  assign _T_956 = _T_952 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@21760.4]
  assign _T_957 = x549_number[31:2]; // @[FixedPoint.scala 18:52:@21761.4]
  assign _T_979 = RetimeWrapper_48_io_out; // @[package.scala 96:25:@21802.4 package.scala 96:25:@21803.4]
  assign _T_981 = io_rr ? _T_979 : 1'h0; // @[implicits.scala 55:10:@21804.4]
  assign _T_982 = _T_366 & _T_981; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 374:194:@21805.4]
  assign x588_x396_D1 = RetimeWrapper_47_io_out; // @[package.scala 96:25:@21790.4 package.scala 96:25:@21791.4]
  assign _T_983 = _T_982 & x588_x396_D1; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 374:281:@21806.4]
  assign _T_984 = _T_983 & x568_b281_D6; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 374:289:@21807.4]
  assign x405 = x394 | x582_x326_D1; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 378:24:@21818.4]
  assign _T_1008 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@21851.4 package.scala 96:25:@21852.4]
  assign _T_1010 = io_rr ? _T_1008 : 1'h0; // @[implicits.scala 55:10:@21853.4]
  assign _T_1011 = _T_366 & _T_1010; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 389:194:@21854.4]
  assign x589_x406_D1 = RetimeWrapper_49_io_out; // @[package.scala 96:25:@21839.4 package.scala 96:25:@21840.4]
  assign _T_1012 = _T_1011 & x589_x406_D1; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 389:281:@21855.4]
  assign _T_1013 = _T_1012 & x568_b281_D6; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 389:289:@21856.4]
  assign x412 = x394 | x335; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 393:24:@21867.4]
  assign _T_1037 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@21900.4 package.scala 96:25:@21901.4]
  assign _T_1039 = io_rr ? _T_1037 : 1'h0; // @[implicits.scala 55:10:@21902.4]
  assign _T_1040 = _T_366 & _T_1039; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 404:194:@21903.4]
  assign x590_x413_D1 = RetimeWrapper_51_io_out; // @[package.scala 96:25:@21888.4 package.scala 96:25:@21889.4]
  assign _T_1041 = _T_1040 & x590_x413_D1; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 404:281:@21904.4]
  assign _T_1042 = _T_1041 & x568_b281_D6; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 404:289:@21905.4]
  assign x419 = x394 | x347; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 408:24:@21916.4]
  assign _T_1066 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@21949.4 package.scala 96:25:@21950.4]
  assign _T_1068 = io_rr ? _T_1066 : 1'h0; // @[implicits.scala 55:10:@21951.4]
  assign _T_1069 = _T_366 & _T_1068; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 419:194:@21952.4]
  assign x591_x420_D1 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@21937.4 package.scala 96:25:@21938.4]
  assign _T_1070 = _T_1069 & x591_x420_D1; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 419:281:@21953.4]
  assign _T_1071 = _T_1070 & x568_b281_D6; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 419:289:@21954.4]
  assign x332_rd_0_number = x283_lb_0_io_rPort_10_output_0; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 209:29:@21216.4 sm_x472_inr_Foreach_SAMPLER_BOX.scala 213:371:@21237.4]
  assign _GEN_0 = {{1'd0}, x332_rd_0_number}; // @[Math.scala 450:32:@21968.4]
  assign _T_1079 = _GEN_0 << 1; // @[Math.scala 450:32:@21968.4]
  assign x369_rd_0_number = x283_lb_0_io_rPort_11_output_0; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 286:29:@21518.4 sm_x472_inr_Foreach_SAMPLER_BOX.scala 290:371:@21539.4]
  assign _GEN_1 = {{1'd0}, x369_rd_0_number}; // @[Math.scala 450:32:@21973.4]
  assign _T_1083 = _GEN_1 << 1; // @[Math.scala 450:32:@21973.4]
  assign x376_rd_0_number = x283_lb_0_io_rPort_2_output_0; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 313:29:@21587.4 sm_x472_inr_Foreach_SAMPLER_BOX.scala 317:406:@21608.4]
  assign _GEN_2 = {{2'd0}, x376_rd_0_number}; // @[Math.scala 450:32:@21978.4]
  assign _T_1087 = _GEN_2 << 2; // @[Math.scala 450:32:@21978.4]
  assign x383_rd_0_number = x283_lb_0_io_rPort_8_output_0; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 328:29:@21636.4 sm_x472_inr_Foreach_SAMPLER_BOX.scala 332:406:@21657.4]
  assign _GEN_3 = {{1'd0}, x383_rd_0_number}; // @[Math.scala 450:32:@21983.4]
  assign _T_1091 = _GEN_3 << 1; // @[Math.scala 450:32:@21983.4]
  assign x410_rd_0_number = x283_lb_0_io_rPort_9_output_0; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 385:29:@21842.4 sm_x472_inr_Foreach_SAMPLER_BOX.scala 389:406:@21863.4]
  assign _GEN_4 = {{1'd0}, x410_rd_0_number}; // @[Math.scala 450:32:@21988.4]
  assign _T_1095 = _GEN_4 << 1; // @[Math.scala 450:32:@21988.4]
  assign x438_sum_number = x438_sum_1_io_result; // @[Math.scala 154:22:@22077.4 Math.scala 155:14:@22078.4]
  assign _T_1131 = x438_sum_number[7:4]; // @[FixedPoint.scala 18:52:@22083.4]
  assign x440_sub_number = x440_sub_1_io_result; // @[Math.scala 195:22:@22110.4 Math.scala 196:14:@22111.4]
  assign x441 = 8'hf < x440_sub_number; // @[Math.scala 466:37:@22116.4]
  assign x439_number = RetimeWrapper_56_io_out; // @[package.scala 96:25:@22090.4 package.scala 96:25:@22091.4]
  assign x597_x443_D6 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@22183.4 package.scala 96:25:@22184.4]
  assign x596_x439_D6_number = RetimeWrapper_60_io_out; // @[package.scala 96:25:@22174.4 package.scala 96:25:@22175.4]
  assign x445_sum_number = x445_sum_1_io_result; // @[Math.scala 154:22:@22165.4 Math.scala 155:14:@22166.4]
  assign x446_number = x597_x443_D6 ? x596_x439_D6_number : x445_sum_number; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 483:24:@22187.4]
  assign x344_rd_0_number = x283_lb_0_io_rPort_1_output_0; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 234:29:@21313.4 sm_x472_inr_Foreach_SAMPLER_BOX.scala 238:371:@21334.4]
  assign _GEN_5 = {{1'd0}, x344_rd_0_number}; // @[Math.scala 450:32:@22191.4]
  assign _T_1186 = _GEN_5 << 1; // @[Math.scala 450:32:@22191.4]
  assign _GEN_6 = {{1'd0}, x376_rd_0_number}; // @[Math.scala 450:32:@22196.4]
  assign _T_1190 = _GEN_6 << 1; // @[Math.scala 450:32:@22196.4]
  assign _GEN_7 = {{2'd0}, x383_rd_0_number}; // @[Math.scala 450:32:@22201.4]
  assign _T_1194 = _GEN_7 << 2; // @[Math.scala 450:32:@22201.4]
  assign x390_rd_0_number = x283_lb_0_io_rPort_7_output_0; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 343:29:@21685.4 sm_x472_inr_Foreach_SAMPLER_BOX.scala 347:406:@21706.4]
  assign _GEN_8 = {{1'd0}, x390_rd_0_number}; // @[Math.scala 450:32:@22206.4]
  assign _T_1198 = _GEN_8 << 1; // @[Math.scala 450:32:@22206.4]
  assign x417_rd_0_number = x283_lb_0_io_rPort_0_output_0; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 400:29:@21891.4 sm_x472_inr_Foreach_SAMPLER_BOX.scala 404:406:@21912.4]
  assign _GEN_9 = {{1'd0}, x417_rd_0_number}; // @[Math.scala 450:32:@22211.4]
  assign _T_1202 = _GEN_9 << 1; // @[Math.scala 450:32:@22211.4]
  assign x459_sum_number = x459_sum_1_io_result; // @[Math.scala 154:22:@22300.4 Math.scala 155:14:@22301.4]
  assign _T_1238 = x459_sum_number[7:4]; // @[FixedPoint.scala 18:52:@22306.4]
  assign x461_sub_number = x461_sub_1_io_result; // @[Math.scala 195:22:@22333.4 Math.scala 196:14:@22334.4]
  assign x462 = 8'hf < x461_sub_number; // @[Math.scala 466:37:@22339.4]
  assign x460_number = RetimeWrapper_63_io_out; // @[package.scala 96:25:@22313.4 package.scala 96:25:@22314.4]
  assign x602_x464_D6 = RetimeWrapper_67_io_out; // @[package.scala 96:25:@22399.4 package.scala 96:25:@22400.4]
  assign x603_x460_D6_number = RetimeWrapper_68_io_out; // @[package.scala 96:25:@22408.4 package.scala 96:25:@22409.4]
  assign x466_sum_number = x466_sum_1_io_result; // @[Math.scala 154:22:@22390.4 Math.scala 155:14:@22391.4]
  assign x467_number = x602_x464_D6 ? x603_x460_D6_number : x466_sum_number; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 545:24:@22412.4]
  assign _T_1313 = RetimeWrapper_72_io_out; // @[package.scala 96:25:@22453.4 package.scala 96:25:@22454.4]
  assign _T_1315 = io_rr ? _T_1313 : 1'h0; // @[implicits.scala 55:10:@22455.4]
  assign x605_b281_D19 = RetimeWrapper_71_io_out; // @[package.scala 96:25:@22444.4 package.scala 96:25:@22445.4]
  assign _T_1316 = _T_1315 & x605_b281_D19; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 555:116:@22456.4]
  assign x604_b282_D19 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@22435.4 package.scala 96:25:@22436.4]
  assign _T_1317 = _T_1316 & x604_b282_D19; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 555:122:@22457.4]
  assign x553_x297_sum_D1_number = RetimeWrapper_2_io_out; // @[package.scala 96:25:@20815.4 package.scala 96:25:@20816.4]
  assign x554_x541_D2_number = RetimeWrapper_3_io_out; // @[package.scala 96:25:@20824.4 package.scala 96:25:@20825.4]
  assign x556_x540_D2_number = RetimeWrapper_5_io_out; // @[package.scala 96:25:@20842.4 package.scala 96:25:@20843.4]
  assign x307_sum_number = x307_sum_1_io_result; // @[Math.scala 154:22:@20927.4 Math.scala 155:14:@20928.4]
  assign x559_x542_D1_number = RetimeWrapper_9_io_out; // @[package.scala 96:25:@20936.4 package.scala 96:25:@20937.4]
  assign x320_sum_number = x320_sum_1_io_result; // @[Math.scala 154:22:@21074.4 Math.scala 155:14:@21075.4]
  assign x566_x542_D5_number = RetimeWrapper_17_io_out; // @[package.scala 96:25:@21083.4 package.scala 96:25:@21084.4]
  assign x570_x544_D2_number = RetimeWrapper_21_io_out; // @[package.scala 96:25:@21119.4 package.scala 96:25:@21120.4]
  assign x573_x329_sum_D1_number = RetimeWrapper_25_io_out; // @[package.scala 96:25:@21195.4 package.scala 96:25:@21196.4]
  assign x575_x541_D6_number = RetimeWrapper_27_io_out; // @[package.scala 96:25:@21213.4 package.scala 96:25:@21214.4]
  assign x340_sum_number = x340_sum_1_io_result; // @[Math.scala 154:22:@21292.4 Math.scala 155:14:@21293.4]
  assign x576_x545_D1_number = RetimeWrapper_29_io_out; // @[package.scala 96:25:@21301.4 package.scala 96:25:@21302.4]
  assign x352_sum_number = x352_sum_1_io_result; // @[Math.scala 154:22:@21389.4 Math.scala 155:14:@21390.4]
  assign x578_x546_D1_number = RetimeWrapper_32_io_out; // @[package.scala 96:25:@21398.4 package.scala 96:25:@21399.4]
  assign x365_sum_number = x365_sum_1_io_result; // @[Math.scala 154:22:@21497.4 Math.scala 155:14:@21498.4]
  assign x581_x548_D1_number = RetimeWrapper_36_io_out; // @[package.scala 96:25:@21515.4 package.scala 96:25:@21516.4]
  assign x373_sum_number = x373_sum_1_io_result; // @[Math.scala 154:22:@21575.4 Math.scala 155:14:@21576.4]
  assign x380_sum_number = x380_sum_1_io_result; // @[Math.scala 154:22:@21624.4 Math.scala 155:14:@21625.4]
  assign x387_sum_number = x387_sum_1_io_result; // @[Math.scala 154:22:@21673.4 Math.scala 155:14:@21674.4]
  assign x399_sum_number = x399_sum_1_io_result; // @[Math.scala 154:22:@21772.4 Math.scala 155:14:@21773.4]
  assign x587_x550_D1_number = RetimeWrapper_46_io_out; // @[package.scala 96:25:@21781.4 package.scala 96:25:@21782.4]
  assign x407_sum_number = x407_sum_1_io_result; // @[Math.scala 154:22:@21830.4 Math.scala 155:14:@21831.4]
  assign x414_sum_number = x414_sum_1_io_result; // @[Math.scala 154:22:@21879.4 Math.scala 155:14:@21880.4]
  assign x421_sum_number = x421_sum_1_io_result; // @[Math.scala 154:22:@21928.4 Math.scala 155:14:@21929.4]
  assign io_in_x270_TREADY = _T_212 & _T_214; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 68:22:@20674.4 sm_x472_inr_Foreach_SAMPLER_BOX.scala 70:22:@20682.4]
  assign io_in_x271_TVALID = _T_1317 & io_sigsIn_backpressure; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 555:22:@22459.4]
  assign io_in_x271_TDATA = {{240'd0}, RetimeWrapper_69_io_out}; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 556:24:@22460.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 710:17:@20559.4]
  assign __1_io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_1); // @[Math.scala 710:17:@20571.4]
  assign x283_lb_0_clock = clock; // @[:@20579.4]
  assign x283_lb_0_reset = reset; // @[:@20580.4]
  assign x283_lb_0_io_rPort_11_banks_1 = x566_x542_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@21535.4]
  assign x283_lb_0_io_rPort_11_banks_0 = x581_x548_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@21534.4]
  assign x283_lb_0_io_rPort_11_ofs_0 = x365_sum_number[0]; // @[MemInterfaceType.scala 107:54:@21536.4]
  assign x283_lb_0_io_rPort_11_en_0 = _T_808 & x569_b282_D6; // @[MemInterfaceType.scala 110:79:@21538.4]
  assign x283_lb_0_io_rPort_11_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@21537.4]
  assign x283_lb_0_io_rPort_10_banks_1 = x575_x541_D6_number[2:0]; // @[MemInterfaceType.scala 106:58:@21233.4]
  assign x283_lb_0_io_rPort_10_banks_0 = x570_x544_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@21232.4]
  assign x283_lb_0_io_rPort_10_ofs_0 = x573_x329_sum_D1_number[0]; // @[MemInterfaceType.scala 107:54:@21234.4]
  assign x283_lb_0_io_rPort_10_en_0 = _T_589 & x569_b282_D6; // @[MemInterfaceType.scala 110:79:@21236.4]
  assign x283_lb_0_io_rPort_10_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@21235.4]
  assign x283_lb_0_io_rPort_9_banks_1 = x575_x541_D6_number[2:0]; // @[MemInterfaceType.scala 106:58:@21859.4]
  assign x283_lb_0_io_rPort_9_banks_0 = x587_x550_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@21858.4]
  assign x283_lb_0_io_rPort_9_ofs_0 = x407_sum_number[0]; // @[MemInterfaceType.scala 107:54:@21860.4]
  assign x283_lb_0_io_rPort_9_en_0 = _T_1013 & x569_b282_D6; // @[MemInterfaceType.scala 110:79:@21862.4]
  assign x283_lb_0_io_rPort_9_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@21861.4]
  assign x283_lb_0_io_rPort_8_banks_1 = x576_x545_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@21653.4]
  assign x283_lb_0_io_rPort_8_banks_0 = x581_x548_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@21652.4]
  assign x283_lb_0_io_rPort_8_ofs_0 = x380_sum_number[0]; // @[MemInterfaceType.scala 107:54:@21654.4]
  assign x283_lb_0_io_rPort_8_en_0 = _T_874 & x569_b282_D6; // @[MemInterfaceType.scala 110:79:@21656.4]
  assign x283_lb_0_io_rPort_8_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@21655.4]
  assign x283_lb_0_io_rPort_7_banks_1 = x578_x546_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@21702.4]
  assign x283_lb_0_io_rPort_7_banks_0 = x581_x548_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@21701.4]
  assign x283_lb_0_io_rPort_7_ofs_0 = x387_sum_number[0]; // @[MemInterfaceType.scala 107:54:@21703.4]
  assign x283_lb_0_io_rPort_7_en_0 = _T_903 & x569_b282_D6; // @[MemInterfaceType.scala 110:79:@21705.4]
  assign x283_lb_0_io_rPort_7_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@21704.4]
  assign x283_lb_0_io_rPort_6_banks_1 = x578_x546_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@21427.4]
  assign x283_lb_0_io_rPort_6_banks_0 = x570_x544_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@21426.4]
  assign x283_lb_0_io_rPort_6_ofs_0 = x352_sum_number[0]; // @[MemInterfaceType.scala 107:54:@21428.4]
  assign x283_lb_0_io_rPort_6_en_0 = _T_727 & x569_b282_D6; // @[MemInterfaceType.scala 110:79:@21430.4]
  assign x283_lb_0_io_rPort_6_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@21429.4]
  assign x283_lb_0_io_rPort_5_banks_1 = x566_x542_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@21810.4]
  assign x283_lb_0_io_rPort_5_banks_0 = x587_x550_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@21809.4]
  assign x283_lb_0_io_rPort_5_ofs_0 = x399_sum_number[0]; // @[MemInterfaceType.scala 107:54:@21811.4]
  assign x283_lb_0_io_rPort_5_en_0 = _T_984 & x569_b282_D6; // @[MemInterfaceType.scala 110:79:@21813.4]
  assign x283_lb_0_io_rPort_5_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@21812.4]
  assign x283_lb_0_io_rPort_4_banks_1 = x566_x542_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@21139.4]
  assign x283_lb_0_io_rPort_4_banks_0 = x570_x544_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@21138.4]
  assign x283_lb_0_io_rPort_4_ofs_0 = x320_sum_number[0]; // @[MemInterfaceType.scala 107:54:@21140.4]
  assign x283_lb_0_io_rPort_4_en_0 = _T_538 & x569_b282_D6; // @[MemInterfaceType.scala 110:79:@21142.4]
  assign x283_lb_0_io_rPort_4_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@21141.4]
  assign x283_lb_0_io_rPort_3_banks_1 = x578_x546_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@21957.4]
  assign x283_lb_0_io_rPort_3_banks_0 = x587_x550_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@21956.4]
  assign x283_lb_0_io_rPort_3_ofs_0 = x421_sum_number[0]; // @[MemInterfaceType.scala 107:54:@21958.4]
  assign x283_lb_0_io_rPort_3_en_0 = _T_1071 & x569_b282_D6; // @[MemInterfaceType.scala 110:79:@21960.4]
  assign x283_lb_0_io_rPort_3_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@21959.4]
  assign x283_lb_0_io_rPort_2_banks_1 = x575_x541_D6_number[2:0]; // @[MemInterfaceType.scala 106:58:@21604.4]
  assign x283_lb_0_io_rPort_2_banks_0 = x581_x548_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@21603.4]
  assign x283_lb_0_io_rPort_2_ofs_0 = x373_sum_number[0]; // @[MemInterfaceType.scala 107:54:@21605.4]
  assign x283_lb_0_io_rPort_2_en_0 = _T_845 & x569_b282_D6; // @[MemInterfaceType.scala 110:79:@21607.4]
  assign x283_lb_0_io_rPort_2_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@21606.4]
  assign x283_lb_0_io_rPort_1_banks_1 = x576_x545_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@21330.4]
  assign x283_lb_0_io_rPort_1_banks_0 = x570_x544_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@21329.4]
  assign x283_lb_0_io_rPort_1_ofs_0 = x340_sum_number[0]; // @[MemInterfaceType.scala 107:54:@21331.4]
  assign x283_lb_0_io_rPort_1_en_0 = _T_658 & x569_b282_D6; // @[MemInterfaceType.scala 110:79:@21333.4]
  assign x283_lb_0_io_rPort_1_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@21332.4]
  assign x283_lb_0_io_rPort_0_banks_1 = x576_x545_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@21908.4]
  assign x283_lb_0_io_rPort_0_banks_0 = x587_x550_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@21907.4]
  assign x283_lb_0_io_rPort_0_ofs_0 = x414_sum_number[0]; // @[MemInterfaceType.scala 107:54:@21909.4]
  assign x283_lb_0_io_rPort_0_en_0 = _T_1042 & x569_b282_D6; // @[MemInterfaceType.scala 110:79:@21911.4]
  assign x283_lb_0_io_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@21910.4]
  assign x283_lb_0_io_wPort_1_banks_1 = x559_x542_D1_number[2:0]; // @[MemInterfaceType.scala 88:58:@20966.4]
  assign x283_lb_0_io_wPort_1_banks_0 = x556_x540_D2_number[2:0]; // @[MemInterfaceType.scala 88:58:@20965.4]
  assign x283_lb_0_io_wPort_1_ofs_0 = x307_sum_number[0]; // @[MemInterfaceType.scala 89:54:@20967.4]
  assign x283_lb_0_io_wPort_1_data_0 = RetimeWrapper_10_io_out; // @[MemInterfaceType.scala 90:56:@20968.4]
  assign x283_lb_0_io_wPort_1_en_0 = _T_433 & x557_b282_D2; // @[MemInterfaceType.scala 93:57:@20970.4]
  assign x283_lb_0_io_wPort_0_banks_1 = x554_x541_D2_number[2:0]; // @[MemInterfaceType.scala 88:58:@20872.4]
  assign x283_lb_0_io_wPort_0_banks_0 = x556_x540_D2_number[2:0]; // @[MemInterfaceType.scala 88:58:@20871.4]
  assign x283_lb_0_io_wPort_0_ofs_0 = x553_x297_sum_D1_number[0]; // @[MemInterfaceType.scala 89:54:@20873.4]
  assign x283_lb_0_io_wPort_0_data_0 = RetimeWrapper_1_io_out; // @[MemInterfaceType.scala 90:56:@20874.4]
  assign x283_lb_0_io_wPort_0_en_0 = _T_377 & x557_b282_D2; // @[MemInterfaceType.scala 93:57:@20876.4]
  assign RetimeWrapper_clock = clock; // @[:@20685.4]
  assign RetimeWrapper_reset = reset; // @[:@20686.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@20688.4]
  assign RetimeWrapper_io_in = io_in_x270_TDATA[15:0]; // @[package.scala 94:16:@20687.4]
  assign x297_sum_1_clock = clock; // @[:@20792.4]
  assign x297_sum_1_reset = reset; // @[:@20793.4]
  assign x297_sum_1_io_a = {_T_331,_T_332}; // @[Math.scala 151:17:@20794.4]
  assign x297_sum_1_io_b = {_T_341,_T_342}; // @[Math.scala 152:17:@20795.4]
  assign x297_sum_1_io_flow = io_in_x271_TREADY; // @[Math.scala 153:20:@20796.4]
  assign RetimeWrapper_1_clock = clock; // @[:@20802.4]
  assign RetimeWrapper_1_reset = reset; // @[:@20803.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@20805.4]
  assign RetimeWrapper_1_io_in = x551_x284_D1_0_number[7:0]; // @[package.scala 94:16:@20804.4]
  assign RetimeWrapper_2_clock = clock; // @[:@20811.4]
  assign RetimeWrapper_2_reset = reset; // @[:@20812.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@20814.4]
  assign RetimeWrapper_2_io_in = x297_sum_1_io_result; // @[package.scala 94:16:@20813.4]
  assign RetimeWrapper_3_clock = clock; // @[:@20820.4]
  assign RetimeWrapper_3_reset = reset; // @[:@20821.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@20823.4]
  assign RetimeWrapper_3_io_in = $unsigned(_T_322); // @[package.scala 94:16:@20822.4]
  assign RetimeWrapper_4_clock = clock; // @[:@20829.4]
  assign RetimeWrapper_4_reset = reset; // @[:@20830.4]
  assign RetimeWrapper_4_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@20832.4]
  assign RetimeWrapper_4_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@20831.4]
  assign RetimeWrapper_5_clock = clock; // @[:@20838.4]
  assign RetimeWrapper_5_reset = reset; // @[:@20839.4]
  assign RetimeWrapper_5_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@20841.4]
  assign RetimeWrapper_5_io_in = $unsigned(_T_310); // @[package.scala 94:16:@20840.4]
  assign RetimeWrapper_6_clock = clock; // @[:@20847.4]
  assign RetimeWrapper_6_reset = reset; // @[:@20848.4]
  assign RetimeWrapper_6_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@20850.4]
  assign RetimeWrapper_6_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@20849.4]
  assign RetimeWrapper_7_clock = clock; // @[:@20858.4]
  assign RetimeWrapper_7_reset = reset; // @[:@20859.4]
  assign RetimeWrapper_7_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@20861.4]
  assign RetimeWrapper_7_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@20860.4]
  assign x303_rdcol_1_clock = clock; // @[:@20881.4]
  assign x303_rdcol_1_reset = reset; // @[:@20882.4]
  assign x303_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@20883.4]
  assign x303_rdcol_1_io_b = 32'h1; // @[Math.scala 152:17:@20884.4]
  assign x303_rdcol_1_io_flow = io_in_x271_TREADY; // @[Math.scala 153:20:@20885.4]
  assign RetimeWrapper_8_clock = clock; // @[:@20913.4]
  assign RetimeWrapper_8_reset = reset; // @[:@20914.4]
  assign RetimeWrapper_8_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@20916.4]
  assign RetimeWrapper_8_io_in = {_T_331,_T_332}; // @[package.scala 94:16:@20915.4]
  assign x307_sum_1_clock = clock; // @[:@20922.4]
  assign x307_sum_1_reset = reset; // @[:@20923.4]
  assign x307_sum_1_io_a = RetimeWrapper_8_io_out; // @[Math.scala 151:17:@20924.4]
  assign x307_sum_1_io_b = {_T_406,_T_407}; // @[Math.scala 152:17:@20925.4]
  assign x307_sum_1_io_flow = io_in_x271_TREADY; // @[Math.scala 153:20:@20926.4]
  assign RetimeWrapper_9_clock = clock; // @[:@20932.4]
  assign RetimeWrapper_9_reset = reset; // @[:@20933.4]
  assign RetimeWrapper_9_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@20935.4]
  assign RetimeWrapper_9_io_in = $unsigned(_T_397); // @[package.scala 94:16:@20934.4]
  assign RetimeWrapper_10_clock = clock; // @[:@20941.4]
  assign RetimeWrapper_10_reset = reset; // @[:@20942.4]
  assign RetimeWrapper_10_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@20944.4]
  assign RetimeWrapper_10_io_in = x551_x284_D1_0_number[15:8]; // @[package.scala 94:16:@20943.4]
  assign RetimeWrapper_11_clock = clock; // @[:@20952.4]
  assign RetimeWrapper_11_reset = reset; // @[:@20953.4]
  assign RetimeWrapper_11_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@20955.4]
  assign RetimeWrapper_11_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@20954.4]
  assign RetimeWrapper_12_clock = clock; // @[:@20973.4]
  assign RetimeWrapper_12_reset = reset; // @[:@20974.4]
  assign RetimeWrapper_12_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@20976.4]
  assign RetimeWrapper_12_io_in = __io_result; // @[package.scala 94:16:@20975.4]
  assign RetimeWrapper_13_clock = clock; // @[:@21000.4]
  assign RetimeWrapper_13_reset = reset; // @[:@21001.4]
  assign RetimeWrapper_13_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21003.4]
  assign RetimeWrapper_13_io_in = x303_rdcol_1_io_result; // @[package.scala 94:16:@21002.4]
  assign RetimeWrapper_14_clock = clock; // @[:@21016.4]
  assign RetimeWrapper_14_reset = reset; // @[:@21017.4]
  assign RetimeWrapper_14_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21019.4]
  assign RetimeWrapper_14_io_in = $signed(_T_445) < $signed(32'sh0); // @[package.scala 94:16:@21018.4]
  assign RetimeWrapper_15_clock = clock; // @[:@21051.4]
  assign RetimeWrapper_15_reset = reset; // @[:@21052.4]
  assign RetimeWrapper_15_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21054.4]
  assign RetimeWrapper_15_io_in = {_T_495,_T_496}; // @[package.scala 94:16:@21053.4]
  assign RetimeWrapper_16_clock = clock; // @[:@21060.4]
  assign RetimeWrapper_16_reset = reset; // @[:@21061.4]
  assign RetimeWrapper_16_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21063.4]
  assign RetimeWrapper_16_io_in = {_T_406,_T_407}; // @[package.scala 94:16:@21062.4]
  assign x320_sum_1_clock = clock; // @[:@21069.4]
  assign x320_sum_1_reset = reset; // @[:@21070.4]
  assign x320_sum_1_io_a = RetimeWrapper_15_io_out; // @[Math.scala 151:17:@21071.4]
  assign x320_sum_1_io_b = RetimeWrapper_16_io_out; // @[Math.scala 152:17:@21072.4]
  assign x320_sum_1_io_flow = io_in_x271_TREADY; // @[Math.scala 153:20:@21073.4]
  assign RetimeWrapper_17_clock = clock; // @[:@21079.4]
  assign RetimeWrapper_17_reset = reset; // @[:@21080.4]
  assign RetimeWrapper_17_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21082.4]
  assign RetimeWrapper_17_io_in = $unsigned(_T_397); // @[package.scala 94:16:@21081.4]
  assign RetimeWrapper_18_clock = clock; // @[:@21088.4]
  assign RetimeWrapper_18_reset = reset; // @[:@21089.4]
  assign RetimeWrapper_18_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21091.4]
  assign RetimeWrapper_18_io_in = ~ x316; // @[package.scala 94:16:@21090.4]
  assign RetimeWrapper_19_clock = clock; // @[:@21097.4]
  assign RetimeWrapper_19_reset = reset; // @[:@21098.4]
  assign RetimeWrapper_19_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21100.4]
  assign RetimeWrapper_19_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@21099.4]
  assign RetimeWrapper_20_clock = clock; // @[:@21106.4]
  assign RetimeWrapper_20_reset = reset; // @[:@21107.4]
  assign RetimeWrapper_20_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21109.4]
  assign RetimeWrapper_20_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@21108.4]
  assign RetimeWrapper_21_clock = clock; // @[:@21115.4]
  assign RetimeWrapper_21_reset = reset; // @[:@21116.4]
  assign RetimeWrapper_21_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21118.4]
  assign RetimeWrapper_21_io_in = $unsigned(_T_486); // @[package.scala 94:16:@21117.4]
  assign RetimeWrapper_22_clock = clock; // @[:@21127.4]
  assign RetimeWrapper_22_reset = reset; // @[:@21128.4]
  assign RetimeWrapper_22_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21130.4]
  assign RetimeWrapper_22_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@21129.4]
  assign RetimeWrapper_23_clock = clock; // @[:@21148.4]
  assign RetimeWrapper_23_reset = reset; // @[:@21149.4]
  assign RetimeWrapper_23_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21151.4]
  assign RetimeWrapper_23_io_in = __1_io_result; // @[package.scala 94:16:@21150.4]
  assign RetimeWrapper_24_clock = clock; // @[:@21172.4]
  assign RetimeWrapper_24_reset = reset; // @[:@21173.4]
  assign RetimeWrapper_24_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21175.4]
  assign RetimeWrapper_24_io_in = {_T_341,_T_342}; // @[package.scala 94:16:@21174.4]
  assign x329_sum_1_clock = clock; // @[:@21181.4]
  assign x329_sum_1_reset = reset; // @[:@21182.4]
  assign x329_sum_1_io_a = {_T_495,_T_496}; // @[Math.scala 151:17:@21183.4]
  assign x329_sum_1_io_b = RetimeWrapper_24_io_out; // @[Math.scala 152:17:@21184.4]
  assign x329_sum_1_io_flow = io_in_x271_TREADY; // @[Math.scala 153:20:@21185.4]
  assign RetimeWrapper_25_clock = clock; // @[:@21191.4]
  assign RetimeWrapper_25_reset = reset; // @[:@21192.4]
  assign RetimeWrapper_25_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21194.4]
  assign RetimeWrapper_25_io_in = x329_sum_1_io_result; // @[package.scala 94:16:@21193.4]
  assign RetimeWrapper_26_clock = clock; // @[:@21200.4]
  assign RetimeWrapper_26_reset = reset; // @[:@21201.4]
  assign RetimeWrapper_26_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21203.4]
  assign RetimeWrapper_26_io_in = ~ x327; // @[package.scala 94:16:@21202.4]
  assign RetimeWrapper_27_clock = clock; // @[:@21209.4]
  assign RetimeWrapper_27_reset = reset; // @[:@21210.4]
  assign RetimeWrapper_27_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21212.4]
  assign RetimeWrapper_27_io_in = $unsigned(_T_322); // @[package.scala 94:16:@21211.4]
  assign RetimeWrapper_28_clock = clock; // @[:@21221.4]
  assign RetimeWrapper_28_reset = reset; // @[:@21222.4]
  assign RetimeWrapper_28_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21224.4]
  assign RetimeWrapper_28_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@21223.4]
  assign x334_rdcol_1_clock = clock; // @[:@21244.4]
  assign x334_rdcol_1_reset = reset; // @[:@21245.4]
  assign x334_rdcol_1_io_a = RetimeWrapper_23_io_out; // @[Math.scala 151:17:@21246.4]
  assign x334_rdcol_1_io_b = 32'hffffffff; // @[Math.scala 152:17:@21247.4]
  assign x334_rdcol_1_io_flow = io_in_x271_TREADY; // @[Math.scala 153:20:@21248.4]
  assign x340_sum_1_clock = clock; // @[:@21287.4]
  assign x340_sum_1_reset = reset; // @[:@21288.4]
  assign x340_sum_1_io_a = RetimeWrapper_15_io_out; // @[Math.scala 151:17:@21289.4]
  assign x340_sum_1_io_b = {_T_630,_T_631}; // @[Math.scala 152:17:@21290.4]
  assign x340_sum_1_io_flow = io_in_x271_TREADY; // @[Math.scala 153:20:@21291.4]
  assign RetimeWrapper_29_clock = clock; // @[:@21297.4]
  assign RetimeWrapper_29_reset = reset; // @[:@21298.4]
  assign RetimeWrapper_29_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21300.4]
  assign RetimeWrapper_29_io_in = $unsigned(_T_621); // @[package.scala 94:16:@21299.4]
  assign RetimeWrapper_30_clock = clock; // @[:@21306.4]
  assign RetimeWrapper_30_reset = reset; // @[:@21307.4]
  assign RetimeWrapper_30_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21309.4]
  assign RetimeWrapper_30_io_in = ~ x336; // @[package.scala 94:16:@21308.4]
  assign RetimeWrapper_31_clock = clock; // @[:@21318.4]
  assign RetimeWrapper_31_reset = reset; // @[:@21319.4]
  assign RetimeWrapper_31_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21321.4]
  assign RetimeWrapper_31_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@21320.4]
  assign x346_rdcol_1_clock = clock; // @[:@21341.4]
  assign x346_rdcol_1_reset = reset; // @[:@21342.4]
  assign x346_rdcol_1_io_a = RetimeWrapper_23_io_out; // @[Math.scala 151:17:@21343.4]
  assign x346_rdcol_1_io_b = 32'hfffffffe; // @[Math.scala 152:17:@21344.4]
  assign x346_rdcol_1_io_flow = io_in_x271_TREADY; // @[Math.scala 153:20:@21345.4]
  assign x352_sum_1_clock = clock; // @[:@21384.4]
  assign x352_sum_1_reset = reset; // @[:@21385.4]
  assign x352_sum_1_io_a = RetimeWrapper_15_io_out; // @[Math.scala 151:17:@21386.4]
  assign x352_sum_1_io_b = {_T_699,_T_700}; // @[Math.scala 152:17:@21387.4]
  assign x352_sum_1_io_flow = io_in_x271_TREADY; // @[Math.scala 153:20:@21388.4]
  assign RetimeWrapper_32_clock = clock; // @[:@21394.4]
  assign RetimeWrapper_32_reset = reset; // @[:@21395.4]
  assign RetimeWrapper_32_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21397.4]
  assign RetimeWrapper_32_io_in = $unsigned(_T_690); // @[package.scala 94:16:@21396.4]
  assign RetimeWrapper_33_clock = clock; // @[:@21403.4]
  assign RetimeWrapper_33_reset = reset; // @[:@21404.4]
  assign RetimeWrapper_33_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21406.4]
  assign RetimeWrapper_33_io_in = ~ x348; // @[package.scala 94:16:@21405.4]
  assign RetimeWrapper_34_clock = clock; // @[:@21415.4]
  assign RetimeWrapper_34_reset = reset; // @[:@21416.4]
  assign RetimeWrapper_34_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21418.4]
  assign RetimeWrapper_34_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@21417.4]
  assign x358_rdrow_1_clock = clock; // @[:@21438.4]
  assign x358_rdrow_1_reset = reset; // @[:@21439.4]
  assign x358_rdrow_1_io_a = RetimeWrapper_12_io_out; // @[Math.scala 192:17:@21440.4]
  assign x358_rdrow_1_io_b = 32'h1; // @[Math.scala 193:17:@21441.4]
  assign x358_rdrow_1_io_flow = io_in_x271_TREADY; // @[Math.scala 194:20:@21442.4]
  assign x365_sum_1_clock = clock; // @[:@21492.4]
  assign x365_sum_1_reset = reset; // @[:@21493.4]
  assign x365_sum_1_io_a = {_T_780,_T_781}; // @[Math.scala 151:17:@21494.4]
  assign x365_sum_1_io_b = RetimeWrapper_16_io_out; // @[Math.scala 152:17:@21495.4]
  assign x365_sum_1_io_flow = io_in_x271_TREADY; // @[Math.scala 153:20:@21496.4]
  assign RetimeWrapper_35_clock = clock; // @[:@21502.4]
  assign RetimeWrapper_35_reset = reset; // @[:@21503.4]
  assign RetimeWrapper_35_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21505.4]
  assign RetimeWrapper_35_io_in = ~ x361; // @[package.scala 94:16:@21504.4]
  assign RetimeWrapper_36_clock = clock; // @[:@21511.4]
  assign RetimeWrapper_36_reset = reset; // @[:@21512.4]
  assign RetimeWrapper_36_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21514.4]
  assign RetimeWrapper_36_io_in = $unsigned(_T_771); // @[package.scala 94:16:@21513.4]
  assign RetimeWrapper_37_clock = clock; // @[:@21523.4]
  assign RetimeWrapper_37_reset = reset; // @[:@21524.4]
  assign RetimeWrapper_37_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21526.4]
  assign RetimeWrapper_37_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@21525.4]
  assign RetimeWrapper_38_clock = clock; // @[:@21544.4]
  assign RetimeWrapper_38_reset = reset; // @[:@21545.4]
  assign RetimeWrapper_38_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21547.4]
  assign RetimeWrapper_38_io_in = $signed(_T_551) < $signed(32'sh0); // @[package.scala 94:16:@21546.4]
  assign RetimeWrapper_39_clock = clock; // @[:@21559.4]
  assign RetimeWrapper_39_reset = reset; // @[:@21560.4]
  assign RetimeWrapper_39_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21562.4]
  assign RetimeWrapper_39_io_in = {_T_341,_T_342}; // @[package.scala 94:16:@21561.4]
  assign x373_sum_1_clock = clock; // @[:@21570.4]
  assign x373_sum_1_reset = reset; // @[:@21571.4]
  assign x373_sum_1_io_a = {_T_780,_T_781}; // @[Math.scala 151:17:@21572.4]
  assign x373_sum_1_io_b = RetimeWrapper_39_io_out; // @[Math.scala 152:17:@21573.4]
  assign x373_sum_1_io_flow = io_in_x271_TREADY; // @[Math.scala 153:20:@21574.4]
  assign RetimeWrapper_40_clock = clock; // @[:@21580.4]
  assign RetimeWrapper_40_reset = reset; // @[:@21581.4]
  assign RetimeWrapper_40_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21583.4]
  assign RetimeWrapper_40_io_in = ~ x371; // @[package.scala 94:16:@21582.4]
  assign RetimeWrapper_41_clock = clock; // @[:@21592.4]
  assign RetimeWrapper_41_reset = reset; // @[:@21593.4]
  assign RetimeWrapper_41_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21595.4]
  assign RetimeWrapper_41_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@21594.4]
  assign x380_sum_1_clock = clock; // @[:@21619.4]
  assign x380_sum_1_reset = reset; // @[:@21620.4]
  assign x380_sum_1_io_a = {_T_780,_T_781}; // @[Math.scala 151:17:@21621.4]
  assign x380_sum_1_io_b = {_T_630,_T_631}; // @[Math.scala 152:17:@21622.4]
  assign x380_sum_1_io_flow = io_in_x271_TREADY; // @[Math.scala 153:20:@21623.4]
  assign RetimeWrapper_42_clock = clock; // @[:@21629.4]
  assign RetimeWrapper_42_reset = reset; // @[:@21630.4]
  assign RetimeWrapper_42_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21632.4]
  assign RetimeWrapper_42_io_in = ~ x378; // @[package.scala 94:16:@21631.4]
  assign RetimeWrapper_43_clock = clock; // @[:@21641.4]
  assign RetimeWrapper_43_reset = reset; // @[:@21642.4]
  assign RetimeWrapper_43_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21644.4]
  assign RetimeWrapper_43_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@21643.4]
  assign x387_sum_1_clock = clock; // @[:@21668.4]
  assign x387_sum_1_reset = reset; // @[:@21669.4]
  assign x387_sum_1_io_a = {_T_780,_T_781}; // @[Math.scala 151:17:@21670.4]
  assign x387_sum_1_io_b = {_T_699,_T_700}; // @[Math.scala 152:17:@21671.4]
  assign x387_sum_1_io_flow = io_in_x271_TREADY; // @[Math.scala 153:20:@21672.4]
  assign RetimeWrapper_44_clock = clock; // @[:@21678.4]
  assign RetimeWrapper_44_reset = reset; // @[:@21679.4]
  assign RetimeWrapper_44_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21681.4]
  assign RetimeWrapper_44_io_in = ~ x385; // @[package.scala 94:16:@21680.4]
  assign RetimeWrapper_45_clock = clock; // @[:@21690.4]
  assign RetimeWrapper_45_reset = reset; // @[:@21691.4]
  assign RetimeWrapper_45_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21693.4]
  assign RetimeWrapper_45_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@21692.4]
  assign x392_rdrow_1_clock = clock; // @[:@21713.4]
  assign x392_rdrow_1_reset = reset; // @[:@21714.4]
  assign x392_rdrow_1_io_a = RetimeWrapper_12_io_out; // @[Math.scala 192:17:@21715.4]
  assign x392_rdrow_1_io_b = 32'h2; // @[Math.scala 193:17:@21716.4]
  assign x392_rdrow_1_io_flow = io_in_x271_TREADY; // @[Math.scala 194:20:@21717.4]
  assign x399_sum_1_clock = clock; // @[:@21767.4]
  assign x399_sum_1_reset = reset; // @[:@21768.4]
  assign x399_sum_1_io_a = {_T_956,_T_957}; // @[Math.scala 151:17:@21769.4]
  assign x399_sum_1_io_b = RetimeWrapper_16_io_out; // @[Math.scala 152:17:@21770.4]
  assign x399_sum_1_io_flow = io_in_x271_TREADY; // @[Math.scala 153:20:@21771.4]
  assign RetimeWrapper_46_clock = clock; // @[:@21777.4]
  assign RetimeWrapper_46_reset = reset; // @[:@21778.4]
  assign RetimeWrapper_46_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21780.4]
  assign RetimeWrapper_46_io_in = $unsigned(_T_947); // @[package.scala 94:16:@21779.4]
  assign RetimeWrapper_47_clock = clock; // @[:@21786.4]
  assign RetimeWrapper_47_reset = reset; // @[:@21787.4]
  assign RetimeWrapper_47_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21789.4]
  assign RetimeWrapper_47_io_in = ~ x395; // @[package.scala 94:16:@21788.4]
  assign RetimeWrapper_48_clock = clock; // @[:@21798.4]
  assign RetimeWrapper_48_reset = reset; // @[:@21799.4]
  assign RetimeWrapper_48_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21801.4]
  assign RetimeWrapper_48_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@21800.4]
  assign x407_sum_1_clock = clock; // @[:@21825.4]
  assign x407_sum_1_reset = reset; // @[:@21826.4]
  assign x407_sum_1_io_a = {_T_956,_T_957}; // @[Math.scala 151:17:@21827.4]
  assign x407_sum_1_io_b = RetimeWrapper_39_io_out; // @[Math.scala 152:17:@21828.4]
  assign x407_sum_1_io_flow = io_in_x271_TREADY; // @[Math.scala 153:20:@21829.4]
  assign RetimeWrapper_49_clock = clock; // @[:@21835.4]
  assign RetimeWrapper_49_reset = reset; // @[:@21836.4]
  assign RetimeWrapper_49_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21838.4]
  assign RetimeWrapper_49_io_in = ~ x405; // @[package.scala 94:16:@21837.4]
  assign RetimeWrapper_50_clock = clock; // @[:@21847.4]
  assign RetimeWrapper_50_reset = reset; // @[:@21848.4]
  assign RetimeWrapper_50_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21850.4]
  assign RetimeWrapper_50_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@21849.4]
  assign x414_sum_1_clock = clock; // @[:@21874.4]
  assign x414_sum_1_reset = reset; // @[:@21875.4]
  assign x414_sum_1_io_a = {_T_956,_T_957}; // @[Math.scala 151:17:@21876.4]
  assign x414_sum_1_io_b = {_T_630,_T_631}; // @[Math.scala 152:17:@21877.4]
  assign x414_sum_1_io_flow = io_in_x271_TREADY; // @[Math.scala 153:20:@21878.4]
  assign RetimeWrapper_51_clock = clock; // @[:@21884.4]
  assign RetimeWrapper_51_reset = reset; // @[:@21885.4]
  assign RetimeWrapper_51_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21887.4]
  assign RetimeWrapper_51_io_in = ~ x412; // @[package.scala 94:16:@21886.4]
  assign RetimeWrapper_52_clock = clock; // @[:@21896.4]
  assign RetimeWrapper_52_reset = reset; // @[:@21897.4]
  assign RetimeWrapper_52_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21899.4]
  assign RetimeWrapper_52_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@21898.4]
  assign x421_sum_1_clock = clock; // @[:@21923.4]
  assign x421_sum_1_reset = reset; // @[:@21924.4]
  assign x421_sum_1_io_a = {_T_956,_T_957}; // @[Math.scala 151:17:@21925.4]
  assign x421_sum_1_io_b = {_T_699,_T_700}; // @[Math.scala 152:17:@21926.4]
  assign x421_sum_1_io_flow = io_in_x271_TREADY; // @[Math.scala 153:20:@21927.4]
  assign RetimeWrapper_53_clock = clock; // @[:@21933.4]
  assign RetimeWrapper_53_reset = reset; // @[:@21934.4]
  assign RetimeWrapper_53_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21936.4]
  assign RetimeWrapper_53_io_in = ~ x419; // @[package.scala 94:16:@21935.4]
  assign RetimeWrapper_54_clock = clock; // @[:@21945.4]
  assign RetimeWrapper_54_reset = reset; // @[:@21946.4]
  assign RetimeWrapper_54_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@21948.4]
  assign RetimeWrapper_54_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@21947.4]
  assign x431_x17_1_clock = clock; // @[:@21993.4]
  assign x431_x17_1_reset = reset; // @[:@21994.4]
  assign x431_x17_1_io_a = x283_lb_0_io_rPort_4_output_0; // @[Math.scala 151:17:@21995.4]
  assign x431_x17_1_io_b = _T_1079[7:0]; // @[Math.scala 152:17:@21996.4]
  assign x431_x17_1_io_flow = io_in_x271_TREADY; // @[Math.scala 153:20:@21997.4]
  assign x432_x18_1_clock = clock; // @[:@22003.4]
  assign x432_x18_1_reset = reset; // @[:@22004.4]
  assign x432_x18_1_io_a = x283_lb_0_io_rPort_1_output_0; // @[Math.scala 151:17:@22005.4]
  assign x432_x18_1_io_b = _T_1083[7:0]; // @[Math.scala 152:17:@22006.4]
  assign x432_x18_1_io_flow = io_in_x271_TREADY; // @[Math.scala 153:20:@22007.4]
  assign x433_x17_1_clock = clock; // @[:@22013.4]
  assign x433_x17_1_reset = reset; // @[:@22014.4]
  assign x433_x17_1_io_a = _T_1087[7:0]; // @[Math.scala 151:17:@22015.4]
  assign x433_x17_1_io_b = _T_1091[7:0]; // @[Math.scala 152:17:@22016.4]
  assign x433_x17_1_io_flow = io_in_x271_TREADY; // @[Math.scala 153:20:@22017.4]
  assign x434_x18_1_clock = clock; // @[:@22023.4]
  assign x434_x18_1_reset = reset; // @[:@22024.4]
  assign x434_x18_1_io_a = x283_lb_0_io_rPort_5_output_0; // @[Math.scala 151:17:@22025.4]
  assign x434_x18_1_io_b = _T_1095[7:0]; // @[Math.scala 152:17:@22026.4]
  assign x434_x18_1_io_flow = io_in_x271_TREADY; // @[Math.scala 153:20:@22027.4]
  assign x435_x17_1_io_a = x431_x17_1_io_result; // @[Math.scala 151:17:@22035.4]
  assign x435_x17_1_io_b = x432_x18_1_io_result; // @[Math.scala 152:17:@22036.4]
  assign x436_x18_1_io_a = x433_x17_1_io_result; // @[Math.scala 151:17:@22045.4]
  assign x436_x18_1_io_b = x434_x18_1_io_result; // @[Math.scala 152:17:@22046.4]
  assign x437_x17_1_io_a = x435_x17_1_io_result; // @[Math.scala 151:17:@22055.4]
  assign x437_x17_1_io_b = x436_x18_1_io_result; // @[Math.scala 152:17:@22056.4]
  assign RetimeWrapper_55_clock = clock; // @[:@22063.4]
  assign RetimeWrapper_55_reset = reset; // @[:@22064.4]
  assign RetimeWrapper_55_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22066.4]
  assign RetimeWrapper_55_io_in = x283_lb_0_io_rPort_0_output_0; // @[package.scala 94:16:@22065.4]
  assign x438_sum_1_io_a = x437_x17_1_io_result; // @[Math.scala 151:17:@22074.4]
  assign x438_sum_1_io_b = RetimeWrapper_55_io_out; // @[Math.scala 152:17:@22075.4]
  assign RetimeWrapper_56_clock = clock; // @[:@22086.4]
  assign RetimeWrapper_56_reset = reset; // @[:@22087.4]
  assign RetimeWrapper_56_io_flow = io_in_x271_TREADY; // @[package.scala 95:18:@22089.4]
  assign RetimeWrapper_56_io_in = {4'h0,_T_1131}; // @[package.scala 94:16:@22088.4]
  assign RetimeWrapper_57_clock = clock; // @[:@22096.4]
  assign RetimeWrapper_57_reset = reset; // @[:@22097.4]
  assign RetimeWrapper_57_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22099.4]
  assign RetimeWrapper_57_io_in = x283_lb_0_io_rPort_4_output_0; // @[package.scala 94:16:@22098.4]
  assign x440_sub_1_io_a = RetimeWrapper_57_io_out; // @[Math.scala 192:17:@22107.4]
  assign x440_sub_1_io_b = RetimeWrapper_56_io_out; // @[Math.scala 193:17:@22108.4]
  assign RetimeWrapper_58_clock = clock; // @[:@22130.4]
  assign RetimeWrapper_58_reset = reset; // @[:@22131.4]
  assign RetimeWrapper_58_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22133.4]
  assign RetimeWrapper_58_io_in = x441 ? x440_sub_number : 8'h0; // @[package.scala 94:16:@22132.4]
  assign x444_div_1_clock = clock; // @[:@22141.4]
  assign x444_div_1_reset = reset; // @[:@22142.4]
  assign x444_div_1_io_a = RetimeWrapper_58_io_out; // @[Math.scala 328:17:@22143.4]
  assign x444_div_1_io_flow = io_in_x271_TREADY; // @[Math.scala 330:20:@22145.4]
  assign RetimeWrapper_59_clock = clock; // @[:@22151.4]
  assign RetimeWrapper_59_reset = reset; // @[:@22152.4]
  assign RetimeWrapper_59_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22154.4]
  assign RetimeWrapper_59_io_in = x283_lb_0_io_rPort_4_output_0; // @[package.scala 94:16:@22153.4]
  assign x445_sum_1_io_a = RetimeWrapper_59_io_out; // @[Math.scala 151:17:@22162.4]
  assign x445_sum_1_io_b = x444_div_1_io_result; // @[Math.scala 152:17:@22163.4]
  assign RetimeWrapper_60_clock = clock; // @[:@22170.4]
  assign RetimeWrapper_60_reset = reset; // @[:@22171.4]
  assign RetimeWrapper_60_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22173.4]
  assign RetimeWrapper_60_io_in = RetimeWrapper_56_io_out; // @[package.scala 94:16:@22172.4]
  assign RetimeWrapper_61_clock = clock; // @[:@22179.4]
  assign RetimeWrapper_61_reset = reset; // @[:@22180.4]
  assign RetimeWrapper_61_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22182.4]
  assign RetimeWrapper_61_io_in = x439_number == 8'h0; // @[package.scala 94:16:@22181.4]
  assign x452_x17_1_clock = clock; // @[:@22216.4]
  assign x452_x17_1_reset = reset; // @[:@22217.4]
  assign x452_x17_1_io_a = x283_lb_0_io_rPort_10_output_0; // @[Math.scala 151:17:@22218.4]
  assign x452_x17_1_io_b = _T_1186[7:0]; // @[Math.scala 152:17:@22219.4]
  assign x452_x17_1_io_flow = io_in_x271_TREADY; // @[Math.scala 153:20:@22220.4]
  assign x453_x18_1_clock = clock; // @[:@22226.4]
  assign x453_x18_1_reset = reset; // @[:@22227.4]
  assign x453_x18_1_io_a = x283_lb_0_io_rPort_6_output_0; // @[Math.scala 151:17:@22228.4]
  assign x453_x18_1_io_b = _T_1190[7:0]; // @[Math.scala 152:17:@22229.4]
  assign x453_x18_1_io_flow = io_in_x271_TREADY; // @[Math.scala 153:20:@22230.4]
  assign x454_x17_1_clock = clock; // @[:@22236.4]
  assign x454_x17_1_reset = reset; // @[:@22237.4]
  assign x454_x17_1_io_a = _T_1194[7:0]; // @[Math.scala 151:17:@22238.4]
  assign x454_x17_1_io_b = _T_1198[7:0]; // @[Math.scala 152:17:@22239.4]
  assign x454_x17_1_io_flow = io_in_x271_TREADY; // @[Math.scala 153:20:@22240.4]
  assign x455_x18_1_clock = clock; // @[:@22246.4]
  assign x455_x18_1_reset = reset; // @[:@22247.4]
  assign x455_x18_1_io_a = x283_lb_0_io_rPort_9_output_0; // @[Math.scala 151:17:@22248.4]
  assign x455_x18_1_io_b = _T_1202[7:0]; // @[Math.scala 152:17:@22249.4]
  assign x455_x18_1_io_flow = io_in_x271_TREADY; // @[Math.scala 153:20:@22250.4]
  assign x456_x17_1_io_a = x452_x17_1_io_result; // @[Math.scala 151:17:@22258.4]
  assign x456_x17_1_io_b = x453_x18_1_io_result; // @[Math.scala 152:17:@22259.4]
  assign x457_x18_1_io_a = x454_x17_1_io_result; // @[Math.scala 151:17:@22268.4]
  assign x457_x18_1_io_b = x455_x18_1_io_result; // @[Math.scala 152:17:@22269.4]
  assign x458_x17_1_io_a = x456_x17_1_io_result; // @[Math.scala 151:17:@22278.4]
  assign x458_x17_1_io_b = x457_x18_1_io_result; // @[Math.scala 152:17:@22279.4]
  assign RetimeWrapper_62_clock = clock; // @[:@22286.4]
  assign RetimeWrapper_62_reset = reset; // @[:@22287.4]
  assign RetimeWrapper_62_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22289.4]
  assign RetimeWrapper_62_io_in = x283_lb_0_io_rPort_3_output_0; // @[package.scala 94:16:@22288.4]
  assign x459_sum_1_io_a = x458_x17_1_io_result; // @[Math.scala 151:17:@22297.4]
  assign x459_sum_1_io_b = RetimeWrapper_62_io_out; // @[Math.scala 152:17:@22298.4]
  assign RetimeWrapper_63_clock = clock; // @[:@22309.4]
  assign RetimeWrapper_63_reset = reset; // @[:@22310.4]
  assign RetimeWrapper_63_io_flow = io_in_x271_TREADY; // @[package.scala 95:18:@22312.4]
  assign RetimeWrapper_63_io_in = {4'h0,_T_1238}; // @[package.scala 94:16:@22311.4]
  assign RetimeWrapper_64_clock = clock; // @[:@22319.4]
  assign RetimeWrapper_64_reset = reset; // @[:@22320.4]
  assign RetimeWrapper_64_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22322.4]
  assign RetimeWrapper_64_io_in = x283_lb_0_io_rPort_10_output_0; // @[package.scala 94:16:@22321.4]
  assign x461_sub_1_io_a = RetimeWrapper_64_io_out; // @[Math.scala 192:17:@22330.4]
  assign x461_sub_1_io_b = RetimeWrapper_63_io_out; // @[Math.scala 193:17:@22331.4]
  assign RetimeWrapper_65_clock = clock; // @[:@22353.4]
  assign RetimeWrapper_65_reset = reset; // @[:@22354.4]
  assign RetimeWrapper_65_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22356.4]
  assign RetimeWrapper_65_io_in = x462 ? x461_sub_number : 8'h0; // @[package.scala 94:16:@22355.4]
  assign x465_div_1_clock = clock; // @[:@22366.4]
  assign x465_div_1_reset = reset; // @[:@22367.4]
  assign x465_div_1_io_a = RetimeWrapper_65_io_out; // @[Math.scala 328:17:@22368.4]
  assign x465_div_1_io_flow = io_in_x271_TREADY; // @[Math.scala 330:20:@22370.4]
  assign RetimeWrapper_66_clock = clock; // @[:@22376.4]
  assign RetimeWrapper_66_reset = reset; // @[:@22377.4]
  assign RetimeWrapper_66_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22379.4]
  assign RetimeWrapper_66_io_in = x283_lb_0_io_rPort_10_output_0; // @[package.scala 94:16:@22378.4]
  assign x466_sum_1_io_a = RetimeWrapper_66_io_out; // @[Math.scala 151:17:@22387.4]
  assign x466_sum_1_io_b = x465_div_1_io_result; // @[Math.scala 152:17:@22388.4]
  assign RetimeWrapper_67_clock = clock; // @[:@22395.4]
  assign RetimeWrapper_67_reset = reset; // @[:@22396.4]
  assign RetimeWrapper_67_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22398.4]
  assign RetimeWrapper_67_io_in = x460_number == 8'h0; // @[package.scala 94:16:@22397.4]
  assign RetimeWrapper_68_clock = clock; // @[:@22404.4]
  assign RetimeWrapper_68_reset = reset; // @[:@22405.4]
  assign RetimeWrapper_68_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22407.4]
  assign RetimeWrapper_68_io_in = RetimeWrapper_63_io_out; // @[package.scala 94:16:@22406.4]
  assign RetimeWrapper_69_clock = clock; // @[:@22422.4]
  assign RetimeWrapper_69_reset = reset; // @[:@22423.4]
  assign RetimeWrapper_69_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22425.4]
  assign RetimeWrapper_69_io_in = {x446_number,x467_number}; // @[package.scala 94:16:@22424.4]
  assign RetimeWrapper_70_clock = clock; // @[:@22431.4]
  assign RetimeWrapper_70_reset = reset; // @[:@22432.4]
  assign RetimeWrapper_70_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22434.4]
  assign RetimeWrapper_70_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@22433.4]
  assign RetimeWrapper_71_clock = clock; // @[:@22440.4]
  assign RetimeWrapper_71_reset = reset; // @[:@22441.4]
  assign RetimeWrapper_71_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22443.4]
  assign RetimeWrapper_71_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@22442.4]
  assign RetimeWrapper_72_clock = clock; // @[:@22449.4]
  assign RetimeWrapper_72_reset = reset; // @[:@22450.4]
  assign RetimeWrapper_72_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@22452.4]
  assign RetimeWrapper_72_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@22451.4]
endmodule
module x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1( // @[:@22470.2]
  input          clock, // @[:@22471.4]
  input          reset, // @[:@22472.4]
  input          io_in_x270_TVALID, // @[:@22473.4]
  output         io_in_x270_TREADY, // @[:@22473.4]
  input  [255:0] io_in_x270_TDATA, // @[:@22473.4]
  input  [7:0]   io_in_x270_TID, // @[:@22473.4]
  input  [7:0]   io_in_x270_TDEST, // @[:@22473.4]
  output         io_in_x271_TVALID, // @[:@22473.4]
  input          io_in_x271_TREADY, // @[:@22473.4]
  output [255:0] io_in_x271_TDATA, // @[:@22473.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@22473.4]
  input          io_sigsIn_smChildAcks_0, // @[:@22473.4]
  output         io_sigsOut_smDoneIn_0, // @[:@22473.4]
  output         io_sigsOut_smCtrCopyDone_0, // @[:@22473.4]
  input          io_rr // @[:@22473.4]
);
  wire  x278_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@22483.4]
  wire  x278_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@22483.4]
  wire  x278_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@22483.4]
  wire  x278_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@22483.4]
  wire [31:0] x278_ctrchain_io_output_counts_1; // @[SpatialBlocks.scala 37:22:@22483.4]
  wire [31:0] x278_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@22483.4]
  wire  x278_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@22483.4]
  wire  x278_ctrchain_io_output_oobs_1; // @[SpatialBlocks.scala 37:22:@22483.4]
  wire  x278_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@22483.4]
  wire  x472_inr_Foreach_SAMPLER_BOX_sm_clock; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 32:18:@22542.4]
  wire  x472_inr_Foreach_SAMPLER_BOX_sm_reset; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 32:18:@22542.4]
  wire  x472_inr_Foreach_SAMPLER_BOX_sm_io_enable; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 32:18:@22542.4]
  wire  x472_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 32:18:@22542.4]
  wire  x472_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 32:18:@22542.4]
  wire  x472_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 32:18:@22542.4]
  wire  x472_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 32:18:@22542.4]
  wire  x472_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 32:18:@22542.4]
  wire  x472_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 32:18:@22542.4]
  wire  x472_inr_Foreach_SAMPLER_BOX_sm_io_parentAck; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 32:18:@22542.4]
  wire  x472_inr_Foreach_SAMPLER_BOX_sm_io_backpressure; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 32:18:@22542.4]
  wire  x472_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 32:18:@22542.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@22570.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@22570.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@22570.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@22570.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@22570.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@22612.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@22612.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@22612.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@22612.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@22612.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@22620.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@22620.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@22620.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@22620.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@22620.4]
  wire  x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_clock; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 568:24:@22652.4]
  wire  x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_reset; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 568:24:@22652.4]
  wire  x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x270_TREADY; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 568:24:@22652.4]
  wire [255:0] x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x270_TDATA; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 568:24:@22652.4]
  wire [7:0] x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x270_TID; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 568:24:@22652.4]
  wire [7:0] x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x270_TDEST; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 568:24:@22652.4]
  wire  x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x271_TVALID; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 568:24:@22652.4]
  wire  x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x271_TREADY; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 568:24:@22652.4]
  wire [255:0] x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x271_TDATA; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 568:24:@22652.4]
  wire  x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 568:24:@22652.4]
  wire  x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 568:24:@22652.4]
  wire  x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 568:24:@22652.4]
  wire [31:0] x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 568:24:@22652.4]
  wire [31:0] x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 568:24:@22652.4]
  wire  x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 568:24:@22652.4]
  wire  x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 568:24:@22652.4]
  wire  x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_rr; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 568:24:@22652.4]
  wire  _T_239; // @[package.scala 96:25:@22575.4 package.scala 96:25:@22576.4]
  wire  x472_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[sm_x473_outr_UnitPipe.scala 68:66:@22581.4]
  wire  _T_252; // @[package.scala 96:25:@22617.4 package.scala 96:25:@22618.4]
  wire  _T_258; // @[package.scala 96:25:@22625.4 package.scala 96:25:@22626.4]
  wire  _T_261; // @[SpatialBlocks.scala 110:93:@22628.4]
  wire  x472_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn; // @[SpatialBlocks.scala 110:90:@22629.4]
  wire  _T_263; // @[SpatialBlocks.scala 128:36:@22637.4]
  wire  _T_264; // @[SpatialBlocks.scala 128:78:@22638.4]
  wire  _T_269; // @[SpatialBlocks.scala 130:61:@22647.4]
  x278_ctrchain x278_ctrchain ( // @[SpatialBlocks.scala 37:22:@22483.4]
    .clock(x278_ctrchain_clock),
    .reset(x278_ctrchain_reset),
    .io_input_reset(x278_ctrchain_io_input_reset),
    .io_input_enable(x278_ctrchain_io_input_enable),
    .io_output_counts_1(x278_ctrchain_io_output_counts_1),
    .io_output_counts_0(x278_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x278_ctrchain_io_output_oobs_0),
    .io_output_oobs_1(x278_ctrchain_io_output_oobs_1),
    .io_output_done(x278_ctrchain_io_output_done)
  );
  x472_inr_Foreach_SAMPLER_BOX_sm x472_inr_Foreach_SAMPLER_BOX_sm ( // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 32:18:@22542.4]
    .clock(x472_inr_Foreach_SAMPLER_BOX_sm_clock),
    .reset(x472_inr_Foreach_SAMPLER_BOX_sm_reset),
    .io_enable(x472_inr_Foreach_SAMPLER_BOX_sm_io_enable),
    .io_done(x472_inr_Foreach_SAMPLER_BOX_sm_io_done),
    .io_doneLatch(x472_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch),
    .io_ctrDone(x472_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone),
    .io_datapathEn(x472_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn),
    .io_ctrInc(x472_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc),
    .io_ctrRst(x472_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst),
    .io_parentAck(x472_inr_Foreach_SAMPLER_BOX_sm_io_parentAck),
    .io_backpressure(x472_inr_Foreach_SAMPLER_BOX_sm_io_backpressure),
    .io_break(x472_inr_Foreach_SAMPLER_BOX_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@22570.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@22612.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@22620.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1 x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1 ( // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 568:24:@22652.4]
    .clock(x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_clock),
    .reset(x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_reset),
    .io_in_x270_TREADY(x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x270_TREADY),
    .io_in_x270_TDATA(x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x270_TDATA),
    .io_in_x270_TID(x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x270_TID),
    .io_in_x270_TDEST(x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x270_TDEST),
    .io_in_x271_TVALID(x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x271_TVALID),
    .io_in_x271_TREADY(x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x271_TREADY),
    .io_in_x271_TDATA(x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x271_TDATA),
    .io_sigsIn_backpressure(x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_1(x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsIn_cchainOutputs_0_oobs_1(x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1),
    .io_rr(x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_rr)
  );
  assign _T_239 = RetimeWrapper_io_out; // @[package.scala 96:25:@22575.4 package.scala 96:25:@22576.4]
  assign x472_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure = io_in_x270_TVALID | x472_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x473_outr_UnitPipe.scala 68:66:@22581.4]
  assign _T_252 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@22617.4 package.scala 96:25:@22618.4]
  assign _T_258 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@22625.4 package.scala 96:25:@22626.4]
  assign _T_261 = ~ _T_258; // @[SpatialBlocks.scala 110:93:@22628.4]
  assign x472_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn = _T_252 & _T_261; // @[SpatialBlocks.scala 110:90:@22629.4]
  assign _T_263 = x472_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[SpatialBlocks.scala 128:36:@22637.4]
  assign _T_264 = ~ x472_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[SpatialBlocks.scala 128:78:@22638.4]
  assign _T_269 = x472_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[SpatialBlocks.scala 130:61:@22647.4]
  assign io_in_x270_TREADY = x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x270_TREADY; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 48:23:@22709.4]
  assign io_in_x271_TVALID = x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x271_TVALID; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 49:23:@22719.4]
  assign io_in_x271_TDATA = x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x271_TDATA; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 49:23:@22717.4]
  assign io_sigsOut_smDoneIn_0 = x472_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[SpatialBlocks.scala 127:53:@22635.4]
  assign io_sigsOut_smCtrCopyDone_0 = x472_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[SpatialBlocks.scala 139:125:@22651.4]
  assign x278_ctrchain_clock = clock; // @[:@22484.4]
  assign x278_ctrchain_reset = reset; // @[:@22485.4]
  assign x278_ctrchain_io_input_reset = x472_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[SpatialBlocks.scala 130:103:@22650.4]
  assign x278_ctrchain_io_input_enable = _T_269 & x472_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 104:75:@22605.4 SpatialBlocks.scala 130:45:@22649.4]
  assign x472_inr_Foreach_SAMPLER_BOX_sm_clock = clock; // @[:@22543.4]
  assign x472_inr_Foreach_SAMPLER_BOX_sm_reset = reset; // @[:@22544.4]
  assign x472_inr_Foreach_SAMPLER_BOX_sm_io_enable = x472_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn & x472_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 112:18:@22632.4]
  assign x472_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone = io_rr ? _T_239 : 1'h0; // @[sm_x473_outr_UnitPipe.scala 66:50:@22578.4]
  assign x472_inr_Foreach_SAMPLER_BOX_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 114:21:@22634.4]
  assign x472_inr_Foreach_SAMPLER_BOX_sm_io_backpressure = io_in_x271_TREADY | x472_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[SpatialBlocks.scala 105:24:@22606.4]
  assign x472_inr_Foreach_SAMPLER_BOX_sm_io_break = 1'h0; // @[sm_x473_outr_UnitPipe.scala 70:48:@22584.4]
  assign RetimeWrapper_clock = clock; // @[:@22571.4]
  assign RetimeWrapper_reset = reset; // @[:@22572.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@22574.4]
  assign RetimeWrapper_io_in = x278_ctrchain_io_output_done; // @[package.scala 94:16:@22573.4]
  assign RetimeWrapper_1_clock = clock; // @[:@22613.4]
  assign RetimeWrapper_1_reset = reset; // @[:@22614.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@22616.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@22615.4]
  assign RetimeWrapper_2_clock = clock; // @[:@22621.4]
  assign RetimeWrapper_2_reset = reset; // @[:@22622.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@22624.4]
  assign RetimeWrapper_2_io_in = x472_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[package.scala 94:16:@22623.4]
  assign x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_clock = clock; // @[:@22653.4]
  assign x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_reset = reset; // @[:@22654.4]
  assign x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x270_TDATA = io_in_x270_TDATA; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 48:23:@22708.4]
  assign x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x270_TID = io_in_x270_TID; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 48:23:@22704.4]
  assign x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x270_TDEST = io_in_x270_TDEST; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 48:23:@22703.4]
  assign x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x271_TREADY = io_in_x271_TREADY; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 49:23:@22718.4]
  assign x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure = io_in_x271_TREADY | x472_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 572:22:@22736.4]
  assign x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn = _T_263 & _T_264; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 572:22:@22734.4]
  assign x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break = x472_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 572:22:@22732.4]
  assign x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1 = x278_ctrchain_io_output_counts_1; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 572:22:@22727.4]
  assign x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = x278_ctrchain_io_output_counts_0; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 572:22:@22726.4]
  assign x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x278_ctrchain_io_output_oobs_0; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 572:22:@22724.4]
  assign x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1 = x278_ctrchain_io_output_oobs_1; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 572:22:@22725.4]
  assign x472_inr_Foreach_SAMPLER_BOX_kernelx472_inr_Foreach_SAMPLER_BOX_concrete1_io_rr = io_rr; // @[sm_x472_inr_Foreach_SAMPLER_BOX.scala 571:18:@22720.4]
endmodule
module RootController_kernelRootController_concrete1( // @[:@22749.2]
  input          clock, // @[:@22750.4]
  input          reset, // @[:@22751.4]
  input          io_in_x270_TVALID, // @[:@22752.4]
  output         io_in_x270_TREADY, // @[:@22752.4]
  input  [255:0] io_in_x270_TDATA, // @[:@22752.4]
  input  [7:0]   io_in_x270_TID, // @[:@22752.4]
  input  [7:0]   io_in_x270_TDEST, // @[:@22752.4]
  output         io_in_x271_TVALID, // @[:@22752.4]
  input          io_in_x271_TREADY, // @[:@22752.4]
  output [255:0] io_in_x271_TDATA, // @[:@22752.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@22752.4]
  input          io_sigsIn_smChildAcks_0, // @[:@22752.4]
  output         io_sigsOut_smDoneIn_0, // @[:@22752.4]
  input          io_rr // @[:@22752.4]
);
  wire  x473_outr_UnitPipe_sm_clock; // @[sm_x473_outr_UnitPipe.scala 32:18:@22893.4]
  wire  x473_outr_UnitPipe_sm_reset; // @[sm_x473_outr_UnitPipe.scala 32:18:@22893.4]
  wire  x473_outr_UnitPipe_sm_io_enable; // @[sm_x473_outr_UnitPipe.scala 32:18:@22893.4]
  wire  x473_outr_UnitPipe_sm_io_done; // @[sm_x473_outr_UnitPipe.scala 32:18:@22893.4]
  wire  x473_outr_UnitPipe_sm_io_parentAck; // @[sm_x473_outr_UnitPipe.scala 32:18:@22893.4]
  wire  x473_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x473_outr_UnitPipe.scala 32:18:@22893.4]
  wire  x473_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x473_outr_UnitPipe.scala 32:18:@22893.4]
  wire  x473_outr_UnitPipe_sm_io_childAck_0; // @[sm_x473_outr_UnitPipe.scala 32:18:@22893.4]
  wire  x473_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x473_outr_UnitPipe.scala 32:18:@22893.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@22945.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@22945.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@22945.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@22945.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@22945.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@22953.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@22953.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@22953.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@22953.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@22953.4]
  wire  x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_clock; // @[sm_x473_outr_UnitPipe.scala 75:24:@22980.4]
  wire  x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_reset; // @[sm_x473_outr_UnitPipe.scala 75:24:@22980.4]
  wire  x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_io_in_x270_TVALID; // @[sm_x473_outr_UnitPipe.scala 75:24:@22980.4]
  wire  x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_io_in_x270_TREADY; // @[sm_x473_outr_UnitPipe.scala 75:24:@22980.4]
  wire [255:0] x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_io_in_x270_TDATA; // @[sm_x473_outr_UnitPipe.scala 75:24:@22980.4]
  wire [7:0] x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_io_in_x270_TID; // @[sm_x473_outr_UnitPipe.scala 75:24:@22980.4]
  wire [7:0] x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_io_in_x270_TDEST; // @[sm_x473_outr_UnitPipe.scala 75:24:@22980.4]
  wire  x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_io_in_x271_TVALID; // @[sm_x473_outr_UnitPipe.scala 75:24:@22980.4]
  wire  x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_io_in_x271_TREADY; // @[sm_x473_outr_UnitPipe.scala 75:24:@22980.4]
  wire [255:0] x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_io_in_x271_TDATA; // @[sm_x473_outr_UnitPipe.scala 75:24:@22980.4]
  wire  x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x473_outr_UnitPipe.scala 75:24:@22980.4]
  wire  x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x473_outr_UnitPipe.scala 75:24:@22980.4]
  wire  x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x473_outr_UnitPipe.scala 75:24:@22980.4]
  wire  x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x473_outr_UnitPipe.scala 75:24:@22980.4]
  wire  x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_io_rr; // @[sm_x473_outr_UnitPipe.scala 75:24:@22980.4]
  wire  _T_246; // @[package.scala 96:25:@22950.4 package.scala 96:25:@22951.4]
  wire  _T_252; // @[package.scala 96:25:@22958.4 package.scala 96:25:@22959.4]
  wire  _T_255; // @[SpatialBlocks.scala 110:93:@22961.4]
  x473_outr_UnitPipe_sm x473_outr_UnitPipe_sm ( // @[sm_x473_outr_UnitPipe.scala 32:18:@22893.4]
    .clock(x473_outr_UnitPipe_sm_clock),
    .reset(x473_outr_UnitPipe_sm_reset),
    .io_enable(x473_outr_UnitPipe_sm_io_enable),
    .io_done(x473_outr_UnitPipe_sm_io_done),
    .io_parentAck(x473_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x473_outr_UnitPipe_sm_io_doneIn_0),
    .io_enableOut_0(x473_outr_UnitPipe_sm_io_enableOut_0),
    .io_childAck_0(x473_outr_UnitPipe_sm_io_childAck_0),
    .io_ctrCopyDone_0(x473_outr_UnitPipe_sm_io_ctrCopyDone_0)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@22945.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@22953.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1 x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1 ( // @[sm_x473_outr_UnitPipe.scala 75:24:@22980.4]
    .clock(x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_clock),
    .reset(x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_reset),
    .io_in_x270_TVALID(x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_io_in_x270_TVALID),
    .io_in_x270_TREADY(x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_io_in_x270_TREADY),
    .io_in_x270_TDATA(x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_io_in_x270_TDATA),
    .io_in_x270_TID(x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_io_in_x270_TID),
    .io_in_x270_TDEST(x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_io_in_x270_TDEST),
    .io_in_x271_TVALID(x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_io_in_x271_TVALID),
    .io_in_x271_TREADY(x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_io_in_x271_TREADY),
    .io_in_x271_TDATA(x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_io_in_x271_TDATA),
    .io_sigsIn_smEnableOuts_0(x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smCtrCopyDone_0(x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_rr(x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_246 = RetimeWrapper_io_out; // @[package.scala 96:25:@22950.4 package.scala 96:25:@22951.4]
  assign _T_252 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@22958.4 package.scala 96:25:@22959.4]
  assign _T_255 = ~ _T_252; // @[SpatialBlocks.scala 110:93:@22961.4]
  assign io_in_x270_TREADY = x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_io_in_x270_TREADY; // @[sm_x473_outr_UnitPipe.scala 48:23:@23035.4]
  assign io_in_x271_TVALID = x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_io_in_x271_TVALID; // @[sm_x473_outr_UnitPipe.scala 49:23:@23045.4]
  assign io_in_x271_TDATA = x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_io_in_x271_TDATA; // @[sm_x473_outr_UnitPipe.scala 49:23:@23043.4]
  assign io_sigsOut_smDoneIn_0 = x473_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 127:53:@22968.4]
  assign x473_outr_UnitPipe_sm_clock = clock; // @[:@22894.4]
  assign x473_outr_UnitPipe_sm_reset = reset; // @[:@22895.4]
  assign x473_outr_UnitPipe_sm_io_enable = _T_246 & _T_255; // @[SpatialBlocks.scala 112:18:@22965.4]
  assign x473_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 114:21:@22967.4]
  assign x473_outr_UnitPipe_sm_io_doneIn_0 = x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 102:67:@22937.4]
  assign x473_outr_UnitPipe_sm_io_ctrCopyDone_0 = x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 132:80:@22979.4]
  assign RetimeWrapper_clock = clock; // @[:@22946.4]
  assign RetimeWrapper_reset = reset; // @[:@22947.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@22949.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@22948.4]
  assign RetimeWrapper_1_clock = clock; // @[:@22954.4]
  assign RetimeWrapper_1_reset = reset; // @[:@22955.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@22957.4]
  assign RetimeWrapper_1_io_in = x473_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@22956.4]
  assign x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_clock = clock; // @[:@22981.4]
  assign x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_reset = reset; // @[:@22982.4]
  assign x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_io_in_x270_TVALID = io_in_x270_TVALID; // @[sm_x473_outr_UnitPipe.scala 48:23:@23036.4]
  assign x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_io_in_x270_TDATA = io_in_x270_TDATA; // @[sm_x473_outr_UnitPipe.scala 48:23:@23034.4]
  assign x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_io_in_x270_TID = io_in_x270_TID; // @[sm_x473_outr_UnitPipe.scala 48:23:@23030.4]
  assign x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_io_in_x270_TDEST = io_in_x270_TDEST; // @[sm_x473_outr_UnitPipe.scala 48:23:@23029.4]
  assign x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_io_in_x271_TREADY = io_in_x271_TREADY; // @[sm_x473_outr_UnitPipe.scala 49:23:@23044.4]
  assign x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x473_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x473_outr_UnitPipe.scala 79:22:@23054.4]
  assign x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x473_outr_UnitPipe_sm_io_childAck_0; // @[sm_x473_outr_UnitPipe.scala 79:22:@23052.4]
  assign x473_outr_UnitPipe_kernelx473_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x473_outr_UnitPipe.scala 78:18:@23046.4]
endmodule
module AccelUnit( // @[:@23073.2]
  input          clock, // @[:@23074.4]
  input          reset, // @[:@23075.4]
  input          io_enable, // @[:@23076.4]
  output         io_done, // @[:@23076.4]
  input          io_reset, // @[:@23076.4]
  input          io_memStreams_loads_0_cmd_ready, // @[:@23076.4]
  output         io_memStreams_loads_0_cmd_valid, // @[:@23076.4]
  output [63:0]  io_memStreams_loads_0_cmd_bits_addr, // @[:@23076.4]
  output [31:0]  io_memStreams_loads_0_cmd_bits_size, // @[:@23076.4]
  output         io_memStreams_loads_0_data_ready, // @[:@23076.4]
  input          io_memStreams_loads_0_data_valid, // @[:@23076.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_0, // @[:@23076.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_1, // @[:@23076.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_2, // @[:@23076.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_3, // @[:@23076.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_4, // @[:@23076.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_5, // @[:@23076.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_6, // @[:@23076.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_7, // @[:@23076.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_8, // @[:@23076.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_9, // @[:@23076.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_10, // @[:@23076.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_11, // @[:@23076.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_12, // @[:@23076.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_13, // @[:@23076.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_14, // @[:@23076.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_15, // @[:@23076.4]
  input          io_memStreams_stores_0_cmd_ready, // @[:@23076.4]
  output         io_memStreams_stores_0_cmd_valid, // @[:@23076.4]
  output [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@23076.4]
  output [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@23076.4]
  input          io_memStreams_stores_0_data_ready, // @[:@23076.4]
  output         io_memStreams_stores_0_data_valid, // @[:@23076.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_0, // @[:@23076.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_1, // @[:@23076.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_2, // @[:@23076.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_3, // @[:@23076.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_4, // @[:@23076.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_5, // @[:@23076.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_6, // @[:@23076.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_7, // @[:@23076.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_8, // @[:@23076.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_9, // @[:@23076.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_10, // @[:@23076.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_11, // @[:@23076.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_12, // @[:@23076.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_13, // @[:@23076.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_14, // @[:@23076.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_15, // @[:@23076.4]
  output [15:0]  io_memStreams_stores_0_data_bits_wstrb, // @[:@23076.4]
  output         io_memStreams_stores_0_wresp_ready, // @[:@23076.4]
  input          io_memStreams_stores_0_wresp_valid, // @[:@23076.4]
  input          io_memStreams_stores_0_wresp_bits, // @[:@23076.4]
  input          io_memStreams_gathers_0_cmd_ready, // @[:@23076.4]
  output         io_memStreams_gathers_0_cmd_valid, // @[:@23076.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_0, // @[:@23076.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_1, // @[:@23076.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_2, // @[:@23076.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_3, // @[:@23076.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_4, // @[:@23076.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_5, // @[:@23076.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_6, // @[:@23076.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_7, // @[:@23076.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_8, // @[:@23076.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_9, // @[:@23076.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_10, // @[:@23076.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_11, // @[:@23076.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_12, // @[:@23076.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_13, // @[:@23076.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_14, // @[:@23076.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_15, // @[:@23076.4]
  output         io_memStreams_gathers_0_data_ready, // @[:@23076.4]
  input          io_memStreams_gathers_0_data_valid, // @[:@23076.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_0, // @[:@23076.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_1, // @[:@23076.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_2, // @[:@23076.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_3, // @[:@23076.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_4, // @[:@23076.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_5, // @[:@23076.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_6, // @[:@23076.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_7, // @[:@23076.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_8, // @[:@23076.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_9, // @[:@23076.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_10, // @[:@23076.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_11, // @[:@23076.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_12, // @[:@23076.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_13, // @[:@23076.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_14, // @[:@23076.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_15, // @[:@23076.4]
  input          io_memStreams_scatters_0_cmd_ready, // @[:@23076.4]
  output         io_memStreams_scatters_0_cmd_valid, // @[:@23076.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_0, // @[:@23076.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_1, // @[:@23076.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_2, // @[:@23076.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_3, // @[:@23076.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_4, // @[:@23076.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_5, // @[:@23076.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_6, // @[:@23076.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_7, // @[:@23076.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_8, // @[:@23076.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_9, // @[:@23076.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_10, // @[:@23076.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_11, // @[:@23076.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_12, // @[:@23076.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_13, // @[:@23076.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_14, // @[:@23076.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_15, // @[:@23076.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_0, // @[:@23076.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_1, // @[:@23076.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_2, // @[:@23076.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_3, // @[:@23076.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_4, // @[:@23076.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_5, // @[:@23076.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_6, // @[:@23076.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_7, // @[:@23076.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_8, // @[:@23076.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_9, // @[:@23076.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_10, // @[:@23076.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_11, // @[:@23076.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_12, // @[:@23076.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_13, // @[:@23076.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_14, // @[:@23076.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_15, // @[:@23076.4]
  output         io_memStreams_scatters_0_wresp_ready, // @[:@23076.4]
  input          io_memStreams_scatters_0_wresp_valid, // @[:@23076.4]
  input          io_memStreams_scatters_0_wresp_bits, // @[:@23076.4]
  input          io_axiStreamsIn_0_TVALID, // @[:@23076.4]
  output         io_axiStreamsIn_0_TREADY, // @[:@23076.4]
  input  [255:0] io_axiStreamsIn_0_TDATA, // @[:@23076.4]
  input  [31:0]  io_axiStreamsIn_0_TSTRB, // @[:@23076.4]
  input  [31:0]  io_axiStreamsIn_0_TKEEP, // @[:@23076.4]
  input          io_axiStreamsIn_0_TLAST, // @[:@23076.4]
  input  [7:0]   io_axiStreamsIn_0_TID, // @[:@23076.4]
  input  [7:0]   io_axiStreamsIn_0_TDEST, // @[:@23076.4]
  input  [31:0]  io_axiStreamsIn_0_TUSER, // @[:@23076.4]
  output         io_axiStreamsOut_0_TVALID, // @[:@23076.4]
  input          io_axiStreamsOut_0_TREADY, // @[:@23076.4]
  output [255:0] io_axiStreamsOut_0_TDATA, // @[:@23076.4]
  output [31:0]  io_axiStreamsOut_0_TSTRB, // @[:@23076.4]
  output [31:0]  io_axiStreamsOut_0_TKEEP, // @[:@23076.4]
  output         io_axiStreamsOut_0_TLAST, // @[:@23076.4]
  output [7:0]   io_axiStreamsOut_0_TID, // @[:@23076.4]
  output [7:0]   io_axiStreamsOut_0_TDEST, // @[:@23076.4]
  output [31:0]  io_axiStreamsOut_0_TUSER, // @[:@23076.4]
  output         io_heap_0_req_valid, // @[:@23076.4]
  output         io_heap_0_req_bits_allocDealloc, // @[:@23076.4]
  output [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@23076.4]
  input          io_heap_0_resp_valid, // @[:@23076.4]
  input          io_heap_0_resp_bits_allocDealloc, // @[:@23076.4]
  input  [63:0]  io_heap_0_resp_bits_sizeAddr, // @[:@23076.4]
  input  [63:0]  io_argIns_0, // @[:@23076.4]
  input  [63:0]  io_argIns_1, // @[:@23076.4]
  input          io_argOuts_0_port_ready, // @[:@23076.4]
  output         io_argOuts_0_port_valid, // @[:@23076.4]
  output [63:0]  io_argOuts_0_port_bits, // @[:@23076.4]
  input  [63:0]  io_argOuts_0_echo // @[:@23076.4]
);
  wire  SingleCounter_clock; // @[Main.scala 35:32:@23239.4]
  wire  SingleCounter_reset; // @[Main.scala 35:32:@23239.4]
  wire  SingleCounter_io_input_reset; // @[Main.scala 35:32:@23239.4]
  wire  SingleCounter_io_output_done; // @[Main.scala 35:32:@23239.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@23257.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@23257.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@23257.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@23257.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@23257.4]
  wire  SRFF_clock; // @[Main.scala 39:28:@23266.4]
  wire  SRFF_reset; // @[Main.scala 39:28:@23266.4]
  wire  SRFF_io_input_set; // @[Main.scala 39:28:@23266.4]
  wire  SRFF_io_input_reset; // @[Main.scala 39:28:@23266.4]
  wire  SRFF_io_input_asyn_reset; // @[Main.scala 39:28:@23266.4]
  wire  SRFF_io_output; // @[Main.scala 39:28:@23266.4]
  wire  RootController_sm_clock; // @[sm_RootController.scala 32:18:@23304.4]
  wire  RootController_sm_reset; // @[sm_RootController.scala 32:18:@23304.4]
  wire  RootController_sm_io_enable; // @[sm_RootController.scala 32:18:@23304.4]
  wire  RootController_sm_io_done; // @[sm_RootController.scala 32:18:@23304.4]
  wire  RootController_sm_io_rst; // @[sm_RootController.scala 32:18:@23304.4]
  wire  RootController_sm_io_ctrDone; // @[sm_RootController.scala 32:18:@23304.4]
  wire  RootController_sm_io_ctrInc; // @[sm_RootController.scala 32:18:@23304.4]
  wire  RootController_sm_io_doneIn_0; // @[sm_RootController.scala 32:18:@23304.4]
  wire  RootController_sm_io_enableOut_0; // @[sm_RootController.scala 32:18:@23304.4]
  wire  RootController_sm_io_childAck_0; // @[sm_RootController.scala 32:18:@23304.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@23336.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@23336.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@23336.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@23336.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@23336.4]
  wire  RootController_kernelRootController_concrete1_clock; // @[sm_RootController.scala 73:24:@23395.4]
  wire  RootController_kernelRootController_concrete1_reset; // @[sm_RootController.scala 73:24:@23395.4]
  wire  RootController_kernelRootController_concrete1_io_in_x270_TVALID; // @[sm_RootController.scala 73:24:@23395.4]
  wire  RootController_kernelRootController_concrete1_io_in_x270_TREADY; // @[sm_RootController.scala 73:24:@23395.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x270_TDATA; // @[sm_RootController.scala 73:24:@23395.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x270_TID; // @[sm_RootController.scala 73:24:@23395.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x270_TDEST; // @[sm_RootController.scala 73:24:@23395.4]
  wire  RootController_kernelRootController_concrete1_io_in_x271_TVALID; // @[sm_RootController.scala 73:24:@23395.4]
  wire  RootController_kernelRootController_concrete1_io_in_x271_TREADY; // @[sm_RootController.scala 73:24:@23395.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x271_TDATA; // @[sm_RootController.scala 73:24:@23395.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_RootController.scala 73:24:@23395.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0; // @[sm_RootController.scala 73:24:@23395.4]
  wire  RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[sm_RootController.scala 73:24:@23395.4]
  wire  RootController_kernelRootController_concrete1_io_rr; // @[sm_RootController.scala 73:24:@23395.4]
  wire  _T_599; // @[package.scala 96:25:@23262.4 package.scala 96:25:@23263.4]
  wire  _T_664; // @[Main.scala 41:50:@23332.4]
  wire  _T_665; // @[Main.scala 41:59:@23333.4]
  wire  _T_677; // @[package.scala 100:49:@23353.4]
  reg  _T_680; // @[package.scala 48:56:@23354.4]
  reg [31:0] _RAND_0;
  SingleCounter SingleCounter ( // @[Main.scala 35:32:@23239.4]
    .clock(SingleCounter_clock),
    .reset(SingleCounter_reset),
    .io_input_reset(SingleCounter_io_input_reset),
    .io_output_done(SingleCounter_io_output_done)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@23257.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  SRFF SRFF ( // @[Main.scala 39:28:@23266.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  RootController_sm RootController_sm ( // @[sm_RootController.scala 32:18:@23304.4]
    .clock(RootController_sm_clock),
    .reset(RootController_sm_reset),
    .io_enable(RootController_sm_io_enable),
    .io_done(RootController_sm_io_done),
    .io_rst(RootController_sm_io_rst),
    .io_ctrDone(RootController_sm_io_ctrDone),
    .io_ctrInc(RootController_sm_io_ctrInc),
    .io_doneIn_0(RootController_sm_io_doneIn_0),
    .io_enableOut_0(RootController_sm_io_enableOut_0),
    .io_childAck_0(RootController_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@23336.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RootController_kernelRootController_concrete1 RootController_kernelRootController_concrete1 ( // @[sm_RootController.scala 73:24:@23395.4]
    .clock(RootController_kernelRootController_concrete1_clock),
    .reset(RootController_kernelRootController_concrete1_reset),
    .io_in_x270_TVALID(RootController_kernelRootController_concrete1_io_in_x270_TVALID),
    .io_in_x270_TREADY(RootController_kernelRootController_concrete1_io_in_x270_TREADY),
    .io_in_x270_TDATA(RootController_kernelRootController_concrete1_io_in_x270_TDATA),
    .io_in_x270_TID(RootController_kernelRootController_concrete1_io_in_x270_TID),
    .io_in_x270_TDEST(RootController_kernelRootController_concrete1_io_in_x270_TDEST),
    .io_in_x271_TVALID(RootController_kernelRootController_concrete1_io_in_x271_TVALID),
    .io_in_x271_TREADY(RootController_kernelRootController_concrete1_io_in_x271_TREADY),
    .io_in_x271_TDATA(RootController_kernelRootController_concrete1_io_in_x271_TDATA),
    .io_sigsIn_smEnableOuts_0(RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(RootController_kernelRootController_concrete1_io_rr)
  );
  assign _T_599 = RetimeWrapper_io_out; // @[package.scala 96:25:@23262.4 package.scala 96:25:@23263.4]
  assign _T_664 = io_enable & _T_599; // @[Main.scala 41:50:@23332.4]
  assign _T_665 = ~ SRFF_io_output; // @[Main.scala 41:59:@23333.4]
  assign _T_677 = RootController_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@23353.4]
  assign io_done = SRFF_io_output; // @[Main.scala 48:23:@23352.4]
  assign io_memStreams_loads_0_cmd_valid = 1'h0;
  assign io_memStreams_loads_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_loads_0_cmd_bits_size = 32'h0;
  assign io_memStreams_loads_0_data_ready = 1'h0;
  assign io_memStreams_stores_0_cmd_valid = 1'h0;
  assign io_memStreams_stores_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_stores_0_cmd_bits_size = 32'h0;
  assign io_memStreams_stores_0_data_valid = 1'h0;
  assign io_memStreams_stores_0_data_bits_wdata_0 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_1 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_2 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_3 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_4 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_5 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_6 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_7 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_8 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_9 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_10 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_11 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_12 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_13 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_14 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_15 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wstrb = 16'h0;
  assign io_memStreams_stores_0_wresp_ready = 1'h0;
  assign io_memStreams_gathers_0_cmd_valid = 1'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_0 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_1 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_2 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_3 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_4 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_5 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_6 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_7 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_8 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_9 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_10 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_11 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_12 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_13 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_14 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_15 = 64'h0;
  assign io_memStreams_gathers_0_data_ready = 1'h0;
  assign io_memStreams_scatters_0_cmd_valid = 1'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_0 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_1 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_2 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_3 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_4 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_5 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_6 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_7 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_8 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_9 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_10 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_11 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_12 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_13 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_14 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_15 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_0 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_1 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_2 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_3 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_4 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_5 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_6 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_7 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_8 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_9 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_10 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_11 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_12 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_13 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_14 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_15 = 32'h0;
  assign io_memStreams_scatters_0_wresp_ready = 1'h0;
  assign io_axiStreamsIn_0_TREADY = RootController_kernelRootController_concrete1_io_in_x270_TREADY; // @[sm_RootController.scala 48:23:@23450.4]
  assign io_axiStreamsOut_0_TVALID = RootController_kernelRootController_concrete1_io_in_x271_TVALID; // @[sm_RootController.scala 49:23:@23460.4]
  assign io_axiStreamsOut_0_TDATA = RootController_kernelRootController_concrete1_io_in_x271_TDATA; // @[sm_RootController.scala 49:23:@23458.4]
  assign io_axiStreamsOut_0_TSTRB = 32'hffffffff; // @[sm_RootController.scala 49:23:@23457.4]
  assign io_axiStreamsOut_0_TKEEP = 32'hffffffff; // @[sm_RootController.scala 49:23:@23456.4]
  assign io_axiStreamsOut_0_TLAST = 1'h0; // @[sm_RootController.scala 49:23:@23455.4]
  assign io_axiStreamsOut_0_TID = 8'h0; // @[sm_RootController.scala 49:23:@23454.4]
  assign io_axiStreamsOut_0_TDEST = 8'h0; // @[sm_RootController.scala 49:23:@23453.4]
  assign io_axiStreamsOut_0_TUSER = 32'h4; // @[sm_RootController.scala 49:23:@23452.4]
  assign io_heap_0_req_valid = 1'h0;
  assign io_heap_0_req_bits_allocDealloc = 1'h0;
  assign io_heap_0_req_bits_sizeAddr = 64'h0;
  assign io_argOuts_0_port_valid = 1'h0;
  assign io_argOuts_0_port_bits = 64'h0;
  assign SingleCounter_clock = clock; // @[:@23240.4]
  assign SingleCounter_reset = reset; // @[:@23241.4]
  assign SingleCounter_io_input_reset = reset; // @[Main.scala 36:79:@23255.4]
  assign RetimeWrapper_clock = clock; // @[:@23258.4]
  assign RetimeWrapper_reset = reset; // @[:@23259.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@23261.4]
  assign RetimeWrapper_io_in = SingleCounter_io_output_done; // @[package.scala 94:16:@23260.4]
  assign SRFF_clock = clock; // @[:@23267.4]
  assign SRFF_reset = reset; // @[:@23268.4]
  assign SRFF_io_input_set = RootController_sm_io_done; // @[Main.scala 57:29:@23487.4]
  assign SRFF_io_input_reset = RetimeWrapper_1_io_out; // @[Main.scala 46:31:@23350.4]
  assign SRFF_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[Main.scala 47:36:@23351.4]
  assign RootController_sm_clock = clock; // @[:@23305.4]
  assign RootController_sm_reset = reset; // @[:@23306.4]
  assign RootController_sm_io_enable = _T_664 & _T_665; // @[Main.scala 45:33:@23349.4 SpatialBlocks.scala 112:18:@23383.4]
  assign RootController_sm_io_rst = RetimeWrapper_1_io_out; // @[SpatialBlocks.scala 106:15:@23377.4]
  assign RootController_sm_io_ctrDone = RootController_sm_io_ctrInc & _T_680; // @[Main.scala 49:34:@23357.4]
  assign RootController_sm_io_doneIn_0 = RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 102:67:@23374.4]
  assign RetimeWrapper_1_clock = clock; // @[:@23337.4]
  assign RetimeWrapper_1_reset = reset; // @[:@23338.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@23340.4]
  assign RetimeWrapper_1_io_in = reset | io_reset; // @[package.scala 94:16:@23339.4]
  assign RootController_kernelRootController_concrete1_clock = clock; // @[:@23396.4]
  assign RootController_kernelRootController_concrete1_reset = reset; // @[:@23397.4]
  assign RootController_kernelRootController_concrete1_io_in_x270_TVALID = io_axiStreamsIn_0_TVALID; // @[sm_RootController.scala 48:23:@23451.4]
  assign RootController_kernelRootController_concrete1_io_in_x270_TDATA = io_axiStreamsIn_0_TDATA; // @[sm_RootController.scala 48:23:@23449.4]
  assign RootController_kernelRootController_concrete1_io_in_x270_TID = io_axiStreamsIn_0_TID; // @[sm_RootController.scala 48:23:@23445.4]
  assign RootController_kernelRootController_concrete1_io_in_x270_TDEST = io_axiStreamsIn_0_TDEST; // @[sm_RootController.scala 48:23:@23444.4]
  assign RootController_kernelRootController_concrete1_io_in_x271_TREADY = io_axiStreamsOut_0_TREADY; // @[sm_RootController.scala 49:23:@23459.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0 = RootController_sm_io_enableOut_0; // @[sm_RootController.scala 77:22:@23469.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0 = RootController_sm_io_childAck_0; // @[sm_RootController.scala 77:22:@23467.4]
  assign RootController_kernelRootController_concrete1_io_rr = RetimeWrapper_io_out; // @[sm_RootController.scala 76:18:@23461.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_680 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_680 <= 1'h0;
    end else begin
      _T_680 <= _T_677;
    end
  end
endmodule
module SpatialIP( // @[:@23489.2]
  input         clock, // @[:@23490.4]
  input         reset, // @[:@23491.4]
  input  [31:0] io_raddr, // @[:@23492.4]
  input         io_wen, // @[:@23492.4]
  input  [31:0] io_waddr, // @[:@23492.4]
  input  [63:0] io_wdata, // @[:@23492.4]
  output [63:0] io_rdata // @[:@23492.4]
);
  wire  accel_clock; // @[Instantiator.scala 53:44:@23494.4]
  wire  accel_reset; // @[Instantiator.scala 53:44:@23494.4]
  wire  accel_io_enable; // @[Instantiator.scala 53:44:@23494.4]
  wire  accel_io_done; // @[Instantiator.scala 53:44:@23494.4]
  wire  accel_io_reset; // @[Instantiator.scala 53:44:@23494.4]
  wire  accel_io_memStreams_loads_0_cmd_ready; // @[Instantiator.scala 53:44:@23494.4]
  wire  accel_io_memStreams_loads_0_cmd_valid; // @[Instantiator.scala 53:44:@23494.4]
  wire [63:0] accel_io_memStreams_loads_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_loads_0_cmd_bits_size; // @[Instantiator.scala 53:44:@23494.4]
  wire  accel_io_memStreams_loads_0_data_ready; // @[Instantiator.scala 53:44:@23494.4]
  wire  accel_io_memStreams_loads_0_data_valid; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_0; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_1; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_2; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_3; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_4; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_5; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_6; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_7; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_8; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_9; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_10; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_11; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_12; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_13; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_14; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_15; // @[Instantiator.scala 53:44:@23494.4]
  wire  accel_io_memStreams_stores_0_cmd_ready; // @[Instantiator.scala 53:44:@23494.4]
  wire  accel_io_memStreams_stores_0_cmd_valid; // @[Instantiator.scala 53:44:@23494.4]
  wire [63:0] accel_io_memStreams_stores_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_stores_0_cmd_bits_size; // @[Instantiator.scala 53:44:@23494.4]
  wire  accel_io_memStreams_stores_0_data_ready; // @[Instantiator.scala 53:44:@23494.4]
  wire  accel_io_memStreams_stores_0_data_valid; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_1; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_2; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_3; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_4; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_5; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_6; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_7; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_8; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_9; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_10; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_11; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_12; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_13; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_14; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_15; // @[Instantiator.scala 53:44:@23494.4]
  wire [15:0] accel_io_memStreams_stores_0_data_bits_wstrb; // @[Instantiator.scala 53:44:@23494.4]
  wire  accel_io_memStreams_stores_0_wresp_ready; // @[Instantiator.scala 53:44:@23494.4]
  wire  accel_io_memStreams_stores_0_wresp_valid; // @[Instantiator.scala 53:44:@23494.4]
  wire  accel_io_memStreams_stores_0_wresp_bits; // @[Instantiator.scala 53:44:@23494.4]
  wire  accel_io_memStreams_gathers_0_cmd_ready; // @[Instantiator.scala 53:44:@23494.4]
  wire  accel_io_memStreams_gathers_0_cmd_valid; // @[Instantiator.scala 53:44:@23494.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_0; // @[Instantiator.scala 53:44:@23494.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_1; // @[Instantiator.scala 53:44:@23494.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_2; // @[Instantiator.scala 53:44:@23494.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_3; // @[Instantiator.scala 53:44:@23494.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_4; // @[Instantiator.scala 53:44:@23494.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_5; // @[Instantiator.scala 53:44:@23494.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_6; // @[Instantiator.scala 53:44:@23494.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_7; // @[Instantiator.scala 53:44:@23494.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_8; // @[Instantiator.scala 53:44:@23494.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_9; // @[Instantiator.scala 53:44:@23494.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_10; // @[Instantiator.scala 53:44:@23494.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_11; // @[Instantiator.scala 53:44:@23494.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_12; // @[Instantiator.scala 53:44:@23494.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_13; // @[Instantiator.scala 53:44:@23494.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_14; // @[Instantiator.scala 53:44:@23494.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_15; // @[Instantiator.scala 53:44:@23494.4]
  wire  accel_io_memStreams_gathers_0_data_ready; // @[Instantiator.scala 53:44:@23494.4]
  wire  accel_io_memStreams_gathers_0_data_valid; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_0; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_1; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_2; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_3; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_4; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_5; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_6; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_7; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_8; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_9; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_10; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_11; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_12; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_13; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_14; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_15; // @[Instantiator.scala 53:44:@23494.4]
  wire  accel_io_memStreams_scatters_0_cmd_ready; // @[Instantiator.scala 53:44:@23494.4]
  wire  accel_io_memStreams_scatters_0_cmd_valid; // @[Instantiator.scala 53:44:@23494.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0; // @[Instantiator.scala 53:44:@23494.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1; // @[Instantiator.scala 53:44:@23494.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2; // @[Instantiator.scala 53:44:@23494.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3; // @[Instantiator.scala 53:44:@23494.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4; // @[Instantiator.scala 53:44:@23494.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5; // @[Instantiator.scala 53:44:@23494.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6; // @[Instantiator.scala 53:44:@23494.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7; // @[Instantiator.scala 53:44:@23494.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8; // @[Instantiator.scala 53:44:@23494.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9; // @[Instantiator.scala 53:44:@23494.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10; // @[Instantiator.scala 53:44:@23494.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11; // @[Instantiator.scala 53:44:@23494.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12; // @[Instantiator.scala 53:44:@23494.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13; // @[Instantiator.scala 53:44:@23494.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14; // @[Instantiator.scala 53:44:@23494.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_0; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_1; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_2; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_3; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_4; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_5; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_6; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_7; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_8; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_9; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_10; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_11; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_12; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_13; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_14; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_15; // @[Instantiator.scala 53:44:@23494.4]
  wire  accel_io_memStreams_scatters_0_wresp_ready; // @[Instantiator.scala 53:44:@23494.4]
  wire  accel_io_memStreams_scatters_0_wresp_valid; // @[Instantiator.scala 53:44:@23494.4]
  wire  accel_io_memStreams_scatters_0_wresp_bits; // @[Instantiator.scala 53:44:@23494.4]
  wire  accel_io_axiStreamsIn_0_TVALID; // @[Instantiator.scala 53:44:@23494.4]
  wire  accel_io_axiStreamsIn_0_TREADY; // @[Instantiator.scala 53:44:@23494.4]
  wire [255:0] accel_io_axiStreamsIn_0_TDATA; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_axiStreamsIn_0_TSTRB; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_axiStreamsIn_0_TKEEP; // @[Instantiator.scala 53:44:@23494.4]
  wire  accel_io_axiStreamsIn_0_TLAST; // @[Instantiator.scala 53:44:@23494.4]
  wire [7:0] accel_io_axiStreamsIn_0_TID; // @[Instantiator.scala 53:44:@23494.4]
  wire [7:0] accel_io_axiStreamsIn_0_TDEST; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_axiStreamsIn_0_TUSER; // @[Instantiator.scala 53:44:@23494.4]
  wire  accel_io_axiStreamsOut_0_TVALID; // @[Instantiator.scala 53:44:@23494.4]
  wire  accel_io_axiStreamsOut_0_TREADY; // @[Instantiator.scala 53:44:@23494.4]
  wire [255:0] accel_io_axiStreamsOut_0_TDATA; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_axiStreamsOut_0_TSTRB; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_axiStreamsOut_0_TKEEP; // @[Instantiator.scala 53:44:@23494.4]
  wire  accel_io_axiStreamsOut_0_TLAST; // @[Instantiator.scala 53:44:@23494.4]
  wire [7:0] accel_io_axiStreamsOut_0_TID; // @[Instantiator.scala 53:44:@23494.4]
  wire [7:0] accel_io_axiStreamsOut_0_TDEST; // @[Instantiator.scala 53:44:@23494.4]
  wire [31:0] accel_io_axiStreamsOut_0_TUSER; // @[Instantiator.scala 53:44:@23494.4]
  wire  accel_io_heap_0_req_valid; // @[Instantiator.scala 53:44:@23494.4]
  wire  accel_io_heap_0_req_bits_allocDealloc; // @[Instantiator.scala 53:44:@23494.4]
  wire [63:0] accel_io_heap_0_req_bits_sizeAddr; // @[Instantiator.scala 53:44:@23494.4]
  wire  accel_io_heap_0_resp_valid; // @[Instantiator.scala 53:44:@23494.4]
  wire  accel_io_heap_0_resp_bits_allocDealloc; // @[Instantiator.scala 53:44:@23494.4]
  wire [63:0] accel_io_heap_0_resp_bits_sizeAddr; // @[Instantiator.scala 53:44:@23494.4]
  wire [63:0] accel_io_argIns_0; // @[Instantiator.scala 53:44:@23494.4]
  wire [63:0] accel_io_argIns_1; // @[Instantiator.scala 53:44:@23494.4]
  wire  accel_io_argOuts_0_port_ready; // @[Instantiator.scala 53:44:@23494.4]
  wire  accel_io_argOuts_0_port_valid; // @[Instantiator.scala 53:44:@23494.4]
  wire [63:0] accel_io_argOuts_0_port_bits; // @[Instantiator.scala 53:44:@23494.4]
  wire [63:0] accel_io_argOuts_0_echo; // @[Instantiator.scala 53:44:@23494.4]
  AccelUnit accel ( // @[Instantiator.scala 53:44:@23494.4]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_enable(accel_io_enable),
    .io_done(accel_io_done),
    .io_reset(accel_io_reset),
    .io_memStreams_loads_0_cmd_ready(accel_io_memStreams_loads_0_cmd_ready),
    .io_memStreams_loads_0_cmd_valid(accel_io_memStreams_loads_0_cmd_valid),
    .io_memStreams_loads_0_cmd_bits_addr(accel_io_memStreams_loads_0_cmd_bits_addr),
    .io_memStreams_loads_0_cmd_bits_size(accel_io_memStreams_loads_0_cmd_bits_size),
    .io_memStreams_loads_0_data_ready(accel_io_memStreams_loads_0_data_ready),
    .io_memStreams_loads_0_data_valid(accel_io_memStreams_loads_0_data_valid),
    .io_memStreams_loads_0_data_bits_rdata_0(accel_io_memStreams_loads_0_data_bits_rdata_0),
    .io_memStreams_loads_0_data_bits_rdata_1(accel_io_memStreams_loads_0_data_bits_rdata_1),
    .io_memStreams_loads_0_data_bits_rdata_2(accel_io_memStreams_loads_0_data_bits_rdata_2),
    .io_memStreams_loads_0_data_bits_rdata_3(accel_io_memStreams_loads_0_data_bits_rdata_3),
    .io_memStreams_loads_0_data_bits_rdata_4(accel_io_memStreams_loads_0_data_bits_rdata_4),
    .io_memStreams_loads_0_data_bits_rdata_5(accel_io_memStreams_loads_0_data_bits_rdata_5),
    .io_memStreams_loads_0_data_bits_rdata_6(accel_io_memStreams_loads_0_data_bits_rdata_6),
    .io_memStreams_loads_0_data_bits_rdata_7(accel_io_memStreams_loads_0_data_bits_rdata_7),
    .io_memStreams_loads_0_data_bits_rdata_8(accel_io_memStreams_loads_0_data_bits_rdata_8),
    .io_memStreams_loads_0_data_bits_rdata_9(accel_io_memStreams_loads_0_data_bits_rdata_9),
    .io_memStreams_loads_0_data_bits_rdata_10(accel_io_memStreams_loads_0_data_bits_rdata_10),
    .io_memStreams_loads_0_data_bits_rdata_11(accel_io_memStreams_loads_0_data_bits_rdata_11),
    .io_memStreams_loads_0_data_bits_rdata_12(accel_io_memStreams_loads_0_data_bits_rdata_12),
    .io_memStreams_loads_0_data_bits_rdata_13(accel_io_memStreams_loads_0_data_bits_rdata_13),
    .io_memStreams_loads_0_data_bits_rdata_14(accel_io_memStreams_loads_0_data_bits_rdata_14),
    .io_memStreams_loads_0_data_bits_rdata_15(accel_io_memStreams_loads_0_data_bits_rdata_15),
    .io_memStreams_stores_0_cmd_ready(accel_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(accel_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(accel_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(accel_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(accel_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(accel_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(accel_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wdata_1(accel_io_memStreams_stores_0_data_bits_wdata_1),
    .io_memStreams_stores_0_data_bits_wdata_2(accel_io_memStreams_stores_0_data_bits_wdata_2),
    .io_memStreams_stores_0_data_bits_wdata_3(accel_io_memStreams_stores_0_data_bits_wdata_3),
    .io_memStreams_stores_0_data_bits_wdata_4(accel_io_memStreams_stores_0_data_bits_wdata_4),
    .io_memStreams_stores_0_data_bits_wdata_5(accel_io_memStreams_stores_0_data_bits_wdata_5),
    .io_memStreams_stores_0_data_bits_wdata_6(accel_io_memStreams_stores_0_data_bits_wdata_6),
    .io_memStreams_stores_0_data_bits_wdata_7(accel_io_memStreams_stores_0_data_bits_wdata_7),
    .io_memStreams_stores_0_data_bits_wdata_8(accel_io_memStreams_stores_0_data_bits_wdata_8),
    .io_memStreams_stores_0_data_bits_wdata_9(accel_io_memStreams_stores_0_data_bits_wdata_9),
    .io_memStreams_stores_0_data_bits_wdata_10(accel_io_memStreams_stores_0_data_bits_wdata_10),
    .io_memStreams_stores_0_data_bits_wdata_11(accel_io_memStreams_stores_0_data_bits_wdata_11),
    .io_memStreams_stores_0_data_bits_wdata_12(accel_io_memStreams_stores_0_data_bits_wdata_12),
    .io_memStreams_stores_0_data_bits_wdata_13(accel_io_memStreams_stores_0_data_bits_wdata_13),
    .io_memStreams_stores_0_data_bits_wdata_14(accel_io_memStreams_stores_0_data_bits_wdata_14),
    .io_memStreams_stores_0_data_bits_wdata_15(accel_io_memStreams_stores_0_data_bits_wdata_15),
    .io_memStreams_stores_0_data_bits_wstrb(accel_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(accel_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(accel_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(accel_io_memStreams_stores_0_wresp_bits),
    .io_memStreams_gathers_0_cmd_ready(accel_io_memStreams_gathers_0_cmd_ready),
    .io_memStreams_gathers_0_cmd_valid(accel_io_memStreams_gathers_0_cmd_valid),
    .io_memStreams_gathers_0_cmd_bits_addr_0(accel_io_memStreams_gathers_0_cmd_bits_addr_0),
    .io_memStreams_gathers_0_cmd_bits_addr_1(accel_io_memStreams_gathers_0_cmd_bits_addr_1),
    .io_memStreams_gathers_0_cmd_bits_addr_2(accel_io_memStreams_gathers_0_cmd_bits_addr_2),
    .io_memStreams_gathers_0_cmd_bits_addr_3(accel_io_memStreams_gathers_0_cmd_bits_addr_3),
    .io_memStreams_gathers_0_cmd_bits_addr_4(accel_io_memStreams_gathers_0_cmd_bits_addr_4),
    .io_memStreams_gathers_0_cmd_bits_addr_5(accel_io_memStreams_gathers_0_cmd_bits_addr_5),
    .io_memStreams_gathers_0_cmd_bits_addr_6(accel_io_memStreams_gathers_0_cmd_bits_addr_6),
    .io_memStreams_gathers_0_cmd_bits_addr_7(accel_io_memStreams_gathers_0_cmd_bits_addr_7),
    .io_memStreams_gathers_0_cmd_bits_addr_8(accel_io_memStreams_gathers_0_cmd_bits_addr_8),
    .io_memStreams_gathers_0_cmd_bits_addr_9(accel_io_memStreams_gathers_0_cmd_bits_addr_9),
    .io_memStreams_gathers_0_cmd_bits_addr_10(accel_io_memStreams_gathers_0_cmd_bits_addr_10),
    .io_memStreams_gathers_0_cmd_bits_addr_11(accel_io_memStreams_gathers_0_cmd_bits_addr_11),
    .io_memStreams_gathers_0_cmd_bits_addr_12(accel_io_memStreams_gathers_0_cmd_bits_addr_12),
    .io_memStreams_gathers_0_cmd_bits_addr_13(accel_io_memStreams_gathers_0_cmd_bits_addr_13),
    .io_memStreams_gathers_0_cmd_bits_addr_14(accel_io_memStreams_gathers_0_cmd_bits_addr_14),
    .io_memStreams_gathers_0_cmd_bits_addr_15(accel_io_memStreams_gathers_0_cmd_bits_addr_15),
    .io_memStreams_gathers_0_data_ready(accel_io_memStreams_gathers_0_data_ready),
    .io_memStreams_gathers_0_data_valid(accel_io_memStreams_gathers_0_data_valid),
    .io_memStreams_gathers_0_data_bits_0(accel_io_memStreams_gathers_0_data_bits_0),
    .io_memStreams_gathers_0_data_bits_1(accel_io_memStreams_gathers_0_data_bits_1),
    .io_memStreams_gathers_0_data_bits_2(accel_io_memStreams_gathers_0_data_bits_2),
    .io_memStreams_gathers_0_data_bits_3(accel_io_memStreams_gathers_0_data_bits_3),
    .io_memStreams_gathers_0_data_bits_4(accel_io_memStreams_gathers_0_data_bits_4),
    .io_memStreams_gathers_0_data_bits_5(accel_io_memStreams_gathers_0_data_bits_5),
    .io_memStreams_gathers_0_data_bits_6(accel_io_memStreams_gathers_0_data_bits_6),
    .io_memStreams_gathers_0_data_bits_7(accel_io_memStreams_gathers_0_data_bits_7),
    .io_memStreams_gathers_0_data_bits_8(accel_io_memStreams_gathers_0_data_bits_8),
    .io_memStreams_gathers_0_data_bits_9(accel_io_memStreams_gathers_0_data_bits_9),
    .io_memStreams_gathers_0_data_bits_10(accel_io_memStreams_gathers_0_data_bits_10),
    .io_memStreams_gathers_0_data_bits_11(accel_io_memStreams_gathers_0_data_bits_11),
    .io_memStreams_gathers_0_data_bits_12(accel_io_memStreams_gathers_0_data_bits_12),
    .io_memStreams_gathers_0_data_bits_13(accel_io_memStreams_gathers_0_data_bits_13),
    .io_memStreams_gathers_0_data_bits_14(accel_io_memStreams_gathers_0_data_bits_14),
    .io_memStreams_gathers_0_data_bits_15(accel_io_memStreams_gathers_0_data_bits_15),
    .io_memStreams_scatters_0_cmd_ready(accel_io_memStreams_scatters_0_cmd_ready),
    .io_memStreams_scatters_0_cmd_valid(accel_io_memStreams_scatters_0_cmd_valid),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_0(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_1(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_2(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_3(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_4(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_5(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_6(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_7(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_8(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_9(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_10(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_11(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_12(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_13(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_14(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_15(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15),
    .io_memStreams_scatters_0_cmd_bits_wdata_0(accel_io_memStreams_scatters_0_cmd_bits_wdata_0),
    .io_memStreams_scatters_0_cmd_bits_wdata_1(accel_io_memStreams_scatters_0_cmd_bits_wdata_1),
    .io_memStreams_scatters_0_cmd_bits_wdata_2(accel_io_memStreams_scatters_0_cmd_bits_wdata_2),
    .io_memStreams_scatters_0_cmd_bits_wdata_3(accel_io_memStreams_scatters_0_cmd_bits_wdata_3),
    .io_memStreams_scatters_0_cmd_bits_wdata_4(accel_io_memStreams_scatters_0_cmd_bits_wdata_4),
    .io_memStreams_scatters_0_cmd_bits_wdata_5(accel_io_memStreams_scatters_0_cmd_bits_wdata_5),
    .io_memStreams_scatters_0_cmd_bits_wdata_6(accel_io_memStreams_scatters_0_cmd_bits_wdata_6),
    .io_memStreams_scatters_0_cmd_bits_wdata_7(accel_io_memStreams_scatters_0_cmd_bits_wdata_7),
    .io_memStreams_scatters_0_cmd_bits_wdata_8(accel_io_memStreams_scatters_0_cmd_bits_wdata_8),
    .io_memStreams_scatters_0_cmd_bits_wdata_9(accel_io_memStreams_scatters_0_cmd_bits_wdata_9),
    .io_memStreams_scatters_0_cmd_bits_wdata_10(accel_io_memStreams_scatters_0_cmd_bits_wdata_10),
    .io_memStreams_scatters_0_cmd_bits_wdata_11(accel_io_memStreams_scatters_0_cmd_bits_wdata_11),
    .io_memStreams_scatters_0_cmd_bits_wdata_12(accel_io_memStreams_scatters_0_cmd_bits_wdata_12),
    .io_memStreams_scatters_0_cmd_bits_wdata_13(accel_io_memStreams_scatters_0_cmd_bits_wdata_13),
    .io_memStreams_scatters_0_cmd_bits_wdata_14(accel_io_memStreams_scatters_0_cmd_bits_wdata_14),
    .io_memStreams_scatters_0_cmd_bits_wdata_15(accel_io_memStreams_scatters_0_cmd_bits_wdata_15),
    .io_memStreams_scatters_0_wresp_ready(accel_io_memStreams_scatters_0_wresp_ready),
    .io_memStreams_scatters_0_wresp_valid(accel_io_memStreams_scatters_0_wresp_valid),
    .io_memStreams_scatters_0_wresp_bits(accel_io_memStreams_scatters_0_wresp_bits),
    .io_axiStreamsIn_0_TVALID(accel_io_axiStreamsIn_0_TVALID),
    .io_axiStreamsIn_0_TREADY(accel_io_axiStreamsIn_0_TREADY),
    .io_axiStreamsIn_0_TDATA(accel_io_axiStreamsIn_0_TDATA),
    .io_axiStreamsIn_0_TSTRB(accel_io_axiStreamsIn_0_TSTRB),
    .io_axiStreamsIn_0_TKEEP(accel_io_axiStreamsIn_0_TKEEP),
    .io_axiStreamsIn_0_TLAST(accel_io_axiStreamsIn_0_TLAST),
    .io_axiStreamsIn_0_TID(accel_io_axiStreamsIn_0_TID),
    .io_axiStreamsIn_0_TDEST(accel_io_axiStreamsIn_0_TDEST),
    .io_axiStreamsIn_0_TUSER(accel_io_axiStreamsIn_0_TUSER),
    .io_axiStreamsOut_0_TVALID(accel_io_axiStreamsOut_0_TVALID),
    .io_axiStreamsOut_0_TREADY(accel_io_axiStreamsOut_0_TREADY),
    .io_axiStreamsOut_0_TDATA(accel_io_axiStreamsOut_0_TDATA),
    .io_axiStreamsOut_0_TSTRB(accel_io_axiStreamsOut_0_TSTRB),
    .io_axiStreamsOut_0_TKEEP(accel_io_axiStreamsOut_0_TKEEP),
    .io_axiStreamsOut_0_TLAST(accel_io_axiStreamsOut_0_TLAST),
    .io_axiStreamsOut_0_TID(accel_io_axiStreamsOut_0_TID),
    .io_axiStreamsOut_0_TDEST(accel_io_axiStreamsOut_0_TDEST),
    .io_axiStreamsOut_0_TUSER(accel_io_axiStreamsOut_0_TUSER),
    .io_heap_0_req_valid(accel_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(accel_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(accel_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(accel_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(accel_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(accel_io_heap_0_resp_bits_sizeAddr),
    .io_argIns_0(accel_io_argIns_0),
    .io_argIns_1(accel_io_argIns_1),
    .io_argOuts_0_port_ready(accel_io_argOuts_0_port_ready),
    .io_argOuts_0_port_valid(accel_io_argOuts_0_port_valid),
    .io_argOuts_0_port_bits(accel_io_argOuts_0_port_bits),
    .io_argOuts_0_echo(accel_io_argOuts_0_echo)
  );
  assign io_rdata = 64'h0;
  assign accel_clock = clock; // @[:@23495.4]
  assign accel_reset = reset; // @[:@23496.4]
  assign accel_io_enable = 1'h0;
  assign accel_io_reset = 1'h0;
  assign accel_io_memStreams_loads_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_loads_0_data_valid = 1'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_0 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_1 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_2 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_3 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_4 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_5 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_6 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_7 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_8 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_9 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_10 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_11 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_12 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_13 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_14 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_15 = 32'h0;
  assign accel_io_memStreams_stores_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_stores_0_data_ready = 1'h0;
  assign accel_io_memStreams_stores_0_wresp_valid = 1'h0;
  assign accel_io_memStreams_stores_0_wresp_bits = 1'h0;
  assign accel_io_memStreams_gathers_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_gathers_0_data_valid = 1'h0;
  assign accel_io_memStreams_gathers_0_data_bits_0 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_1 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_2 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_3 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_4 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_5 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_6 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_7 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_8 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_9 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_10 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_11 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_12 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_13 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_14 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_15 = 32'h0;
  assign accel_io_memStreams_scatters_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_scatters_0_wresp_valid = 1'h0;
  assign accel_io_memStreams_scatters_0_wresp_bits = 1'h0;
  assign accel_io_axiStreamsIn_0_TVALID = 1'h0;
  assign accel_io_axiStreamsIn_0_TDATA = 256'h0;
  assign accel_io_axiStreamsIn_0_TSTRB = 32'h0;
  assign accel_io_axiStreamsIn_0_TKEEP = 32'h0;
  assign accel_io_axiStreamsIn_0_TLAST = 1'h0;
  assign accel_io_axiStreamsIn_0_TID = 8'h0;
  assign accel_io_axiStreamsIn_0_TDEST = 8'h0;
  assign accel_io_axiStreamsIn_0_TUSER = 32'h0;
  assign accel_io_axiStreamsOut_0_TREADY = 1'h0;
  assign accel_io_heap_0_resp_valid = 1'h0;
  assign accel_io_heap_0_resp_bits_allocDealloc = 1'h0;
  assign accel_io_heap_0_resp_bits_sizeAddr = 64'h0;
  assign accel_io_argIns_0 = 64'h0;
  assign accel_io_argIns_1 = 64'h0;
  assign accel_io_argOuts_0_port_ready = 1'h0;
  assign accel_io_argOuts_0_echo = 64'h0;
endmodule
