module stupleToSSeq_tInt_n3 (input [7:0] I_0, input [7:0] I_1, input [7:0] I_2, output [7:0] O_0, output [7:0] O_1, output [7:0] O_2, output valid_down, input valid_up);
assign O_0 = I_0;
assign O_1 = I_1;
assign O_2 = I_2;
assign valid_down = valid_up;
endmodule

module sseqTupleCreator_tInt (input [7:0] I0, input [7:0] I1, output [7:0] O_0, output [7:0] O_1, output valid_down, input valid_up);
assign O_0 = I0;
assign O_1 = I1;
assign valid_down = valid_up;
endmodule

module sseqTupleAppender_tInt_n2 (input [7:0] I0_0, input [7:0] I0_1, input [7:0] I1, output [7:0] O_0, output [7:0] O_1, output [7:0] O_2, output valid_down, input valid_up);
assign O_0 = I0_0;
assign O_1 = I0_1;
assign O_2 = I1;
assign valid_down = valid_up;
endmodule

module corebit_and (input in0, input in1, output out);
  assign out = in0 & in1;
endmodule

module atomTupleCreator_t0Int_t1Int (input [7:0] I0, input [7:0] I1, output [7:0] O__0, output [7:0] O__1, output valid_down, input valid_up);
assign O__0 = I0;
assign O__1 = I1;
assign valid_down = valid_up;
endmodule

module coreir_ult #(parameter width = 1) (input [width-1:0] in0, input [width-1:0] in1, output out);
  assign out = in0 < in1;
endmodule

module coreir_term #(parameter width = 1) (input [width-1:0] in);

endmodule

module coreir_shl #(parameter width = 1) (input [width-1:0] in0, input [width-1:0] in1, output [width-1:0] out);
  assign out = in0 << in1;
endmodule

module coreir_reg #(parameter width = 1, parameter clk_posedge = 1, parameter init = 1) (input clk, input [width-1:0] in, output [width-1:0] out);
  reg [width-1:0] outReg=init;
  wire real_clk;
  assign real_clk = clk_posedge ? clk : ~clk;
  always @(posedge real_clk) begin
    outReg <= in;
  end
  assign out = outReg;
endmodule

module coreir_mux #(parameter width = 1) (input [width-1:0] in0, input [width-1:0] in1, input sel, output [width-1:0] out);
  assign out = sel ? in1 : in0;
endmodule

module coreir_lshr #(parameter width = 1) (input [width-1:0] in0, input [width-1:0] in1, output [width-1:0] out);
  assign out = in0 >> in1;
endmodule

module coreir_eq #(parameter width = 1) (input [width-1:0] in0, input [width-1:0] in1, output out);
  assign out = in0 == in1;
endmodule

module coreir_const #(parameter width = 1, parameter value = 1) (output [width-1:0] out);
  assign out = value;
endmodule

module coreir_add #(parameter width = 1) (input [width-1:0] in0, input [width-1:0] in1, output [width-1:0] out);
  assign out = in0 + in1;
endmodule

module \commonlib_muxn__N2__width2 (input [1:0] in_data_0, input [1:0] in_data_1, input [0:0] in_sel, output [1:0] out);
wire [1:0] _join_out;
coreir_mux #(.width(2)) _join(.in0(in_data_0), .in1(in_data_1), .out(_join_out), .sel(in_sel[0]));
assign out = _join_out;
endmodule

module \commonlib_muxn__N2__width1 (input [0:0] in_data_0, input [0:0] in_data_1, input [0:0] in_sel, output [0:0] out);
wire [0:0] _join_out;
coreir_mux #(.width(1)) _join(.in0(in_data_0), .in1(in_data_1), .out(_join_out), .sel(in_sel[0]));
assign out = _join_out;
endmodule

module lutN #(parameter N = 1, parameter init = 1) (input [N-1:0] in, output out);
  assign out = init[in];
endmodule

module \aetherlinglib_hydrate__hydratedTypeBit83 (input [23:0] in, output [7:0] out_0, output [7:0] out_1, output [7:0] out_2);
assign out_0 = {in[7],in[6],in[5],in[4],in[3],in[2],in[1],in[0]};
assign out_1 = {in[15],in[14],in[13],in[12],in[11],in[10],in[9],in[8]};
assign out_2 = {in[23],in[22],in[21],in[20],in[19],in[18],in[17],in[16]};
endmodule

module \aetherlinglib_hydrate__hydratedTypeBit81 (input [7:0] in, output [7:0] out_0);
assign out_0 = {in[7],in[6],in[5],in[4],in[3],in[2],in[1],in[0]};
endmodule

module \aetherlinglib_dehydrate__hydratedTypeBit812 (input [7:0] in_0_0, input [7:0] in_1_0, output [15:0] out);
assign out = {in_1_0[7],in_1_0[6],in_1_0[5],in_1_0[4],in_1_0[3],in_1_0[2],in_1_0[1],in_1_0[0],in_0_0[7],in_0_0[6],in_0_0[5],in_0_0[4],in_0_0[3],in_0_0[2],in_0_0[1],in_0_0[0]};
endmodule

module \aetherlinglib_dehydrate__hydratedTypeBit (input in, output [0:0] out);
assign out = in;
endmodule

module Term_Bitt (input I);
wire [0:0] dehydrate_tBit_inst0_out;
\aetherlinglib_dehydrate__hydratedTypeBit dehydrate_tBit_inst0(.in(I), .out(dehydrate_tBit_inst0_out));
coreir_term #(.width(1)) term_w1_inst0(.in(dehydrate_tBit_inst0_out));
endmodule

module Term_Array_2_Array_1_Array_8_Bit___t (input [7:0] I_0_0, input [7:0] I_1_0);
wire [15:0] dehydrate_tArray_2_Array_1_Array_8_Bit____inst0_out;
\aetherlinglib_dehydrate__hydratedTypeBit812 dehydrate_tArray_2_Array_1_Array_8_Bit____inst0(.in_0_0(I_0_0), .in_1_0(I_1_0), .out(dehydrate_tArray_2_Array_1_Array_8_Bit____inst0_out));
coreir_term #(.width(16)) term_w16_inst0(.in(dehydrate_tArray_2_Array_1_Array_8_Bit____inst0_out));
endmodule

module SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse (input CE, input CLK, output [0:0] O);
wire [0:0] const_0_1_out;
Term_Bitt Term_Bitt_inst0(.I(CE));
coreir_const #(.value(1'h0), .width(1)) const_0_1(.out(const_0_1_out));
assign O = const_0_1_out;
endmodule

module Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue (input CLK, input [7:0] I_0_0, input [7:0] I_1_0, input [7:0] I_2_0, input [7:0] I_3_0, input [7:0] I_4_0, input [7:0] I_5_0, input [7:0] I_6_0, input [7:0] I_7_0, input [7:0] I_8_0, output [7:0] O_0_0, output [7:0] O_1_0, output [7:0] O_2_0, output [7:0] O_3_0, output [7:0] O_4_0, output [7:0] O_5_0, output [7:0] O_6_0, output [7:0] O_7_0, output [7:0] O_8_0, output valid_down, input valid_up);
assign O_0_0 = I_8_0;
assign O_1_0 = I_0_0;
assign O_2_0 = I_1_0;
assign O_3_0 = I_2_0;
assign O_4_0 = I_3_0;
assign O_5_0 = I_4_0;
assign O_6_0 = I_5_0;
assign O_7_0 = I_6_0;
assign O_8_0 = I_7_0;
assign valid_down = valid_up;
endmodule

module Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue (input CLK, input [7:0] I_0_0, input [7:0] I_10_0, input [7:0] I_11_0, input [7:0] I_12_0, input [7:0] I_13_0, input [7:0] I_14_0, input [7:0] I_15_0, input [7:0] I_16_0, input [7:0] I_17_0, input [7:0] I_18_0, input [7:0] I_19_0, input [7:0] I_1_0, input [7:0] I_20_0, input [7:0] I_21_0, input [7:0] I_22_0, input [7:0] I_23_0, input [7:0] I_24_0, input [7:0] I_25_0, input [7:0] I_26_0, input [7:0] I_2_0, input [7:0] I_3_0, input [7:0] I_4_0, input [7:0] I_5_0, input [7:0] I_6_0, input [7:0] I_7_0, input [7:0] I_8_0, input [7:0] I_9_0, output [7:0] O_0_0, output [7:0] O_10_0, output [7:0] O_11_0, output [7:0] O_12_0, output [7:0] O_13_0, output [7:0] O_14_0, output [7:0] O_15_0, output [7:0] O_16_0, output [7:0] O_17_0, output [7:0] O_18_0, output [7:0] O_19_0, output [7:0] O_1_0, output [7:0] O_20_0, output [7:0] O_21_0, output [7:0] O_22_0, output [7:0] O_23_0, output [7:0] O_24_0, output [7:0] O_25_0, output [7:0] O_26_0, output [7:0] O_2_0, output [7:0] O_3_0, output [7:0] O_4_0, output [7:0] O_5_0, output [7:0] O_6_0, output [7:0] O_7_0, output [7:0] O_8_0, output [7:0] O_9_0, output valid_down, input valid_up);
assign O_0_0 = I_26_0;
assign O_10_0 = I_9_0;
assign O_11_0 = I_10_0;
assign O_12_0 = I_11_0;
assign O_13_0 = I_12_0;
assign O_14_0 = I_13_0;
assign O_15_0 = I_14_0;
assign O_16_0 = I_15_0;
assign O_17_0 = I_16_0;
assign O_18_0 = I_17_0;
assign O_19_0 = I_18_0;
assign O_1_0 = I_0_0;
assign O_20_0 = I_19_0;
assign O_21_0 = I_20_0;
assign O_22_0 = I_21_0;
assign O_23_0 = I_22_0;
assign O_24_0 = I_23_0;
assign O_25_0 = I_24_0;
assign O_26_0 = I_25_0;
assign O_2_0 = I_1_0;
assign O_3_0 = I_2_0;
assign O_4_0 = I_3_0;
assign O_5_0 = I_4_0;
assign O_6_0 = I_5_0;
assign O_7_0 = I_6_0;
assign O_8_0 = I_7_0;
assign O_9_0 = I_8_0;
assign valid_down = valid_up;
endmodule

module Remove_1_S (input [7:0] I_0_0, input [7:0] I_0_1, input [7:0] I_0_2, output [7:0] O_0, output [7:0] O_1, output [7:0] O_2, output valid_down, input valid_up);
wire [7:0] stupleToSSeq_tInt_n3_inst0_O_0;
wire [7:0] stupleToSSeq_tInt_n3_inst0_O_1;
wire [7:0] stupleToSSeq_tInt_n3_inst0_O_2;
wire stupleToSSeq_tInt_n3_inst0_valid_down;
stupleToSSeq_tInt_n3 stupleToSSeq_tInt_n3_inst0(.I_0(I_0_0), .I_1(I_0_1), .I_2(I_0_2), .O_0(stupleToSSeq_tInt_n3_inst0_O_0), .O_1(stupleToSSeq_tInt_n3_inst0_O_1), .O_2(stupleToSSeq_tInt_n3_inst0_O_2), .valid_down(stupleToSSeq_tInt_n3_inst0_valid_down), .valid_up(valid_up));
assign O_0 = stupleToSSeq_tInt_n3_inst0_O_0;
assign O_1 = stupleToSSeq_tInt_n3_inst0_O_1;
assign O_2 = stupleToSSeq_tInt_n3_inst0_O_2;
assign valid_down = stupleToSSeq_tInt_n3_inst0_valid_down;
endmodule

module RShift_Atom (input [7:0] I__0, input [7:0] I__1, output [7:0] O, output valid_down, input valid_up);
wire [7:0] lshr8_inst0_out;
coreir_lshr #(.width(8)) lshr8_inst0(.in0(I__0), .in1(I__1), .out(lshr8_inst0_out));
assign O = lshr8_inst0_out;
assign valid_down = valid_up;
endmodule

module Partition_S_no9_ni3_tElSSeq_1_Int__vTrue (input CLK, input [7:0] I_0_0, input [7:0] I_10_0, input [7:0] I_11_0, input [7:0] I_12_0, input [7:0] I_13_0, input [7:0] I_14_0, input [7:0] I_15_0, input [7:0] I_16_0, input [7:0] I_17_0, input [7:0] I_18_0, input [7:0] I_19_0, input [7:0] I_1_0, input [7:0] I_20_0, input [7:0] I_21_0, input [7:0] I_22_0, input [7:0] I_23_0, input [7:0] I_24_0, input [7:0] I_25_0, input [7:0] I_26_0, input [7:0] I_2_0, input [7:0] I_3_0, input [7:0] I_4_0, input [7:0] I_5_0, input [7:0] I_6_0, input [7:0] I_7_0, input [7:0] I_8_0, input [7:0] I_9_0, output [7:0] O_0_0_0, output [7:0] O_0_1_0, output [7:0] O_0_2_0, output [7:0] O_1_0_0, output [7:0] O_1_1_0, output [7:0] O_1_2_0, output [7:0] O_2_0_0, output [7:0] O_2_1_0, output [7:0] O_2_2_0, output [7:0] O_3_0_0, output [7:0] O_3_1_0, output [7:0] O_3_2_0, output [7:0] O_4_0_0, output [7:0] O_4_1_0, output [7:0] O_4_2_0, output [7:0] O_5_0_0, output [7:0] O_5_1_0, output [7:0] O_5_2_0, output [7:0] O_6_0_0, output [7:0] O_6_1_0, output [7:0] O_6_2_0, output [7:0] O_7_0_0, output [7:0] O_7_1_0, output [7:0] O_7_2_0, output [7:0] O_8_0_0, output [7:0] O_8_1_0, output [7:0] O_8_2_0, output valid_down, input valid_up);
assign O_0_0_0 = I_0_0;
assign O_0_1_0 = I_1_0;
assign O_0_2_0 = I_2_0;
assign O_1_0_0 = I_3_0;
assign O_1_1_0 = I_4_0;
assign O_1_2_0 = I_5_0;
assign O_2_0_0 = I_6_0;
assign O_2_1_0 = I_7_0;
assign O_2_2_0 = I_8_0;
assign O_3_0_0 = I_9_0;
assign O_3_1_0 = I_10_0;
assign O_3_2_0 = I_11_0;
assign O_4_0_0 = I_12_0;
assign O_4_1_0 = I_13_0;
assign O_4_2_0 = I_14_0;
assign O_5_0_0 = I_15_0;
assign O_5_1_0 = I_16_0;
assign O_5_2_0 = I_17_0;
assign O_6_0_0 = I_18_0;
assign O_6_1_0 = I_19_0;
assign O_6_2_0 = I_20_0;
assign O_7_0_0 = I_21_0;
assign O_7_1_0 = I_22_0;
assign O_7_2_0 = I_23_0;
assign O_8_0_0 = I_24_0;
assign O_8_1_0 = I_25_0;
assign O_8_2_0 = I_26_0;
assign valid_down = valid_up;
endmodule

module Partition_S_no9_ni1_tElSSeq_1_Int__vTrue (input CLK, input [7:0] I_0_0_0, input [7:0] I_1_0_0, input [7:0] I_2_0_0, input [7:0] I_3_0_0, input [7:0] I_4_0_0, input [7:0] I_5_0_0, input [7:0] I_6_0_0, input [7:0] I_7_0_0, input [7:0] I_8_0_0, output [7:0] O_0_0, output [7:0] O_1_0, output [7:0] O_2_0, output [7:0] O_3_0, output [7:0] O_4_0, output [7:0] O_5_0, output [7:0] O_6_0, output [7:0] O_7_0, output [7:0] O_8_0, output valid_down, input valid_up);
assign O_0_0 = I_0_0_0;
assign O_1_0 = I_1_0_0;
assign O_2_0 = I_2_0_0;
assign O_3_0 = I_3_0_0;
assign O_4_0 = I_4_0_0;
assign O_5_0 = I_5_0_0;
assign O_6_0 = I_6_0_0;
assign O_7_0 = I_7_0_0;
assign O_8_0 = I_8_0_0;
assign valid_down = valid_up;
endmodule

module Partition_S_no3_ni3_tElSSeq_1_Int__vTrue (input CLK, input [7:0] I_0_0, input [7:0] I_1_0, input [7:0] I_2_0, input [7:0] I_3_0, input [7:0] I_4_0, input [7:0] I_5_0, input [7:0] I_6_0, input [7:0] I_7_0, input [7:0] I_8_0, output [7:0] O_0_0_0, output [7:0] O_0_1_0, output [7:0] O_0_2_0, output [7:0] O_1_0_0, output [7:0] O_1_1_0, output [7:0] O_1_2_0, output [7:0] O_2_0_0, output [7:0] O_2_1_0, output [7:0] O_2_2_0, output valid_down, input valid_up);
assign O_0_0_0 = I_0_0;
assign O_0_1_0 = I_1_0;
assign O_0_2_0 = I_2_0;
assign O_1_0_0 = I_3_0;
assign O_1_1_0 = I_4_0;
assign O_1_2_0 = I_5_0;
assign O_2_0_0 = I_6_0;
assign O_2_1_0 = I_7_0;
assign O_2_2_0 = I_8_0;
assign valid_down = valid_up;
endmodule

module Partition_S_no3_ni1_tElSSeq_1_Int__vTrue (input CLK, input [7:0] I_0_0_0, input [7:0] I_1_0_0, input [7:0] I_2_0_0, output [7:0] O_0_0, output [7:0] O_1_0, output [7:0] O_2_0, output valid_down, input valid_up);
assign O_0_0 = I_0_0_0;
assign O_1_0 = I_1_0_0;
assign O_2_0 = I_2_0_0;
assign valid_down = valid_up;
endmodule

module NativeMapParallel_n9_unq3 (input [7:0] I_0_0_0, input [7:0] I_0_0_1, input [7:0] I_0_0_2, input [7:0] I_1_0_0, input [7:0] I_1_0_1, input [7:0] I_1_0_2, input [7:0] I_2_0_0, input [7:0] I_2_0_1, input [7:0] I_2_0_2, input [7:0] I_3_0_0, input [7:0] I_3_0_1, input [7:0] I_3_0_2, input [7:0] I_4_0_0, input [7:0] I_4_0_1, input [7:0] I_4_0_2, input [7:0] I_5_0_0, input [7:0] I_5_0_1, input [7:0] I_5_0_2, input [7:0] I_6_0_0, input [7:0] I_6_0_1, input [7:0] I_6_0_2, input [7:0] I_7_0_0, input [7:0] I_7_0_1, input [7:0] I_7_0_2, input [7:0] I_8_0_0, input [7:0] I_8_0_1, input [7:0] I_8_0_2, output [7:0] O_0_0, output [7:0] O_0_1, output [7:0] O_0_2, output [7:0] O_1_0, output [7:0] O_1_1, output [7:0] O_1_2, output [7:0] O_2_0, output [7:0] O_2_1, output [7:0] O_2_2, output [7:0] O_3_0, output [7:0] O_3_1, output [7:0] O_3_2, output [7:0] O_4_0, output [7:0] O_4_1, output [7:0] O_4_2, output [7:0] O_5_0, output [7:0] O_5_1, output [7:0] O_5_2, output [7:0] O_6_0, output [7:0] O_6_1, output [7:0] O_6_2, output [7:0] O_7_0, output [7:0] O_7_1, output [7:0] O_7_2, output [7:0] O_8_0, output [7:0] O_8_1, output [7:0] O_8_2, output valid_down, input valid_up);
wire [7:0] Remove_1_S_inst0_O_0;
wire [7:0] Remove_1_S_inst0_O_1;
wire [7:0] Remove_1_S_inst0_O_2;
wire Remove_1_S_inst0_valid_down;
wire [7:0] Remove_1_S_inst1_O_0;
wire [7:0] Remove_1_S_inst1_O_1;
wire [7:0] Remove_1_S_inst1_O_2;
wire Remove_1_S_inst1_valid_down;
wire [7:0] Remove_1_S_inst2_O_0;
wire [7:0] Remove_1_S_inst2_O_1;
wire [7:0] Remove_1_S_inst2_O_2;
wire Remove_1_S_inst2_valid_down;
wire [7:0] Remove_1_S_inst3_O_0;
wire [7:0] Remove_1_S_inst3_O_1;
wire [7:0] Remove_1_S_inst3_O_2;
wire Remove_1_S_inst3_valid_down;
wire [7:0] Remove_1_S_inst4_O_0;
wire [7:0] Remove_1_S_inst4_O_1;
wire [7:0] Remove_1_S_inst4_O_2;
wire Remove_1_S_inst4_valid_down;
wire [7:0] Remove_1_S_inst5_O_0;
wire [7:0] Remove_1_S_inst5_O_1;
wire [7:0] Remove_1_S_inst5_O_2;
wire Remove_1_S_inst5_valid_down;
wire [7:0] Remove_1_S_inst6_O_0;
wire [7:0] Remove_1_S_inst6_O_1;
wire [7:0] Remove_1_S_inst6_O_2;
wire Remove_1_S_inst6_valid_down;
wire [7:0] Remove_1_S_inst7_O_0;
wire [7:0] Remove_1_S_inst7_O_1;
wire [7:0] Remove_1_S_inst7_O_2;
wire Remove_1_S_inst7_valid_down;
wire [7:0] Remove_1_S_inst8_O_0;
wire [7:0] Remove_1_S_inst8_O_1;
wire [7:0] Remove_1_S_inst8_O_2;
wire Remove_1_S_inst8_valid_down;
wire and_inst0_out;
wire and_inst1_out;
wire and_inst2_out;
wire and_inst3_out;
wire and_inst4_out;
wire and_inst5_out;
wire and_inst6_out;
wire and_inst7_out;
Remove_1_S Remove_1_S_inst0(.I_0_0(I_0_0_0), .I_0_1(I_0_0_1), .I_0_2(I_0_0_2), .O_0(Remove_1_S_inst0_O_0), .O_1(Remove_1_S_inst0_O_1), .O_2(Remove_1_S_inst0_O_2), .valid_down(Remove_1_S_inst0_valid_down), .valid_up(valid_up));
Remove_1_S Remove_1_S_inst1(.I_0_0(I_1_0_0), .I_0_1(I_1_0_1), .I_0_2(I_1_0_2), .O_0(Remove_1_S_inst1_O_0), .O_1(Remove_1_S_inst1_O_1), .O_2(Remove_1_S_inst1_O_2), .valid_down(Remove_1_S_inst1_valid_down), .valid_up(valid_up));
Remove_1_S Remove_1_S_inst2(.I_0_0(I_2_0_0), .I_0_1(I_2_0_1), .I_0_2(I_2_0_2), .O_0(Remove_1_S_inst2_O_0), .O_1(Remove_1_S_inst2_O_1), .O_2(Remove_1_S_inst2_O_2), .valid_down(Remove_1_S_inst2_valid_down), .valid_up(valid_up));
Remove_1_S Remove_1_S_inst3(.I_0_0(I_3_0_0), .I_0_1(I_3_0_1), .I_0_2(I_3_0_2), .O_0(Remove_1_S_inst3_O_0), .O_1(Remove_1_S_inst3_O_1), .O_2(Remove_1_S_inst3_O_2), .valid_down(Remove_1_S_inst3_valid_down), .valid_up(valid_up));
Remove_1_S Remove_1_S_inst4(.I_0_0(I_4_0_0), .I_0_1(I_4_0_1), .I_0_2(I_4_0_2), .O_0(Remove_1_S_inst4_O_0), .O_1(Remove_1_S_inst4_O_1), .O_2(Remove_1_S_inst4_O_2), .valid_down(Remove_1_S_inst4_valid_down), .valid_up(valid_up));
Remove_1_S Remove_1_S_inst5(.I_0_0(I_5_0_0), .I_0_1(I_5_0_1), .I_0_2(I_5_0_2), .O_0(Remove_1_S_inst5_O_0), .O_1(Remove_1_S_inst5_O_1), .O_2(Remove_1_S_inst5_O_2), .valid_down(Remove_1_S_inst5_valid_down), .valid_up(valid_up));
Remove_1_S Remove_1_S_inst6(.I_0_0(I_6_0_0), .I_0_1(I_6_0_1), .I_0_2(I_6_0_2), .O_0(Remove_1_S_inst6_O_0), .O_1(Remove_1_S_inst6_O_1), .O_2(Remove_1_S_inst6_O_2), .valid_down(Remove_1_S_inst6_valid_down), .valid_up(valid_up));
Remove_1_S Remove_1_S_inst7(.I_0_0(I_7_0_0), .I_0_1(I_7_0_1), .I_0_2(I_7_0_2), .O_0(Remove_1_S_inst7_O_0), .O_1(Remove_1_S_inst7_O_1), .O_2(Remove_1_S_inst7_O_2), .valid_down(Remove_1_S_inst7_valid_down), .valid_up(valid_up));
Remove_1_S Remove_1_S_inst8(.I_0_0(I_8_0_0), .I_0_1(I_8_0_1), .I_0_2(I_8_0_2), .O_0(Remove_1_S_inst8_O_0), .O_1(Remove_1_S_inst8_O_1), .O_2(Remove_1_S_inst8_O_2), .valid_down(Remove_1_S_inst8_valid_down), .valid_up(valid_up));
corebit_and and_inst0(.in0(Remove_1_S_inst0_valid_down), .in1(Remove_1_S_inst1_valid_down), .out(and_inst0_out));
corebit_and and_inst1(.in0(and_inst0_out), .in1(Remove_1_S_inst2_valid_down), .out(and_inst1_out));
corebit_and and_inst2(.in0(and_inst1_out), .in1(Remove_1_S_inst3_valid_down), .out(and_inst2_out));
corebit_and and_inst3(.in0(and_inst2_out), .in1(Remove_1_S_inst4_valid_down), .out(and_inst3_out));
corebit_and and_inst4(.in0(and_inst3_out), .in1(Remove_1_S_inst5_valid_down), .out(and_inst4_out));
corebit_and and_inst5(.in0(and_inst4_out), .in1(Remove_1_S_inst6_valid_down), .out(and_inst5_out));
corebit_and and_inst6(.in0(and_inst5_out), .in1(Remove_1_S_inst7_valid_down), .out(and_inst6_out));
corebit_and and_inst7(.in0(and_inst6_out), .in1(Remove_1_S_inst8_valid_down), .out(and_inst7_out));
assign O_0_0 = Remove_1_S_inst0_O_0;
assign O_0_1 = Remove_1_S_inst0_O_1;
assign O_0_2 = Remove_1_S_inst0_O_2;
assign O_1_0 = Remove_1_S_inst1_O_0;
assign O_1_1 = Remove_1_S_inst1_O_1;
assign O_1_2 = Remove_1_S_inst1_O_2;
assign O_2_0 = Remove_1_S_inst2_O_0;
assign O_2_1 = Remove_1_S_inst2_O_1;
assign O_2_2 = Remove_1_S_inst2_O_2;
assign O_3_0 = Remove_1_S_inst3_O_0;
assign O_3_1 = Remove_1_S_inst3_O_1;
assign O_3_2 = Remove_1_S_inst3_O_2;
assign O_4_0 = Remove_1_S_inst4_O_0;
assign O_4_1 = Remove_1_S_inst4_O_1;
assign O_4_2 = Remove_1_S_inst4_O_2;
assign O_5_0 = Remove_1_S_inst5_O_0;
assign O_5_1 = Remove_1_S_inst5_O_1;
assign O_5_2 = Remove_1_S_inst5_O_2;
assign O_6_0 = Remove_1_S_inst6_O_0;
assign O_6_1 = Remove_1_S_inst6_O_1;
assign O_6_2 = Remove_1_S_inst6_O_2;
assign O_7_0 = Remove_1_S_inst7_O_0;
assign O_7_1 = Remove_1_S_inst7_O_1;
assign O_7_2 = Remove_1_S_inst7_O_2;
assign O_8_0 = Remove_1_S_inst8_O_0;
assign O_8_1 = Remove_1_S_inst8_O_1;
assign O_8_2 = Remove_1_S_inst8_O_2;
assign valid_down = and_inst7_out;
endmodule

module NativeMapParallel_n3 (input [7:0] I0_0, input [7:0] I0_1, input [7:0] I0_2, input [7:0] I1_0, input [7:0] I1_1, input [7:0] I1_2, output [7:0] O_0__0, output [7:0] O_0__1, output [7:0] O_1__0, output [7:0] O_1__1, output [7:0] O_2__0, output [7:0] O_2__1, output valid_down, input valid_up);
wire and_inst0_out;
wire and_inst1_out;
wire [7:0] atomTupleCreator_t0Int_t1Int_inst0_O__0;
wire [7:0] atomTupleCreator_t0Int_t1Int_inst0_O__1;
wire atomTupleCreator_t0Int_t1Int_inst0_valid_down;
wire [7:0] atomTupleCreator_t0Int_t1Int_inst1_O__0;
wire [7:0] atomTupleCreator_t0Int_t1Int_inst1_O__1;
wire atomTupleCreator_t0Int_t1Int_inst1_valid_down;
wire [7:0] atomTupleCreator_t0Int_t1Int_inst2_O__0;
wire [7:0] atomTupleCreator_t0Int_t1Int_inst2_O__1;
wire atomTupleCreator_t0Int_t1Int_inst2_valid_down;
corebit_and and_inst0(.in0(atomTupleCreator_t0Int_t1Int_inst0_valid_down), .in1(atomTupleCreator_t0Int_t1Int_inst1_valid_down), .out(and_inst0_out));
corebit_and and_inst1(.in0(and_inst0_out), .in1(atomTupleCreator_t0Int_t1Int_inst2_valid_down), .out(and_inst1_out));
atomTupleCreator_t0Int_t1Int atomTupleCreator_t0Int_t1Int_inst0(.I0(I0_0), .I1(I1_0), .O__0(atomTupleCreator_t0Int_t1Int_inst0_O__0), .O__1(atomTupleCreator_t0Int_t1Int_inst0_O__1), .valid_down(atomTupleCreator_t0Int_t1Int_inst0_valid_down), .valid_up(valid_up));
atomTupleCreator_t0Int_t1Int atomTupleCreator_t0Int_t1Int_inst1(.I0(I0_1), .I1(I1_1), .O__0(atomTupleCreator_t0Int_t1Int_inst1_O__0), .O__1(atomTupleCreator_t0Int_t1Int_inst1_O__1), .valid_down(atomTupleCreator_t0Int_t1Int_inst1_valid_down), .valid_up(valid_up));
atomTupleCreator_t0Int_t1Int atomTupleCreator_t0Int_t1Int_inst2(.I0(I0_2), .I1(I1_2), .O__0(atomTupleCreator_t0Int_t1Int_inst2_O__0), .O__1(atomTupleCreator_t0Int_t1Int_inst2_O__1), .valid_down(atomTupleCreator_t0Int_t1Int_inst2_valid_down), .valid_up(valid_up));
assign O_0__0 = atomTupleCreator_t0Int_t1Int_inst0_O__0;
assign O_0__1 = atomTupleCreator_t0Int_t1Int_inst0_O__1;
assign O_1__0 = atomTupleCreator_t0Int_t1Int_inst1_O__0;
assign O_1__1 = atomTupleCreator_t0Int_t1Int_inst1_O__1;
assign O_2__0 = atomTupleCreator_t0Int_t1Int_inst2_O__0;
assign O_2__1 = atomTupleCreator_t0Int_t1Int_inst2_O__1;
assign valid_down = and_inst1_out;
endmodule

module NativeMapParallel_n27_unq2 (input [7:0] I_0_0_0, input [7:0] I_0_0_1, input [7:0] I_0_0_2, input [7:0] I_10_0_0, input [7:0] I_10_0_1, input [7:0] I_10_0_2, input [7:0] I_11_0_0, input [7:0] I_11_0_1, input [7:0] I_11_0_2, input [7:0] I_12_0_0, input [7:0] I_12_0_1, input [7:0] I_12_0_2, input [7:0] I_13_0_0, input [7:0] I_13_0_1, input [7:0] I_13_0_2, input [7:0] I_14_0_0, input [7:0] I_14_0_1, input [7:0] I_14_0_2, input [7:0] I_15_0_0, input [7:0] I_15_0_1, input [7:0] I_15_0_2, input [7:0] I_16_0_0, input [7:0] I_16_0_1, input [7:0] I_16_0_2, input [7:0] I_17_0_0, input [7:0] I_17_0_1, input [7:0] I_17_0_2, input [7:0] I_18_0_0, input [7:0] I_18_0_1, input [7:0] I_18_0_2, input [7:0] I_19_0_0, input [7:0] I_19_0_1, input [7:0] I_19_0_2, input [7:0] I_1_0_0, input [7:0] I_1_0_1, input [7:0] I_1_0_2, input [7:0] I_20_0_0, input [7:0] I_20_0_1, input [7:0] I_20_0_2, input [7:0] I_21_0_0, input [7:0] I_21_0_1, input [7:0] I_21_0_2, input [7:0] I_22_0_0, input [7:0] I_22_0_1, input [7:0] I_22_0_2, input [7:0] I_23_0_0, input [7:0] I_23_0_1, input [7:0] I_23_0_2, input [7:0] I_24_0_0, input [7:0] I_24_0_1, input [7:0] I_24_0_2, input [7:0] I_25_0_0, input [7:0] I_25_0_1, input [7:0] I_25_0_2, input [7:0] I_26_0_0, input [7:0] I_26_0_1, input [7:0] I_26_0_2, input [7:0] I_2_0_0, input [7:0] I_2_0_1, input [7:0] I_2_0_2, input [7:0] I_3_0_0, input [7:0] I_3_0_1, input [7:0] I_3_0_2, input [7:0] I_4_0_0, input [7:0] I_4_0_1, input [7:0] I_4_0_2, input [7:0] I_5_0_0, input [7:0] I_5_0_1, input [7:0] I_5_0_2, input [7:0] I_6_0_0, input [7:0] I_6_0_1, input [7:0] I_6_0_2, input [7:0] I_7_0_0, input [7:0] I_7_0_1, input [7:0] I_7_0_2, input [7:0] I_8_0_0, input [7:0] I_8_0_1, input [7:0] I_8_0_2, input [7:0] I_9_0_0, input [7:0] I_9_0_1, input [7:0] I_9_0_2, output [7:0] O_0_0, output [7:0] O_0_1, output [7:0] O_0_2, output [7:0] O_10_0, output [7:0] O_10_1, output [7:0] O_10_2, output [7:0] O_11_0, output [7:0] O_11_1, output [7:0] O_11_2, output [7:0] O_12_0, output [7:0] O_12_1, output [7:0] O_12_2, output [7:0] O_13_0, output [7:0] O_13_1, output [7:0] O_13_2, output [7:0] O_14_0, output [7:0] O_14_1, output [7:0] O_14_2, output [7:0] O_15_0, output [7:0] O_15_1, output [7:0] O_15_2, output [7:0] O_16_0, output [7:0] O_16_1, output [7:0] O_16_2, output [7:0] O_17_0, output [7:0] O_17_1, output [7:0] O_17_2, output [7:0] O_18_0, output [7:0] O_18_1, output [7:0] O_18_2, output [7:0] O_19_0, output [7:0] O_19_1, output [7:0] O_19_2, output [7:0] O_1_0, output [7:0] O_1_1, output [7:0] O_1_2, output [7:0] O_20_0, output [7:0] O_20_1, output [7:0] O_20_2, output [7:0] O_21_0, output [7:0] O_21_1, output [7:0] O_21_2, output [7:0] O_22_0, output [7:0] O_22_1, output [7:0] O_22_2, output [7:0] O_23_0, output [7:0] O_23_1, output [7:0] O_23_2, output [7:0] O_24_0, output [7:0] O_24_1, output [7:0] O_24_2, output [7:0] O_25_0, output [7:0] O_25_1, output [7:0] O_25_2, output [7:0] O_26_0, output [7:0] O_26_1, output [7:0] O_26_2, output [7:0] O_2_0, output [7:0] O_2_1, output [7:0] O_2_2, output [7:0] O_3_0, output [7:0] O_3_1, output [7:0] O_3_2, output [7:0] O_4_0, output [7:0] O_4_1, output [7:0] O_4_2, output [7:0] O_5_0, output [7:0] O_5_1, output [7:0] O_5_2, output [7:0] O_6_0, output [7:0] O_6_1, output [7:0] O_6_2, output [7:0] O_7_0, output [7:0] O_7_1, output [7:0] O_7_2, output [7:0] O_8_0, output [7:0] O_8_1, output [7:0] O_8_2, output [7:0] O_9_0, output [7:0] O_9_1, output [7:0] O_9_2, output valid_down, input valid_up);
wire [7:0] Remove_1_S_inst0_O_0;
wire [7:0] Remove_1_S_inst0_O_1;
wire [7:0] Remove_1_S_inst0_O_2;
wire Remove_1_S_inst0_valid_down;
wire [7:0] Remove_1_S_inst1_O_0;
wire [7:0] Remove_1_S_inst1_O_1;
wire [7:0] Remove_1_S_inst1_O_2;
wire Remove_1_S_inst1_valid_down;
wire [7:0] Remove_1_S_inst10_O_0;
wire [7:0] Remove_1_S_inst10_O_1;
wire [7:0] Remove_1_S_inst10_O_2;
wire Remove_1_S_inst10_valid_down;
wire [7:0] Remove_1_S_inst11_O_0;
wire [7:0] Remove_1_S_inst11_O_1;
wire [7:0] Remove_1_S_inst11_O_2;
wire Remove_1_S_inst11_valid_down;
wire [7:0] Remove_1_S_inst12_O_0;
wire [7:0] Remove_1_S_inst12_O_1;
wire [7:0] Remove_1_S_inst12_O_2;
wire Remove_1_S_inst12_valid_down;
wire [7:0] Remove_1_S_inst13_O_0;
wire [7:0] Remove_1_S_inst13_O_1;
wire [7:0] Remove_1_S_inst13_O_2;
wire Remove_1_S_inst13_valid_down;
wire [7:0] Remove_1_S_inst14_O_0;
wire [7:0] Remove_1_S_inst14_O_1;
wire [7:0] Remove_1_S_inst14_O_2;
wire Remove_1_S_inst14_valid_down;
wire [7:0] Remove_1_S_inst15_O_0;
wire [7:0] Remove_1_S_inst15_O_1;
wire [7:0] Remove_1_S_inst15_O_2;
wire Remove_1_S_inst15_valid_down;
wire [7:0] Remove_1_S_inst16_O_0;
wire [7:0] Remove_1_S_inst16_O_1;
wire [7:0] Remove_1_S_inst16_O_2;
wire Remove_1_S_inst16_valid_down;
wire [7:0] Remove_1_S_inst17_O_0;
wire [7:0] Remove_1_S_inst17_O_1;
wire [7:0] Remove_1_S_inst17_O_2;
wire Remove_1_S_inst17_valid_down;
wire [7:0] Remove_1_S_inst18_O_0;
wire [7:0] Remove_1_S_inst18_O_1;
wire [7:0] Remove_1_S_inst18_O_2;
wire Remove_1_S_inst18_valid_down;
wire [7:0] Remove_1_S_inst19_O_0;
wire [7:0] Remove_1_S_inst19_O_1;
wire [7:0] Remove_1_S_inst19_O_2;
wire Remove_1_S_inst19_valid_down;
wire [7:0] Remove_1_S_inst2_O_0;
wire [7:0] Remove_1_S_inst2_O_1;
wire [7:0] Remove_1_S_inst2_O_2;
wire Remove_1_S_inst2_valid_down;
wire [7:0] Remove_1_S_inst20_O_0;
wire [7:0] Remove_1_S_inst20_O_1;
wire [7:0] Remove_1_S_inst20_O_2;
wire Remove_1_S_inst20_valid_down;
wire [7:0] Remove_1_S_inst21_O_0;
wire [7:0] Remove_1_S_inst21_O_1;
wire [7:0] Remove_1_S_inst21_O_2;
wire Remove_1_S_inst21_valid_down;
wire [7:0] Remove_1_S_inst22_O_0;
wire [7:0] Remove_1_S_inst22_O_1;
wire [7:0] Remove_1_S_inst22_O_2;
wire Remove_1_S_inst22_valid_down;
wire [7:0] Remove_1_S_inst23_O_0;
wire [7:0] Remove_1_S_inst23_O_1;
wire [7:0] Remove_1_S_inst23_O_2;
wire Remove_1_S_inst23_valid_down;
wire [7:0] Remove_1_S_inst24_O_0;
wire [7:0] Remove_1_S_inst24_O_1;
wire [7:0] Remove_1_S_inst24_O_2;
wire Remove_1_S_inst24_valid_down;
wire [7:0] Remove_1_S_inst25_O_0;
wire [7:0] Remove_1_S_inst25_O_1;
wire [7:0] Remove_1_S_inst25_O_2;
wire Remove_1_S_inst25_valid_down;
wire [7:0] Remove_1_S_inst26_O_0;
wire [7:0] Remove_1_S_inst26_O_1;
wire [7:0] Remove_1_S_inst26_O_2;
wire Remove_1_S_inst26_valid_down;
wire [7:0] Remove_1_S_inst3_O_0;
wire [7:0] Remove_1_S_inst3_O_1;
wire [7:0] Remove_1_S_inst3_O_2;
wire Remove_1_S_inst3_valid_down;
wire [7:0] Remove_1_S_inst4_O_0;
wire [7:0] Remove_1_S_inst4_O_1;
wire [7:0] Remove_1_S_inst4_O_2;
wire Remove_1_S_inst4_valid_down;
wire [7:0] Remove_1_S_inst5_O_0;
wire [7:0] Remove_1_S_inst5_O_1;
wire [7:0] Remove_1_S_inst5_O_2;
wire Remove_1_S_inst5_valid_down;
wire [7:0] Remove_1_S_inst6_O_0;
wire [7:0] Remove_1_S_inst6_O_1;
wire [7:0] Remove_1_S_inst6_O_2;
wire Remove_1_S_inst6_valid_down;
wire [7:0] Remove_1_S_inst7_O_0;
wire [7:0] Remove_1_S_inst7_O_1;
wire [7:0] Remove_1_S_inst7_O_2;
wire Remove_1_S_inst7_valid_down;
wire [7:0] Remove_1_S_inst8_O_0;
wire [7:0] Remove_1_S_inst8_O_1;
wire [7:0] Remove_1_S_inst8_O_2;
wire Remove_1_S_inst8_valid_down;
wire [7:0] Remove_1_S_inst9_O_0;
wire [7:0] Remove_1_S_inst9_O_1;
wire [7:0] Remove_1_S_inst9_O_2;
wire Remove_1_S_inst9_valid_down;
wire and_inst0_out;
wire and_inst1_out;
wire and_inst10_out;
wire and_inst11_out;
wire and_inst12_out;
wire and_inst13_out;
wire and_inst14_out;
wire and_inst15_out;
wire and_inst16_out;
wire and_inst17_out;
wire and_inst18_out;
wire and_inst19_out;
wire and_inst2_out;
wire and_inst20_out;
wire and_inst21_out;
wire and_inst22_out;
wire and_inst23_out;
wire and_inst24_out;
wire and_inst25_out;
wire and_inst3_out;
wire and_inst4_out;
wire and_inst5_out;
wire and_inst6_out;
wire and_inst7_out;
wire and_inst8_out;
wire and_inst9_out;
Remove_1_S Remove_1_S_inst0(.I_0_0(I_0_0_0), .I_0_1(I_0_0_1), .I_0_2(I_0_0_2), .O_0(Remove_1_S_inst0_O_0), .O_1(Remove_1_S_inst0_O_1), .O_2(Remove_1_S_inst0_O_2), .valid_down(Remove_1_S_inst0_valid_down), .valid_up(valid_up));
Remove_1_S Remove_1_S_inst1(.I_0_0(I_1_0_0), .I_0_1(I_1_0_1), .I_0_2(I_1_0_2), .O_0(Remove_1_S_inst1_O_0), .O_1(Remove_1_S_inst1_O_1), .O_2(Remove_1_S_inst1_O_2), .valid_down(Remove_1_S_inst1_valid_down), .valid_up(valid_up));
Remove_1_S Remove_1_S_inst10(.I_0_0(I_10_0_0), .I_0_1(I_10_0_1), .I_0_2(I_10_0_2), .O_0(Remove_1_S_inst10_O_0), .O_1(Remove_1_S_inst10_O_1), .O_2(Remove_1_S_inst10_O_2), .valid_down(Remove_1_S_inst10_valid_down), .valid_up(valid_up));
Remove_1_S Remove_1_S_inst11(.I_0_0(I_11_0_0), .I_0_1(I_11_0_1), .I_0_2(I_11_0_2), .O_0(Remove_1_S_inst11_O_0), .O_1(Remove_1_S_inst11_O_1), .O_2(Remove_1_S_inst11_O_2), .valid_down(Remove_1_S_inst11_valid_down), .valid_up(valid_up));
Remove_1_S Remove_1_S_inst12(.I_0_0(I_12_0_0), .I_0_1(I_12_0_1), .I_0_2(I_12_0_2), .O_0(Remove_1_S_inst12_O_0), .O_1(Remove_1_S_inst12_O_1), .O_2(Remove_1_S_inst12_O_2), .valid_down(Remove_1_S_inst12_valid_down), .valid_up(valid_up));
Remove_1_S Remove_1_S_inst13(.I_0_0(I_13_0_0), .I_0_1(I_13_0_1), .I_0_2(I_13_0_2), .O_0(Remove_1_S_inst13_O_0), .O_1(Remove_1_S_inst13_O_1), .O_2(Remove_1_S_inst13_O_2), .valid_down(Remove_1_S_inst13_valid_down), .valid_up(valid_up));
Remove_1_S Remove_1_S_inst14(.I_0_0(I_14_0_0), .I_0_1(I_14_0_1), .I_0_2(I_14_0_2), .O_0(Remove_1_S_inst14_O_0), .O_1(Remove_1_S_inst14_O_1), .O_2(Remove_1_S_inst14_O_2), .valid_down(Remove_1_S_inst14_valid_down), .valid_up(valid_up));
Remove_1_S Remove_1_S_inst15(.I_0_0(I_15_0_0), .I_0_1(I_15_0_1), .I_0_2(I_15_0_2), .O_0(Remove_1_S_inst15_O_0), .O_1(Remove_1_S_inst15_O_1), .O_2(Remove_1_S_inst15_O_2), .valid_down(Remove_1_S_inst15_valid_down), .valid_up(valid_up));
Remove_1_S Remove_1_S_inst16(.I_0_0(I_16_0_0), .I_0_1(I_16_0_1), .I_0_2(I_16_0_2), .O_0(Remove_1_S_inst16_O_0), .O_1(Remove_1_S_inst16_O_1), .O_2(Remove_1_S_inst16_O_2), .valid_down(Remove_1_S_inst16_valid_down), .valid_up(valid_up));
Remove_1_S Remove_1_S_inst17(.I_0_0(I_17_0_0), .I_0_1(I_17_0_1), .I_0_2(I_17_0_2), .O_0(Remove_1_S_inst17_O_0), .O_1(Remove_1_S_inst17_O_1), .O_2(Remove_1_S_inst17_O_2), .valid_down(Remove_1_S_inst17_valid_down), .valid_up(valid_up));
Remove_1_S Remove_1_S_inst18(.I_0_0(I_18_0_0), .I_0_1(I_18_0_1), .I_0_2(I_18_0_2), .O_0(Remove_1_S_inst18_O_0), .O_1(Remove_1_S_inst18_O_1), .O_2(Remove_1_S_inst18_O_2), .valid_down(Remove_1_S_inst18_valid_down), .valid_up(valid_up));
Remove_1_S Remove_1_S_inst19(.I_0_0(I_19_0_0), .I_0_1(I_19_0_1), .I_0_2(I_19_0_2), .O_0(Remove_1_S_inst19_O_0), .O_1(Remove_1_S_inst19_O_1), .O_2(Remove_1_S_inst19_O_2), .valid_down(Remove_1_S_inst19_valid_down), .valid_up(valid_up));
Remove_1_S Remove_1_S_inst2(.I_0_0(I_2_0_0), .I_0_1(I_2_0_1), .I_0_2(I_2_0_2), .O_0(Remove_1_S_inst2_O_0), .O_1(Remove_1_S_inst2_O_1), .O_2(Remove_1_S_inst2_O_2), .valid_down(Remove_1_S_inst2_valid_down), .valid_up(valid_up));
Remove_1_S Remove_1_S_inst20(.I_0_0(I_20_0_0), .I_0_1(I_20_0_1), .I_0_2(I_20_0_2), .O_0(Remove_1_S_inst20_O_0), .O_1(Remove_1_S_inst20_O_1), .O_2(Remove_1_S_inst20_O_2), .valid_down(Remove_1_S_inst20_valid_down), .valid_up(valid_up));
Remove_1_S Remove_1_S_inst21(.I_0_0(I_21_0_0), .I_0_1(I_21_0_1), .I_0_2(I_21_0_2), .O_0(Remove_1_S_inst21_O_0), .O_1(Remove_1_S_inst21_O_1), .O_2(Remove_1_S_inst21_O_2), .valid_down(Remove_1_S_inst21_valid_down), .valid_up(valid_up));
Remove_1_S Remove_1_S_inst22(.I_0_0(I_22_0_0), .I_0_1(I_22_0_1), .I_0_2(I_22_0_2), .O_0(Remove_1_S_inst22_O_0), .O_1(Remove_1_S_inst22_O_1), .O_2(Remove_1_S_inst22_O_2), .valid_down(Remove_1_S_inst22_valid_down), .valid_up(valid_up));
Remove_1_S Remove_1_S_inst23(.I_0_0(I_23_0_0), .I_0_1(I_23_0_1), .I_0_2(I_23_0_2), .O_0(Remove_1_S_inst23_O_0), .O_1(Remove_1_S_inst23_O_1), .O_2(Remove_1_S_inst23_O_2), .valid_down(Remove_1_S_inst23_valid_down), .valid_up(valid_up));
Remove_1_S Remove_1_S_inst24(.I_0_0(I_24_0_0), .I_0_1(I_24_0_1), .I_0_2(I_24_0_2), .O_0(Remove_1_S_inst24_O_0), .O_1(Remove_1_S_inst24_O_1), .O_2(Remove_1_S_inst24_O_2), .valid_down(Remove_1_S_inst24_valid_down), .valid_up(valid_up));
Remove_1_S Remove_1_S_inst25(.I_0_0(I_25_0_0), .I_0_1(I_25_0_1), .I_0_2(I_25_0_2), .O_0(Remove_1_S_inst25_O_0), .O_1(Remove_1_S_inst25_O_1), .O_2(Remove_1_S_inst25_O_2), .valid_down(Remove_1_S_inst25_valid_down), .valid_up(valid_up));
Remove_1_S Remove_1_S_inst26(.I_0_0(I_26_0_0), .I_0_1(I_26_0_1), .I_0_2(I_26_0_2), .O_0(Remove_1_S_inst26_O_0), .O_1(Remove_1_S_inst26_O_1), .O_2(Remove_1_S_inst26_O_2), .valid_down(Remove_1_S_inst26_valid_down), .valid_up(valid_up));
Remove_1_S Remove_1_S_inst3(.I_0_0(I_3_0_0), .I_0_1(I_3_0_1), .I_0_2(I_3_0_2), .O_0(Remove_1_S_inst3_O_0), .O_1(Remove_1_S_inst3_O_1), .O_2(Remove_1_S_inst3_O_2), .valid_down(Remove_1_S_inst3_valid_down), .valid_up(valid_up));
Remove_1_S Remove_1_S_inst4(.I_0_0(I_4_0_0), .I_0_1(I_4_0_1), .I_0_2(I_4_0_2), .O_0(Remove_1_S_inst4_O_0), .O_1(Remove_1_S_inst4_O_1), .O_2(Remove_1_S_inst4_O_2), .valid_down(Remove_1_S_inst4_valid_down), .valid_up(valid_up));
Remove_1_S Remove_1_S_inst5(.I_0_0(I_5_0_0), .I_0_1(I_5_0_1), .I_0_2(I_5_0_2), .O_0(Remove_1_S_inst5_O_0), .O_1(Remove_1_S_inst5_O_1), .O_2(Remove_1_S_inst5_O_2), .valid_down(Remove_1_S_inst5_valid_down), .valid_up(valid_up));
Remove_1_S Remove_1_S_inst6(.I_0_0(I_6_0_0), .I_0_1(I_6_0_1), .I_0_2(I_6_0_2), .O_0(Remove_1_S_inst6_O_0), .O_1(Remove_1_S_inst6_O_1), .O_2(Remove_1_S_inst6_O_2), .valid_down(Remove_1_S_inst6_valid_down), .valid_up(valid_up));
Remove_1_S Remove_1_S_inst7(.I_0_0(I_7_0_0), .I_0_1(I_7_0_1), .I_0_2(I_7_0_2), .O_0(Remove_1_S_inst7_O_0), .O_1(Remove_1_S_inst7_O_1), .O_2(Remove_1_S_inst7_O_2), .valid_down(Remove_1_S_inst7_valid_down), .valid_up(valid_up));
Remove_1_S Remove_1_S_inst8(.I_0_0(I_8_0_0), .I_0_1(I_8_0_1), .I_0_2(I_8_0_2), .O_0(Remove_1_S_inst8_O_0), .O_1(Remove_1_S_inst8_O_1), .O_2(Remove_1_S_inst8_O_2), .valid_down(Remove_1_S_inst8_valid_down), .valid_up(valid_up));
Remove_1_S Remove_1_S_inst9(.I_0_0(I_9_0_0), .I_0_1(I_9_0_1), .I_0_2(I_9_0_2), .O_0(Remove_1_S_inst9_O_0), .O_1(Remove_1_S_inst9_O_1), .O_2(Remove_1_S_inst9_O_2), .valid_down(Remove_1_S_inst9_valid_down), .valid_up(valid_up));
corebit_and and_inst0(.in0(Remove_1_S_inst0_valid_down), .in1(Remove_1_S_inst1_valid_down), .out(and_inst0_out));
corebit_and and_inst1(.in0(and_inst0_out), .in1(Remove_1_S_inst2_valid_down), .out(and_inst1_out));
corebit_and and_inst10(.in0(and_inst9_out), .in1(Remove_1_S_inst11_valid_down), .out(and_inst10_out));
corebit_and and_inst11(.in0(and_inst10_out), .in1(Remove_1_S_inst12_valid_down), .out(and_inst11_out));
corebit_and and_inst12(.in0(and_inst11_out), .in1(Remove_1_S_inst13_valid_down), .out(and_inst12_out));
corebit_and and_inst13(.in0(and_inst12_out), .in1(Remove_1_S_inst14_valid_down), .out(and_inst13_out));
corebit_and and_inst14(.in0(and_inst13_out), .in1(Remove_1_S_inst15_valid_down), .out(and_inst14_out));
corebit_and and_inst15(.in0(and_inst14_out), .in1(Remove_1_S_inst16_valid_down), .out(and_inst15_out));
corebit_and and_inst16(.in0(and_inst15_out), .in1(Remove_1_S_inst17_valid_down), .out(and_inst16_out));
corebit_and and_inst17(.in0(and_inst16_out), .in1(Remove_1_S_inst18_valid_down), .out(and_inst17_out));
corebit_and and_inst18(.in0(and_inst17_out), .in1(Remove_1_S_inst19_valid_down), .out(and_inst18_out));
corebit_and and_inst19(.in0(and_inst18_out), .in1(Remove_1_S_inst20_valid_down), .out(and_inst19_out));
corebit_and and_inst2(.in0(and_inst1_out), .in1(Remove_1_S_inst3_valid_down), .out(and_inst2_out));
corebit_and and_inst20(.in0(and_inst19_out), .in1(Remove_1_S_inst21_valid_down), .out(and_inst20_out));
corebit_and and_inst21(.in0(and_inst20_out), .in1(Remove_1_S_inst22_valid_down), .out(and_inst21_out));
corebit_and and_inst22(.in0(and_inst21_out), .in1(Remove_1_S_inst23_valid_down), .out(and_inst22_out));
corebit_and and_inst23(.in0(and_inst22_out), .in1(Remove_1_S_inst24_valid_down), .out(and_inst23_out));
corebit_and and_inst24(.in0(and_inst23_out), .in1(Remove_1_S_inst25_valid_down), .out(and_inst24_out));
corebit_and and_inst25(.in0(and_inst24_out), .in1(Remove_1_S_inst26_valid_down), .out(and_inst25_out));
corebit_and and_inst3(.in0(and_inst2_out), .in1(Remove_1_S_inst4_valid_down), .out(and_inst3_out));
corebit_and and_inst4(.in0(and_inst3_out), .in1(Remove_1_S_inst5_valid_down), .out(and_inst4_out));
corebit_and and_inst5(.in0(and_inst4_out), .in1(Remove_1_S_inst6_valid_down), .out(and_inst5_out));
corebit_and and_inst6(.in0(and_inst5_out), .in1(Remove_1_S_inst7_valid_down), .out(and_inst6_out));
corebit_and and_inst7(.in0(and_inst6_out), .in1(Remove_1_S_inst8_valid_down), .out(and_inst7_out));
corebit_and and_inst8(.in0(and_inst7_out), .in1(Remove_1_S_inst9_valid_down), .out(and_inst8_out));
corebit_and and_inst9(.in0(and_inst8_out), .in1(Remove_1_S_inst10_valid_down), .out(and_inst9_out));
assign O_0_0 = Remove_1_S_inst0_O_0;
assign O_0_1 = Remove_1_S_inst0_O_1;
assign O_0_2 = Remove_1_S_inst0_O_2;
assign O_10_0 = Remove_1_S_inst10_O_0;
assign O_10_1 = Remove_1_S_inst10_O_1;
assign O_10_2 = Remove_1_S_inst10_O_2;
assign O_11_0 = Remove_1_S_inst11_O_0;
assign O_11_1 = Remove_1_S_inst11_O_1;
assign O_11_2 = Remove_1_S_inst11_O_2;
assign O_12_0 = Remove_1_S_inst12_O_0;
assign O_12_1 = Remove_1_S_inst12_O_1;
assign O_12_2 = Remove_1_S_inst12_O_2;
assign O_13_0 = Remove_1_S_inst13_O_0;
assign O_13_1 = Remove_1_S_inst13_O_1;
assign O_13_2 = Remove_1_S_inst13_O_2;
assign O_14_0 = Remove_1_S_inst14_O_0;
assign O_14_1 = Remove_1_S_inst14_O_1;
assign O_14_2 = Remove_1_S_inst14_O_2;
assign O_15_0 = Remove_1_S_inst15_O_0;
assign O_15_1 = Remove_1_S_inst15_O_1;
assign O_15_2 = Remove_1_S_inst15_O_2;
assign O_16_0 = Remove_1_S_inst16_O_0;
assign O_16_1 = Remove_1_S_inst16_O_1;
assign O_16_2 = Remove_1_S_inst16_O_2;
assign O_17_0 = Remove_1_S_inst17_O_0;
assign O_17_1 = Remove_1_S_inst17_O_1;
assign O_17_2 = Remove_1_S_inst17_O_2;
assign O_18_0 = Remove_1_S_inst18_O_0;
assign O_18_1 = Remove_1_S_inst18_O_1;
assign O_18_2 = Remove_1_S_inst18_O_2;
assign O_19_0 = Remove_1_S_inst19_O_0;
assign O_19_1 = Remove_1_S_inst19_O_1;
assign O_19_2 = Remove_1_S_inst19_O_2;
assign O_1_0 = Remove_1_S_inst1_O_0;
assign O_1_1 = Remove_1_S_inst1_O_1;
assign O_1_2 = Remove_1_S_inst1_O_2;
assign O_20_0 = Remove_1_S_inst20_O_0;
assign O_20_1 = Remove_1_S_inst20_O_1;
assign O_20_2 = Remove_1_S_inst20_O_2;
assign O_21_0 = Remove_1_S_inst21_O_0;
assign O_21_1 = Remove_1_S_inst21_O_1;
assign O_21_2 = Remove_1_S_inst21_O_2;
assign O_22_0 = Remove_1_S_inst22_O_0;
assign O_22_1 = Remove_1_S_inst22_O_1;
assign O_22_2 = Remove_1_S_inst22_O_2;
assign O_23_0 = Remove_1_S_inst23_O_0;
assign O_23_1 = Remove_1_S_inst23_O_1;
assign O_23_2 = Remove_1_S_inst23_O_2;
assign O_24_0 = Remove_1_S_inst24_O_0;
assign O_24_1 = Remove_1_S_inst24_O_1;
assign O_24_2 = Remove_1_S_inst24_O_2;
assign O_25_0 = Remove_1_S_inst25_O_0;
assign O_25_1 = Remove_1_S_inst25_O_1;
assign O_25_2 = Remove_1_S_inst25_O_2;
assign O_26_0 = Remove_1_S_inst26_O_0;
assign O_26_1 = Remove_1_S_inst26_O_1;
assign O_26_2 = Remove_1_S_inst26_O_2;
assign O_2_0 = Remove_1_S_inst2_O_0;
assign O_2_1 = Remove_1_S_inst2_O_1;
assign O_2_2 = Remove_1_S_inst2_O_2;
assign O_3_0 = Remove_1_S_inst3_O_0;
assign O_3_1 = Remove_1_S_inst3_O_1;
assign O_3_2 = Remove_1_S_inst3_O_2;
assign O_4_0 = Remove_1_S_inst4_O_0;
assign O_4_1 = Remove_1_S_inst4_O_1;
assign O_4_2 = Remove_1_S_inst4_O_2;
assign O_5_0 = Remove_1_S_inst5_O_0;
assign O_5_1 = Remove_1_S_inst5_O_1;
assign O_5_2 = Remove_1_S_inst5_O_2;
assign O_6_0 = Remove_1_S_inst6_O_0;
assign O_6_1 = Remove_1_S_inst6_O_1;
assign O_6_2 = Remove_1_S_inst6_O_2;
assign O_7_0 = Remove_1_S_inst7_O_0;
assign O_7_1 = Remove_1_S_inst7_O_1;
assign O_7_2 = Remove_1_S_inst7_O_2;
assign O_8_0 = Remove_1_S_inst8_O_0;
assign O_8_1 = Remove_1_S_inst8_O_1;
assign O_8_2 = Remove_1_S_inst8_O_2;
assign O_9_0 = Remove_1_S_inst9_O_0;
assign O_9_1 = Remove_1_S_inst9_O_1;
assign O_9_2 = Remove_1_S_inst9_O_2;
assign valid_down = and_inst25_out;
endmodule

module NativeMapParallel_n1_unq3 (input [7:0] I_0__0, input [7:0] I_0__1, output [7:0] O_0, output valid_down, input valid_up);
wire [7:0] RShift_Atom_inst0_O;
wire RShift_Atom_inst0_valid_down;
RShift_Atom RShift_Atom_inst0(.I__0(I_0__0), .I__1(I_0__1), .O(RShift_Atom_inst0_O), .valid_down(RShift_Atom_inst0_valid_down), .valid_up(valid_up));
assign O_0 = RShift_Atom_inst0_O;
assign valid_down = RShift_Atom_inst0_valid_down;
endmodule

module NativeMapParallel_n1_unq2 (input [7:0] I0_0, input [7:0] I1_0, output [7:0] O_0__0, output [7:0] O_0__1, output valid_down, input valid_up);
wire [7:0] atomTupleCreator_t0Int_t1Int_inst0_O__0;
wire [7:0] atomTupleCreator_t0Int_t1Int_inst0_O__1;
wire atomTupleCreator_t0Int_t1Int_inst0_valid_down;
atomTupleCreator_t0Int_t1Int atomTupleCreator_t0Int_t1Int_inst0(.I0(I0_0), .I1(I1_0), .O__0(atomTupleCreator_t0Int_t1Int_inst0_O__0), .O__1(atomTupleCreator_t0Int_t1Int_inst0_O__1), .valid_down(atomTupleCreator_t0Int_t1Int_inst0_valid_down), .valid_up(valid_up));
assign O_0__0 = atomTupleCreator_t0Int_t1Int_inst0_O__0;
assign O_0__1 = atomTupleCreator_t0Int_t1Int_inst0_O__1;
assign valid_down = atomTupleCreator_t0Int_t1Int_inst0_valid_down;
endmodule

module NativeMapParallel_n1_unq1 (input [7:0] I0_0_0, input [7:0] I0_0_1, input [7:0] I1_0, output [7:0] O_0_0, output [7:0] O_0_1, output [7:0] O_0_2, output valid_down, input valid_up);
wire [7:0] sseqTupleAppender_tInt_n2_inst0_O_0;
wire [7:0] sseqTupleAppender_tInt_n2_inst0_O_1;
wire [7:0] sseqTupleAppender_tInt_n2_inst0_O_2;
wire sseqTupleAppender_tInt_n2_inst0_valid_down;
sseqTupleAppender_tInt_n2 sseqTupleAppender_tInt_n2_inst0(.I0_0(I0_0_0), .I0_1(I0_0_1), .I1(I1_0), .O_0(sseqTupleAppender_tInt_n2_inst0_O_0), .O_1(sseqTupleAppender_tInt_n2_inst0_O_1), .O_2(sseqTupleAppender_tInt_n2_inst0_O_2), .valid_down(sseqTupleAppender_tInt_n2_inst0_valid_down), .valid_up(valid_up));
assign O_0_0 = sseqTupleAppender_tInt_n2_inst0_O_0;
assign O_0_1 = sseqTupleAppender_tInt_n2_inst0_O_1;
assign O_0_2 = sseqTupleAppender_tInt_n2_inst0_O_2;
assign valid_down = sseqTupleAppender_tInt_n2_inst0_valid_down;
endmodule

module NativeMapParallel_n9_unq2 (input [7:0] I0_0_0_0, input [7:0] I0_0_0_1, input [7:0] I0_1_0_0, input [7:0] I0_1_0_1, input [7:0] I0_2_0_0, input [7:0] I0_2_0_1, input [7:0] I0_3_0_0, input [7:0] I0_3_0_1, input [7:0] I0_4_0_0, input [7:0] I0_4_0_1, input [7:0] I0_5_0_0, input [7:0] I0_5_0_1, input [7:0] I0_6_0_0, input [7:0] I0_6_0_1, input [7:0] I0_7_0_0, input [7:0] I0_7_0_1, input [7:0] I0_8_0_0, input [7:0] I0_8_0_1, input [7:0] I1_0_0, input [7:0] I1_1_0, input [7:0] I1_2_0, input [7:0] I1_3_0, input [7:0] I1_4_0, input [7:0] I1_5_0, input [7:0] I1_6_0, input [7:0] I1_7_0, input [7:0] I1_8_0, output [7:0] O_0_0_0, output [7:0] O_0_0_1, output [7:0] O_0_0_2, output [7:0] O_1_0_0, output [7:0] O_1_0_1, output [7:0] O_1_0_2, output [7:0] O_2_0_0, output [7:0] O_2_0_1, output [7:0] O_2_0_2, output [7:0] O_3_0_0, output [7:0] O_3_0_1, output [7:0] O_3_0_2, output [7:0] O_4_0_0, output [7:0] O_4_0_1, output [7:0] O_4_0_2, output [7:0] O_5_0_0, output [7:0] O_5_0_1, output [7:0] O_5_0_2, output [7:0] O_6_0_0, output [7:0] O_6_0_1, output [7:0] O_6_0_2, output [7:0] O_7_0_0, output [7:0] O_7_0_1, output [7:0] O_7_0_2, output [7:0] O_8_0_0, output [7:0] O_8_0_1, output [7:0] O_8_0_2, output valid_down, input valid_up);
wire [7:0] NativeMapParallel_n1_inst0_O_0_0;
wire [7:0] NativeMapParallel_n1_inst0_O_0_1;
wire [7:0] NativeMapParallel_n1_inst0_O_0_2;
wire NativeMapParallel_n1_inst0_valid_down;
wire [7:0] NativeMapParallel_n1_inst1_O_0_0;
wire [7:0] NativeMapParallel_n1_inst1_O_0_1;
wire [7:0] NativeMapParallel_n1_inst1_O_0_2;
wire NativeMapParallel_n1_inst1_valid_down;
wire [7:0] NativeMapParallel_n1_inst2_O_0_0;
wire [7:0] NativeMapParallel_n1_inst2_O_0_1;
wire [7:0] NativeMapParallel_n1_inst2_O_0_2;
wire NativeMapParallel_n1_inst2_valid_down;
wire [7:0] NativeMapParallel_n1_inst3_O_0_0;
wire [7:0] NativeMapParallel_n1_inst3_O_0_1;
wire [7:0] NativeMapParallel_n1_inst3_O_0_2;
wire NativeMapParallel_n1_inst3_valid_down;
wire [7:0] NativeMapParallel_n1_inst4_O_0_0;
wire [7:0] NativeMapParallel_n1_inst4_O_0_1;
wire [7:0] NativeMapParallel_n1_inst4_O_0_2;
wire NativeMapParallel_n1_inst4_valid_down;
wire [7:0] NativeMapParallel_n1_inst5_O_0_0;
wire [7:0] NativeMapParallel_n1_inst5_O_0_1;
wire [7:0] NativeMapParallel_n1_inst5_O_0_2;
wire NativeMapParallel_n1_inst5_valid_down;
wire [7:0] NativeMapParallel_n1_inst6_O_0_0;
wire [7:0] NativeMapParallel_n1_inst6_O_0_1;
wire [7:0] NativeMapParallel_n1_inst6_O_0_2;
wire NativeMapParallel_n1_inst6_valid_down;
wire [7:0] NativeMapParallel_n1_inst7_O_0_0;
wire [7:0] NativeMapParallel_n1_inst7_O_0_1;
wire [7:0] NativeMapParallel_n1_inst7_O_0_2;
wire NativeMapParallel_n1_inst7_valid_down;
wire [7:0] NativeMapParallel_n1_inst8_O_0_0;
wire [7:0] NativeMapParallel_n1_inst8_O_0_1;
wire [7:0] NativeMapParallel_n1_inst8_O_0_2;
wire NativeMapParallel_n1_inst8_valid_down;
wire and_inst0_out;
wire and_inst1_out;
wire and_inst2_out;
wire and_inst3_out;
wire and_inst4_out;
wire and_inst5_out;
wire and_inst6_out;
wire and_inst7_out;
NativeMapParallel_n1_unq1 NativeMapParallel_n1_inst0(.I0_0_0(I0_0_0_0), .I0_0_1(I0_0_0_1), .I1_0(I1_0_0), .O_0_0(NativeMapParallel_n1_inst0_O_0_0), .O_0_1(NativeMapParallel_n1_inst0_O_0_1), .O_0_2(NativeMapParallel_n1_inst0_O_0_2), .valid_down(NativeMapParallel_n1_inst0_valid_down), .valid_up(valid_up));
NativeMapParallel_n1_unq1 NativeMapParallel_n1_inst1(.I0_0_0(I0_1_0_0), .I0_0_1(I0_1_0_1), .I1_0(I1_1_0), .O_0_0(NativeMapParallel_n1_inst1_O_0_0), .O_0_1(NativeMapParallel_n1_inst1_O_0_1), .O_0_2(NativeMapParallel_n1_inst1_O_0_2), .valid_down(NativeMapParallel_n1_inst1_valid_down), .valid_up(valid_up));
NativeMapParallel_n1_unq1 NativeMapParallel_n1_inst2(.I0_0_0(I0_2_0_0), .I0_0_1(I0_2_0_1), .I1_0(I1_2_0), .O_0_0(NativeMapParallel_n1_inst2_O_0_0), .O_0_1(NativeMapParallel_n1_inst2_O_0_1), .O_0_2(NativeMapParallel_n1_inst2_O_0_2), .valid_down(NativeMapParallel_n1_inst2_valid_down), .valid_up(valid_up));
NativeMapParallel_n1_unq1 NativeMapParallel_n1_inst3(.I0_0_0(I0_3_0_0), .I0_0_1(I0_3_0_1), .I1_0(I1_3_0), .O_0_0(NativeMapParallel_n1_inst3_O_0_0), .O_0_1(NativeMapParallel_n1_inst3_O_0_1), .O_0_2(NativeMapParallel_n1_inst3_O_0_2), .valid_down(NativeMapParallel_n1_inst3_valid_down), .valid_up(valid_up));
NativeMapParallel_n1_unq1 NativeMapParallel_n1_inst4(.I0_0_0(I0_4_0_0), .I0_0_1(I0_4_0_1), .I1_0(I1_4_0), .O_0_0(NativeMapParallel_n1_inst4_O_0_0), .O_0_1(NativeMapParallel_n1_inst4_O_0_1), .O_0_2(NativeMapParallel_n1_inst4_O_0_2), .valid_down(NativeMapParallel_n1_inst4_valid_down), .valid_up(valid_up));
NativeMapParallel_n1_unq1 NativeMapParallel_n1_inst5(.I0_0_0(I0_5_0_0), .I0_0_1(I0_5_0_1), .I1_0(I1_5_0), .O_0_0(NativeMapParallel_n1_inst5_O_0_0), .O_0_1(NativeMapParallel_n1_inst5_O_0_1), .O_0_2(NativeMapParallel_n1_inst5_O_0_2), .valid_down(NativeMapParallel_n1_inst5_valid_down), .valid_up(valid_up));
NativeMapParallel_n1_unq1 NativeMapParallel_n1_inst6(.I0_0_0(I0_6_0_0), .I0_0_1(I0_6_0_1), .I1_0(I1_6_0), .O_0_0(NativeMapParallel_n1_inst6_O_0_0), .O_0_1(NativeMapParallel_n1_inst6_O_0_1), .O_0_2(NativeMapParallel_n1_inst6_O_0_2), .valid_down(NativeMapParallel_n1_inst6_valid_down), .valid_up(valid_up));
NativeMapParallel_n1_unq1 NativeMapParallel_n1_inst7(.I0_0_0(I0_7_0_0), .I0_0_1(I0_7_0_1), .I1_0(I1_7_0), .O_0_0(NativeMapParallel_n1_inst7_O_0_0), .O_0_1(NativeMapParallel_n1_inst7_O_0_1), .O_0_2(NativeMapParallel_n1_inst7_O_0_2), .valid_down(NativeMapParallel_n1_inst7_valid_down), .valid_up(valid_up));
NativeMapParallel_n1_unq1 NativeMapParallel_n1_inst8(.I0_0_0(I0_8_0_0), .I0_0_1(I0_8_0_1), .I1_0(I1_8_0), .O_0_0(NativeMapParallel_n1_inst8_O_0_0), .O_0_1(NativeMapParallel_n1_inst8_O_0_1), .O_0_2(NativeMapParallel_n1_inst8_O_0_2), .valid_down(NativeMapParallel_n1_inst8_valid_down), .valid_up(valid_up));
corebit_and and_inst0(.in0(NativeMapParallel_n1_inst0_valid_down), .in1(NativeMapParallel_n1_inst1_valid_down), .out(and_inst0_out));
corebit_and and_inst1(.in0(and_inst0_out), .in1(NativeMapParallel_n1_inst2_valid_down), .out(and_inst1_out));
corebit_and and_inst2(.in0(and_inst1_out), .in1(NativeMapParallel_n1_inst3_valid_down), .out(and_inst2_out));
corebit_and and_inst3(.in0(and_inst2_out), .in1(NativeMapParallel_n1_inst4_valid_down), .out(and_inst3_out));
corebit_and and_inst4(.in0(and_inst3_out), .in1(NativeMapParallel_n1_inst5_valid_down), .out(and_inst4_out));
corebit_and and_inst5(.in0(and_inst4_out), .in1(NativeMapParallel_n1_inst6_valid_down), .out(and_inst5_out));
corebit_and and_inst6(.in0(and_inst5_out), .in1(NativeMapParallel_n1_inst7_valid_down), .out(and_inst6_out));
corebit_and and_inst7(.in0(and_inst6_out), .in1(NativeMapParallel_n1_inst8_valid_down), .out(and_inst7_out));
assign O_0_0_0 = NativeMapParallel_n1_inst0_O_0_0;
assign O_0_0_1 = NativeMapParallel_n1_inst0_O_0_1;
assign O_0_0_2 = NativeMapParallel_n1_inst0_O_0_2;
assign O_1_0_0 = NativeMapParallel_n1_inst1_O_0_0;
assign O_1_0_1 = NativeMapParallel_n1_inst1_O_0_1;
assign O_1_0_2 = NativeMapParallel_n1_inst1_O_0_2;
assign O_2_0_0 = NativeMapParallel_n1_inst2_O_0_0;
assign O_2_0_1 = NativeMapParallel_n1_inst2_O_0_1;
assign O_2_0_2 = NativeMapParallel_n1_inst2_O_0_2;
assign O_3_0_0 = NativeMapParallel_n1_inst3_O_0_0;
assign O_3_0_1 = NativeMapParallel_n1_inst3_O_0_1;
assign O_3_0_2 = NativeMapParallel_n1_inst3_O_0_2;
assign O_4_0_0 = NativeMapParallel_n1_inst4_O_0_0;
assign O_4_0_1 = NativeMapParallel_n1_inst4_O_0_1;
assign O_4_0_2 = NativeMapParallel_n1_inst4_O_0_2;
assign O_5_0_0 = NativeMapParallel_n1_inst5_O_0_0;
assign O_5_0_1 = NativeMapParallel_n1_inst5_O_0_1;
assign O_5_0_2 = NativeMapParallel_n1_inst5_O_0_2;
assign O_6_0_0 = NativeMapParallel_n1_inst6_O_0_0;
assign O_6_0_1 = NativeMapParallel_n1_inst6_O_0_1;
assign O_6_0_2 = NativeMapParallel_n1_inst6_O_0_2;
assign O_7_0_0 = NativeMapParallel_n1_inst7_O_0_0;
assign O_7_0_1 = NativeMapParallel_n1_inst7_O_0_1;
assign O_7_0_2 = NativeMapParallel_n1_inst7_O_0_2;
assign O_8_0_0 = NativeMapParallel_n1_inst8_O_0_0;
assign O_8_0_1 = NativeMapParallel_n1_inst8_O_0_1;
assign O_8_0_2 = NativeMapParallel_n1_inst8_O_0_2;
assign valid_down = and_inst7_out;
endmodule

module NativeMapParallel_n27_unq1 (input [7:0] I0_0_0_0, input [7:0] I0_0_0_1, input [7:0] I0_10_0_0, input [7:0] I0_10_0_1, input [7:0] I0_11_0_0, input [7:0] I0_11_0_1, input [7:0] I0_12_0_0, input [7:0] I0_12_0_1, input [7:0] I0_13_0_0, input [7:0] I0_13_0_1, input [7:0] I0_14_0_0, input [7:0] I0_14_0_1, input [7:0] I0_15_0_0, input [7:0] I0_15_0_1, input [7:0] I0_16_0_0, input [7:0] I0_16_0_1, input [7:0] I0_17_0_0, input [7:0] I0_17_0_1, input [7:0] I0_18_0_0, input [7:0] I0_18_0_1, input [7:0] I0_19_0_0, input [7:0] I0_19_0_1, input [7:0] I0_1_0_0, input [7:0] I0_1_0_1, input [7:0] I0_20_0_0, input [7:0] I0_20_0_1, input [7:0] I0_21_0_0, input [7:0] I0_21_0_1, input [7:0] I0_22_0_0, input [7:0] I0_22_0_1, input [7:0] I0_23_0_0, input [7:0] I0_23_0_1, input [7:0] I0_24_0_0, input [7:0] I0_24_0_1, input [7:0] I0_25_0_0, input [7:0] I0_25_0_1, input [7:0] I0_26_0_0, input [7:0] I0_26_0_1, input [7:0] I0_2_0_0, input [7:0] I0_2_0_1, input [7:0] I0_3_0_0, input [7:0] I0_3_0_1, input [7:0] I0_4_0_0, input [7:0] I0_4_0_1, input [7:0] I0_5_0_0, input [7:0] I0_5_0_1, input [7:0] I0_6_0_0, input [7:0] I0_6_0_1, input [7:0] I0_7_0_0, input [7:0] I0_7_0_1, input [7:0] I0_8_0_0, input [7:0] I0_8_0_1, input [7:0] I0_9_0_0, input [7:0] I0_9_0_1, input [7:0] I1_0_0, input [7:0] I1_10_0, input [7:0] I1_11_0, input [7:0] I1_12_0, input [7:0] I1_13_0, input [7:0] I1_14_0, input [7:0] I1_15_0, input [7:0] I1_16_0, input [7:0] I1_17_0, input [7:0] I1_18_0, input [7:0] I1_19_0, input [7:0] I1_1_0, input [7:0] I1_20_0, input [7:0] I1_21_0, input [7:0] I1_22_0, input [7:0] I1_23_0, input [7:0] I1_24_0, input [7:0] I1_25_0, input [7:0] I1_26_0, input [7:0] I1_2_0, input [7:0] I1_3_0, input [7:0] I1_4_0, input [7:0] I1_5_0, input [7:0] I1_6_0, input [7:0] I1_7_0, input [7:0] I1_8_0, input [7:0] I1_9_0, output [7:0] O_0_0_0, output [7:0] O_0_0_1, output [7:0] O_0_0_2, output [7:0] O_10_0_0, output [7:0] O_10_0_1, output [7:0] O_10_0_2, output [7:0] O_11_0_0, output [7:0] O_11_0_1, output [7:0] O_11_0_2, output [7:0] O_12_0_0, output [7:0] O_12_0_1, output [7:0] O_12_0_2, output [7:0] O_13_0_0, output [7:0] O_13_0_1, output [7:0] O_13_0_2, output [7:0] O_14_0_0, output [7:0] O_14_0_1, output [7:0] O_14_0_2, output [7:0] O_15_0_0, output [7:0] O_15_0_1, output [7:0] O_15_0_2, output [7:0] O_16_0_0, output [7:0] O_16_0_1, output [7:0] O_16_0_2, output [7:0] O_17_0_0, output [7:0] O_17_0_1, output [7:0] O_17_0_2, output [7:0] O_18_0_0, output [7:0] O_18_0_1, output [7:0] O_18_0_2, output [7:0] O_19_0_0, output [7:0] O_19_0_1, output [7:0] O_19_0_2, output [7:0] O_1_0_0, output [7:0] O_1_0_1, output [7:0] O_1_0_2, output [7:0] O_20_0_0, output [7:0] O_20_0_1, output [7:0] O_20_0_2, output [7:0] O_21_0_0, output [7:0] O_21_0_1, output [7:0] O_21_0_2, output [7:0] O_22_0_0, output [7:0] O_22_0_1, output [7:0] O_22_0_2, output [7:0] O_23_0_0, output [7:0] O_23_0_1, output [7:0] O_23_0_2, output [7:0] O_24_0_0, output [7:0] O_24_0_1, output [7:0] O_24_0_2, output [7:0] O_25_0_0, output [7:0] O_25_0_1, output [7:0] O_25_0_2, output [7:0] O_26_0_0, output [7:0] O_26_0_1, output [7:0] O_26_0_2, output [7:0] O_2_0_0, output [7:0] O_2_0_1, output [7:0] O_2_0_2, output [7:0] O_3_0_0, output [7:0] O_3_0_1, output [7:0] O_3_0_2, output [7:0] O_4_0_0, output [7:0] O_4_0_1, output [7:0] O_4_0_2, output [7:0] O_5_0_0, output [7:0] O_5_0_1, output [7:0] O_5_0_2, output [7:0] O_6_0_0, output [7:0] O_6_0_1, output [7:0] O_6_0_2, output [7:0] O_7_0_0, output [7:0] O_7_0_1, output [7:0] O_7_0_2, output [7:0] O_8_0_0, output [7:0] O_8_0_1, output [7:0] O_8_0_2, output [7:0] O_9_0_0, output [7:0] O_9_0_1, output [7:0] O_9_0_2, output valid_down, input valid_up);
wire [7:0] NativeMapParallel_n1_inst0_O_0_0;
wire [7:0] NativeMapParallel_n1_inst0_O_0_1;
wire [7:0] NativeMapParallel_n1_inst0_O_0_2;
wire NativeMapParallel_n1_inst0_valid_down;
wire [7:0] NativeMapParallel_n1_inst1_O_0_0;
wire [7:0] NativeMapParallel_n1_inst1_O_0_1;
wire [7:0] NativeMapParallel_n1_inst1_O_0_2;
wire NativeMapParallel_n1_inst1_valid_down;
wire [7:0] NativeMapParallel_n1_inst10_O_0_0;
wire [7:0] NativeMapParallel_n1_inst10_O_0_1;
wire [7:0] NativeMapParallel_n1_inst10_O_0_2;
wire NativeMapParallel_n1_inst10_valid_down;
wire [7:0] NativeMapParallel_n1_inst11_O_0_0;
wire [7:0] NativeMapParallel_n1_inst11_O_0_1;
wire [7:0] NativeMapParallel_n1_inst11_O_0_2;
wire NativeMapParallel_n1_inst11_valid_down;
wire [7:0] NativeMapParallel_n1_inst12_O_0_0;
wire [7:0] NativeMapParallel_n1_inst12_O_0_1;
wire [7:0] NativeMapParallel_n1_inst12_O_0_2;
wire NativeMapParallel_n1_inst12_valid_down;
wire [7:0] NativeMapParallel_n1_inst13_O_0_0;
wire [7:0] NativeMapParallel_n1_inst13_O_0_1;
wire [7:0] NativeMapParallel_n1_inst13_O_0_2;
wire NativeMapParallel_n1_inst13_valid_down;
wire [7:0] NativeMapParallel_n1_inst14_O_0_0;
wire [7:0] NativeMapParallel_n1_inst14_O_0_1;
wire [7:0] NativeMapParallel_n1_inst14_O_0_2;
wire NativeMapParallel_n1_inst14_valid_down;
wire [7:0] NativeMapParallel_n1_inst15_O_0_0;
wire [7:0] NativeMapParallel_n1_inst15_O_0_1;
wire [7:0] NativeMapParallel_n1_inst15_O_0_2;
wire NativeMapParallel_n1_inst15_valid_down;
wire [7:0] NativeMapParallel_n1_inst16_O_0_0;
wire [7:0] NativeMapParallel_n1_inst16_O_0_1;
wire [7:0] NativeMapParallel_n1_inst16_O_0_2;
wire NativeMapParallel_n1_inst16_valid_down;
wire [7:0] NativeMapParallel_n1_inst17_O_0_0;
wire [7:0] NativeMapParallel_n1_inst17_O_0_1;
wire [7:0] NativeMapParallel_n1_inst17_O_0_2;
wire NativeMapParallel_n1_inst17_valid_down;
wire [7:0] NativeMapParallel_n1_inst18_O_0_0;
wire [7:0] NativeMapParallel_n1_inst18_O_0_1;
wire [7:0] NativeMapParallel_n1_inst18_O_0_2;
wire NativeMapParallel_n1_inst18_valid_down;
wire [7:0] NativeMapParallel_n1_inst19_O_0_0;
wire [7:0] NativeMapParallel_n1_inst19_O_0_1;
wire [7:0] NativeMapParallel_n1_inst19_O_0_2;
wire NativeMapParallel_n1_inst19_valid_down;
wire [7:0] NativeMapParallel_n1_inst2_O_0_0;
wire [7:0] NativeMapParallel_n1_inst2_O_0_1;
wire [7:0] NativeMapParallel_n1_inst2_O_0_2;
wire NativeMapParallel_n1_inst2_valid_down;
wire [7:0] NativeMapParallel_n1_inst20_O_0_0;
wire [7:0] NativeMapParallel_n1_inst20_O_0_1;
wire [7:0] NativeMapParallel_n1_inst20_O_0_2;
wire NativeMapParallel_n1_inst20_valid_down;
wire [7:0] NativeMapParallel_n1_inst21_O_0_0;
wire [7:0] NativeMapParallel_n1_inst21_O_0_1;
wire [7:0] NativeMapParallel_n1_inst21_O_0_2;
wire NativeMapParallel_n1_inst21_valid_down;
wire [7:0] NativeMapParallel_n1_inst22_O_0_0;
wire [7:0] NativeMapParallel_n1_inst22_O_0_1;
wire [7:0] NativeMapParallel_n1_inst22_O_0_2;
wire NativeMapParallel_n1_inst22_valid_down;
wire [7:0] NativeMapParallel_n1_inst23_O_0_0;
wire [7:0] NativeMapParallel_n1_inst23_O_0_1;
wire [7:0] NativeMapParallel_n1_inst23_O_0_2;
wire NativeMapParallel_n1_inst23_valid_down;
wire [7:0] NativeMapParallel_n1_inst24_O_0_0;
wire [7:0] NativeMapParallel_n1_inst24_O_0_1;
wire [7:0] NativeMapParallel_n1_inst24_O_0_2;
wire NativeMapParallel_n1_inst24_valid_down;
wire [7:0] NativeMapParallel_n1_inst25_O_0_0;
wire [7:0] NativeMapParallel_n1_inst25_O_0_1;
wire [7:0] NativeMapParallel_n1_inst25_O_0_2;
wire NativeMapParallel_n1_inst25_valid_down;
wire [7:0] NativeMapParallel_n1_inst26_O_0_0;
wire [7:0] NativeMapParallel_n1_inst26_O_0_1;
wire [7:0] NativeMapParallel_n1_inst26_O_0_2;
wire NativeMapParallel_n1_inst26_valid_down;
wire [7:0] NativeMapParallel_n1_inst3_O_0_0;
wire [7:0] NativeMapParallel_n1_inst3_O_0_1;
wire [7:0] NativeMapParallel_n1_inst3_O_0_2;
wire NativeMapParallel_n1_inst3_valid_down;
wire [7:0] NativeMapParallel_n1_inst4_O_0_0;
wire [7:0] NativeMapParallel_n1_inst4_O_0_1;
wire [7:0] NativeMapParallel_n1_inst4_O_0_2;
wire NativeMapParallel_n1_inst4_valid_down;
wire [7:0] NativeMapParallel_n1_inst5_O_0_0;
wire [7:0] NativeMapParallel_n1_inst5_O_0_1;
wire [7:0] NativeMapParallel_n1_inst5_O_0_2;
wire NativeMapParallel_n1_inst5_valid_down;
wire [7:0] NativeMapParallel_n1_inst6_O_0_0;
wire [7:0] NativeMapParallel_n1_inst6_O_0_1;
wire [7:0] NativeMapParallel_n1_inst6_O_0_2;
wire NativeMapParallel_n1_inst6_valid_down;
wire [7:0] NativeMapParallel_n1_inst7_O_0_0;
wire [7:0] NativeMapParallel_n1_inst7_O_0_1;
wire [7:0] NativeMapParallel_n1_inst7_O_0_2;
wire NativeMapParallel_n1_inst7_valid_down;
wire [7:0] NativeMapParallel_n1_inst8_O_0_0;
wire [7:0] NativeMapParallel_n1_inst8_O_0_1;
wire [7:0] NativeMapParallel_n1_inst8_O_0_2;
wire NativeMapParallel_n1_inst8_valid_down;
wire [7:0] NativeMapParallel_n1_inst9_O_0_0;
wire [7:0] NativeMapParallel_n1_inst9_O_0_1;
wire [7:0] NativeMapParallel_n1_inst9_O_0_2;
wire NativeMapParallel_n1_inst9_valid_down;
wire and_inst0_out;
wire and_inst1_out;
wire and_inst10_out;
wire and_inst11_out;
wire and_inst12_out;
wire and_inst13_out;
wire and_inst14_out;
wire and_inst15_out;
wire and_inst16_out;
wire and_inst17_out;
wire and_inst18_out;
wire and_inst19_out;
wire and_inst2_out;
wire and_inst20_out;
wire and_inst21_out;
wire and_inst22_out;
wire and_inst23_out;
wire and_inst24_out;
wire and_inst25_out;
wire and_inst3_out;
wire and_inst4_out;
wire and_inst5_out;
wire and_inst6_out;
wire and_inst7_out;
wire and_inst8_out;
wire and_inst9_out;
NativeMapParallel_n1_unq1 NativeMapParallel_n1_inst0(.I0_0_0(I0_0_0_0), .I0_0_1(I0_0_0_1), .I1_0(I1_0_0), .O_0_0(NativeMapParallel_n1_inst0_O_0_0), .O_0_1(NativeMapParallel_n1_inst0_O_0_1), .O_0_2(NativeMapParallel_n1_inst0_O_0_2), .valid_down(NativeMapParallel_n1_inst0_valid_down), .valid_up(valid_up));
NativeMapParallel_n1_unq1 NativeMapParallel_n1_inst1(.I0_0_0(I0_1_0_0), .I0_0_1(I0_1_0_1), .I1_0(I1_1_0), .O_0_0(NativeMapParallel_n1_inst1_O_0_0), .O_0_1(NativeMapParallel_n1_inst1_O_0_1), .O_0_2(NativeMapParallel_n1_inst1_O_0_2), .valid_down(NativeMapParallel_n1_inst1_valid_down), .valid_up(valid_up));
NativeMapParallel_n1_unq1 NativeMapParallel_n1_inst10(.I0_0_0(I0_10_0_0), .I0_0_1(I0_10_0_1), .I1_0(I1_10_0), .O_0_0(NativeMapParallel_n1_inst10_O_0_0), .O_0_1(NativeMapParallel_n1_inst10_O_0_1), .O_0_2(NativeMapParallel_n1_inst10_O_0_2), .valid_down(NativeMapParallel_n1_inst10_valid_down), .valid_up(valid_up));
NativeMapParallel_n1_unq1 NativeMapParallel_n1_inst11(.I0_0_0(I0_11_0_0), .I0_0_1(I0_11_0_1), .I1_0(I1_11_0), .O_0_0(NativeMapParallel_n1_inst11_O_0_0), .O_0_1(NativeMapParallel_n1_inst11_O_0_1), .O_0_2(NativeMapParallel_n1_inst11_O_0_2), .valid_down(NativeMapParallel_n1_inst11_valid_down), .valid_up(valid_up));
NativeMapParallel_n1_unq1 NativeMapParallel_n1_inst12(.I0_0_0(I0_12_0_0), .I0_0_1(I0_12_0_1), .I1_0(I1_12_0), .O_0_0(NativeMapParallel_n1_inst12_O_0_0), .O_0_1(NativeMapParallel_n1_inst12_O_0_1), .O_0_2(NativeMapParallel_n1_inst12_O_0_2), .valid_down(NativeMapParallel_n1_inst12_valid_down), .valid_up(valid_up));
NativeMapParallel_n1_unq1 NativeMapParallel_n1_inst13(.I0_0_0(I0_13_0_0), .I0_0_1(I0_13_0_1), .I1_0(I1_13_0), .O_0_0(NativeMapParallel_n1_inst13_O_0_0), .O_0_1(NativeMapParallel_n1_inst13_O_0_1), .O_0_2(NativeMapParallel_n1_inst13_O_0_2), .valid_down(NativeMapParallel_n1_inst13_valid_down), .valid_up(valid_up));
NativeMapParallel_n1_unq1 NativeMapParallel_n1_inst14(.I0_0_0(I0_14_0_0), .I0_0_1(I0_14_0_1), .I1_0(I1_14_0), .O_0_0(NativeMapParallel_n1_inst14_O_0_0), .O_0_1(NativeMapParallel_n1_inst14_O_0_1), .O_0_2(NativeMapParallel_n1_inst14_O_0_2), .valid_down(NativeMapParallel_n1_inst14_valid_down), .valid_up(valid_up));
NativeMapParallel_n1_unq1 NativeMapParallel_n1_inst15(.I0_0_0(I0_15_0_0), .I0_0_1(I0_15_0_1), .I1_0(I1_15_0), .O_0_0(NativeMapParallel_n1_inst15_O_0_0), .O_0_1(NativeMapParallel_n1_inst15_O_0_1), .O_0_2(NativeMapParallel_n1_inst15_O_0_2), .valid_down(NativeMapParallel_n1_inst15_valid_down), .valid_up(valid_up));
NativeMapParallel_n1_unq1 NativeMapParallel_n1_inst16(.I0_0_0(I0_16_0_0), .I0_0_1(I0_16_0_1), .I1_0(I1_16_0), .O_0_0(NativeMapParallel_n1_inst16_O_0_0), .O_0_1(NativeMapParallel_n1_inst16_O_0_1), .O_0_2(NativeMapParallel_n1_inst16_O_0_2), .valid_down(NativeMapParallel_n1_inst16_valid_down), .valid_up(valid_up));
NativeMapParallel_n1_unq1 NativeMapParallel_n1_inst17(.I0_0_0(I0_17_0_0), .I0_0_1(I0_17_0_1), .I1_0(I1_17_0), .O_0_0(NativeMapParallel_n1_inst17_O_0_0), .O_0_1(NativeMapParallel_n1_inst17_O_0_1), .O_0_2(NativeMapParallel_n1_inst17_O_0_2), .valid_down(NativeMapParallel_n1_inst17_valid_down), .valid_up(valid_up));
NativeMapParallel_n1_unq1 NativeMapParallel_n1_inst18(.I0_0_0(I0_18_0_0), .I0_0_1(I0_18_0_1), .I1_0(I1_18_0), .O_0_0(NativeMapParallel_n1_inst18_O_0_0), .O_0_1(NativeMapParallel_n1_inst18_O_0_1), .O_0_2(NativeMapParallel_n1_inst18_O_0_2), .valid_down(NativeMapParallel_n1_inst18_valid_down), .valid_up(valid_up));
NativeMapParallel_n1_unq1 NativeMapParallel_n1_inst19(.I0_0_0(I0_19_0_0), .I0_0_1(I0_19_0_1), .I1_0(I1_19_0), .O_0_0(NativeMapParallel_n1_inst19_O_0_0), .O_0_1(NativeMapParallel_n1_inst19_O_0_1), .O_0_2(NativeMapParallel_n1_inst19_O_0_2), .valid_down(NativeMapParallel_n1_inst19_valid_down), .valid_up(valid_up));
NativeMapParallel_n1_unq1 NativeMapParallel_n1_inst2(.I0_0_0(I0_2_0_0), .I0_0_1(I0_2_0_1), .I1_0(I1_2_0), .O_0_0(NativeMapParallel_n1_inst2_O_0_0), .O_0_1(NativeMapParallel_n1_inst2_O_0_1), .O_0_2(NativeMapParallel_n1_inst2_O_0_2), .valid_down(NativeMapParallel_n1_inst2_valid_down), .valid_up(valid_up));
NativeMapParallel_n1_unq1 NativeMapParallel_n1_inst20(.I0_0_0(I0_20_0_0), .I0_0_1(I0_20_0_1), .I1_0(I1_20_0), .O_0_0(NativeMapParallel_n1_inst20_O_0_0), .O_0_1(NativeMapParallel_n1_inst20_O_0_1), .O_0_2(NativeMapParallel_n1_inst20_O_0_2), .valid_down(NativeMapParallel_n1_inst20_valid_down), .valid_up(valid_up));
NativeMapParallel_n1_unq1 NativeMapParallel_n1_inst21(.I0_0_0(I0_21_0_0), .I0_0_1(I0_21_0_1), .I1_0(I1_21_0), .O_0_0(NativeMapParallel_n1_inst21_O_0_0), .O_0_1(NativeMapParallel_n1_inst21_O_0_1), .O_0_2(NativeMapParallel_n1_inst21_O_0_2), .valid_down(NativeMapParallel_n1_inst21_valid_down), .valid_up(valid_up));
NativeMapParallel_n1_unq1 NativeMapParallel_n1_inst22(.I0_0_0(I0_22_0_0), .I0_0_1(I0_22_0_1), .I1_0(I1_22_0), .O_0_0(NativeMapParallel_n1_inst22_O_0_0), .O_0_1(NativeMapParallel_n1_inst22_O_0_1), .O_0_2(NativeMapParallel_n1_inst22_O_0_2), .valid_down(NativeMapParallel_n1_inst22_valid_down), .valid_up(valid_up));
NativeMapParallel_n1_unq1 NativeMapParallel_n1_inst23(.I0_0_0(I0_23_0_0), .I0_0_1(I0_23_0_1), .I1_0(I1_23_0), .O_0_0(NativeMapParallel_n1_inst23_O_0_0), .O_0_1(NativeMapParallel_n1_inst23_O_0_1), .O_0_2(NativeMapParallel_n1_inst23_O_0_2), .valid_down(NativeMapParallel_n1_inst23_valid_down), .valid_up(valid_up));
NativeMapParallel_n1_unq1 NativeMapParallel_n1_inst24(.I0_0_0(I0_24_0_0), .I0_0_1(I0_24_0_1), .I1_0(I1_24_0), .O_0_0(NativeMapParallel_n1_inst24_O_0_0), .O_0_1(NativeMapParallel_n1_inst24_O_0_1), .O_0_2(NativeMapParallel_n1_inst24_O_0_2), .valid_down(NativeMapParallel_n1_inst24_valid_down), .valid_up(valid_up));
NativeMapParallel_n1_unq1 NativeMapParallel_n1_inst25(.I0_0_0(I0_25_0_0), .I0_0_1(I0_25_0_1), .I1_0(I1_25_0), .O_0_0(NativeMapParallel_n1_inst25_O_0_0), .O_0_1(NativeMapParallel_n1_inst25_O_0_1), .O_0_2(NativeMapParallel_n1_inst25_O_0_2), .valid_down(NativeMapParallel_n1_inst25_valid_down), .valid_up(valid_up));
NativeMapParallel_n1_unq1 NativeMapParallel_n1_inst26(.I0_0_0(I0_26_0_0), .I0_0_1(I0_26_0_1), .I1_0(I1_26_0), .O_0_0(NativeMapParallel_n1_inst26_O_0_0), .O_0_1(NativeMapParallel_n1_inst26_O_0_1), .O_0_2(NativeMapParallel_n1_inst26_O_0_2), .valid_down(NativeMapParallel_n1_inst26_valid_down), .valid_up(valid_up));
NativeMapParallel_n1_unq1 NativeMapParallel_n1_inst3(.I0_0_0(I0_3_0_0), .I0_0_1(I0_3_0_1), .I1_0(I1_3_0), .O_0_0(NativeMapParallel_n1_inst3_O_0_0), .O_0_1(NativeMapParallel_n1_inst3_O_0_1), .O_0_2(NativeMapParallel_n1_inst3_O_0_2), .valid_down(NativeMapParallel_n1_inst3_valid_down), .valid_up(valid_up));
NativeMapParallel_n1_unq1 NativeMapParallel_n1_inst4(.I0_0_0(I0_4_0_0), .I0_0_1(I0_4_0_1), .I1_0(I1_4_0), .O_0_0(NativeMapParallel_n1_inst4_O_0_0), .O_0_1(NativeMapParallel_n1_inst4_O_0_1), .O_0_2(NativeMapParallel_n1_inst4_O_0_2), .valid_down(NativeMapParallel_n1_inst4_valid_down), .valid_up(valid_up));
NativeMapParallel_n1_unq1 NativeMapParallel_n1_inst5(.I0_0_0(I0_5_0_0), .I0_0_1(I0_5_0_1), .I1_0(I1_5_0), .O_0_0(NativeMapParallel_n1_inst5_O_0_0), .O_0_1(NativeMapParallel_n1_inst5_O_0_1), .O_0_2(NativeMapParallel_n1_inst5_O_0_2), .valid_down(NativeMapParallel_n1_inst5_valid_down), .valid_up(valid_up));
NativeMapParallel_n1_unq1 NativeMapParallel_n1_inst6(.I0_0_0(I0_6_0_0), .I0_0_1(I0_6_0_1), .I1_0(I1_6_0), .O_0_0(NativeMapParallel_n1_inst6_O_0_0), .O_0_1(NativeMapParallel_n1_inst6_O_0_1), .O_0_2(NativeMapParallel_n1_inst6_O_0_2), .valid_down(NativeMapParallel_n1_inst6_valid_down), .valid_up(valid_up));
NativeMapParallel_n1_unq1 NativeMapParallel_n1_inst7(.I0_0_0(I0_7_0_0), .I0_0_1(I0_7_0_1), .I1_0(I1_7_0), .O_0_0(NativeMapParallel_n1_inst7_O_0_0), .O_0_1(NativeMapParallel_n1_inst7_O_0_1), .O_0_2(NativeMapParallel_n1_inst7_O_0_2), .valid_down(NativeMapParallel_n1_inst7_valid_down), .valid_up(valid_up));
NativeMapParallel_n1_unq1 NativeMapParallel_n1_inst8(.I0_0_0(I0_8_0_0), .I0_0_1(I0_8_0_1), .I1_0(I1_8_0), .O_0_0(NativeMapParallel_n1_inst8_O_0_0), .O_0_1(NativeMapParallel_n1_inst8_O_0_1), .O_0_2(NativeMapParallel_n1_inst8_O_0_2), .valid_down(NativeMapParallel_n1_inst8_valid_down), .valid_up(valid_up));
NativeMapParallel_n1_unq1 NativeMapParallel_n1_inst9(.I0_0_0(I0_9_0_0), .I0_0_1(I0_9_0_1), .I1_0(I1_9_0), .O_0_0(NativeMapParallel_n1_inst9_O_0_0), .O_0_1(NativeMapParallel_n1_inst9_O_0_1), .O_0_2(NativeMapParallel_n1_inst9_O_0_2), .valid_down(NativeMapParallel_n1_inst9_valid_down), .valid_up(valid_up));
corebit_and and_inst0(.in0(NativeMapParallel_n1_inst0_valid_down), .in1(NativeMapParallel_n1_inst1_valid_down), .out(and_inst0_out));
corebit_and and_inst1(.in0(and_inst0_out), .in1(NativeMapParallel_n1_inst2_valid_down), .out(and_inst1_out));
corebit_and and_inst10(.in0(and_inst9_out), .in1(NativeMapParallel_n1_inst11_valid_down), .out(and_inst10_out));
corebit_and and_inst11(.in0(and_inst10_out), .in1(NativeMapParallel_n1_inst12_valid_down), .out(and_inst11_out));
corebit_and and_inst12(.in0(and_inst11_out), .in1(NativeMapParallel_n1_inst13_valid_down), .out(and_inst12_out));
corebit_and and_inst13(.in0(and_inst12_out), .in1(NativeMapParallel_n1_inst14_valid_down), .out(and_inst13_out));
corebit_and and_inst14(.in0(and_inst13_out), .in1(NativeMapParallel_n1_inst15_valid_down), .out(and_inst14_out));
corebit_and and_inst15(.in0(and_inst14_out), .in1(NativeMapParallel_n1_inst16_valid_down), .out(and_inst15_out));
corebit_and and_inst16(.in0(and_inst15_out), .in1(NativeMapParallel_n1_inst17_valid_down), .out(and_inst16_out));
corebit_and and_inst17(.in0(and_inst16_out), .in1(NativeMapParallel_n1_inst18_valid_down), .out(and_inst17_out));
corebit_and and_inst18(.in0(and_inst17_out), .in1(NativeMapParallel_n1_inst19_valid_down), .out(and_inst18_out));
corebit_and and_inst19(.in0(and_inst18_out), .in1(NativeMapParallel_n1_inst20_valid_down), .out(and_inst19_out));
corebit_and and_inst2(.in0(and_inst1_out), .in1(NativeMapParallel_n1_inst3_valid_down), .out(and_inst2_out));
corebit_and and_inst20(.in0(and_inst19_out), .in1(NativeMapParallel_n1_inst21_valid_down), .out(and_inst20_out));
corebit_and and_inst21(.in0(and_inst20_out), .in1(NativeMapParallel_n1_inst22_valid_down), .out(and_inst21_out));
corebit_and and_inst22(.in0(and_inst21_out), .in1(NativeMapParallel_n1_inst23_valid_down), .out(and_inst22_out));
corebit_and and_inst23(.in0(and_inst22_out), .in1(NativeMapParallel_n1_inst24_valid_down), .out(and_inst23_out));
corebit_and and_inst24(.in0(and_inst23_out), .in1(NativeMapParallel_n1_inst25_valid_down), .out(and_inst24_out));
corebit_and and_inst25(.in0(and_inst24_out), .in1(NativeMapParallel_n1_inst26_valid_down), .out(and_inst25_out));
corebit_and and_inst3(.in0(and_inst2_out), .in1(NativeMapParallel_n1_inst4_valid_down), .out(and_inst3_out));
corebit_and and_inst4(.in0(and_inst3_out), .in1(NativeMapParallel_n1_inst5_valid_down), .out(and_inst4_out));
corebit_and and_inst5(.in0(and_inst4_out), .in1(NativeMapParallel_n1_inst6_valid_down), .out(and_inst5_out));
corebit_and and_inst6(.in0(and_inst5_out), .in1(NativeMapParallel_n1_inst7_valid_down), .out(and_inst6_out));
corebit_and and_inst7(.in0(and_inst6_out), .in1(NativeMapParallel_n1_inst8_valid_down), .out(and_inst7_out));
corebit_and and_inst8(.in0(and_inst7_out), .in1(NativeMapParallel_n1_inst9_valid_down), .out(and_inst8_out));
corebit_and and_inst9(.in0(and_inst8_out), .in1(NativeMapParallel_n1_inst10_valid_down), .out(and_inst9_out));
assign O_0_0_0 = NativeMapParallel_n1_inst0_O_0_0;
assign O_0_0_1 = NativeMapParallel_n1_inst0_O_0_1;
assign O_0_0_2 = NativeMapParallel_n1_inst0_O_0_2;
assign O_10_0_0 = NativeMapParallel_n1_inst10_O_0_0;
assign O_10_0_1 = NativeMapParallel_n1_inst10_O_0_1;
assign O_10_0_2 = NativeMapParallel_n1_inst10_O_0_2;
assign O_11_0_0 = NativeMapParallel_n1_inst11_O_0_0;
assign O_11_0_1 = NativeMapParallel_n1_inst11_O_0_1;
assign O_11_0_2 = NativeMapParallel_n1_inst11_O_0_2;
assign O_12_0_0 = NativeMapParallel_n1_inst12_O_0_0;
assign O_12_0_1 = NativeMapParallel_n1_inst12_O_0_1;
assign O_12_0_2 = NativeMapParallel_n1_inst12_O_0_2;
assign O_13_0_0 = NativeMapParallel_n1_inst13_O_0_0;
assign O_13_0_1 = NativeMapParallel_n1_inst13_O_0_1;
assign O_13_0_2 = NativeMapParallel_n1_inst13_O_0_2;
assign O_14_0_0 = NativeMapParallel_n1_inst14_O_0_0;
assign O_14_0_1 = NativeMapParallel_n1_inst14_O_0_1;
assign O_14_0_2 = NativeMapParallel_n1_inst14_O_0_2;
assign O_15_0_0 = NativeMapParallel_n1_inst15_O_0_0;
assign O_15_0_1 = NativeMapParallel_n1_inst15_O_0_1;
assign O_15_0_2 = NativeMapParallel_n1_inst15_O_0_2;
assign O_16_0_0 = NativeMapParallel_n1_inst16_O_0_0;
assign O_16_0_1 = NativeMapParallel_n1_inst16_O_0_1;
assign O_16_0_2 = NativeMapParallel_n1_inst16_O_0_2;
assign O_17_0_0 = NativeMapParallel_n1_inst17_O_0_0;
assign O_17_0_1 = NativeMapParallel_n1_inst17_O_0_1;
assign O_17_0_2 = NativeMapParallel_n1_inst17_O_0_2;
assign O_18_0_0 = NativeMapParallel_n1_inst18_O_0_0;
assign O_18_0_1 = NativeMapParallel_n1_inst18_O_0_1;
assign O_18_0_2 = NativeMapParallel_n1_inst18_O_0_2;
assign O_19_0_0 = NativeMapParallel_n1_inst19_O_0_0;
assign O_19_0_1 = NativeMapParallel_n1_inst19_O_0_1;
assign O_19_0_2 = NativeMapParallel_n1_inst19_O_0_2;
assign O_1_0_0 = NativeMapParallel_n1_inst1_O_0_0;
assign O_1_0_1 = NativeMapParallel_n1_inst1_O_0_1;
assign O_1_0_2 = NativeMapParallel_n1_inst1_O_0_2;
assign O_20_0_0 = NativeMapParallel_n1_inst20_O_0_0;
assign O_20_0_1 = NativeMapParallel_n1_inst20_O_0_1;
assign O_20_0_2 = NativeMapParallel_n1_inst20_O_0_2;
assign O_21_0_0 = NativeMapParallel_n1_inst21_O_0_0;
assign O_21_0_1 = NativeMapParallel_n1_inst21_O_0_1;
assign O_21_0_2 = NativeMapParallel_n1_inst21_O_0_2;
assign O_22_0_0 = NativeMapParallel_n1_inst22_O_0_0;
assign O_22_0_1 = NativeMapParallel_n1_inst22_O_0_1;
assign O_22_0_2 = NativeMapParallel_n1_inst22_O_0_2;
assign O_23_0_0 = NativeMapParallel_n1_inst23_O_0_0;
assign O_23_0_1 = NativeMapParallel_n1_inst23_O_0_1;
assign O_23_0_2 = NativeMapParallel_n1_inst23_O_0_2;
assign O_24_0_0 = NativeMapParallel_n1_inst24_O_0_0;
assign O_24_0_1 = NativeMapParallel_n1_inst24_O_0_1;
assign O_24_0_2 = NativeMapParallel_n1_inst24_O_0_2;
assign O_25_0_0 = NativeMapParallel_n1_inst25_O_0_0;
assign O_25_0_1 = NativeMapParallel_n1_inst25_O_0_1;
assign O_25_0_2 = NativeMapParallel_n1_inst25_O_0_2;
assign O_26_0_0 = NativeMapParallel_n1_inst26_O_0_0;
assign O_26_0_1 = NativeMapParallel_n1_inst26_O_0_1;
assign O_26_0_2 = NativeMapParallel_n1_inst26_O_0_2;
assign O_2_0_0 = NativeMapParallel_n1_inst2_O_0_0;
assign O_2_0_1 = NativeMapParallel_n1_inst2_O_0_1;
assign O_2_0_2 = NativeMapParallel_n1_inst2_O_0_2;
assign O_3_0_0 = NativeMapParallel_n1_inst3_O_0_0;
assign O_3_0_1 = NativeMapParallel_n1_inst3_O_0_1;
assign O_3_0_2 = NativeMapParallel_n1_inst3_O_0_2;
assign O_4_0_0 = NativeMapParallel_n1_inst4_O_0_0;
assign O_4_0_1 = NativeMapParallel_n1_inst4_O_0_1;
assign O_4_0_2 = NativeMapParallel_n1_inst4_O_0_2;
assign O_5_0_0 = NativeMapParallel_n1_inst5_O_0_0;
assign O_5_0_1 = NativeMapParallel_n1_inst5_O_0_1;
assign O_5_0_2 = NativeMapParallel_n1_inst5_O_0_2;
assign O_6_0_0 = NativeMapParallel_n1_inst6_O_0_0;
assign O_6_0_1 = NativeMapParallel_n1_inst6_O_0_1;
assign O_6_0_2 = NativeMapParallel_n1_inst6_O_0_2;
assign O_7_0_0 = NativeMapParallel_n1_inst7_O_0_0;
assign O_7_0_1 = NativeMapParallel_n1_inst7_O_0_1;
assign O_7_0_2 = NativeMapParallel_n1_inst7_O_0_2;
assign O_8_0_0 = NativeMapParallel_n1_inst8_O_0_0;
assign O_8_0_1 = NativeMapParallel_n1_inst8_O_0_1;
assign O_8_0_2 = NativeMapParallel_n1_inst8_O_0_2;
assign O_9_0_0 = NativeMapParallel_n1_inst9_O_0_0;
assign O_9_0_1 = NativeMapParallel_n1_inst9_O_0_1;
assign O_9_0_2 = NativeMapParallel_n1_inst9_O_0_2;
assign valid_down = and_inst25_out;
endmodule

module NativeMapParallel_n1 (input [7:0] I0_0, input [7:0] I1_0, output [7:0] O_0_0, output [7:0] O_0_1, output valid_down, input valid_up);
wire [7:0] sseqTupleCreator_tInt_inst0_O_0;
wire [7:0] sseqTupleCreator_tInt_inst0_O_1;
wire sseqTupleCreator_tInt_inst0_valid_down;
sseqTupleCreator_tInt sseqTupleCreator_tInt_inst0(.I0(I0_0), .I1(I1_0), .O_0(sseqTupleCreator_tInt_inst0_O_0), .O_1(sseqTupleCreator_tInt_inst0_O_1), .valid_down(sseqTupleCreator_tInt_inst0_valid_down), .valid_up(valid_up));
assign O_0_0 = sseqTupleCreator_tInt_inst0_O_0;
assign O_0_1 = sseqTupleCreator_tInt_inst0_O_1;
assign valid_down = sseqTupleCreator_tInt_inst0_valid_down;
endmodule

module NativeMapParallel_n9_unq1 (input [7:0] I0_0_0, input [7:0] I0_1_0, input [7:0] I0_2_0, input [7:0] I0_3_0, input [7:0] I0_4_0, input [7:0] I0_5_0, input [7:0] I0_6_0, input [7:0] I0_7_0, input [7:0] I0_8_0, input [7:0] I1_0_0, input [7:0] I1_1_0, input [7:0] I1_2_0, input [7:0] I1_3_0, input [7:0] I1_4_0, input [7:0] I1_5_0, input [7:0] I1_6_0, input [7:0] I1_7_0, input [7:0] I1_8_0, output [7:0] O_0_0_0, output [7:0] O_0_0_1, output [7:0] O_1_0_0, output [7:0] O_1_0_1, output [7:0] O_2_0_0, output [7:0] O_2_0_1, output [7:0] O_3_0_0, output [7:0] O_3_0_1, output [7:0] O_4_0_0, output [7:0] O_4_0_1, output [7:0] O_5_0_0, output [7:0] O_5_0_1, output [7:0] O_6_0_0, output [7:0] O_6_0_1, output [7:0] O_7_0_0, output [7:0] O_7_0_1, output [7:0] O_8_0_0, output [7:0] O_8_0_1, output valid_down, input valid_up);
wire [7:0] NativeMapParallel_n1_inst0_O_0_0;
wire [7:0] NativeMapParallel_n1_inst0_O_0_1;
wire NativeMapParallel_n1_inst0_valid_down;
wire [7:0] NativeMapParallel_n1_inst1_O_0_0;
wire [7:0] NativeMapParallel_n1_inst1_O_0_1;
wire NativeMapParallel_n1_inst1_valid_down;
wire [7:0] NativeMapParallel_n1_inst2_O_0_0;
wire [7:0] NativeMapParallel_n1_inst2_O_0_1;
wire NativeMapParallel_n1_inst2_valid_down;
wire [7:0] NativeMapParallel_n1_inst3_O_0_0;
wire [7:0] NativeMapParallel_n1_inst3_O_0_1;
wire NativeMapParallel_n1_inst3_valid_down;
wire [7:0] NativeMapParallel_n1_inst4_O_0_0;
wire [7:0] NativeMapParallel_n1_inst4_O_0_1;
wire NativeMapParallel_n1_inst4_valid_down;
wire [7:0] NativeMapParallel_n1_inst5_O_0_0;
wire [7:0] NativeMapParallel_n1_inst5_O_0_1;
wire NativeMapParallel_n1_inst5_valid_down;
wire [7:0] NativeMapParallel_n1_inst6_O_0_0;
wire [7:0] NativeMapParallel_n1_inst6_O_0_1;
wire NativeMapParallel_n1_inst6_valid_down;
wire [7:0] NativeMapParallel_n1_inst7_O_0_0;
wire [7:0] NativeMapParallel_n1_inst7_O_0_1;
wire NativeMapParallel_n1_inst7_valid_down;
wire [7:0] NativeMapParallel_n1_inst8_O_0_0;
wire [7:0] NativeMapParallel_n1_inst8_O_0_1;
wire NativeMapParallel_n1_inst8_valid_down;
wire and_inst0_out;
wire and_inst1_out;
wire and_inst2_out;
wire and_inst3_out;
wire and_inst4_out;
wire and_inst5_out;
wire and_inst6_out;
wire and_inst7_out;
NativeMapParallel_n1 NativeMapParallel_n1_inst0(.I0_0(I0_0_0), .I1_0(I1_0_0), .O_0_0(NativeMapParallel_n1_inst0_O_0_0), .O_0_1(NativeMapParallel_n1_inst0_O_0_1), .valid_down(NativeMapParallel_n1_inst0_valid_down), .valid_up(valid_up));
NativeMapParallel_n1 NativeMapParallel_n1_inst1(.I0_0(I0_1_0), .I1_0(I1_1_0), .O_0_0(NativeMapParallel_n1_inst1_O_0_0), .O_0_1(NativeMapParallel_n1_inst1_O_0_1), .valid_down(NativeMapParallel_n1_inst1_valid_down), .valid_up(valid_up));
NativeMapParallel_n1 NativeMapParallel_n1_inst2(.I0_0(I0_2_0), .I1_0(I1_2_0), .O_0_0(NativeMapParallel_n1_inst2_O_0_0), .O_0_1(NativeMapParallel_n1_inst2_O_0_1), .valid_down(NativeMapParallel_n1_inst2_valid_down), .valid_up(valid_up));
NativeMapParallel_n1 NativeMapParallel_n1_inst3(.I0_0(I0_3_0), .I1_0(I1_3_0), .O_0_0(NativeMapParallel_n1_inst3_O_0_0), .O_0_1(NativeMapParallel_n1_inst3_O_0_1), .valid_down(NativeMapParallel_n1_inst3_valid_down), .valid_up(valid_up));
NativeMapParallel_n1 NativeMapParallel_n1_inst4(.I0_0(I0_4_0), .I1_0(I1_4_0), .O_0_0(NativeMapParallel_n1_inst4_O_0_0), .O_0_1(NativeMapParallel_n1_inst4_O_0_1), .valid_down(NativeMapParallel_n1_inst4_valid_down), .valid_up(valid_up));
NativeMapParallel_n1 NativeMapParallel_n1_inst5(.I0_0(I0_5_0), .I1_0(I1_5_0), .O_0_0(NativeMapParallel_n1_inst5_O_0_0), .O_0_1(NativeMapParallel_n1_inst5_O_0_1), .valid_down(NativeMapParallel_n1_inst5_valid_down), .valid_up(valid_up));
NativeMapParallel_n1 NativeMapParallel_n1_inst6(.I0_0(I0_6_0), .I1_0(I1_6_0), .O_0_0(NativeMapParallel_n1_inst6_O_0_0), .O_0_1(NativeMapParallel_n1_inst6_O_0_1), .valid_down(NativeMapParallel_n1_inst6_valid_down), .valid_up(valid_up));
NativeMapParallel_n1 NativeMapParallel_n1_inst7(.I0_0(I0_7_0), .I1_0(I1_7_0), .O_0_0(NativeMapParallel_n1_inst7_O_0_0), .O_0_1(NativeMapParallel_n1_inst7_O_0_1), .valid_down(NativeMapParallel_n1_inst7_valid_down), .valid_up(valid_up));
NativeMapParallel_n1 NativeMapParallel_n1_inst8(.I0_0(I0_8_0), .I1_0(I1_8_0), .O_0_0(NativeMapParallel_n1_inst8_O_0_0), .O_0_1(NativeMapParallel_n1_inst8_O_0_1), .valid_down(NativeMapParallel_n1_inst8_valid_down), .valid_up(valid_up));
corebit_and and_inst0(.in0(NativeMapParallel_n1_inst0_valid_down), .in1(NativeMapParallel_n1_inst1_valid_down), .out(and_inst0_out));
corebit_and and_inst1(.in0(and_inst0_out), .in1(NativeMapParallel_n1_inst2_valid_down), .out(and_inst1_out));
corebit_and and_inst2(.in0(and_inst1_out), .in1(NativeMapParallel_n1_inst3_valid_down), .out(and_inst2_out));
corebit_and and_inst3(.in0(and_inst2_out), .in1(NativeMapParallel_n1_inst4_valid_down), .out(and_inst3_out));
corebit_and and_inst4(.in0(and_inst3_out), .in1(NativeMapParallel_n1_inst5_valid_down), .out(and_inst4_out));
corebit_and and_inst5(.in0(and_inst4_out), .in1(NativeMapParallel_n1_inst6_valid_down), .out(and_inst5_out));
corebit_and and_inst6(.in0(and_inst5_out), .in1(NativeMapParallel_n1_inst7_valid_down), .out(and_inst6_out));
corebit_and and_inst7(.in0(and_inst6_out), .in1(NativeMapParallel_n1_inst8_valid_down), .out(and_inst7_out));
assign O_0_0_0 = NativeMapParallel_n1_inst0_O_0_0;
assign O_0_0_1 = NativeMapParallel_n1_inst0_O_0_1;
assign O_1_0_0 = NativeMapParallel_n1_inst1_O_0_0;
assign O_1_0_1 = NativeMapParallel_n1_inst1_O_0_1;
assign O_2_0_0 = NativeMapParallel_n1_inst2_O_0_0;
assign O_2_0_1 = NativeMapParallel_n1_inst2_O_0_1;
assign O_3_0_0 = NativeMapParallel_n1_inst3_O_0_0;
assign O_3_0_1 = NativeMapParallel_n1_inst3_O_0_1;
assign O_4_0_0 = NativeMapParallel_n1_inst4_O_0_0;
assign O_4_0_1 = NativeMapParallel_n1_inst4_O_0_1;
assign O_5_0_0 = NativeMapParallel_n1_inst5_O_0_0;
assign O_5_0_1 = NativeMapParallel_n1_inst5_O_0_1;
assign O_6_0_0 = NativeMapParallel_n1_inst6_O_0_0;
assign O_6_0_1 = NativeMapParallel_n1_inst6_O_0_1;
assign O_7_0_0 = NativeMapParallel_n1_inst7_O_0_0;
assign O_7_0_1 = NativeMapParallel_n1_inst7_O_0_1;
assign O_8_0_0 = NativeMapParallel_n1_inst8_O_0_0;
assign O_8_0_1 = NativeMapParallel_n1_inst8_O_0_1;
assign valid_down = and_inst7_out;
endmodule

module NativeMapParallel_n27 (input [7:0] I0_0_0, input [7:0] I0_10_0, input [7:0] I0_11_0, input [7:0] I0_12_0, input [7:0] I0_13_0, input [7:0] I0_14_0, input [7:0] I0_15_0, input [7:0] I0_16_0, input [7:0] I0_17_0, input [7:0] I0_18_0, input [7:0] I0_19_0, input [7:0] I0_1_0, input [7:0] I0_20_0, input [7:0] I0_21_0, input [7:0] I0_22_0, input [7:0] I0_23_0, input [7:0] I0_24_0, input [7:0] I0_25_0, input [7:0] I0_26_0, input [7:0] I0_2_0, input [7:0] I0_3_0, input [7:0] I0_4_0, input [7:0] I0_5_0, input [7:0] I0_6_0, input [7:0] I0_7_0, input [7:0] I0_8_0, input [7:0] I0_9_0, input [7:0] I1_0_0, input [7:0] I1_10_0, input [7:0] I1_11_0, input [7:0] I1_12_0, input [7:0] I1_13_0, input [7:0] I1_14_0, input [7:0] I1_15_0, input [7:0] I1_16_0, input [7:0] I1_17_0, input [7:0] I1_18_0, input [7:0] I1_19_0, input [7:0] I1_1_0, input [7:0] I1_20_0, input [7:0] I1_21_0, input [7:0] I1_22_0, input [7:0] I1_23_0, input [7:0] I1_24_0, input [7:0] I1_25_0, input [7:0] I1_26_0, input [7:0] I1_2_0, input [7:0] I1_3_0, input [7:0] I1_4_0, input [7:0] I1_5_0, input [7:0] I1_6_0, input [7:0] I1_7_0, input [7:0] I1_8_0, input [7:0] I1_9_0, output [7:0] O_0_0_0, output [7:0] O_0_0_1, output [7:0] O_10_0_0, output [7:0] O_10_0_1, output [7:0] O_11_0_0, output [7:0] O_11_0_1, output [7:0] O_12_0_0, output [7:0] O_12_0_1, output [7:0] O_13_0_0, output [7:0] O_13_0_1, output [7:0] O_14_0_0, output [7:0] O_14_0_1, output [7:0] O_15_0_0, output [7:0] O_15_0_1, output [7:0] O_16_0_0, output [7:0] O_16_0_1, output [7:0] O_17_0_0, output [7:0] O_17_0_1, output [7:0] O_18_0_0, output [7:0] O_18_0_1, output [7:0] O_19_0_0, output [7:0] O_19_0_1, output [7:0] O_1_0_0, output [7:0] O_1_0_1, output [7:0] O_20_0_0, output [7:0] O_20_0_1, output [7:0] O_21_0_0, output [7:0] O_21_0_1, output [7:0] O_22_0_0, output [7:0] O_22_0_1, output [7:0] O_23_0_0, output [7:0] O_23_0_1, output [7:0] O_24_0_0, output [7:0] O_24_0_1, output [7:0] O_25_0_0, output [7:0] O_25_0_1, output [7:0] O_26_0_0, output [7:0] O_26_0_1, output [7:0] O_2_0_0, output [7:0] O_2_0_1, output [7:0] O_3_0_0, output [7:0] O_3_0_1, output [7:0] O_4_0_0, output [7:0] O_4_0_1, output [7:0] O_5_0_0, output [7:0] O_5_0_1, output [7:0] O_6_0_0, output [7:0] O_6_0_1, output [7:0] O_7_0_0, output [7:0] O_7_0_1, output [7:0] O_8_0_0, output [7:0] O_8_0_1, output [7:0] O_9_0_0, output [7:0] O_9_0_1, output valid_down, input valid_up);
wire [7:0] NativeMapParallel_n1_inst0_O_0_0;
wire [7:0] NativeMapParallel_n1_inst0_O_0_1;
wire NativeMapParallel_n1_inst0_valid_down;
wire [7:0] NativeMapParallel_n1_inst1_O_0_0;
wire [7:0] NativeMapParallel_n1_inst1_O_0_1;
wire NativeMapParallel_n1_inst1_valid_down;
wire [7:0] NativeMapParallel_n1_inst10_O_0_0;
wire [7:0] NativeMapParallel_n1_inst10_O_0_1;
wire NativeMapParallel_n1_inst10_valid_down;
wire [7:0] NativeMapParallel_n1_inst11_O_0_0;
wire [7:0] NativeMapParallel_n1_inst11_O_0_1;
wire NativeMapParallel_n1_inst11_valid_down;
wire [7:0] NativeMapParallel_n1_inst12_O_0_0;
wire [7:0] NativeMapParallel_n1_inst12_O_0_1;
wire NativeMapParallel_n1_inst12_valid_down;
wire [7:0] NativeMapParallel_n1_inst13_O_0_0;
wire [7:0] NativeMapParallel_n1_inst13_O_0_1;
wire NativeMapParallel_n1_inst13_valid_down;
wire [7:0] NativeMapParallel_n1_inst14_O_0_0;
wire [7:0] NativeMapParallel_n1_inst14_O_0_1;
wire NativeMapParallel_n1_inst14_valid_down;
wire [7:0] NativeMapParallel_n1_inst15_O_0_0;
wire [7:0] NativeMapParallel_n1_inst15_O_0_1;
wire NativeMapParallel_n1_inst15_valid_down;
wire [7:0] NativeMapParallel_n1_inst16_O_0_0;
wire [7:0] NativeMapParallel_n1_inst16_O_0_1;
wire NativeMapParallel_n1_inst16_valid_down;
wire [7:0] NativeMapParallel_n1_inst17_O_0_0;
wire [7:0] NativeMapParallel_n1_inst17_O_0_1;
wire NativeMapParallel_n1_inst17_valid_down;
wire [7:0] NativeMapParallel_n1_inst18_O_0_0;
wire [7:0] NativeMapParallel_n1_inst18_O_0_1;
wire NativeMapParallel_n1_inst18_valid_down;
wire [7:0] NativeMapParallel_n1_inst19_O_0_0;
wire [7:0] NativeMapParallel_n1_inst19_O_0_1;
wire NativeMapParallel_n1_inst19_valid_down;
wire [7:0] NativeMapParallel_n1_inst2_O_0_0;
wire [7:0] NativeMapParallel_n1_inst2_O_0_1;
wire NativeMapParallel_n1_inst2_valid_down;
wire [7:0] NativeMapParallel_n1_inst20_O_0_0;
wire [7:0] NativeMapParallel_n1_inst20_O_0_1;
wire NativeMapParallel_n1_inst20_valid_down;
wire [7:0] NativeMapParallel_n1_inst21_O_0_0;
wire [7:0] NativeMapParallel_n1_inst21_O_0_1;
wire NativeMapParallel_n1_inst21_valid_down;
wire [7:0] NativeMapParallel_n1_inst22_O_0_0;
wire [7:0] NativeMapParallel_n1_inst22_O_0_1;
wire NativeMapParallel_n1_inst22_valid_down;
wire [7:0] NativeMapParallel_n1_inst23_O_0_0;
wire [7:0] NativeMapParallel_n1_inst23_O_0_1;
wire NativeMapParallel_n1_inst23_valid_down;
wire [7:0] NativeMapParallel_n1_inst24_O_0_0;
wire [7:0] NativeMapParallel_n1_inst24_O_0_1;
wire NativeMapParallel_n1_inst24_valid_down;
wire [7:0] NativeMapParallel_n1_inst25_O_0_0;
wire [7:0] NativeMapParallel_n1_inst25_O_0_1;
wire NativeMapParallel_n1_inst25_valid_down;
wire [7:0] NativeMapParallel_n1_inst26_O_0_0;
wire [7:0] NativeMapParallel_n1_inst26_O_0_1;
wire NativeMapParallel_n1_inst26_valid_down;
wire [7:0] NativeMapParallel_n1_inst3_O_0_0;
wire [7:0] NativeMapParallel_n1_inst3_O_0_1;
wire NativeMapParallel_n1_inst3_valid_down;
wire [7:0] NativeMapParallel_n1_inst4_O_0_0;
wire [7:0] NativeMapParallel_n1_inst4_O_0_1;
wire NativeMapParallel_n1_inst4_valid_down;
wire [7:0] NativeMapParallel_n1_inst5_O_0_0;
wire [7:0] NativeMapParallel_n1_inst5_O_0_1;
wire NativeMapParallel_n1_inst5_valid_down;
wire [7:0] NativeMapParallel_n1_inst6_O_0_0;
wire [7:0] NativeMapParallel_n1_inst6_O_0_1;
wire NativeMapParallel_n1_inst6_valid_down;
wire [7:0] NativeMapParallel_n1_inst7_O_0_0;
wire [7:0] NativeMapParallel_n1_inst7_O_0_1;
wire NativeMapParallel_n1_inst7_valid_down;
wire [7:0] NativeMapParallel_n1_inst8_O_0_0;
wire [7:0] NativeMapParallel_n1_inst8_O_0_1;
wire NativeMapParallel_n1_inst8_valid_down;
wire [7:0] NativeMapParallel_n1_inst9_O_0_0;
wire [7:0] NativeMapParallel_n1_inst9_O_0_1;
wire NativeMapParallel_n1_inst9_valid_down;
wire and_inst0_out;
wire and_inst1_out;
wire and_inst10_out;
wire and_inst11_out;
wire and_inst12_out;
wire and_inst13_out;
wire and_inst14_out;
wire and_inst15_out;
wire and_inst16_out;
wire and_inst17_out;
wire and_inst18_out;
wire and_inst19_out;
wire and_inst2_out;
wire and_inst20_out;
wire and_inst21_out;
wire and_inst22_out;
wire and_inst23_out;
wire and_inst24_out;
wire and_inst25_out;
wire and_inst3_out;
wire and_inst4_out;
wire and_inst5_out;
wire and_inst6_out;
wire and_inst7_out;
wire and_inst8_out;
wire and_inst9_out;
NativeMapParallel_n1 NativeMapParallel_n1_inst0(.I0_0(I0_0_0), .I1_0(I1_0_0), .O_0_0(NativeMapParallel_n1_inst0_O_0_0), .O_0_1(NativeMapParallel_n1_inst0_O_0_1), .valid_down(NativeMapParallel_n1_inst0_valid_down), .valid_up(valid_up));
NativeMapParallel_n1 NativeMapParallel_n1_inst1(.I0_0(I0_1_0), .I1_0(I1_1_0), .O_0_0(NativeMapParallel_n1_inst1_O_0_0), .O_0_1(NativeMapParallel_n1_inst1_O_0_1), .valid_down(NativeMapParallel_n1_inst1_valid_down), .valid_up(valid_up));
NativeMapParallel_n1 NativeMapParallel_n1_inst10(.I0_0(I0_10_0), .I1_0(I1_10_0), .O_0_0(NativeMapParallel_n1_inst10_O_0_0), .O_0_1(NativeMapParallel_n1_inst10_O_0_1), .valid_down(NativeMapParallel_n1_inst10_valid_down), .valid_up(valid_up));
NativeMapParallel_n1 NativeMapParallel_n1_inst11(.I0_0(I0_11_0), .I1_0(I1_11_0), .O_0_0(NativeMapParallel_n1_inst11_O_0_0), .O_0_1(NativeMapParallel_n1_inst11_O_0_1), .valid_down(NativeMapParallel_n1_inst11_valid_down), .valid_up(valid_up));
NativeMapParallel_n1 NativeMapParallel_n1_inst12(.I0_0(I0_12_0), .I1_0(I1_12_0), .O_0_0(NativeMapParallel_n1_inst12_O_0_0), .O_0_1(NativeMapParallel_n1_inst12_O_0_1), .valid_down(NativeMapParallel_n1_inst12_valid_down), .valid_up(valid_up));
NativeMapParallel_n1 NativeMapParallel_n1_inst13(.I0_0(I0_13_0), .I1_0(I1_13_0), .O_0_0(NativeMapParallel_n1_inst13_O_0_0), .O_0_1(NativeMapParallel_n1_inst13_O_0_1), .valid_down(NativeMapParallel_n1_inst13_valid_down), .valid_up(valid_up));
NativeMapParallel_n1 NativeMapParallel_n1_inst14(.I0_0(I0_14_0), .I1_0(I1_14_0), .O_0_0(NativeMapParallel_n1_inst14_O_0_0), .O_0_1(NativeMapParallel_n1_inst14_O_0_1), .valid_down(NativeMapParallel_n1_inst14_valid_down), .valid_up(valid_up));
NativeMapParallel_n1 NativeMapParallel_n1_inst15(.I0_0(I0_15_0), .I1_0(I1_15_0), .O_0_0(NativeMapParallel_n1_inst15_O_0_0), .O_0_1(NativeMapParallel_n1_inst15_O_0_1), .valid_down(NativeMapParallel_n1_inst15_valid_down), .valid_up(valid_up));
NativeMapParallel_n1 NativeMapParallel_n1_inst16(.I0_0(I0_16_0), .I1_0(I1_16_0), .O_0_0(NativeMapParallel_n1_inst16_O_0_0), .O_0_1(NativeMapParallel_n1_inst16_O_0_1), .valid_down(NativeMapParallel_n1_inst16_valid_down), .valid_up(valid_up));
NativeMapParallel_n1 NativeMapParallel_n1_inst17(.I0_0(I0_17_0), .I1_0(I1_17_0), .O_0_0(NativeMapParallel_n1_inst17_O_0_0), .O_0_1(NativeMapParallel_n1_inst17_O_0_1), .valid_down(NativeMapParallel_n1_inst17_valid_down), .valid_up(valid_up));
NativeMapParallel_n1 NativeMapParallel_n1_inst18(.I0_0(I0_18_0), .I1_0(I1_18_0), .O_0_0(NativeMapParallel_n1_inst18_O_0_0), .O_0_1(NativeMapParallel_n1_inst18_O_0_1), .valid_down(NativeMapParallel_n1_inst18_valid_down), .valid_up(valid_up));
NativeMapParallel_n1 NativeMapParallel_n1_inst19(.I0_0(I0_19_0), .I1_0(I1_19_0), .O_0_0(NativeMapParallel_n1_inst19_O_0_0), .O_0_1(NativeMapParallel_n1_inst19_O_0_1), .valid_down(NativeMapParallel_n1_inst19_valid_down), .valid_up(valid_up));
NativeMapParallel_n1 NativeMapParallel_n1_inst2(.I0_0(I0_2_0), .I1_0(I1_2_0), .O_0_0(NativeMapParallel_n1_inst2_O_0_0), .O_0_1(NativeMapParallel_n1_inst2_O_0_1), .valid_down(NativeMapParallel_n1_inst2_valid_down), .valid_up(valid_up));
NativeMapParallel_n1 NativeMapParallel_n1_inst20(.I0_0(I0_20_0), .I1_0(I1_20_0), .O_0_0(NativeMapParallel_n1_inst20_O_0_0), .O_0_1(NativeMapParallel_n1_inst20_O_0_1), .valid_down(NativeMapParallel_n1_inst20_valid_down), .valid_up(valid_up));
NativeMapParallel_n1 NativeMapParallel_n1_inst21(.I0_0(I0_21_0), .I1_0(I1_21_0), .O_0_0(NativeMapParallel_n1_inst21_O_0_0), .O_0_1(NativeMapParallel_n1_inst21_O_0_1), .valid_down(NativeMapParallel_n1_inst21_valid_down), .valid_up(valid_up));
NativeMapParallel_n1 NativeMapParallel_n1_inst22(.I0_0(I0_22_0), .I1_0(I1_22_0), .O_0_0(NativeMapParallel_n1_inst22_O_0_0), .O_0_1(NativeMapParallel_n1_inst22_O_0_1), .valid_down(NativeMapParallel_n1_inst22_valid_down), .valid_up(valid_up));
NativeMapParallel_n1 NativeMapParallel_n1_inst23(.I0_0(I0_23_0), .I1_0(I1_23_0), .O_0_0(NativeMapParallel_n1_inst23_O_0_0), .O_0_1(NativeMapParallel_n1_inst23_O_0_1), .valid_down(NativeMapParallel_n1_inst23_valid_down), .valid_up(valid_up));
NativeMapParallel_n1 NativeMapParallel_n1_inst24(.I0_0(I0_24_0), .I1_0(I1_24_0), .O_0_0(NativeMapParallel_n1_inst24_O_0_0), .O_0_1(NativeMapParallel_n1_inst24_O_0_1), .valid_down(NativeMapParallel_n1_inst24_valid_down), .valid_up(valid_up));
NativeMapParallel_n1 NativeMapParallel_n1_inst25(.I0_0(I0_25_0), .I1_0(I1_25_0), .O_0_0(NativeMapParallel_n1_inst25_O_0_0), .O_0_1(NativeMapParallel_n1_inst25_O_0_1), .valid_down(NativeMapParallel_n1_inst25_valid_down), .valid_up(valid_up));
NativeMapParallel_n1 NativeMapParallel_n1_inst26(.I0_0(I0_26_0), .I1_0(I1_26_0), .O_0_0(NativeMapParallel_n1_inst26_O_0_0), .O_0_1(NativeMapParallel_n1_inst26_O_0_1), .valid_down(NativeMapParallel_n1_inst26_valid_down), .valid_up(valid_up));
NativeMapParallel_n1 NativeMapParallel_n1_inst3(.I0_0(I0_3_0), .I1_0(I1_3_0), .O_0_0(NativeMapParallel_n1_inst3_O_0_0), .O_0_1(NativeMapParallel_n1_inst3_O_0_1), .valid_down(NativeMapParallel_n1_inst3_valid_down), .valid_up(valid_up));
NativeMapParallel_n1 NativeMapParallel_n1_inst4(.I0_0(I0_4_0), .I1_0(I1_4_0), .O_0_0(NativeMapParallel_n1_inst4_O_0_0), .O_0_1(NativeMapParallel_n1_inst4_O_0_1), .valid_down(NativeMapParallel_n1_inst4_valid_down), .valid_up(valid_up));
NativeMapParallel_n1 NativeMapParallel_n1_inst5(.I0_0(I0_5_0), .I1_0(I1_5_0), .O_0_0(NativeMapParallel_n1_inst5_O_0_0), .O_0_1(NativeMapParallel_n1_inst5_O_0_1), .valid_down(NativeMapParallel_n1_inst5_valid_down), .valid_up(valid_up));
NativeMapParallel_n1 NativeMapParallel_n1_inst6(.I0_0(I0_6_0), .I1_0(I1_6_0), .O_0_0(NativeMapParallel_n1_inst6_O_0_0), .O_0_1(NativeMapParallel_n1_inst6_O_0_1), .valid_down(NativeMapParallel_n1_inst6_valid_down), .valid_up(valid_up));
NativeMapParallel_n1 NativeMapParallel_n1_inst7(.I0_0(I0_7_0), .I1_0(I1_7_0), .O_0_0(NativeMapParallel_n1_inst7_O_0_0), .O_0_1(NativeMapParallel_n1_inst7_O_0_1), .valid_down(NativeMapParallel_n1_inst7_valid_down), .valid_up(valid_up));
NativeMapParallel_n1 NativeMapParallel_n1_inst8(.I0_0(I0_8_0), .I1_0(I1_8_0), .O_0_0(NativeMapParallel_n1_inst8_O_0_0), .O_0_1(NativeMapParallel_n1_inst8_O_0_1), .valid_down(NativeMapParallel_n1_inst8_valid_down), .valid_up(valid_up));
NativeMapParallel_n1 NativeMapParallel_n1_inst9(.I0_0(I0_9_0), .I1_0(I1_9_0), .O_0_0(NativeMapParallel_n1_inst9_O_0_0), .O_0_1(NativeMapParallel_n1_inst9_O_0_1), .valid_down(NativeMapParallel_n1_inst9_valid_down), .valid_up(valid_up));
corebit_and and_inst0(.in0(NativeMapParallel_n1_inst0_valid_down), .in1(NativeMapParallel_n1_inst1_valid_down), .out(and_inst0_out));
corebit_and and_inst1(.in0(and_inst0_out), .in1(NativeMapParallel_n1_inst2_valid_down), .out(and_inst1_out));
corebit_and and_inst10(.in0(and_inst9_out), .in1(NativeMapParallel_n1_inst11_valid_down), .out(and_inst10_out));
corebit_and and_inst11(.in0(and_inst10_out), .in1(NativeMapParallel_n1_inst12_valid_down), .out(and_inst11_out));
corebit_and and_inst12(.in0(and_inst11_out), .in1(NativeMapParallel_n1_inst13_valid_down), .out(and_inst12_out));
corebit_and and_inst13(.in0(and_inst12_out), .in1(NativeMapParallel_n1_inst14_valid_down), .out(and_inst13_out));
corebit_and and_inst14(.in0(and_inst13_out), .in1(NativeMapParallel_n1_inst15_valid_down), .out(and_inst14_out));
corebit_and and_inst15(.in0(and_inst14_out), .in1(NativeMapParallel_n1_inst16_valid_down), .out(and_inst15_out));
corebit_and and_inst16(.in0(and_inst15_out), .in1(NativeMapParallel_n1_inst17_valid_down), .out(and_inst16_out));
corebit_and and_inst17(.in0(and_inst16_out), .in1(NativeMapParallel_n1_inst18_valid_down), .out(and_inst17_out));
corebit_and and_inst18(.in0(and_inst17_out), .in1(NativeMapParallel_n1_inst19_valid_down), .out(and_inst18_out));
corebit_and and_inst19(.in0(and_inst18_out), .in1(NativeMapParallel_n1_inst20_valid_down), .out(and_inst19_out));
corebit_and and_inst2(.in0(and_inst1_out), .in1(NativeMapParallel_n1_inst3_valid_down), .out(and_inst2_out));
corebit_and and_inst20(.in0(and_inst19_out), .in1(NativeMapParallel_n1_inst21_valid_down), .out(and_inst20_out));
corebit_and and_inst21(.in0(and_inst20_out), .in1(NativeMapParallel_n1_inst22_valid_down), .out(and_inst21_out));
corebit_and and_inst22(.in0(and_inst21_out), .in1(NativeMapParallel_n1_inst23_valid_down), .out(and_inst22_out));
corebit_and and_inst23(.in0(and_inst22_out), .in1(NativeMapParallel_n1_inst24_valid_down), .out(and_inst23_out));
corebit_and and_inst24(.in0(and_inst23_out), .in1(NativeMapParallel_n1_inst25_valid_down), .out(and_inst24_out));
corebit_and and_inst25(.in0(and_inst24_out), .in1(NativeMapParallel_n1_inst26_valid_down), .out(and_inst25_out));
corebit_and and_inst3(.in0(and_inst2_out), .in1(NativeMapParallel_n1_inst4_valid_down), .out(and_inst3_out));
corebit_and and_inst4(.in0(and_inst3_out), .in1(NativeMapParallel_n1_inst5_valid_down), .out(and_inst4_out));
corebit_and and_inst5(.in0(and_inst4_out), .in1(NativeMapParallel_n1_inst6_valid_down), .out(and_inst5_out));
corebit_and and_inst6(.in0(and_inst5_out), .in1(NativeMapParallel_n1_inst7_valid_down), .out(and_inst6_out));
corebit_and and_inst7(.in0(and_inst6_out), .in1(NativeMapParallel_n1_inst8_valid_down), .out(and_inst7_out));
corebit_and and_inst8(.in0(and_inst7_out), .in1(NativeMapParallel_n1_inst9_valid_down), .out(and_inst8_out));
corebit_and and_inst9(.in0(and_inst8_out), .in1(NativeMapParallel_n1_inst10_valid_down), .out(and_inst9_out));
assign O_0_0_0 = NativeMapParallel_n1_inst0_O_0_0;
assign O_0_0_1 = NativeMapParallel_n1_inst0_O_0_1;
assign O_10_0_0 = NativeMapParallel_n1_inst10_O_0_0;
assign O_10_0_1 = NativeMapParallel_n1_inst10_O_0_1;
assign O_11_0_0 = NativeMapParallel_n1_inst11_O_0_0;
assign O_11_0_1 = NativeMapParallel_n1_inst11_O_0_1;
assign O_12_0_0 = NativeMapParallel_n1_inst12_O_0_0;
assign O_12_0_1 = NativeMapParallel_n1_inst12_O_0_1;
assign O_13_0_0 = NativeMapParallel_n1_inst13_O_0_0;
assign O_13_0_1 = NativeMapParallel_n1_inst13_O_0_1;
assign O_14_0_0 = NativeMapParallel_n1_inst14_O_0_0;
assign O_14_0_1 = NativeMapParallel_n1_inst14_O_0_1;
assign O_15_0_0 = NativeMapParallel_n1_inst15_O_0_0;
assign O_15_0_1 = NativeMapParallel_n1_inst15_O_0_1;
assign O_16_0_0 = NativeMapParallel_n1_inst16_O_0_0;
assign O_16_0_1 = NativeMapParallel_n1_inst16_O_0_1;
assign O_17_0_0 = NativeMapParallel_n1_inst17_O_0_0;
assign O_17_0_1 = NativeMapParallel_n1_inst17_O_0_1;
assign O_18_0_0 = NativeMapParallel_n1_inst18_O_0_0;
assign O_18_0_1 = NativeMapParallel_n1_inst18_O_0_1;
assign O_19_0_0 = NativeMapParallel_n1_inst19_O_0_0;
assign O_19_0_1 = NativeMapParallel_n1_inst19_O_0_1;
assign O_1_0_0 = NativeMapParallel_n1_inst1_O_0_0;
assign O_1_0_1 = NativeMapParallel_n1_inst1_O_0_1;
assign O_20_0_0 = NativeMapParallel_n1_inst20_O_0_0;
assign O_20_0_1 = NativeMapParallel_n1_inst20_O_0_1;
assign O_21_0_0 = NativeMapParallel_n1_inst21_O_0_0;
assign O_21_0_1 = NativeMapParallel_n1_inst21_O_0_1;
assign O_22_0_0 = NativeMapParallel_n1_inst22_O_0_0;
assign O_22_0_1 = NativeMapParallel_n1_inst22_O_0_1;
assign O_23_0_0 = NativeMapParallel_n1_inst23_O_0_0;
assign O_23_0_1 = NativeMapParallel_n1_inst23_O_0_1;
assign O_24_0_0 = NativeMapParallel_n1_inst24_O_0_0;
assign O_24_0_1 = NativeMapParallel_n1_inst24_O_0_1;
assign O_25_0_0 = NativeMapParallel_n1_inst25_O_0_0;
assign O_25_0_1 = NativeMapParallel_n1_inst25_O_0_1;
assign O_26_0_0 = NativeMapParallel_n1_inst26_O_0_0;
assign O_26_0_1 = NativeMapParallel_n1_inst26_O_0_1;
assign O_2_0_0 = NativeMapParallel_n1_inst2_O_0_0;
assign O_2_0_1 = NativeMapParallel_n1_inst2_O_0_1;
assign O_3_0_0 = NativeMapParallel_n1_inst3_O_0_0;
assign O_3_0_1 = NativeMapParallel_n1_inst3_O_0_1;
assign O_4_0_0 = NativeMapParallel_n1_inst4_O_0_0;
assign O_4_0_1 = NativeMapParallel_n1_inst4_O_0_1;
assign O_5_0_0 = NativeMapParallel_n1_inst5_O_0_0;
assign O_5_0_1 = NativeMapParallel_n1_inst5_O_0_1;
assign O_6_0_0 = NativeMapParallel_n1_inst6_O_0_0;
assign O_6_0_1 = NativeMapParallel_n1_inst6_O_0_1;
assign O_7_0_0 = NativeMapParallel_n1_inst7_O_0_0;
assign O_7_0_1 = NativeMapParallel_n1_inst7_O_0_1;
assign O_8_0_0 = NativeMapParallel_n1_inst8_O_0_0;
assign O_8_0_1 = NativeMapParallel_n1_inst8_O_0_1;
assign O_9_0_0 = NativeMapParallel_n1_inst9_O_0_0;
assign O_9_0_1 = NativeMapParallel_n1_inst9_O_0_1;
assign valid_down = and_inst25_out;
endmodule

module Mux2xOutBits2 (input [1:0] I0, input [1:0] I1, output [1:0] O, input S);
wire [1:0] coreir_commonlib_mux2x2_inst0_out;
\commonlib_muxn__N2__width2 coreir_commonlib_mux2x2_inst0(.in_data_0(I0), .in_data_1(I1), .in_sel(S), .out(coreir_commonlib_mux2x2_inst0_out));
assign O = coreir_commonlib_mux2x2_inst0_out;
endmodule

module Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2 (input CE, input CLK, input [1:0] I, output [1:0] O, input RESET);
wire [1:0] Mux2xOutBits2_inst0_O;
wire [1:0] const_0_2_out;
wire [1:0] enable_mux_O;
wire [1:0] value_out;
Mux2xOutBits2 Mux2xOutBits2_inst0(.I0(enable_mux_O), .I1(const_0_2_out), .O(Mux2xOutBits2_inst0_O), .S(RESET));
coreir_const #(.value(2'h0), .width(2)) const_0_2(.out(const_0_2_out));
Mux2xOutBits2 enable_mux(.I0(value_out), .I1(I), .O(enable_mux_O), .S(CE));
coreir_reg #(.clk_posedge(1), .init(2'h0), .width(2)) value(.clk(CLK), .in(Mux2xOutBits2_inst0_O), .out(value_out));
assign O = value_out;
endmodule

module Mux2xOutBits1 (input [0:0] I0, input [0:0] I1, output [0:0] O, input S);
wire [0:0] coreir_commonlib_mux2x1_inst0_out;
\commonlib_muxn__N2__width1 coreir_commonlib_mux2x1_inst0(.in_data_0(I0), .in_data_1(I1), .in_sel(S), .out(coreir_commonlib_mux2x1_inst0_out));
assign O = coreir_commonlib_mux2x1_inst0_out;
endmodule

module Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1 (input CE, input CLK, input [0:0] I, output [0:0] O, input RESET);
wire [0:0] Mux2xOutBits1_inst0_O;
wire [0:0] const_0_1_out;
wire [0:0] enable_mux_O;
wire [0:0] value_out;
Mux2xOutBits1 Mux2xOutBits1_inst0(.I0(enable_mux_O), .I1(const_0_1_out), .O(Mux2xOutBits1_inst0_O), .S(RESET));
coreir_const #(.value(1'h0), .width(1)) const_0_1(.out(const_0_1_out));
Mux2xOutBits1 enable_mux(.I0(value_out), .I1(I), .O(enable_mux_O), .S(CE));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) value(.clk(CLK), .in(Mux2xOutBits1_inst0_O), .out(value_out));
assign O = value_out;
endmodule

module LUT2_8 (input I0, input I1, output O);
wire coreir_lut2_inst0_out;
lutN #(.init(4'h8), .N(2)) coreir_lut2_inst0(.in({I1,I0}), .out(coreir_lut2_inst0_out));
assign O = coreir_lut2_inst0_out;
endmodule

module LUT2_4 (input I0, input I1, output O);
wire coreir_lut2_inst0_out;
lutN #(.init(4'h4), .N(2)) coreir_lut2_inst0(.in({I1,I0}), .out(coreir_lut2_inst0_out));
assign O = coreir_lut2_inst0_out;
endmodule

module LUT1_2 (input I0, output O);
wire coreir_lut1_inst0_out;
lutN #(.init(2'h2), .N(1)) coreir_lut1_inst0(.in(I0), .out(coreir_lut1_inst0_out));
assign O = coreir_lut1_inst0_out;
endmodule

module LUT1_1 (input I0, output O);
wire coreir_lut1_inst0_out;
lutN #(.init(2'h1), .N(1)) coreir_lut1_inst0(.in(I0), .out(coreir_lut1_inst0_out));
assign O = coreir_lut1_inst0_out;
endmodule

module LUT1_0 (input I0, output O);
wire coreir_lut1_inst0_out;
lutN #(.init(2'h0), .N(1)) coreir_lut1_inst0(.in(I0), .out(coreir_lut1_inst0_out));
assign O = coreir_lut1_inst0_out;
endmodule

module LUT_Array_3_Array_8_Bit__t_1n (input CLK, input [0:0] addr, output [7:0] data_0, output [7:0] data_1, output [7:0] data_2);
wire LUT1_0_inst0_O;
wire LUT1_0_inst1_O;
wire LUT1_0_inst10_O;
wire LUT1_0_inst11_O;
wire LUT1_0_inst12_O;
wire LUT1_0_inst13_O;
wire LUT1_0_inst14_O;
wire LUT1_0_inst15_O;
wire LUT1_0_inst16_O;
wire LUT1_0_inst17_O;
wire LUT1_0_inst18_O;
wire LUT1_0_inst19_O;
wire LUT1_0_inst2_O;
wire LUT1_0_inst20_O;
wire LUT1_0_inst21_O;
wire LUT1_0_inst22_O;
wire LUT1_0_inst3_O;
wire LUT1_0_inst4_O;
wire LUT1_0_inst5_O;
wire LUT1_0_inst6_O;
wire LUT1_0_inst7_O;
wire LUT1_0_inst8_O;
wire LUT1_0_inst9_O;
wire LUT1_1_inst0_O;
wire [7:0] hydrate_tArray_3_Array_8_Bit___inst0_out_0;
wire [7:0] hydrate_tArray_3_Array_8_Bit___inst0_out_1;
wire [7:0] hydrate_tArray_3_Array_8_Bit___inst0_out_2;
LUT1_0 LUT1_0_inst0(.I0(addr[0]), .O(LUT1_0_inst0_O));
LUT1_0 LUT1_0_inst1(.I0(addr[0]), .O(LUT1_0_inst1_O));
LUT1_0 LUT1_0_inst10(.I0(addr[0]), .O(LUT1_0_inst10_O));
LUT1_0 LUT1_0_inst11(.I0(addr[0]), .O(LUT1_0_inst11_O));
LUT1_0 LUT1_0_inst12(.I0(addr[0]), .O(LUT1_0_inst12_O));
LUT1_0 LUT1_0_inst13(.I0(addr[0]), .O(LUT1_0_inst13_O));
LUT1_0 LUT1_0_inst14(.I0(addr[0]), .O(LUT1_0_inst14_O));
LUT1_0 LUT1_0_inst15(.I0(addr[0]), .O(LUT1_0_inst15_O));
LUT1_0 LUT1_0_inst16(.I0(addr[0]), .O(LUT1_0_inst16_O));
LUT1_0 LUT1_0_inst17(.I0(addr[0]), .O(LUT1_0_inst17_O));
LUT1_0 LUT1_0_inst18(.I0(addr[0]), .O(LUT1_0_inst18_O));
LUT1_0 LUT1_0_inst19(.I0(addr[0]), .O(LUT1_0_inst19_O));
LUT1_0 LUT1_0_inst2(.I0(addr[0]), .O(LUT1_0_inst2_O));
LUT1_0 LUT1_0_inst20(.I0(addr[0]), .O(LUT1_0_inst20_O));
LUT1_0 LUT1_0_inst21(.I0(addr[0]), .O(LUT1_0_inst21_O));
LUT1_0 LUT1_0_inst22(.I0(addr[0]), .O(LUT1_0_inst22_O));
LUT1_0 LUT1_0_inst3(.I0(addr[0]), .O(LUT1_0_inst3_O));
LUT1_0 LUT1_0_inst4(.I0(addr[0]), .O(LUT1_0_inst4_O));
LUT1_0 LUT1_0_inst5(.I0(addr[0]), .O(LUT1_0_inst5_O));
LUT1_0 LUT1_0_inst6(.I0(addr[0]), .O(LUT1_0_inst6_O));
LUT1_0 LUT1_0_inst7(.I0(addr[0]), .O(LUT1_0_inst7_O));
LUT1_0 LUT1_0_inst8(.I0(addr[0]), .O(LUT1_0_inst8_O));
LUT1_0 LUT1_0_inst9(.I0(addr[0]), .O(LUT1_0_inst9_O));
LUT1_1 LUT1_1_inst0(.I0(addr[0]), .O(LUT1_1_inst0_O));
\aetherlinglib_hydrate__hydratedTypeBit83 hydrate_tArray_3_Array_8_Bit___inst0(.in({LUT1_0_inst22_O,LUT1_0_inst21_O,LUT1_0_inst20_O,LUT1_0_inst19_O,LUT1_0_inst18_O,LUT1_0_inst17_O,LUT1_0_inst16_O,LUT1_0_inst15_O,LUT1_0_inst14_O,LUT1_0_inst13_O,LUT1_0_inst12_O,LUT1_0_inst11_O,LUT1_0_inst10_O,LUT1_0_inst9_O,LUT1_0_inst8_O,LUT1_1_inst0_O,LUT1_0_inst7_O,LUT1_0_inst6_O,LUT1_0_inst5_O,LUT1_0_inst4_O,LUT1_0_inst3_O,LUT1_0_inst2_O,LUT1_0_inst1_O,LUT1_0_inst0_O}), .out_0(hydrate_tArray_3_Array_8_Bit___inst0_out_0), .out_1(hydrate_tArray_3_Array_8_Bit___inst0_out_1), .out_2(hydrate_tArray_3_Array_8_Bit___inst0_out_2));
assign data_0 = hydrate_tArray_3_Array_8_Bit___inst0_out_0;
assign data_1 = hydrate_tArray_3_Array_8_Bit___inst0_out_1;
assign data_2 = hydrate_tArray_3_Array_8_Bit___inst0_out_2;
endmodule

module LUT_Array_1_Array_8_Bit__t_1n (input CLK, input [0:0] addr, output [7:0] data_0);
wire LUT1_0_inst0_O;
wire LUT1_0_inst1_O;
wire LUT1_0_inst2_O;
wire LUT1_0_inst3_O;
wire LUT1_0_inst4_O;
wire LUT1_0_inst5_O;
wire LUT1_0_inst6_O;
wire LUT1_1_inst0_O;
wire [7:0] hydrate_tArray_1_Array_8_Bit___inst0_out_0;
LUT1_0 LUT1_0_inst0(.I0(addr[0]), .O(LUT1_0_inst0_O));
LUT1_0 LUT1_0_inst1(.I0(addr[0]), .O(LUT1_0_inst1_O));
LUT1_0 LUT1_0_inst2(.I0(addr[0]), .O(LUT1_0_inst2_O));
LUT1_0 LUT1_0_inst3(.I0(addr[0]), .O(LUT1_0_inst3_O));
LUT1_0 LUT1_0_inst4(.I0(addr[0]), .O(LUT1_0_inst4_O));
LUT1_0 LUT1_0_inst5(.I0(addr[0]), .O(LUT1_0_inst5_O));
LUT1_0 LUT1_0_inst6(.I0(addr[0]), .O(LUT1_0_inst6_O));
LUT1_1 LUT1_1_inst0(.I0(addr[0]), .O(LUT1_1_inst0_O));
\aetherlinglib_hydrate__hydratedTypeBit81 hydrate_tArray_1_Array_8_Bit___inst0(.in({LUT1_0_inst6_O,LUT1_0_inst5_O,LUT1_0_inst4_O,LUT1_0_inst3_O,LUT1_0_inst2_O,LUT1_0_inst1_O,LUT1_1_inst0_O,LUT1_0_inst0_O}), .out_0(hydrate_tArray_1_Array_8_Bit___inst0_out_0));
assign data_0 = hydrate_tArray_1_Array_8_Bit___inst0_out_0;
endmodule

module LShift_Atom (input [7:0] I__0, input [7:0] I__1, output [7:0] O, output valid_down, input valid_up);
wire [7:0] shl8_inst0_out;
coreir_shl #(.width(8)) shl8_inst0(.in0(I__0), .in1(I__1), .out(shl8_inst0_out));
assign O = shl8_inst0_out;
assign valid_down = valid_up;
endmodule

module NativeMapParallel_n3_unq1 (input [7:0] I_0__0, input [7:0] I_0__1, input [7:0] I_1__0, input [7:0] I_1__1, input [7:0] I_2__0, input [7:0] I_2__1, output [7:0] O_0, output [7:0] O_1, output [7:0] O_2, output valid_down, input valid_up);
wire [7:0] LShift_Atom_inst0_O;
wire LShift_Atom_inst0_valid_down;
wire [7:0] LShift_Atom_inst1_O;
wire LShift_Atom_inst1_valid_down;
wire [7:0] LShift_Atom_inst2_O;
wire LShift_Atom_inst2_valid_down;
wire and_inst0_out;
wire and_inst1_out;
LShift_Atom LShift_Atom_inst0(.I__0(I_0__0), .I__1(I_0__1), .O(LShift_Atom_inst0_O), .valid_down(LShift_Atom_inst0_valid_down), .valid_up(valid_up));
LShift_Atom LShift_Atom_inst1(.I__0(I_1__0), .I__1(I_1__1), .O(LShift_Atom_inst1_O), .valid_down(LShift_Atom_inst1_valid_down), .valid_up(valid_up));
LShift_Atom LShift_Atom_inst2(.I__0(I_2__0), .I__1(I_2__1), .O(LShift_Atom_inst2_O), .valid_down(LShift_Atom_inst2_valid_down), .valid_up(valid_up));
corebit_and and_inst0(.in0(LShift_Atom_inst0_valid_down), .in1(LShift_Atom_inst1_valid_down), .out(and_inst0_out));
corebit_and and_inst1(.in0(and_inst0_out), .in1(LShift_Atom_inst2_valid_down), .out(and_inst1_out));
assign O_0 = LShift_Atom_inst0_O;
assign O_1 = LShift_Atom_inst1_O;
assign O_2 = LShift_Atom_inst2_O;
assign valid_down = and_inst1_out;
endmodule

module Down_S_n3_sel2_tElSSeq_1_Int__vTrue (input CLK, input [7:0] I_0_0, input [7:0] I_1_0, input [7:0] I_2_0, output [7:0] O_0_0, output valid_down, input valid_up);
Term_Array_2_Array_1_Array_8_Bit___t Term_Array_2_Array_1_Array_8_Bit___t_inst0(.I_0_0(I_0_0), .I_1_0(I_1_0));
assign O_0_0 = I_2_0;
assign valid_down = valid_up;
endmodule

module NativeMapParallel_n9 (input CLK, input [7:0] I_0_0_0, input [7:0] I_0_1_0, input [7:0] I_0_2_0, input [7:0] I_1_0_0, input [7:0] I_1_1_0, input [7:0] I_1_2_0, input [7:0] I_2_0_0, input [7:0] I_2_1_0, input [7:0] I_2_2_0, input [7:0] I_3_0_0, input [7:0] I_3_1_0, input [7:0] I_3_2_0, input [7:0] I_4_0_0, input [7:0] I_4_1_0, input [7:0] I_4_2_0, input [7:0] I_5_0_0, input [7:0] I_5_1_0, input [7:0] I_5_2_0, input [7:0] I_6_0_0, input [7:0] I_6_1_0, input [7:0] I_6_2_0, input [7:0] I_7_0_0, input [7:0] I_7_1_0, input [7:0] I_7_2_0, input [7:0] I_8_0_0, input [7:0] I_8_1_0, input [7:0] I_8_2_0, output [7:0] O_0_0_0, output [7:0] O_1_0_0, output [7:0] O_2_0_0, output [7:0] O_3_0_0, output [7:0] O_4_0_0, output [7:0] O_5_0_0, output [7:0] O_6_0_0, output [7:0] O_7_0_0, output [7:0] O_8_0_0, output valid_down, input valid_up);
wire [7:0] Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst0_O_0_0;
wire Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst0_valid_down;
wire [7:0] Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst1_O_0_0;
wire Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst1_valid_down;
wire [7:0] Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst2_O_0_0;
wire Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst2_valid_down;
wire [7:0] Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst3_O_0_0;
wire Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst3_valid_down;
wire [7:0] Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst4_O_0_0;
wire Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst4_valid_down;
wire [7:0] Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst5_O_0_0;
wire Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst5_valid_down;
wire [7:0] Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst6_O_0_0;
wire Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst6_valid_down;
wire [7:0] Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst7_O_0_0;
wire Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst7_valid_down;
wire [7:0] Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst8_O_0_0;
wire Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst8_valid_down;
wire and_inst0_out;
wire and_inst1_out;
wire and_inst2_out;
wire and_inst3_out;
wire and_inst4_out;
wire and_inst5_out;
wire and_inst6_out;
wire and_inst7_out;
Down_S_n3_sel2_tElSSeq_1_Int__vTrue Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst0(.CLK(CLK), .I_0_0(I_0_0_0), .I_1_0(I_0_1_0), .I_2_0(I_0_2_0), .O_0_0(Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst0_O_0_0), .valid_down(Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst0_valid_down), .valid_up(valid_up));
Down_S_n3_sel2_tElSSeq_1_Int__vTrue Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst1(.CLK(CLK), .I_0_0(I_1_0_0), .I_1_0(I_1_1_0), .I_2_0(I_1_2_0), .O_0_0(Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst1_O_0_0), .valid_down(Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst1_valid_down), .valid_up(valid_up));
Down_S_n3_sel2_tElSSeq_1_Int__vTrue Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst2(.CLK(CLK), .I_0_0(I_2_0_0), .I_1_0(I_2_1_0), .I_2_0(I_2_2_0), .O_0_0(Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst2_O_0_0), .valid_down(Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst2_valid_down), .valid_up(valid_up));
Down_S_n3_sel2_tElSSeq_1_Int__vTrue Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst3(.CLK(CLK), .I_0_0(I_3_0_0), .I_1_0(I_3_1_0), .I_2_0(I_3_2_0), .O_0_0(Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst3_O_0_0), .valid_down(Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst3_valid_down), .valid_up(valid_up));
Down_S_n3_sel2_tElSSeq_1_Int__vTrue Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst4(.CLK(CLK), .I_0_0(I_4_0_0), .I_1_0(I_4_1_0), .I_2_0(I_4_2_0), .O_0_0(Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst4_O_0_0), .valid_down(Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst4_valid_down), .valid_up(valid_up));
Down_S_n3_sel2_tElSSeq_1_Int__vTrue Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst5(.CLK(CLK), .I_0_0(I_5_0_0), .I_1_0(I_5_1_0), .I_2_0(I_5_2_0), .O_0_0(Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst5_O_0_0), .valid_down(Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst5_valid_down), .valid_up(valid_up));
Down_S_n3_sel2_tElSSeq_1_Int__vTrue Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst6(.CLK(CLK), .I_0_0(I_6_0_0), .I_1_0(I_6_1_0), .I_2_0(I_6_2_0), .O_0_0(Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst6_O_0_0), .valid_down(Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst6_valid_down), .valid_up(valid_up));
Down_S_n3_sel2_tElSSeq_1_Int__vTrue Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst7(.CLK(CLK), .I_0_0(I_7_0_0), .I_1_0(I_7_1_0), .I_2_0(I_7_2_0), .O_0_0(Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst7_O_0_0), .valid_down(Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst7_valid_down), .valid_up(valid_up));
Down_S_n3_sel2_tElSSeq_1_Int__vTrue Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst8(.CLK(CLK), .I_0_0(I_8_0_0), .I_1_0(I_8_1_0), .I_2_0(I_8_2_0), .O_0_0(Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst8_O_0_0), .valid_down(Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst8_valid_down), .valid_up(valid_up));
corebit_and and_inst0(.in0(Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst0_valid_down), .in1(Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst1_valid_down), .out(and_inst0_out));
corebit_and and_inst1(.in0(and_inst0_out), .in1(Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst2_valid_down), .out(and_inst1_out));
corebit_and and_inst2(.in0(and_inst1_out), .in1(Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst3_valid_down), .out(and_inst2_out));
corebit_and and_inst3(.in0(and_inst2_out), .in1(Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst4_valid_down), .out(and_inst3_out));
corebit_and and_inst4(.in0(and_inst3_out), .in1(Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst5_valid_down), .out(and_inst4_out));
corebit_and and_inst5(.in0(and_inst4_out), .in1(Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst6_valid_down), .out(and_inst5_out));
corebit_and and_inst6(.in0(and_inst5_out), .in1(Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst7_valid_down), .out(and_inst6_out));
corebit_and and_inst7(.in0(and_inst6_out), .in1(Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst8_valid_down), .out(and_inst7_out));
assign O_0_0_0 = Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst0_O_0_0;
assign O_1_0_0 = Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst1_O_0_0;
assign O_2_0_0 = Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst2_O_0_0;
assign O_3_0_0 = Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst3_O_0_0;
assign O_4_0_0 = Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst4_O_0_0;
assign O_5_0_0 = Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst5_O_0_0;
assign O_6_0_0 = Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst6_O_0_0;
assign O_7_0_0 = Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst7_O_0_0;
assign O_8_0_0 = Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst8_O_0_0;
assign valid_down = and_inst7_out;
endmodule

module NativeMapParallel_n3_unq2 (input CLK, input [7:0] I_0_0_0, input [7:0] I_0_1_0, input [7:0] I_0_2_0, input [7:0] I_1_0_0, input [7:0] I_1_1_0, input [7:0] I_1_2_0, input [7:0] I_2_0_0, input [7:0] I_2_1_0, input [7:0] I_2_2_0, output [7:0] O_0_0_0, output [7:0] O_1_0_0, output [7:0] O_2_0_0, output valid_down, input valid_up);
wire [7:0] Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst0_O_0_0;
wire Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst0_valid_down;
wire [7:0] Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst1_O_0_0;
wire Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst1_valid_down;
wire [7:0] Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst2_O_0_0;
wire Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst2_valid_down;
wire and_inst0_out;
wire and_inst1_out;
Down_S_n3_sel2_tElSSeq_1_Int__vTrue Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst0(.CLK(CLK), .I_0_0(I_0_0_0), .I_1_0(I_0_1_0), .I_2_0(I_0_2_0), .O_0_0(Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst0_O_0_0), .valid_down(Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst0_valid_down), .valid_up(valid_up));
Down_S_n3_sel2_tElSSeq_1_Int__vTrue Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst1(.CLK(CLK), .I_0_0(I_1_0_0), .I_1_0(I_1_1_0), .I_2_0(I_1_2_0), .O_0_0(Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst1_O_0_0), .valid_down(Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst1_valid_down), .valid_up(valid_up));
Down_S_n3_sel2_tElSSeq_1_Int__vTrue Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst2(.CLK(CLK), .I_0_0(I_2_0_0), .I_1_0(I_2_1_0), .I_2_0(I_2_2_0), .O_0_0(Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst2_O_0_0), .valid_down(Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst2_valid_down), .valid_up(valid_up));
corebit_and and_inst0(.in0(Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst0_valid_down), .in1(Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst1_valid_down), .out(and_inst0_out));
corebit_and and_inst1(.in0(and_inst0_out), .in1(Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst2_valid_down), .out(and_inst1_out));
assign O_0_0_0 = Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst0_O_0_0;
assign O_1_0_0 = Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst1_O_0_0;
assign O_2_0_0 = Down_S_n3_sel2_tElSSeq_1_Int__vTrue_inst2_O_0_0;
assign valid_down = and_inst1_out;
endmodule

module DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse (input CLK, input I, output O);
wire [0:0] reg_P_inst0_out;
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) reg_P_inst0(.clk(CLK), .in(I), .out(reg_P_inst0_out));
assign O = reg_P_inst0_out[0];
endmodule

module Register8 (input CLK, input [7:0] I, output [7:0] O);
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7_O;
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0(.CLK(CLK), .I(I[0]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1(.CLK(CLK), .I(I[1]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2(.CLK(CLK), .I(I[2]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3(.CLK(CLK), .I(I[3]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4(.CLK(CLK), .I(I[4]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5(.CLK(CLK), .I(I[5]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6(.CLK(CLK), .I(I[6]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7(.CLK(CLK), .I(I[7]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7_O));
assign O = {DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O};
endmodule

module Register_Array_8_Bit_t_0init_FalseCE_FalseRESET (input CLK, input [7:0] I, output [7:0] O);
wire [7:0] Register8_inst0_O;
Register8 Register8_inst0(.CLK(CLK), .I(I), .O(Register8_inst0_O));
assign O = Register8_inst0_O;
endmodule

module Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET (input CLK, input [7:0] I_0, output [7:0] O_0);
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst0_O;
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst0(.CLK(CLK), .I(I_0), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst0_O));
assign O_0 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst0_O;
endmodule

module Register_Array_3_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET (input CLK, input [7:0] I_0_0, input [7:0] I_1_0, input [7:0] I_2_0, output [7:0] O_0_0, output [7:0] O_1_0, output [7:0] O_2_0);
wire [7:0] Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_0;
wire [7:0] Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst1_O_0;
wire [7:0] Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst2_O_0;
Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0(.CLK(CLK), .I_0(I_0_0), .O_0(Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_0));
Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst1(.CLK(CLK), .I_0(I_1_0), .O_0(Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst1_O_0));
Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst2(.CLK(CLK), .I_0(I_2_0), .O_0(Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst2_O_0));
assign O_0_0 = Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_0;
assign O_1_0 = Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst1_O_0;
assign O_2_0 = Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst2_O_0;
endmodule

module Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET (input CLK, input [7:0] I_0_0, input [7:0] I_10_0, input [7:0] I_11_0, input [7:0] I_12_0, input [7:0] I_13_0, input [7:0] I_14_0, input [7:0] I_15_0, input [7:0] I_16_0, input [7:0] I_17_0, input [7:0] I_18_0, input [7:0] I_19_0, input [7:0] I_1_0, input [7:0] I_20_0, input [7:0] I_21_0, input [7:0] I_22_0, input [7:0] I_23_0, input [7:0] I_24_0, input [7:0] I_25_0, input [7:0] I_26_0, input [7:0] I_2_0, input [7:0] I_3_0, input [7:0] I_4_0, input [7:0] I_5_0, input [7:0] I_6_0, input [7:0] I_7_0, input [7:0] I_8_0, input [7:0] I_9_0, output [7:0] O_0_0, output [7:0] O_10_0, output [7:0] O_11_0, output [7:0] O_12_0, output [7:0] O_13_0, output [7:0] O_14_0, output [7:0] O_15_0, output [7:0] O_16_0, output [7:0] O_17_0, output [7:0] O_18_0, output [7:0] O_19_0, output [7:0] O_1_0, output [7:0] O_20_0, output [7:0] O_21_0, output [7:0] O_22_0, output [7:0] O_23_0, output [7:0] O_24_0, output [7:0] O_25_0, output [7:0] O_26_0, output [7:0] O_2_0, output [7:0] O_3_0, output [7:0] O_4_0, output [7:0] O_5_0, output [7:0] O_6_0, output [7:0] O_7_0, output [7:0] O_8_0, output [7:0] O_9_0);
wire [7:0] Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_0;
wire [7:0] Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst1_O_0;
wire [7:0] Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst10_O_0;
wire [7:0] Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst11_O_0;
wire [7:0] Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst12_O_0;
wire [7:0] Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst13_O_0;
wire [7:0] Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst14_O_0;
wire [7:0] Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst15_O_0;
wire [7:0] Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst16_O_0;
wire [7:0] Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst17_O_0;
wire [7:0] Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst18_O_0;
wire [7:0] Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst19_O_0;
wire [7:0] Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst2_O_0;
wire [7:0] Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst20_O_0;
wire [7:0] Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst21_O_0;
wire [7:0] Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst22_O_0;
wire [7:0] Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst23_O_0;
wire [7:0] Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst24_O_0;
wire [7:0] Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst25_O_0;
wire [7:0] Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst26_O_0;
wire [7:0] Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst3_O_0;
wire [7:0] Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst4_O_0;
wire [7:0] Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst5_O_0;
wire [7:0] Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst6_O_0;
wire [7:0] Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst7_O_0;
wire [7:0] Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst8_O_0;
wire [7:0] Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst9_O_0;
Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0(.CLK(CLK), .I_0(I_0_0), .O_0(Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_0));
Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst1(.CLK(CLK), .I_0(I_1_0), .O_0(Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst1_O_0));
Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst10(.CLK(CLK), .I_0(I_10_0), .O_0(Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst10_O_0));
Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst11(.CLK(CLK), .I_0(I_11_0), .O_0(Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst11_O_0));
Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst12(.CLK(CLK), .I_0(I_12_0), .O_0(Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst12_O_0));
Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst13(.CLK(CLK), .I_0(I_13_0), .O_0(Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst13_O_0));
Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst14(.CLK(CLK), .I_0(I_14_0), .O_0(Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst14_O_0));
Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst15(.CLK(CLK), .I_0(I_15_0), .O_0(Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst15_O_0));
Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst16(.CLK(CLK), .I_0(I_16_0), .O_0(Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst16_O_0));
Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst17(.CLK(CLK), .I_0(I_17_0), .O_0(Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst17_O_0));
Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst18(.CLK(CLK), .I_0(I_18_0), .O_0(Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst18_O_0));
Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst19(.CLK(CLK), .I_0(I_19_0), .O_0(Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst19_O_0));
Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst2(.CLK(CLK), .I_0(I_2_0), .O_0(Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst2_O_0));
Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst20(.CLK(CLK), .I_0(I_20_0), .O_0(Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst20_O_0));
Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst21(.CLK(CLK), .I_0(I_21_0), .O_0(Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst21_O_0));
Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst22(.CLK(CLK), .I_0(I_22_0), .O_0(Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst22_O_0));
Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst23(.CLK(CLK), .I_0(I_23_0), .O_0(Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst23_O_0));
Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst24(.CLK(CLK), .I_0(I_24_0), .O_0(Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst24_O_0));
Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst25(.CLK(CLK), .I_0(I_25_0), .O_0(Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst25_O_0));
Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst26(.CLK(CLK), .I_0(I_26_0), .O_0(Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst26_O_0));
Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst3(.CLK(CLK), .I_0(I_3_0), .O_0(Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst3_O_0));
Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst4(.CLK(CLK), .I_0(I_4_0), .O_0(Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst4_O_0));
Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst5(.CLK(CLK), .I_0(I_5_0), .O_0(Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst5_O_0));
Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst6(.CLK(CLK), .I_0(I_6_0), .O_0(Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst6_O_0));
Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst7(.CLK(CLK), .I_0(I_7_0), .O_0(Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst7_O_0));
Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst8(.CLK(CLK), .I_0(I_8_0), .O_0(Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst8_O_0));
Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst9(.CLK(CLK), .I_0(I_9_0), .O_0(Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst9_O_0));
assign O_0_0 = Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_0;
assign O_10_0 = Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst10_O_0;
assign O_11_0 = Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst11_O_0;
assign O_12_0 = Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst12_O_0;
assign O_13_0 = Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst13_O_0;
assign O_14_0 = Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst14_O_0;
assign O_15_0 = Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst15_O_0;
assign O_16_0 = Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst16_O_0;
assign O_17_0 = Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst17_O_0;
assign O_18_0 = Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst18_O_0;
assign O_19_0 = Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst19_O_0;
assign O_1_0 = Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst1_O_0;
assign O_20_0 = Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst20_O_0;
assign O_21_0 = Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst21_O_0;
assign O_22_0 = Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst22_O_0;
assign O_23_0 = Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst23_O_0;
assign O_24_0 = Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst24_O_0;
assign O_25_0 = Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst25_O_0;
assign O_26_0 = Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst26_O_0;
assign O_2_0 = Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst2_O_0;
assign O_3_0 = Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst3_O_0;
assign O_4_0 = Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst4_O_0;
assign O_5_0 = Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst5_O_0;
assign O_6_0 = Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst6_O_0;
assign O_7_0 = Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst7_O_0;
assign O_8_0 = Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst8_O_0;
assign O_9_0 = Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst9_O_0;
endmodule

module Register1 (input CLK, input [0:0] I, output [0:0] O);
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O;
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0(.CLK(CLK), .I(I[0]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O));
assign O = DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O;
endmodule

module Register_Bitt_0init_FalseCE_FalseRESET (input CLK, input I, output O);
wire [0:0] Register1_inst0_O;
Register1 Register1_inst0(.CLK(CLK), .I(I), .O(Register1_inst0_O));
assign O = Register1_inst0_O[0];
endmodule

module FIFO_tSSeq_3_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue (input CLK, input [7:0] I_0_0, input [7:0] I_1_0, input [7:0] I_2_0, output [7:0] O_0_0, output [7:0] O_1_0, output [7:0] O_2_0, output valid_down, input valid_up);
wire [7:0] Register_Array_3_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_0_0;
wire [7:0] Register_Array_3_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_1_0;
wire [7:0] Register_Array_3_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_2_0;
wire Register_Bitt_0init_FalseCE_FalseRESET_inst0_O;
Register_Array_3_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET Register_Array_3_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0(.CLK(CLK), .I_0_0(I_0_0), .I_1_0(I_1_0), .I_2_0(I_2_0), .O_0_0(Register_Array_3_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_0_0), .O_1_0(Register_Array_3_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_1_0), .O_2_0(Register_Array_3_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_2_0));
Register_Bitt_0init_FalseCE_FalseRESET Register_Bitt_0init_FalseCE_FalseRESET_inst0(.CLK(CLK), .I(valid_up), .O(Register_Bitt_0init_FalseCE_FalseRESET_inst0_O));
assign O_0_0 = Register_Array_3_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_0_0;
assign O_1_0 = Register_Array_3_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_1_0;
assign O_2_0 = Register_Array_3_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_2_0;
assign valid_down = Register_Bitt_0init_FalseCE_FalseRESET_inst0_O;
endmodule

module FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue (input CLK, input [7:0] I_0_0, input [7:0] I_10_0, input [7:0] I_11_0, input [7:0] I_12_0, input [7:0] I_13_0, input [7:0] I_14_0, input [7:0] I_15_0, input [7:0] I_16_0, input [7:0] I_17_0, input [7:0] I_18_0, input [7:0] I_19_0, input [7:0] I_1_0, input [7:0] I_20_0, input [7:0] I_21_0, input [7:0] I_22_0, input [7:0] I_23_0, input [7:0] I_24_0, input [7:0] I_25_0, input [7:0] I_26_0, input [7:0] I_2_0, input [7:0] I_3_0, input [7:0] I_4_0, input [7:0] I_5_0, input [7:0] I_6_0, input [7:0] I_7_0, input [7:0] I_8_0, input [7:0] I_9_0, output [7:0] O_0_0, output [7:0] O_10_0, output [7:0] O_11_0, output [7:0] O_12_0, output [7:0] O_13_0, output [7:0] O_14_0, output [7:0] O_15_0, output [7:0] O_16_0, output [7:0] O_17_0, output [7:0] O_18_0, output [7:0] O_19_0, output [7:0] O_1_0, output [7:0] O_20_0, output [7:0] O_21_0, output [7:0] O_22_0, output [7:0] O_23_0, output [7:0] O_24_0, output [7:0] O_25_0, output [7:0] O_26_0, output [7:0] O_2_0, output [7:0] O_3_0, output [7:0] O_4_0, output [7:0] O_5_0, output [7:0] O_6_0, output [7:0] O_7_0, output [7:0] O_8_0, output [7:0] O_9_0, output valid_down, input valid_up);
wire [7:0] Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_0_0;
wire [7:0] Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_10_0;
wire [7:0] Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_11_0;
wire [7:0] Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_12_0;
wire [7:0] Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_13_0;
wire [7:0] Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_14_0;
wire [7:0] Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_15_0;
wire [7:0] Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_16_0;
wire [7:0] Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_17_0;
wire [7:0] Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_18_0;
wire [7:0] Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_19_0;
wire [7:0] Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_1_0;
wire [7:0] Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_20_0;
wire [7:0] Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_21_0;
wire [7:0] Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_22_0;
wire [7:0] Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_23_0;
wire [7:0] Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_24_0;
wire [7:0] Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_25_0;
wire [7:0] Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_26_0;
wire [7:0] Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_2_0;
wire [7:0] Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_3_0;
wire [7:0] Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_4_0;
wire [7:0] Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_5_0;
wire [7:0] Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_6_0;
wire [7:0] Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_7_0;
wire [7:0] Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_8_0;
wire [7:0] Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_9_0;
wire Register_Bitt_0init_FalseCE_FalseRESET_inst0_O;
Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0(.CLK(CLK), .I_0_0(I_0_0), .I_10_0(I_10_0), .I_11_0(I_11_0), .I_12_0(I_12_0), .I_13_0(I_13_0), .I_14_0(I_14_0), .I_15_0(I_15_0), .I_16_0(I_16_0), .I_17_0(I_17_0), .I_18_0(I_18_0), .I_19_0(I_19_0), .I_1_0(I_1_0), .I_20_0(I_20_0), .I_21_0(I_21_0), .I_22_0(I_22_0), .I_23_0(I_23_0), .I_24_0(I_24_0), .I_25_0(I_25_0), .I_26_0(I_26_0), .I_2_0(I_2_0), .I_3_0(I_3_0), .I_4_0(I_4_0), .I_5_0(I_5_0), .I_6_0(I_6_0), .I_7_0(I_7_0), .I_8_0(I_8_0), .I_9_0(I_9_0), .O_0_0(Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_0_0), .O_10_0(Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_10_0), .O_11_0(Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_11_0), .O_12_0(Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_12_0), .O_13_0(Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_13_0), .O_14_0(Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_14_0), .O_15_0(Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_15_0), .O_16_0(Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_16_0), .O_17_0(Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_17_0), .O_18_0(Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_18_0), .O_19_0(Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_19_0), .O_1_0(Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_1_0), .O_20_0(Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_20_0), .O_21_0(Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_21_0), .O_22_0(Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_22_0), .O_23_0(Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_23_0), .O_24_0(Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_24_0), .O_25_0(Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_25_0), .O_26_0(Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_26_0), .O_2_0(Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_2_0), .O_3_0(Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_3_0), .O_4_0(Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_4_0), .O_5_0(Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_5_0), .O_6_0(Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_6_0), .O_7_0(Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_7_0), .O_8_0(Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_8_0), .O_9_0(Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_9_0));
Register_Bitt_0init_FalseCE_FalseRESET Register_Bitt_0init_FalseCE_FalseRESET_inst0(.CLK(CLK), .I(valid_up), .O(Register_Bitt_0init_FalseCE_FalseRESET_inst0_O));
assign O_0_0 = Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_0_0;
assign O_10_0 = Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_10_0;
assign O_11_0 = Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_11_0;
assign O_12_0 = Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_12_0;
assign O_13_0 = Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_13_0;
assign O_14_0 = Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_14_0;
assign O_15_0 = Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_15_0;
assign O_16_0 = Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_16_0;
assign O_17_0 = Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_17_0;
assign O_18_0 = Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_18_0;
assign O_19_0 = Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_19_0;
assign O_1_0 = Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_1_0;
assign O_20_0 = Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_20_0;
assign O_21_0 = Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_21_0;
assign O_22_0 = Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_22_0;
assign O_23_0 = Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_23_0;
assign O_24_0 = Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_24_0;
assign O_25_0 = Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_25_0;
assign O_26_0 = Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_26_0;
assign O_2_0 = Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_2_0;
assign O_3_0 = Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_3_0;
assign O_4_0 = Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_4_0;
assign O_5_0 = Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_5_0;
assign O_6_0 = Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_6_0;
assign O_7_0 = Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_7_0;
assign O_8_0 = Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_8_0;
assign O_9_0 = Register_Array_27_Array_1_Array_8_Bit___t_0init_FalseCE_FalseRESET_inst0_O_9_0;
assign valid_down = Register_Bitt_0init_FalseCE_FalseRESET_inst0_O;
endmodule

module Counter2CER (input CE, input CLK, output [1:0] O, input RESET);
wire [1:0] Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0_O;
wire [1:0] const_1_2_out;
wire [1:0] coreir_add2_inst0_out;
Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2 Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0(.CE(CE), .CLK(CLK), .I(coreir_add2_inst0_out), .O(Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0_O), .RESET(RESET));
coreir_const #(.value(2'h1), .width(2)) const_1_2(.out(const_1_2_out));
coreir_add #(.width(2)) coreir_add2_inst0(.in0(Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0_O), .in1(const_1_2_out), .out(coreir_add2_inst0_out));
assign O = Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0_O;
endmodule

module Counter2_Mod4CE (input CE, input CLK, output [1:0] O);
wire [1:0] Counter2CER_inst0_O;
wire LUT2_8_inst0_O;
wire and_inst0_out;
Counter2CER Counter2CER_inst0(.CE(CE), .CLK(CLK), .O(Counter2CER_inst0_O), .RESET(and_inst0_out));
LUT2_8 LUT2_8_inst0(.I0(Counter2CER_inst0_O[0]), .I1(Counter2CER_inst0_O[1]), .O(LUT2_8_inst0_O));
corebit_and and_inst0(.in0(LUT2_8_inst0_O), .in1(CE), .out(and_inst0_out));
assign O = Counter2CER_inst0_O;
endmodule

module InitialDelayCounter_3 (input CE, input CLK, output valid);
wire [1:0] Counter2_Mod4CE_inst0_O;
wire and_inst0_out;
wire [1:0] coreir_const23_inst0_out;
wire coreir_eq_2_inst0_out;
wire coreir_ult2_inst0_out;
Counter2_Mod4CE Counter2_Mod4CE_inst0(.CE(and_inst0_out), .CLK(CLK), .O(Counter2_Mod4CE_inst0_O));
corebit_and and_inst0(.in0(CE), .in1(coreir_ult2_inst0_out), .out(and_inst0_out));
coreir_const #(.value(2'h3), .width(2)) coreir_const23_inst0(.out(coreir_const23_inst0_out));
coreir_eq #(.width(2)) coreir_eq_2_inst0(.in0(Counter2_Mod4CE_inst0_O), .in1(coreir_const23_inst0_out), .out(coreir_eq_2_inst0_out));
coreir_ult #(.width(2)) coreir_ult2_inst0(.in0(Counter2_Mod4CE_inst0_O), .in1(coreir_const23_inst0_out), .out(coreir_ult2_inst0_out));
assign valid = coreir_eq_2_inst0_out;
endmodule

module Counter2_Mod3CE (input CE, input CLK, output [1:0] O);
wire [1:0] Counter2CER_inst0_O;
wire LUT2_4_inst0_O;
wire and_inst0_out;
Counter2CER Counter2CER_inst0(.CE(CE), .CLK(CLK), .O(Counter2CER_inst0_O), .RESET(and_inst0_out));
LUT2_4 LUT2_4_inst0(.I0(Counter2CER_inst0_O[0]), .I1(Counter2CER_inst0_O[1]), .O(LUT2_4_inst0_O));
corebit_and and_inst0(.in0(LUT2_4_inst0_O), .in1(CE), .out(and_inst0_out));
assign O = Counter2CER_inst0_O;
endmodule

module InitialDelayCounter_2 (input CE, input CLK, output valid);
wire [1:0] Counter2_Mod3CE_inst0_O;
wire and_inst0_out;
wire [1:0] coreir_const22_inst0_out;
wire coreir_eq_2_inst0_out;
wire coreir_ult2_inst0_out;
Counter2_Mod3CE Counter2_Mod3CE_inst0(.CE(and_inst0_out), .CLK(CLK), .O(Counter2_Mod3CE_inst0_O));
corebit_and and_inst0(.in0(CE), .in1(coreir_ult2_inst0_out), .out(and_inst0_out));
coreir_const #(.value(2'h2), .width(2)) coreir_const22_inst0(.out(coreir_const22_inst0_out));
coreir_eq #(.width(2)) coreir_eq_2_inst0(.in0(Counter2_Mod3CE_inst0_O), .in1(coreir_const22_inst0_out), .out(coreir_eq_2_inst0_out));
coreir_ult #(.width(2)) coreir_ult2_inst0(.in0(Counter2_Mod3CE_inst0_O), .in1(coreir_const22_inst0_out), .out(coreir_ult2_inst0_out));
assign valid = coreir_eq_2_inst0_out;
endmodule

module Counter1CER (input CE, input CLK, output [0:0] O, input RESET);
wire [0:0] Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0_O;
wire [0:0] const_1_1_out;
wire [0:0] coreir_add1_inst0_out;
Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1 Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0(.CE(CE), .CLK(CLK), .I(coreir_add1_inst0_out), .O(Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0_O), .RESET(RESET));
coreir_const #(.value(1'h1), .width(1)) const_1_1(.out(const_1_1_out));
coreir_add #(.width(1)) coreir_add1_inst0(.in0(Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0_O), .in1(const_1_1_out), .out(coreir_add1_inst0_out));
assign O = Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0_O;
endmodule

module Counter1_Mod2CE (input CE, input CLK, output [0:0] O);
wire [0:0] Counter1CER_inst0_O;
wire LUT1_2_inst0_O;
wire and_inst0_out;
Counter1CER Counter1CER_inst0(.CE(CE), .CLK(CLK), .O(Counter1CER_inst0_O), .RESET(and_inst0_out));
LUT1_2 LUT1_2_inst0(.I0(Counter1CER_inst0_O[0]), .O(LUT1_2_inst0_O));
corebit_and and_inst0(.in0(LUT1_2_inst0_O), .in1(CE), .out(and_inst0_out));
assign O = Counter1CER_inst0_O;
endmodule

module InitialDelayCounter_1 (input CE, input CLK, output valid);
wire [0:0] Counter1_Mod2CE_inst0_O;
wire and_inst0_out;
wire [0:0] coreir_const11_inst0_out;
wire coreir_eq_1_inst0_out;
wire coreir_ult1_inst0_out;
Counter1_Mod2CE Counter1_Mod2CE_inst0(.CE(and_inst0_out), .CLK(CLK), .O(Counter1_Mod2CE_inst0_O));
corebit_and and_inst0(.in0(CE), .in1(coreir_ult1_inst0_out), .out(and_inst0_out));
coreir_const #(.value(1'h1), .width(1)) coreir_const11_inst0(.out(coreir_const11_inst0_out));
coreir_eq #(.width(1)) coreir_eq_1_inst0(.in0(Counter1_Mod2CE_inst0_O), .in1(coreir_const11_inst0_out), .out(coreir_eq_1_inst0_out));
coreir_ult #(.width(1)) coreir_ult1_inst0(.in0(Counter1_Mod2CE_inst0_O), .in1(coreir_const11_inst0_out), .out(coreir_ult1_inst0_out));
assign valid = coreir_eq_1_inst0_out;
endmodule

module Const_tSSeq_3_Int__hasCEFalse_hasResetFalse_hasValidTrue_unq1 (input CLK, output [7:0] O_0, output [7:0] O_1, output [7:0] O_2, output valid_down, input valid_up);
wire InitialDelayCounter_2_inst0_valid;
wire [7:0] LUT_Array_3_Array_8_Bit__t_1n_inst0_data_0;
wire [7:0] LUT_Array_3_Array_8_Bit__t_1n_inst0_data_1;
wire [7:0] LUT_Array_3_Array_8_Bit__t_1n_inst0_data_2;
wire [0:0] SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse_inst0_O;
wire [0:0] coreir_const11_inst0_out;
InitialDelayCounter_2 InitialDelayCounter_2_inst0(.CE(coreir_const11_inst0_out[0]), .CLK(CLK), .valid(InitialDelayCounter_2_inst0_valid));
LUT_Array_3_Array_8_Bit__t_1n LUT_Array_3_Array_8_Bit__t_1n_inst0(.CLK(CLK), .addr(SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse_inst0_O), .data_0(LUT_Array_3_Array_8_Bit__t_1n_inst0_data_0), .data_1(LUT_Array_3_Array_8_Bit__t_1n_inst0_data_1), .data_2(LUT_Array_3_Array_8_Bit__t_1n_inst0_data_2));
SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse_inst0(.CE(InitialDelayCounter_2_inst0_valid), .CLK(CLK), .O(SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse_inst0_O));
Term_Bitt Term_Bitt_inst0(.I(valid_up));
coreir_const #(.value(1'h1), .width(1)) coreir_const11_inst0(.out(coreir_const11_inst0_out));
assign O_0 = LUT_Array_3_Array_8_Bit__t_1n_inst0_data_0;
assign O_1 = LUT_Array_3_Array_8_Bit__t_1n_inst0_data_1;
assign O_2 = LUT_Array_3_Array_8_Bit__t_1n_inst0_data_2;
assign valid_down = InitialDelayCounter_2_inst0_valid;
endmodule

module Const_tSSeq_3_Int__hasCEFalse_hasResetFalse_hasValidTrue (input CLK, output [7:0] O_0, output [7:0] O_1, output [7:0] O_2, output valid_down, input valid_up);
wire InitialDelayCounter_1_inst0_valid;
wire [7:0] LUT_Array_3_Array_8_Bit__t_1n_inst0_data_0;
wire [7:0] LUT_Array_3_Array_8_Bit__t_1n_inst0_data_1;
wire [7:0] LUT_Array_3_Array_8_Bit__t_1n_inst0_data_2;
wire [0:0] SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse_inst0_O;
wire [0:0] coreir_const11_inst0_out;
InitialDelayCounter_1 InitialDelayCounter_1_inst0(.CE(coreir_const11_inst0_out[0]), .CLK(CLK), .valid(InitialDelayCounter_1_inst0_valid));
LUT_Array_3_Array_8_Bit__t_1n LUT_Array_3_Array_8_Bit__t_1n_inst0(.CLK(CLK), .addr(SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse_inst0_O), .data_0(LUT_Array_3_Array_8_Bit__t_1n_inst0_data_0), .data_1(LUT_Array_3_Array_8_Bit__t_1n_inst0_data_1), .data_2(LUT_Array_3_Array_8_Bit__t_1n_inst0_data_2));
SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse_inst0(.CE(InitialDelayCounter_1_inst0_valid), .CLK(CLK), .O(SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse_inst0_O));
Term_Bitt Term_Bitt_inst0(.I(valid_up));
coreir_const #(.value(1'h1), .width(1)) coreir_const11_inst0(.out(coreir_const11_inst0_out));
assign O_0 = LUT_Array_3_Array_8_Bit__t_1n_inst0_data_0;
assign O_1 = LUT_Array_3_Array_8_Bit__t_1n_inst0_data_1;
assign O_2 = LUT_Array_3_Array_8_Bit__t_1n_inst0_data_2;
assign valid_down = InitialDelayCounter_1_inst0_valid;
endmodule

module Const_tSSeq_1_Int__hasCEFalse_hasResetFalse_hasValidTrue_unq1 (input CLK, output [7:0] O_0, output valid_down, input valid_up);
wire InitialDelayCounter_3_inst0_valid;
wire [7:0] LUT_Array_1_Array_8_Bit__t_1n_inst0_data_0;
wire [0:0] SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse_inst0_O;
wire [0:0] coreir_const11_inst0_out;
InitialDelayCounter_3 InitialDelayCounter_3_inst0(.CE(coreir_const11_inst0_out[0]), .CLK(CLK), .valid(InitialDelayCounter_3_inst0_valid));
LUT_Array_1_Array_8_Bit__t_1n LUT_Array_1_Array_8_Bit__t_1n_inst0(.CLK(CLK), .addr(SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse_inst0_O), .data_0(LUT_Array_1_Array_8_Bit__t_1n_inst0_data_0));
SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse_inst0(.CE(InitialDelayCounter_3_inst0_valid), .CLK(CLK), .O(SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse_inst0_O));
Term_Bitt Term_Bitt_inst0(.I(valid_up));
coreir_const #(.value(1'h1), .width(1)) coreir_const11_inst0(.out(coreir_const11_inst0_out));
assign O_0 = LUT_Array_1_Array_8_Bit__t_1n_inst0_data_0;
assign valid_down = InitialDelayCounter_3_inst0_valid;
endmodule

module Const_tSSeq_1_Int__hasCEFalse_hasResetFalse_hasValidTrue (input CLK, output [7:0] O_0, output valid_down, input valid_up);
wire InitialDelayCounter_2_inst0_valid;
wire [7:0] LUT_Array_1_Array_8_Bit__t_1n_inst0_data_0;
wire [0:0] SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse_inst0_O;
wire [0:0] coreir_const11_inst0_out;
InitialDelayCounter_2 InitialDelayCounter_2_inst0(.CE(coreir_const11_inst0_out[0]), .CLK(CLK), .valid(InitialDelayCounter_2_inst0_valid));
LUT_Array_1_Array_8_Bit__t_1n LUT_Array_1_Array_8_Bit__t_1n_inst0(.CLK(CLK), .addr(SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse_inst0_O), .data_0(LUT_Array_1_Array_8_Bit__t_1n_inst0_data_0));
SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse_inst0(.CE(InitialDelayCounter_2_inst0_valid), .CLK(CLK), .O(SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse_inst0_O));
Term_Bitt Term_Bitt_inst0(.I(valid_up));
coreir_const #(.value(1'h1), .width(1)) coreir_const11_inst0(.out(coreir_const11_inst0_out));
assign O_0 = LUT_Array_1_Array_8_Bit__t_1n_inst0_data_0;
assign valid_down = InitialDelayCounter_2_inst0_valid;
endmodule

module Add_Atom (input [7:0] I__0, input [7:0] I__1, output [7:0] O);
wire [7:0] coreir_add8_inst0_out;
coreir_add #(.width(8)) coreir_add8_inst0(.in0(I__0), .in1(I__1), .out(coreir_add8_inst0_out));
assign O = coreir_add8_inst0_out;
endmodule

module renamedForReduce (input [7:0] in0, input [7:0] in1, output [7:0] out);
wire [7:0] Add_Atom_inst0_O;
Add_Atom Add_Atom_inst0(.I__0(in0), .I__1(in1), .O(Add_Atom_inst0_O));
assign out = Add_Atom_inst0_O;
endmodule

module ReduceParallel_n3 (input [7:0] I_0, input [7:0] I_1, input [7:0] I_2, output [7:0] O);
wire [7:0] renamedForReduce_inst0_out;
wire [7:0] renamedForReduce_inst1_out;
renamedForReduce renamedForReduce_inst0(.in0(I_2), .in1(renamedForReduce_inst1_out), .out(renamedForReduce_inst0_out));
renamedForReduce renamedForReduce_inst1(.in0(I_1), .in1(I_0), .out(renamedForReduce_inst1_out));
assign O = renamedForReduce_inst0_out;
endmodule

module Reduce_S_n3 (input CLK, input [7:0] I_0, input [7:0] I_1, input [7:0] I_2, output [7:0] O_0, output valid_down, input valid_up);
wire [7:0] ReduceParallel_n3_inst0_O;
wire [7:0] Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_0;
wire [0:0] reg_P_inst0_out;
ReduceParallel_n3 ReduceParallel_n3_inst0(.I_0(I_0), .I_1(I_1), .I_2(I_2), .O(ReduceParallel_n3_inst0_O));
Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0(.CLK(CLK), .I_0(ReduceParallel_n3_inst0_O), .O_0(Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_0));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) reg_P_inst0(.clk(CLK), .in(valid_up), .out(reg_P_inst0_out));
assign O_0 = Register_Array_1_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_0;
assign valid_down = reg_P_inst0_out[0];
endmodule

module Module_1 (input CLK, input [7:0] I_0, input [7:0] I_1, input [7:0] I_2, output [7:0] O_0, output valid_down, input valid_up);
wire [7:0] Const_tSSeq_1_Int__hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0;
wire Const_tSSeq_1_Int__hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down;
wire [7:0] Const_tSSeq_3_Int__hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0;
wire [7:0] Const_tSSeq_3_Int__hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_1;
wire [7:0] Const_tSSeq_3_Int__hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_2;
wire Const_tSSeq_3_Int__hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down;
wire [7:0] NativeMapParallel_n1_inst0_O_0__0;
wire [7:0] NativeMapParallel_n1_inst0_O_0__1;
wire NativeMapParallel_n1_inst0_valid_down;
wire [7:0] NativeMapParallel_n1_inst1_O_0;
wire NativeMapParallel_n1_inst1_valid_down;
wire [7:0] NativeMapParallel_n3_inst0_O_0__0;
wire [7:0] NativeMapParallel_n3_inst0_O_0__1;
wire [7:0] NativeMapParallel_n3_inst0_O_1__0;
wire [7:0] NativeMapParallel_n3_inst0_O_1__1;
wire [7:0] NativeMapParallel_n3_inst0_O_2__0;
wire [7:0] NativeMapParallel_n3_inst0_O_2__1;
wire NativeMapParallel_n3_inst0_valid_down;
wire [7:0] NativeMapParallel_n3_inst1_O_0;
wire [7:0] NativeMapParallel_n3_inst1_O_1;
wire [7:0] NativeMapParallel_n3_inst1_O_2;
wire NativeMapParallel_n3_inst1_valid_down;
wire [7:0] Reduce_S_n3_inst0_O_0;
wire Reduce_S_n3_inst0_valid_down;
wire and_inst0_out;
wire and_inst1_out;
Const_tSSeq_1_Int__hasCEFalse_hasResetFalse_hasValidTrue_unq1 Const_tSSeq_1_Int__hasCEFalse_hasResetFalse_hasValidTrue_inst0(.CLK(CLK), .O_0(Const_tSSeq_1_Int__hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0), .valid_down(Const_tSSeq_1_Int__hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down), .valid_up(valid_up));
Const_tSSeq_3_Int__hasCEFalse_hasResetFalse_hasValidTrue_unq1 Const_tSSeq_3_Int__hasCEFalse_hasResetFalse_hasValidTrue_inst0(.CLK(CLK), .O_0(Const_tSSeq_3_Int__hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0), .O_1(Const_tSSeq_3_Int__hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_1), .O_2(Const_tSSeq_3_Int__hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_2), .valid_down(Const_tSSeq_3_Int__hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down), .valid_up(valid_up));
NativeMapParallel_n1_unq2 NativeMapParallel_n1_inst0(.I0_0(Reduce_S_n3_inst0_O_0), .I1_0(Const_tSSeq_1_Int__hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0), .O_0__0(NativeMapParallel_n1_inst0_O_0__0), .O_0__1(NativeMapParallel_n1_inst0_O_0__1), .valid_down(NativeMapParallel_n1_inst0_valid_down), .valid_up(and_inst1_out));
NativeMapParallel_n1_unq3 NativeMapParallel_n1_inst1(.I_0__0(NativeMapParallel_n1_inst0_O_0__0), .I_0__1(NativeMapParallel_n1_inst0_O_0__1), .O_0(NativeMapParallel_n1_inst1_O_0), .valid_down(NativeMapParallel_n1_inst1_valid_down), .valid_up(NativeMapParallel_n1_inst0_valid_down));
NativeMapParallel_n3 NativeMapParallel_n3_inst0(.I0_0(I_0), .I0_1(I_1), .I0_2(I_2), .I1_0(Const_tSSeq_3_Int__hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0), .I1_1(Const_tSSeq_3_Int__hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_1), .I1_2(Const_tSSeq_3_Int__hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_2), .O_0__0(NativeMapParallel_n3_inst0_O_0__0), .O_0__1(NativeMapParallel_n3_inst0_O_0__1), .O_1__0(NativeMapParallel_n3_inst0_O_1__0), .O_1__1(NativeMapParallel_n3_inst0_O_1__1), .O_2__0(NativeMapParallel_n3_inst0_O_2__0), .O_2__1(NativeMapParallel_n3_inst0_O_2__1), .valid_down(NativeMapParallel_n3_inst0_valid_down), .valid_up(and_inst0_out));
NativeMapParallel_n3_unq1 NativeMapParallel_n3_inst1(.I_0__0(NativeMapParallel_n3_inst0_O_0__0), .I_0__1(NativeMapParallel_n3_inst0_O_0__1), .I_1__0(NativeMapParallel_n3_inst0_O_1__0), .I_1__1(NativeMapParallel_n3_inst0_O_1__1), .I_2__0(NativeMapParallel_n3_inst0_O_2__0), .I_2__1(NativeMapParallel_n3_inst0_O_2__1), .O_0(NativeMapParallel_n3_inst1_O_0), .O_1(NativeMapParallel_n3_inst1_O_1), .O_2(NativeMapParallel_n3_inst1_O_2), .valid_down(NativeMapParallel_n3_inst1_valid_down), .valid_up(NativeMapParallel_n3_inst0_valid_down));
Reduce_S_n3 Reduce_S_n3_inst0(.CLK(CLK), .I_0(NativeMapParallel_n3_inst1_O_0), .I_1(NativeMapParallel_n3_inst1_O_1), .I_2(NativeMapParallel_n3_inst1_O_2), .O_0(Reduce_S_n3_inst0_O_0), .valid_down(Reduce_S_n3_inst0_valid_down), .valid_up(NativeMapParallel_n3_inst1_valid_down));
corebit_and and_inst0(.in0(valid_up), .in1(Const_tSSeq_3_Int__hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down), .out(and_inst0_out));
corebit_and and_inst1(.in0(Reduce_S_n3_inst0_valid_down), .in1(Const_tSSeq_1_Int__hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down), .out(and_inst1_out));
assign O_0 = NativeMapParallel_n1_inst1_O_0;
assign valid_down = NativeMapParallel_n1_inst1_valid_down;
endmodule

module NativeMapParallel_n9_unq4 (input CLK, input [7:0] I_0_0, input [7:0] I_0_1, input [7:0] I_0_2, input [7:0] I_1_0, input [7:0] I_1_1, input [7:0] I_1_2, input [7:0] I_2_0, input [7:0] I_2_1, input [7:0] I_2_2, input [7:0] I_3_0, input [7:0] I_3_1, input [7:0] I_3_2, input [7:0] I_4_0, input [7:0] I_4_1, input [7:0] I_4_2, input [7:0] I_5_0, input [7:0] I_5_1, input [7:0] I_5_2, input [7:0] I_6_0, input [7:0] I_6_1, input [7:0] I_6_2, input [7:0] I_7_0, input [7:0] I_7_1, input [7:0] I_7_2, input [7:0] I_8_0, input [7:0] I_8_1, input [7:0] I_8_2, output [7:0] O_0_0, output [7:0] O_1_0, output [7:0] O_2_0, output [7:0] O_3_0, output [7:0] O_4_0, output [7:0] O_5_0, output [7:0] O_6_0, output [7:0] O_7_0, output [7:0] O_8_0, output valid_down, input valid_up);
wire [7:0] Module_1_inst0_O_0;
wire Module_1_inst0_valid_down;
wire [7:0] Module_1_inst1_O_0;
wire Module_1_inst1_valid_down;
wire [7:0] Module_1_inst2_O_0;
wire Module_1_inst2_valid_down;
wire [7:0] Module_1_inst3_O_0;
wire Module_1_inst3_valid_down;
wire [7:0] Module_1_inst4_O_0;
wire Module_1_inst4_valid_down;
wire [7:0] Module_1_inst5_O_0;
wire Module_1_inst5_valid_down;
wire [7:0] Module_1_inst6_O_0;
wire Module_1_inst6_valid_down;
wire [7:0] Module_1_inst7_O_0;
wire Module_1_inst7_valid_down;
wire [7:0] Module_1_inst8_O_0;
wire Module_1_inst8_valid_down;
wire and_inst0_out;
wire and_inst1_out;
wire and_inst2_out;
wire and_inst3_out;
wire and_inst4_out;
wire and_inst5_out;
wire and_inst6_out;
wire and_inst7_out;
Module_1 Module_1_inst0(.CLK(CLK), .I_0(I_0_0), .I_1(I_0_1), .I_2(I_0_2), .O_0(Module_1_inst0_O_0), .valid_down(Module_1_inst0_valid_down), .valid_up(valid_up));
Module_1 Module_1_inst1(.CLK(CLK), .I_0(I_1_0), .I_1(I_1_1), .I_2(I_1_2), .O_0(Module_1_inst1_O_0), .valid_down(Module_1_inst1_valid_down), .valid_up(valid_up));
Module_1 Module_1_inst2(.CLK(CLK), .I_0(I_2_0), .I_1(I_2_1), .I_2(I_2_2), .O_0(Module_1_inst2_O_0), .valid_down(Module_1_inst2_valid_down), .valid_up(valid_up));
Module_1 Module_1_inst3(.CLK(CLK), .I_0(I_3_0), .I_1(I_3_1), .I_2(I_3_2), .O_0(Module_1_inst3_O_0), .valid_down(Module_1_inst3_valid_down), .valid_up(valid_up));
Module_1 Module_1_inst4(.CLK(CLK), .I_0(I_4_0), .I_1(I_4_1), .I_2(I_4_2), .O_0(Module_1_inst4_O_0), .valid_down(Module_1_inst4_valid_down), .valid_up(valid_up));
Module_1 Module_1_inst5(.CLK(CLK), .I_0(I_5_0), .I_1(I_5_1), .I_2(I_5_2), .O_0(Module_1_inst5_O_0), .valid_down(Module_1_inst5_valid_down), .valid_up(valid_up));
Module_1 Module_1_inst6(.CLK(CLK), .I_0(I_6_0), .I_1(I_6_1), .I_2(I_6_2), .O_0(Module_1_inst6_O_0), .valid_down(Module_1_inst6_valid_down), .valid_up(valid_up));
Module_1 Module_1_inst7(.CLK(CLK), .I_0(I_7_0), .I_1(I_7_1), .I_2(I_7_2), .O_0(Module_1_inst7_O_0), .valid_down(Module_1_inst7_valid_down), .valid_up(valid_up));
Module_1 Module_1_inst8(.CLK(CLK), .I_0(I_8_0), .I_1(I_8_1), .I_2(I_8_2), .O_0(Module_1_inst8_O_0), .valid_down(Module_1_inst8_valid_down), .valid_up(valid_up));
corebit_and and_inst0(.in0(Module_1_inst0_valid_down), .in1(Module_1_inst1_valid_down), .out(and_inst0_out));
corebit_and and_inst1(.in0(and_inst0_out), .in1(Module_1_inst2_valid_down), .out(and_inst1_out));
corebit_and and_inst2(.in0(and_inst1_out), .in1(Module_1_inst3_valid_down), .out(and_inst2_out));
corebit_and and_inst3(.in0(and_inst2_out), .in1(Module_1_inst4_valid_down), .out(and_inst3_out));
corebit_and and_inst4(.in0(and_inst3_out), .in1(Module_1_inst5_valid_down), .out(and_inst4_out));
corebit_and and_inst5(.in0(and_inst4_out), .in1(Module_1_inst6_valid_down), .out(and_inst5_out));
corebit_and and_inst6(.in0(and_inst5_out), .in1(Module_1_inst7_valid_down), .out(and_inst6_out));
corebit_and and_inst7(.in0(and_inst6_out), .in1(Module_1_inst8_valid_down), .out(and_inst7_out));
assign O_0_0 = Module_1_inst0_O_0;
assign O_1_0 = Module_1_inst1_O_0;
assign O_2_0 = Module_1_inst2_O_0;
assign O_3_0 = Module_1_inst3_O_0;
assign O_4_0 = Module_1_inst4_O_0;
assign O_5_0 = Module_1_inst5_O_0;
assign O_6_0 = Module_1_inst6_O_0;
assign O_7_0 = Module_1_inst7_O_0;
assign O_8_0 = Module_1_inst8_O_0;
assign valid_down = and_inst7_out;
endmodule

module Module_0 (input CLK, input [7:0] I_0, input [7:0] I_1, input [7:0] I_2, output [7:0] O_0, output valid_down, input valid_up);
wire [7:0] Const_tSSeq_1_Int__hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0;
wire Const_tSSeq_1_Int__hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down;
wire [7:0] Const_tSSeq_3_Int__hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0;
wire [7:0] Const_tSSeq_3_Int__hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_1;
wire [7:0] Const_tSSeq_3_Int__hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_2;
wire Const_tSSeq_3_Int__hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down;
wire [7:0] NativeMapParallel_n1_inst0_O_0__0;
wire [7:0] NativeMapParallel_n1_inst0_O_0__1;
wire NativeMapParallel_n1_inst0_valid_down;
wire [7:0] NativeMapParallel_n1_inst1_O_0;
wire NativeMapParallel_n1_inst1_valid_down;
wire [7:0] NativeMapParallel_n3_inst0_O_0__0;
wire [7:0] NativeMapParallel_n3_inst0_O_0__1;
wire [7:0] NativeMapParallel_n3_inst0_O_1__0;
wire [7:0] NativeMapParallel_n3_inst0_O_1__1;
wire [7:0] NativeMapParallel_n3_inst0_O_2__0;
wire [7:0] NativeMapParallel_n3_inst0_O_2__1;
wire NativeMapParallel_n3_inst0_valid_down;
wire [7:0] NativeMapParallel_n3_inst1_O_0;
wire [7:0] NativeMapParallel_n3_inst1_O_1;
wire [7:0] NativeMapParallel_n3_inst1_O_2;
wire NativeMapParallel_n3_inst1_valid_down;
wire [7:0] Reduce_S_n3_inst0_O_0;
wire Reduce_S_n3_inst0_valid_down;
wire and_inst0_out;
wire and_inst1_out;
Const_tSSeq_1_Int__hasCEFalse_hasResetFalse_hasValidTrue Const_tSSeq_1_Int__hasCEFalse_hasResetFalse_hasValidTrue_inst0(.CLK(CLK), .O_0(Const_tSSeq_1_Int__hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0), .valid_down(Const_tSSeq_1_Int__hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down), .valid_up(valid_up));
Const_tSSeq_3_Int__hasCEFalse_hasResetFalse_hasValidTrue Const_tSSeq_3_Int__hasCEFalse_hasResetFalse_hasValidTrue_inst0(.CLK(CLK), .O_0(Const_tSSeq_3_Int__hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0), .O_1(Const_tSSeq_3_Int__hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_1), .O_2(Const_tSSeq_3_Int__hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_2), .valid_down(Const_tSSeq_3_Int__hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down), .valid_up(valid_up));
NativeMapParallel_n1_unq2 NativeMapParallel_n1_inst0(.I0_0(Reduce_S_n3_inst0_O_0), .I1_0(Const_tSSeq_1_Int__hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0), .O_0__0(NativeMapParallel_n1_inst0_O_0__0), .O_0__1(NativeMapParallel_n1_inst0_O_0__1), .valid_down(NativeMapParallel_n1_inst0_valid_down), .valid_up(and_inst1_out));
NativeMapParallel_n1_unq3 NativeMapParallel_n1_inst1(.I_0__0(NativeMapParallel_n1_inst0_O_0__0), .I_0__1(NativeMapParallel_n1_inst0_O_0__1), .O_0(NativeMapParallel_n1_inst1_O_0), .valid_down(NativeMapParallel_n1_inst1_valid_down), .valid_up(NativeMapParallel_n1_inst0_valid_down));
NativeMapParallel_n3 NativeMapParallel_n3_inst0(.I0_0(I_0), .I0_1(I_1), .I0_2(I_2), .I1_0(Const_tSSeq_3_Int__hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0), .I1_1(Const_tSSeq_3_Int__hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_1), .I1_2(Const_tSSeq_3_Int__hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_2), .O_0__0(NativeMapParallel_n3_inst0_O_0__0), .O_0__1(NativeMapParallel_n3_inst0_O_0__1), .O_1__0(NativeMapParallel_n3_inst0_O_1__0), .O_1__1(NativeMapParallel_n3_inst0_O_1__1), .O_2__0(NativeMapParallel_n3_inst0_O_2__0), .O_2__1(NativeMapParallel_n3_inst0_O_2__1), .valid_down(NativeMapParallel_n3_inst0_valid_down), .valid_up(and_inst0_out));
NativeMapParallel_n3_unq1 NativeMapParallel_n3_inst1(.I_0__0(NativeMapParallel_n3_inst0_O_0__0), .I_0__1(NativeMapParallel_n3_inst0_O_0__1), .I_1__0(NativeMapParallel_n3_inst0_O_1__0), .I_1__1(NativeMapParallel_n3_inst0_O_1__1), .I_2__0(NativeMapParallel_n3_inst0_O_2__0), .I_2__1(NativeMapParallel_n3_inst0_O_2__1), .O_0(NativeMapParallel_n3_inst1_O_0), .O_1(NativeMapParallel_n3_inst1_O_1), .O_2(NativeMapParallel_n3_inst1_O_2), .valid_down(NativeMapParallel_n3_inst1_valid_down), .valid_up(NativeMapParallel_n3_inst0_valid_down));
Reduce_S_n3 Reduce_S_n3_inst0(.CLK(CLK), .I_0(NativeMapParallel_n3_inst1_O_0), .I_1(NativeMapParallel_n3_inst1_O_1), .I_2(NativeMapParallel_n3_inst1_O_2), .O_0(Reduce_S_n3_inst0_O_0), .valid_down(Reduce_S_n3_inst0_valid_down), .valid_up(NativeMapParallel_n3_inst1_valid_down));
corebit_and and_inst0(.in0(valid_up), .in1(Const_tSSeq_3_Int__hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down), .out(and_inst0_out));
corebit_and and_inst1(.in0(Reduce_S_n3_inst0_valid_down), .in1(Const_tSSeq_1_Int__hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down), .out(and_inst1_out));
assign O_0 = NativeMapParallel_n1_inst1_O_0;
assign valid_down = NativeMapParallel_n1_inst1_valid_down;
endmodule

module NativeMapParallel_n27_unq3 (input CLK, input [7:0] I_0_0, input [7:0] I_0_1, input [7:0] I_0_2, input [7:0] I_10_0, input [7:0] I_10_1, input [7:0] I_10_2, input [7:0] I_11_0, input [7:0] I_11_1, input [7:0] I_11_2, input [7:0] I_12_0, input [7:0] I_12_1, input [7:0] I_12_2, input [7:0] I_13_0, input [7:0] I_13_1, input [7:0] I_13_2, input [7:0] I_14_0, input [7:0] I_14_1, input [7:0] I_14_2, input [7:0] I_15_0, input [7:0] I_15_1, input [7:0] I_15_2, input [7:0] I_16_0, input [7:0] I_16_1, input [7:0] I_16_2, input [7:0] I_17_0, input [7:0] I_17_1, input [7:0] I_17_2, input [7:0] I_18_0, input [7:0] I_18_1, input [7:0] I_18_2, input [7:0] I_19_0, input [7:0] I_19_1, input [7:0] I_19_2, input [7:0] I_1_0, input [7:0] I_1_1, input [7:0] I_1_2, input [7:0] I_20_0, input [7:0] I_20_1, input [7:0] I_20_2, input [7:0] I_21_0, input [7:0] I_21_1, input [7:0] I_21_2, input [7:0] I_22_0, input [7:0] I_22_1, input [7:0] I_22_2, input [7:0] I_23_0, input [7:0] I_23_1, input [7:0] I_23_2, input [7:0] I_24_0, input [7:0] I_24_1, input [7:0] I_24_2, input [7:0] I_25_0, input [7:0] I_25_1, input [7:0] I_25_2, input [7:0] I_26_0, input [7:0] I_26_1, input [7:0] I_26_2, input [7:0] I_2_0, input [7:0] I_2_1, input [7:0] I_2_2, input [7:0] I_3_0, input [7:0] I_3_1, input [7:0] I_3_2, input [7:0] I_4_0, input [7:0] I_4_1, input [7:0] I_4_2, input [7:0] I_5_0, input [7:0] I_5_1, input [7:0] I_5_2, input [7:0] I_6_0, input [7:0] I_6_1, input [7:0] I_6_2, input [7:0] I_7_0, input [7:0] I_7_1, input [7:0] I_7_2, input [7:0] I_8_0, input [7:0] I_8_1, input [7:0] I_8_2, input [7:0] I_9_0, input [7:0] I_9_1, input [7:0] I_9_2, output [7:0] O_0_0, output [7:0] O_10_0, output [7:0] O_11_0, output [7:0] O_12_0, output [7:0] O_13_0, output [7:0] O_14_0, output [7:0] O_15_0, output [7:0] O_16_0, output [7:0] O_17_0, output [7:0] O_18_0, output [7:0] O_19_0, output [7:0] O_1_0, output [7:0] O_20_0, output [7:0] O_21_0, output [7:0] O_22_0, output [7:0] O_23_0, output [7:0] O_24_0, output [7:0] O_25_0, output [7:0] O_26_0, output [7:0] O_2_0, output [7:0] O_3_0, output [7:0] O_4_0, output [7:0] O_5_0, output [7:0] O_6_0, output [7:0] O_7_0, output [7:0] O_8_0, output [7:0] O_9_0, output valid_down, input valid_up);
wire [7:0] Module_0_inst0_O_0;
wire Module_0_inst0_valid_down;
wire [7:0] Module_0_inst1_O_0;
wire Module_0_inst1_valid_down;
wire [7:0] Module_0_inst10_O_0;
wire Module_0_inst10_valid_down;
wire [7:0] Module_0_inst11_O_0;
wire Module_0_inst11_valid_down;
wire [7:0] Module_0_inst12_O_0;
wire Module_0_inst12_valid_down;
wire [7:0] Module_0_inst13_O_0;
wire Module_0_inst13_valid_down;
wire [7:0] Module_0_inst14_O_0;
wire Module_0_inst14_valid_down;
wire [7:0] Module_0_inst15_O_0;
wire Module_0_inst15_valid_down;
wire [7:0] Module_0_inst16_O_0;
wire Module_0_inst16_valid_down;
wire [7:0] Module_0_inst17_O_0;
wire Module_0_inst17_valid_down;
wire [7:0] Module_0_inst18_O_0;
wire Module_0_inst18_valid_down;
wire [7:0] Module_0_inst19_O_0;
wire Module_0_inst19_valid_down;
wire [7:0] Module_0_inst2_O_0;
wire Module_0_inst2_valid_down;
wire [7:0] Module_0_inst20_O_0;
wire Module_0_inst20_valid_down;
wire [7:0] Module_0_inst21_O_0;
wire Module_0_inst21_valid_down;
wire [7:0] Module_0_inst22_O_0;
wire Module_0_inst22_valid_down;
wire [7:0] Module_0_inst23_O_0;
wire Module_0_inst23_valid_down;
wire [7:0] Module_0_inst24_O_0;
wire Module_0_inst24_valid_down;
wire [7:0] Module_0_inst25_O_0;
wire Module_0_inst25_valid_down;
wire [7:0] Module_0_inst26_O_0;
wire Module_0_inst26_valid_down;
wire [7:0] Module_0_inst3_O_0;
wire Module_0_inst3_valid_down;
wire [7:0] Module_0_inst4_O_0;
wire Module_0_inst4_valid_down;
wire [7:0] Module_0_inst5_O_0;
wire Module_0_inst5_valid_down;
wire [7:0] Module_0_inst6_O_0;
wire Module_0_inst6_valid_down;
wire [7:0] Module_0_inst7_O_0;
wire Module_0_inst7_valid_down;
wire [7:0] Module_0_inst8_O_0;
wire Module_0_inst8_valid_down;
wire [7:0] Module_0_inst9_O_0;
wire Module_0_inst9_valid_down;
wire and_inst0_out;
wire and_inst1_out;
wire and_inst10_out;
wire and_inst11_out;
wire and_inst12_out;
wire and_inst13_out;
wire and_inst14_out;
wire and_inst15_out;
wire and_inst16_out;
wire and_inst17_out;
wire and_inst18_out;
wire and_inst19_out;
wire and_inst2_out;
wire and_inst20_out;
wire and_inst21_out;
wire and_inst22_out;
wire and_inst23_out;
wire and_inst24_out;
wire and_inst25_out;
wire and_inst3_out;
wire and_inst4_out;
wire and_inst5_out;
wire and_inst6_out;
wire and_inst7_out;
wire and_inst8_out;
wire and_inst9_out;
Module_0 Module_0_inst0(.CLK(CLK), .I_0(I_0_0), .I_1(I_0_1), .I_2(I_0_2), .O_0(Module_0_inst0_O_0), .valid_down(Module_0_inst0_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst1(.CLK(CLK), .I_0(I_1_0), .I_1(I_1_1), .I_2(I_1_2), .O_0(Module_0_inst1_O_0), .valid_down(Module_0_inst1_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst10(.CLK(CLK), .I_0(I_10_0), .I_1(I_10_1), .I_2(I_10_2), .O_0(Module_0_inst10_O_0), .valid_down(Module_0_inst10_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst11(.CLK(CLK), .I_0(I_11_0), .I_1(I_11_1), .I_2(I_11_2), .O_0(Module_0_inst11_O_0), .valid_down(Module_0_inst11_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst12(.CLK(CLK), .I_0(I_12_0), .I_1(I_12_1), .I_2(I_12_2), .O_0(Module_0_inst12_O_0), .valid_down(Module_0_inst12_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst13(.CLK(CLK), .I_0(I_13_0), .I_1(I_13_1), .I_2(I_13_2), .O_0(Module_0_inst13_O_0), .valid_down(Module_0_inst13_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst14(.CLK(CLK), .I_0(I_14_0), .I_1(I_14_1), .I_2(I_14_2), .O_0(Module_0_inst14_O_0), .valid_down(Module_0_inst14_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst15(.CLK(CLK), .I_0(I_15_0), .I_1(I_15_1), .I_2(I_15_2), .O_0(Module_0_inst15_O_0), .valid_down(Module_0_inst15_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst16(.CLK(CLK), .I_0(I_16_0), .I_1(I_16_1), .I_2(I_16_2), .O_0(Module_0_inst16_O_0), .valid_down(Module_0_inst16_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst17(.CLK(CLK), .I_0(I_17_0), .I_1(I_17_1), .I_2(I_17_2), .O_0(Module_0_inst17_O_0), .valid_down(Module_0_inst17_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst18(.CLK(CLK), .I_0(I_18_0), .I_1(I_18_1), .I_2(I_18_2), .O_0(Module_0_inst18_O_0), .valid_down(Module_0_inst18_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst19(.CLK(CLK), .I_0(I_19_0), .I_1(I_19_1), .I_2(I_19_2), .O_0(Module_0_inst19_O_0), .valid_down(Module_0_inst19_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst2(.CLK(CLK), .I_0(I_2_0), .I_1(I_2_1), .I_2(I_2_2), .O_0(Module_0_inst2_O_0), .valid_down(Module_0_inst2_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst20(.CLK(CLK), .I_0(I_20_0), .I_1(I_20_1), .I_2(I_20_2), .O_0(Module_0_inst20_O_0), .valid_down(Module_0_inst20_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst21(.CLK(CLK), .I_0(I_21_0), .I_1(I_21_1), .I_2(I_21_2), .O_0(Module_0_inst21_O_0), .valid_down(Module_0_inst21_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst22(.CLK(CLK), .I_0(I_22_0), .I_1(I_22_1), .I_2(I_22_2), .O_0(Module_0_inst22_O_0), .valid_down(Module_0_inst22_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst23(.CLK(CLK), .I_0(I_23_0), .I_1(I_23_1), .I_2(I_23_2), .O_0(Module_0_inst23_O_0), .valid_down(Module_0_inst23_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst24(.CLK(CLK), .I_0(I_24_0), .I_1(I_24_1), .I_2(I_24_2), .O_0(Module_0_inst24_O_0), .valid_down(Module_0_inst24_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst25(.CLK(CLK), .I_0(I_25_0), .I_1(I_25_1), .I_2(I_25_2), .O_0(Module_0_inst25_O_0), .valid_down(Module_0_inst25_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst26(.CLK(CLK), .I_0(I_26_0), .I_1(I_26_1), .I_2(I_26_2), .O_0(Module_0_inst26_O_0), .valid_down(Module_0_inst26_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst3(.CLK(CLK), .I_0(I_3_0), .I_1(I_3_1), .I_2(I_3_2), .O_0(Module_0_inst3_O_0), .valid_down(Module_0_inst3_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst4(.CLK(CLK), .I_0(I_4_0), .I_1(I_4_1), .I_2(I_4_2), .O_0(Module_0_inst4_O_0), .valid_down(Module_0_inst4_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst5(.CLK(CLK), .I_0(I_5_0), .I_1(I_5_1), .I_2(I_5_2), .O_0(Module_0_inst5_O_0), .valid_down(Module_0_inst5_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst6(.CLK(CLK), .I_0(I_6_0), .I_1(I_6_1), .I_2(I_6_2), .O_0(Module_0_inst6_O_0), .valid_down(Module_0_inst6_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst7(.CLK(CLK), .I_0(I_7_0), .I_1(I_7_1), .I_2(I_7_2), .O_0(Module_0_inst7_O_0), .valid_down(Module_0_inst7_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst8(.CLK(CLK), .I_0(I_8_0), .I_1(I_8_1), .I_2(I_8_2), .O_0(Module_0_inst8_O_0), .valid_down(Module_0_inst8_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst9(.CLK(CLK), .I_0(I_9_0), .I_1(I_9_1), .I_2(I_9_2), .O_0(Module_0_inst9_O_0), .valid_down(Module_0_inst9_valid_down), .valid_up(valid_up));
corebit_and and_inst0(.in0(Module_0_inst0_valid_down), .in1(Module_0_inst1_valid_down), .out(and_inst0_out));
corebit_and and_inst1(.in0(and_inst0_out), .in1(Module_0_inst2_valid_down), .out(and_inst1_out));
corebit_and and_inst10(.in0(and_inst9_out), .in1(Module_0_inst11_valid_down), .out(and_inst10_out));
corebit_and and_inst11(.in0(and_inst10_out), .in1(Module_0_inst12_valid_down), .out(and_inst11_out));
corebit_and and_inst12(.in0(and_inst11_out), .in1(Module_0_inst13_valid_down), .out(and_inst12_out));
corebit_and and_inst13(.in0(and_inst12_out), .in1(Module_0_inst14_valid_down), .out(and_inst13_out));
corebit_and and_inst14(.in0(and_inst13_out), .in1(Module_0_inst15_valid_down), .out(and_inst14_out));
corebit_and and_inst15(.in0(and_inst14_out), .in1(Module_0_inst16_valid_down), .out(and_inst15_out));
corebit_and and_inst16(.in0(and_inst15_out), .in1(Module_0_inst17_valid_down), .out(and_inst16_out));
corebit_and and_inst17(.in0(and_inst16_out), .in1(Module_0_inst18_valid_down), .out(and_inst17_out));
corebit_and and_inst18(.in0(and_inst17_out), .in1(Module_0_inst19_valid_down), .out(and_inst18_out));
corebit_and and_inst19(.in0(and_inst18_out), .in1(Module_0_inst20_valid_down), .out(and_inst19_out));
corebit_and and_inst2(.in0(and_inst1_out), .in1(Module_0_inst3_valid_down), .out(and_inst2_out));
corebit_and and_inst20(.in0(and_inst19_out), .in1(Module_0_inst21_valid_down), .out(and_inst20_out));
corebit_and and_inst21(.in0(and_inst20_out), .in1(Module_0_inst22_valid_down), .out(and_inst21_out));
corebit_and and_inst22(.in0(and_inst21_out), .in1(Module_0_inst23_valid_down), .out(and_inst22_out));
corebit_and and_inst23(.in0(and_inst22_out), .in1(Module_0_inst24_valid_down), .out(and_inst23_out));
corebit_and and_inst24(.in0(and_inst23_out), .in1(Module_0_inst25_valid_down), .out(and_inst24_out));
corebit_and and_inst25(.in0(and_inst24_out), .in1(Module_0_inst26_valid_down), .out(and_inst25_out));
corebit_and and_inst3(.in0(and_inst2_out), .in1(Module_0_inst4_valid_down), .out(and_inst3_out));
corebit_and and_inst4(.in0(and_inst3_out), .in1(Module_0_inst5_valid_down), .out(and_inst4_out));
corebit_and and_inst5(.in0(and_inst4_out), .in1(Module_0_inst6_valid_down), .out(and_inst5_out));
corebit_and and_inst6(.in0(and_inst5_out), .in1(Module_0_inst7_valid_down), .out(and_inst6_out));
corebit_and and_inst7(.in0(and_inst6_out), .in1(Module_0_inst8_valid_down), .out(and_inst7_out));
corebit_and and_inst8(.in0(and_inst7_out), .in1(Module_0_inst9_valid_down), .out(and_inst8_out));
corebit_and and_inst9(.in0(and_inst8_out), .in1(Module_0_inst10_valid_down), .out(and_inst9_out));
assign O_0_0 = Module_0_inst0_O_0;
assign O_10_0 = Module_0_inst10_O_0;
assign O_11_0 = Module_0_inst11_O_0;
assign O_12_0 = Module_0_inst12_O_0;
assign O_13_0 = Module_0_inst13_O_0;
assign O_14_0 = Module_0_inst14_O_0;
assign O_15_0 = Module_0_inst15_O_0;
assign O_16_0 = Module_0_inst16_O_0;
assign O_17_0 = Module_0_inst17_O_0;
assign O_18_0 = Module_0_inst18_O_0;
assign O_19_0 = Module_0_inst19_O_0;
assign O_1_0 = Module_0_inst1_O_0;
assign O_20_0 = Module_0_inst20_O_0;
assign O_21_0 = Module_0_inst21_O_0;
assign O_22_0 = Module_0_inst22_O_0;
assign O_23_0 = Module_0_inst23_O_0;
assign O_24_0 = Module_0_inst24_O_0;
assign O_25_0 = Module_0_inst25_O_0;
assign O_26_0 = Module_0_inst26_O_0;
assign O_2_0 = Module_0_inst2_O_0;
assign O_3_0 = Module_0_inst3_O_0;
assign O_4_0 = Module_0_inst4_O_0;
assign O_5_0 = Module_0_inst5_O_0;
assign O_6_0 = Module_0_inst6_O_0;
assign O_7_0 = Module_0_inst7_O_0;
assign O_8_0 = Module_0_inst8_O_0;
assign O_9_0 = Module_0_inst9_O_0;
assign valid_down = and_inst25_out;
endmodule

module top (input CLK, input [7:0] I_0_0, input [7:0] I_10_0, input [7:0] I_11_0, input [7:0] I_12_0, input [7:0] I_13_0, input [7:0] I_14_0, input [7:0] I_15_0, input [7:0] I_16_0, input [7:0] I_17_0, input [7:0] I_18_0, input [7:0] I_19_0, input [7:0] I_1_0, input [7:0] I_20_0, input [7:0] I_21_0, input [7:0] I_22_0, input [7:0] I_23_0, input [7:0] I_24_0, input [7:0] I_25_0, input [7:0] I_26_0, input [7:0] I_2_0, input [7:0] I_3_0, input [7:0] I_4_0, input [7:0] I_5_0, input [7:0] I_6_0, input [7:0] I_7_0, input [7:0] I_8_0, input [7:0] I_9_0, output [7:0] O_0_0, output [7:0] O_1_0, output [7:0] O_2_0, output valid_down, input valid_up);
wire [7:0] FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0_0;
wire [7:0] FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_10_0;
wire [7:0] FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_11_0;
wire [7:0] FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_12_0;
wire [7:0] FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_13_0;
wire [7:0] FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_14_0;
wire [7:0] FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_15_0;
wire [7:0] FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_16_0;
wire [7:0] FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_17_0;
wire [7:0] FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_18_0;
wire [7:0] FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_19_0;
wire [7:0] FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_1_0;
wire [7:0] FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_20_0;
wire [7:0] FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_21_0;
wire [7:0] FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_22_0;
wire [7:0] FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_23_0;
wire [7:0] FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_24_0;
wire [7:0] FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_25_0;
wire [7:0] FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_26_0;
wire [7:0] FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_2_0;
wire [7:0] FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_3_0;
wire [7:0] FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_4_0;
wire [7:0] FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_5_0;
wire [7:0] FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_6_0;
wire [7:0] FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_7_0;
wire [7:0] FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_8_0;
wire [7:0] FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_9_0;
wire FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down;
wire [7:0] FIFO_tSSeq_3_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0_0;
wire [7:0] FIFO_tSSeq_3_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_1_0;
wire [7:0] FIFO_tSSeq_3_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_2_0;
wire FIFO_tSSeq_3_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down;
wire [7:0] FIFO_tSSeq_3_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_0_0;
wire [7:0] FIFO_tSSeq_3_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_1_0;
wire [7:0] FIFO_tSSeq_3_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_2_0;
wire FIFO_tSSeq_3_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_valid_down;
wire [7:0] FIFO_tSSeq_3_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_0_0;
wire [7:0] FIFO_tSSeq_3_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_1_0;
wire [7:0] FIFO_tSSeq_3_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_2_0;
wire FIFO_tSSeq_3_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_valid_down;
wire [7:0] NativeMapParallel_n27_inst0_O_0_0_0;
wire [7:0] NativeMapParallel_n27_inst0_O_0_0_1;
wire [7:0] NativeMapParallel_n27_inst0_O_10_0_0;
wire [7:0] NativeMapParallel_n27_inst0_O_10_0_1;
wire [7:0] NativeMapParallel_n27_inst0_O_11_0_0;
wire [7:0] NativeMapParallel_n27_inst0_O_11_0_1;
wire [7:0] NativeMapParallel_n27_inst0_O_12_0_0;
wire [7:0] NativeMapParallel_n27_inst0_O_12_0_1;
wire [7:0] NativeMapParallel_n27_inst0_O_13_0_0;
wire [7:0] NativeMapParallel_n27_inst0_O_13_0_1;
wire [7:0] NativeMapParallel_n27_inst0_O_14_0_0;
wire [7:0] NativeMapParallel_n27_inst0_O_14_0_1;
wire [7:0] NativeMapParallel_n27_inst0_O_15_0_0;
wire [7:0] NativeMapParallel_n27_inst0_O_15_0_1;
wire [7:0] NativeMapParallel_n27_inst0_O_16_0_0;
wire [7:0] NativeMapParallel_n27_inst0_O_16_0_1;
wire [7:0] NativeMapParallel_n27_inst0_O_17_0_0;
wire [7:0] NativeMapParallel_n27_inst0_O_17_0_1;
wire [7:0] NativeMapParallel_n27_inst0_O_18_0_0;
wire [7:0] NativeMapParallel_n27_inst0_O_18_0_1;
wire [7:0] NativeMapParallel_n27_inst0_O_19_0_0;
wire [7:0] NativeMapParallel_n27_inst0_O_19_0_1;
wire [7:0] NativeMapParallel_n27_inst0_O_1_0_0;
wire [7:0] NativeMapParallel_n27_inst0_O_1_0_1;
wire [7:0] NativeMapParallel_n27_inst0_O_20_0_0;
wire [7:0] NativeMapParallel_n27_inst0_O_20_0_1;
wire [7:0] NativeMapParallel_n27_inst0_O_21_0_0;
wire [7:0] NativeMapParallel_n27_inst0_O_21_0_1;
wire [7:0] NativeMapParallel_n27_inst0_O_22_0_0;
wire [7:0] NativeMapParallel_n27_inst0_O_22_0_1;
wire [7:0] NativeMapParallel_n27_inst0_O_23_0_0;
wire [7:0] NativeMapParallel_n27_inst0_O_23_0_1;
wire [7:0] NativeMapParallel_n27_inst0_O_24_0_0;
wire [7:0] NativeMapParallel_n27_inst0_O_24_0_1;
wire [7:0] NativeMapParallel_n27_inst0_O_25_0_0;
wire [7:0] NativeMapParallel_n27_inst0_O_25_0_1;
wire [7:0] NativeMapParallel_n27_inst0_O_26_0_0;
wire [7:0] NativeMapParallel_n27_inst0_O_26_0_1;
wire [7:0] NativeMapParallel_n27_inst0_O_2_0_0;
wire [7:0] NativeMapParallel_n27_inst0_O_2_0_1;
wire [7:0] NativeMapParallel_n27_inst0_O_3_0_0;
wire [7:0] NativeMapParallel_n27_inst0_O_3_0_1;
wire [7:0] NativeMapParallel_n27_inst0_O_4_0_0;
wire [7:0] NativeMapParallel_n27_inst0_O_4_0_1;
wire [7:0] NativeMapParallel_n27_inst0_O_5_0_0;
wire [7:0] NativeMapParallel_n27_inst0_O_5_0_1;
wire [7:0] NativeMapParallel_n27_inst0_O_6_0_0;
wire [7:0] NativeMapParallel_n27_inst0_O_6_0_1;
wire [7:0] NativeMapParallel_n27_inst0_O_7_0_0;
wire [7:0] NativeMapParallel_n27_inst0_O_7_0_1;
wire [7:0] NativeMapParallel_n27_inst0_O_8_0_0;
wire [7:0] NativeMapParallel_n27_inst0_O_8_0_1;
wire [7:0] NativeMapParallel_n27_inst0_O_9_0_0;
wire [7:0] NativeMapParallel_n27_inst0_O_9_0_1;
wire NativeMapParallel_n27_inst0_valid_down;
wire [7:0] NativeMapParallel_n27_inst1_O_0_0_0;
wire [7:0] NativeMapParallel_n27_inst1_O_0_0_1;
wire [7:0] NativeMapParallel_n27_inst1_O_0_0_2;
wire [7:0] NativeMapParallel_n27_inst1_O_10_0_0;
wire [7:0] NativeMapParallel_n27_inst1_O_10_0_1;
wire [7:0] NativeMapParallel_n27_inst1_O_10_0_2;
wire [7:0] NativeMapParallel_n27_inst1_O_11_0_0;
wire [7:0] NativeMapParallel_n27_inst1_O_11_0_1;
wire [7:0] NativeMapParallel_n27_inst1_O_11_0_2;
wire [7:0] NativeMapParallel_n27_inst1_O_12_0_0;
wire [7:0] NativeMapParallel_n27_inst1_O_12_0_1;
wire [7:0] NativeMapParallel_n27_inst1_O_12_0_2;
wire [7:0] NativeMapParallel_n27_inst1_O_13_0_0;
wire [7:0] NativeMapParallel_n27_inst1_O_13_0_1;
wire [7:0] NativeMapParallel_n27_inst1_O_13_0_2;
wire [7:0] NativeMapParallel_n27_inst1_O_14_0_0;
wire [7:0] NativeMapParallel_n27_inst1_O_14_0_1;
wire [7:0] NativeMapParallel_n27_inst1_O_14_0_2;
wire [7:0] NativeMapParallel_n27_inst1_O_15_0_0;
wire [7:0] NativeMapParallel_n27_inst1_O_15_0_1;
wire [7:0] NativeMapParallel_n27_inst1_O_15_0_2;
wire [7:0] NativeMapParallel_n27_inst1_O_16_0_0;
wire [7:0] NativeMapParallel_n27_inst1_O_16_0_1;
wire [7:0] NativeMapParallel_n27_inst1_O_16_0_2;
wire [7:0] NativeMapParallel_n27_inst1_O_17_0_0;
wire [7:0] NativeMapParallel_n27_inst1_O_17_0_1;
wire [7:0] NativeMapParallel_n27_inst1_O_17_0_2;
wire [7:0] NativeMapParallel_n27_inst1_O_18_0_0;
wire [7:0] NativeMapParallel_n27_inst1_O_18_0_1;
wire [7:0] NativeMapParallel_n27_inst1_O_18_0_2;
wire [7:0] NativeMapParallel_n27_inst1_O_19_0_0;
wire [7:0] NativeMapParallel_n27_inst1_O_19_0_1;
wire [7:0] NativeMapParallel_n27_inst1_O_19_0_2;
wire [7:0] NativeMapParallel_n27_inst1_O_1_0_0;
wire [7:0] NativeMapParallel_n27_inst1_O_1_0_1;
wire [7:0] NativeMapParallel_n27_inst1_O_1_0_2;
wire [7:0] NativeMapParallel_n27_inst1_O_20_0_0;
wire [7:0] NativeMapParallel_n27_inst1_O_20_0_1;
wire [7:0] NativeMapParallel_n27_inst1_O_20_0_2;
wire [7:0] NativeMapParallel_n27_inst1_O_21_0_0;
wire [7:0] NativeMapParallel_n27_inst1_O_21_0_1;
wire [7:0] NativeMapParallel_n27_inst1_O_21_0_2;
wire [7:0] NativeMapParallel_n27_inst1_O_22_0_0;
wire [7:0] NativeMapParallel_n27_inst1_O_22_0_1;
wire [7:0] NativeMapParallel_n27_inst1_O_22_0_2;
wire [7:0] NativeMapParallel_n27_inst1_O_23_0_0;
wire [7:0] NativeMapParallel_n27_inst1_O_23_0_1;
wire [7:0] NativeMapParallel_n27_inst1_O_23_0_2;
wire [7:0] NativeMapParallel_n27_inst1_O_24_0_0;
wire [7:0] NativeMapParallel_n27_inst1_O_24_0_1;
wire [7:0] NativeMapParallel_n27_inst1_O_24_0_2;
wire [7:0] NativeMapParallel_n27_inst1_O_25_0_0;
wire [7:0] NativeMapParallel_n27_inst1_O_25_0_1;
wire [7:0] NativeMapParallel_n27_inst1_O_25_0_2;
wire [7:0] NativeMapParallel_n27_inst1_O_26_0_0;
wire [7:0] NativeMapParallel_n27_inst1_O_26_0_1;
wire [7:0] NativeMapParallel_n27_inst1_O_26_0_2;
wire [7:0] NativeMapParallel_n27_inst1_O_2_0_0;
wire [7:0] NativeMapParallel_n27_inst1_O_2_0_1;
wire [7:0] NativeMapParallel_n27_inst1_O_2_0_2;
wire [7:0] NativeMapParallel_n27_inst1_O_3_0_0;
wire [7:0] NativeMapParallel_n27_inst1_O_3_0_1;
wire [7:0] NativeMapParallel_n27_inst1_O_3_0_2;
wire [7:0] NativeMapParallel_n27_inst1_O_4_0_0;
wire [7:0] NativeMapParallel_n27_inst1_O_4_0_1;
wire [7:0] NativeMapParallel_n27_inst1_O_4_0_2;
wire [7:0] NativeMapParallel_n27_inst1_O_5_0_0;
wire [7:0] NativeMapParallel_n27_inst1_O_5_0_1;
wire [7:0] NativeMapParallel_n27_inst1_O_5_0_2;
wire [7:0] NativeMapParallel_n27_inst1_O_6_0_0;
wire [7:0] NativeMapParallel_n27_inst1_O_6_0_1;
wire [7:0] NativeMapParallel_n27_inst1_O_6_0_2;
wire [7:0] NativeMapParallel_n27_inst1_O_7_0_0;
wire [7:0] NativeMapParallel_n27_inst1_O_7_0_1;
wire [7:0] NativeMapParallel_n27_inst1_O_7_0_2;
wire [7:0] NativeMapParallel_n27_inst1_O_8_0_0;
wire [7:0] NativeMapParallel_n27_inst1_O_8_0_1;
wire [7:0] NativeMapParallel_n27_inst1_O_8_0_2;
wire [7:0] NativeMapParallel_n27_inst1_O_9_0_0;
wire [7:0] NativeMapParallel_n27_inst1_O_9_0_1;
wire [7:0] NativeMapParallel_n27_inst1_O_9_0_2;
wire NativeMapParallel_n27_inst1_valid_down;
wire [7:0] NativeMapParallel_n27_inst2_O_0_0;
wire [7:0] NativeMapParallel_n27_inst2_O_0_1;
wire [7:0] NativeMapParallel_n27_inst2_O_0_2;
wire [7:0] NativeMapParallel_n27_inst2_O_10_0;
wire [7:0] NativeMapParallel_n27_inst2_O_10_1;
wire [7:0] NativeMapParallel_n27_inst2_O_10_2;
wire [7:0] NativeMapParallel_n27_inst2_O_11_0;
wire [7:0] NativeMapParallel_n27_inst2_O_11_1;
wire [7:0] NativeMapParallel_n27_inst2_O_11_2;
wire [7:0] NativeMapParallel_n27_inst2_O_12_0;
wire [7:0] NativeMapParallel_n27_inst2_O_12_1;
wire [7:0] NativeMapParallel_n27_inst2_O_12_2;
wire [7:0] NativeMapParallel_n27_inst2_O_13_0;
wire [7:0] NativeMapParallel_n27_inst2_O_13_1;
wire [7:0] NativeMapParallel_n27_inst2_O_13_2;
wire [7:0] NativeMapParallel_n27_inst2_O_14_0;
wire [7:0] NativeMapParallel_n27_inst2_O_14_1;
wire [7:0] NativeMapParallel_n27_inst2_O_14_2;
wire [7:0] NativeMapParallel_n27_inst2_O_15_0;
wire [7:0] NativeMapParallel_n27_inst2_O_15_1;
wire [7:0] NativeMapParallel_n27_inst2_O_15_2;
wire [7:0] NativeMapParallel_n27_inst2_O_16_0;
wire [7:0] NativeMapParallel_n27_inst2_O_16_1;
wire [7:0] NativeMapParallel_n27_inst2_O_16_2;
wire [7:0] NativeMapParallel_n27_inst2_O_17_0;
wire [7:0] NativeMapParallel_n27_inst2_O_17_1;
wire [7:0] NativeMapParallel_n27_inst2_O_17_2;
wire [7:0] NativeMapParallel_n27_inst2_O_18_0;
wire [7:0] NativeMapParallel_n27_inst2_O_18_1;
wire [7:0] NativeMapParallel_n27_inst2_O_18_2;
wire [7:0] NativeMapParallel_n27_inst2_O_19_0;
wire [7:0] NativeMapParallel_n27_inst2_O_19_1;
wire [7:0] NativeMapParallel_n27_inst2_O_19_2;
wire [7:0] NativeMapParallel_n27_inst2_O_1_0;
wire [7:0] NativeMapParallel_n27_inst2_O_1_1;
wire [7:0] NativeMapParallel_n27_inst2_O_1_2;
wire [7:0] NativeMapParallel_n27_inst2_O_20_0;
wire [7:0] NativeMapParallel_n27_inst2_O_20_1;
wire [7:0] NativeMapParallel_n27_inst2_O_20_2;
wire [7:0] NativeMapParallel_n27_inst2_O_21_0;
wire [7:0] NativeMapParallel_n27_inst2_O_21_1;
wire [7:0] NativeMapParallel_n27_inst2_O_21_2;
wire [7:0] NativeMapParallel_n27_inst2_O_22_0;
wire [7:0] NativeMapParallel_n27_inst2_O_22_1;
wire [7:0] NativeMapParallel_n27_inst2_O_22_2;
wire [7:0] NativeMapParallel_n27_inst2_O_23_0;
wire [7:0] NativeMapParallel_n27_inst2_O_23_1;
wire [7:0] NativeMapParallel_n27_inst2_O_23_2;
wire [7:0] NativeMapParallel_n27_inst2_O_24_0;
wire [7:0] NativeMapParallel_n27_inst2_O_24_1;
wire [7:0] NativeMapParallel_n27_inst2_O_24_2;
wire [7:0] NativeMapParallel_n27_inst2_O_25_0;
wire [7:0] NativeMapParallel_n27_inst2_O_25_1;
wire [7:0] NativeMapParallel_n27_inst2_O_25_2;
wire [7:0] NativeMapParallel_n27_inst2_O_26_0;
wire [7:0] NativeMapParallel_n27_inst2_O_26_1;
wire [7:0] NativeMapParallel_n27_inst2_O_26_2;
wire [7:0] NativeMapParallel_n27_inst2_O_2_0;
wire [7:0] NativeMapParallel_n27_inst2_O_2_1;
wire [7:0] NativeMapParallel_n27_inst2_O_2_2;
wire [7:0] NativeMapParallel_n27_inst2_O_3_0;
wire [7:0] NativeMapParallel_n27_inst2_O_3_1;
wire [7:0] NativeMapParallel_n27_inst2_O_3_2;
wire [7:0] NativeMapParallel_n27_inst2_O_4_0;
wire [7:0] NativeMapParallel_n27_inst2_O_4_1;
wire [7:0] NativeMapParallel_n27_inst2_O_4_2;
wire [7:0] NativeMapParallel_n27_inst2_O_5_0;
wire [7:0] NativeMapParallel_n27_inst2_O_5_1;
wire [7:0] NativeMapParallel_n27_inst2_O_5_2;
wire [7:0] NativeMapParallel_n27_inst2_O_6_0;
wire [7:0] NativeMapParallel_n27_inst2_O_6_1;
wire [7:0] NativeMapParallel_n27_inst2_O_6_2;
wire [7:0] NativeMapParallel_n27_inst2_O_7_0;
wire [7:0] NativeMapParallel_n27_inst2_O_7_1;
wire [7:0] NativeMapParallel_n27_inst2_O_7_2;
wire [7:0] NativeMapParallel_n27_inst2_O_8_0;
wire [7:0] NativeMapParallel_n27_inst2_O_8_1;
wire [7:0] NativeMapParallel_n27_inst2_O_8_2;
wire [7:0] NativeMapParallel_n27_inst2_O_9_0;
wire [7:0] NativeMapParallel_n27_inst2_O_9_1;
wire [7:0] NativeMapParallel_n27_inst2_O_9_2;
wire NativeMapParallel_n27_inst2_valid_down;
wire [7:0] NativeMapParallel_n27_inst3_O_0_0;
wire [7:0] NativeMapParallel_n27_inst3_O_10_0;
wire [7:0] NativeMapParallel_n27_inst3_O_11_0;
wire [7:0] NativeMapParallel_n27_inst3_O_12_0;
wire [7:0] NativeMapParallel_n27_inst3_O_13_0;
wire [7:0] NativeMapParallel_n27_inst3_O_14_0;
wire [7:0] NativeMapParallel_n27_inst3_O_15_0;
wire [7:0] NativeMapParallel_n27_inst3_O_16_0;
wire [7:0] NativeMapParallel_n27_inst3_O_17_0;
wire [7:0] NativeMapParallel_n27_inst3_O_18_0;
wire [7:0] NativeMapParallel_n27_inst3_O_19_0;
wire [7:0] NativeMapParallel_n27_inst3_O_1_0;
wire [7:0] NativeMapParallel_n27_inst3_O_20_0;
wire [7:0] NativeMapParallel_n27_inst3_O_21_0;
wire [7:0] NativeMapParallel_n27_inst3_O_22_0;
wire [7:0] NativeMapParallel_n27_inst3_O_23_0;
wire [7:0] NativeMapParallel_n27_inst3_O_24_0;
wire [7:0] NativeMapParallel_n27_inst3_O_25_0;
wire [7:0] NativeMapParallel_n27_inst3_O_26_0;
wire [7:0] NativeMapParallel_n27_inst3_O_2_0;
wire [7:0] NativeMapParallel_n27_inst3_O_3_0;
wire [7:0] NativeMapParallel_n27_inst3_O_4_0;
wire [7:0] NativeMapParallel_n27_inst3_O_5_0;
wire [7:0] NativeMapParallel_n27_inst3_O_6_0;
wire [7:0] NativeMapParallel_n27_inst3_O_7_0;
wire [7:0] NativeMapParallel_n27_inst3_O_8_0;
wire [7:0] NativeMapParallel_n27_inst3_O_9_0;
wire NativeMapParallel_n27_inst3_valid_down;
wire [7:0] NativeMapParallel_n3_inst0_O_0_0_0;
wire [7:0] NativeMapParallel_n3_inst0_O_1_0_0;
wire [7:0] NativeMapParallel_n3_inst0_O_2_0_0;
wire NativeMapParallel_n3_inst0_valid_down;
wire [7:0] NativeMapParallel_n9_inst0_O_0_0_0;
wire [7:0] NativeMapParallel_n9_inst0_O_1_0_0;
wire [7:0] NativeMapParallel_n9_inst0_O_2_0_0;
wire [7:0] NativeMapParallel_n9_inst0_O_3_0_0;
wire [7:0] NativeMapParallel_n9_inst0_O_4_0_0;
wire [7:0] NativeMapParallel_n9_inst0_O_5_0_0;
wire [7:0] NativeMapParallel_n9_inst0_O_6_0_0;
wire [7:0] NativeMapParallel_n9_inst0_O_7_0_0;
wire [7:0] NativeMapParallel_n9_inst0_O_8_0_0;
wire NativeMapParallel_n9_inst0_valid_down;
wire [7:0] NativeMapParallel_n9_inst1_O_0_0_0;
wire [7:0] NativeMapParallel_n9_inst1_O_0_0_1;
wire [7:0] NativeMapParallel_n9_inst1_O_1_0_0;
wire [7:0] NativeMapParallel_n9_inst1_O_1_0_1;
wire [7:0] NativeMapParallel_n9_inst1_O_2_0_0;
wire [7:0] NativeMapParallel_n9_inst1_O_2_0_1;
wire [7:0] NativeMapParallel_n9_inst1_O_3_0_0;
wire [7:0] NativeMapParallel_n9_inst1_O_3_0_1;
wire [7:0] NativeMapParallel_n9_inst1_O_4_0_0;
wire [7:0] NativeMapParallel_n9_inst1_O_4_0_1;
wire [7:0] NativeMapParallel_n9_inst1_O_5_0_0;
wire [7:0] NativeMapParallel_n9_inst1_O_5_0_1;
wire [7:0] NativeMapParallel_n9_inst1_O_6_0_0;
wire [7:0] NativeMapParallel_n9_inst1_O_6_0_1;
wire [7:0] NativeMapParallel_n9_inst1_O_7_0_0;
wire [7:0] NativeMapParallel_n9_inst1_O_7_0_1;
wire [7:0] NativeMapParallel_n9_inst1_O_8_0_0;
wire [7:0] NativeMapParallel_n9_inst1_O_8_0_1;
wire NativeMapParallel_n9_inst1_valid_down;
wire [7:0] NativeMapParallel_n9_inst2_O_0_0_0;
wire [7:0] NativeMapParallel_n9_inst2_O_0_0_1;
wire [7:0] NativeMapParallel_n9_inst2_O_0_0_2;
wire [7:0] NativeMapParallel_n9_inst2_O_1_0_0;
wire [7:0] NativeMapParallel_n9_inst2_O_1_0_1;
wire [7:0] NativeMapParallel_n9_inst2_O_1_0_2;
wire [7:0] NativeMapParallel_n9_inst2_O_2_0_0;
wire [7:0] NativeMapParallel_n9_inst2_O_2_0_1;
wire [7:0] NativeMapParallel_n9_inst2_O_2_0_2;
wire [7:0] NativeMapParallel_n9_inst2_O_3_0_0;
wire [7:0] NativeMapParallel_n9_inst2_O_3_0_1;
wire [7:0] NativeMapParallel_n9_inst2_O_3_0_2;
wire [7:0] NativeMapParallel_n9_inst2_O_4_0_0;
wire [7:0] NativeMapParallel_n9_inst2_O_4_0_1;
wire [7:0] NativeMapParallel_n9_inst2_O_4_0_2;
wire [7:0] NativeMapParallel_n9_inst2_O_5_0_0;
wire [7:0] NativeMapParallel_n9_inst2_O_5_0_1;
wire [7:0] NativeMapParallel_n9_inst2_O_5_0_2;
wire [7:0] NativeMapParallel_n9_inst2_O_6_0_0;
wire [7:0] NativeMapParallel_n9_inst2_O_6_0_1;
wire [7:0] NativeMapParallel_n9_inst2_O_6_0_2;
wire [7:0] NativeMapParallel_n9_inst2_O_7_0_0;
wire [7:0] NativeMapParallel_n9_inst2_O_7_0_1;
wire [7:0] NativeMapParallel_n9_inst2_O_7_0_2;
wire [7:0] NativeMapParallel_n9_inst2_O_8_0_0;
wire [7:0] NativeMapParallel_n9_inst2_O_8_0_1;
wire [7:0] NativeMapParallel_n9_inst2_O_8_0_2;
wire NativeMapParallel_n9_inst2_valid_down;
wire [7:0] NativeMapParallel_n9_inst3_O_0_0;
wire [7:0] NativeMapParallel_n9_inst3_O_0_1;
wire [7:0] NativeMapParallel_n9_inst3_O_0_2;
wire [7:0] NativeMapParallel_n9_inst3_O_1_0;
wire [7:0] NativeMapParallel_n9_inst3_O_1_1;
wire [7:0] NativeMapParallel_n9_inst3_O_1_2;
wire [7:0] NativeMapParallel_n9_inst3_O_2_0;
wire [7:0] NativeMapParallel_n9_inst3_O_2_1;
wire [7:0] NativeMapParallel_n9_inst3_O_2_2;
wire [7:0] NativeMapParallel_n9_inst3_O_3_0;
wire [7:0] NativeMapParallel_n9_inst3_O_3_1;
wire [7:0] NativeMapParallel_n9_inst3_O_3_2;
wire [7:0] NativeMapParallel_n9_inst3_O_4_0;
wire [7:0] NativeMapParallel_n9_inst3_O_4_1;
wire [7:0] NativeMapParallel_n9_inst3_O_4_2;
wire [7:0] NativeMapParallel_n9_inst3_O_5_0;
wire [7:0] NativeMapParallel_n9_inst3_O_5_1;
wire [7:0] NativeMapParallel_n9_inst3_O_5_2;
wire [7:0] NativeMapParallel_n9_inst3_O_6_0;
wire [7:0] NativeMapParallel_n9_inst3_O_6_1;
wire [7:0] NativeMapParallel_n9_inst3_O_6_2;
wire [7:0] NativeMapParallel_n9_inst3_O_7_0;
wire [7:0] NativeMapParallel_n9_inst3_O_7_1;
wire [7:0] NativeMapParallel_n9_inst3_O_7_2;
wire [7:0] NativeMapParallel_n9_inst3_O_8_0;
wire [7:0] NativeMapParallel_n9_inst3_O_8_1;
wire [7:0] NativeMapParallel_n9_inst3_O_8_2;
wire NativeMapParallel_n9_inst3_valid_down;
wire [7:0] NativeMapParallel_n9_inst4_O_0_0;
wire [7:0] NativeMapParallel_n9_inst4_O_1_0;
wire [7:0] NativeMapParallel_n9_inst4_O_2_0;
wire [7:0] NativeMapParallel_n9_inst4_O_3_0;
wire [7:0] NativeMapParallel_n9_inst4_O_4_0;
wire [7:0] NativeMapParallel_n9_inst4_O_5_0;
wire [7:0] NativeMapParallel_n9_inst4_O_6_0;
wire [7:0] NativeMapParallel_n9_inst4_O_7_0;
wire [7:0] NativeMapParallel_n9_inst4_O_8_0;
wire NativeMapParallel_n9_inst4_valid_down;
wire [7:0] Partition_S_no3_ni1_tElSSeq_1_Int__vTrue_inst0_O_0_0;
wire [7:0] Partition_S_no3_ni1_tElSSeq_1_Int__vTrue_inst0_O_1_0;
wire [7:0] Partition_S_no3_ni1_tElSSeq_1_Int__vTrue_inst0_O_2_0;
wire Partition_S_no3_ni1_tElSSeq_1_Int__vTrue_inst0_valid_down;
wire [7:0] Partition_S_no3_ni3_tElSSeq_1_Int__vTrue_inst0_O_0_0_0;
wire [7:0] Partition_S_no3_ni3_tElSSeq_1_Int__vTrue_inst0_O_0_1_0;
wire [7:0] Partition_S_no3_ni3_tElSSeq_1_Int__vTrue_inst0_O_0_2_0;
wire [7:0] Partition_S_no3_ni3_tElSSeq_1_Int__vTrue_inst0_O_1_0_0;
wire [7:0] Partition_S_no3_ni3_tElSSeq_1_Int__vTrue_inst0_O_1_1_0;
wire [7:0] Partition_S_no3_ni3_tElSSeq_1_Int__vTrue_inst0_O_1_2_0;
wire [7:0] Partition_S_no3_ni3_tElSSeq_1_Int__vTrue_inst0_O_2_0_0;
wire [7:0] Partition_S_no3_ni3_tElSSeq_1_Int__vTrue_inst0_O_2_1_0;
wire [7:0] Partition_S_no3_ni3_tElSSeq_1_Int__vTrue_inst0_O_2_2_0;
wire Partition_S_no3_ni3_tElSSeq_1_Int__vTrue_inst0_valid_down;
wire [7:0] Partition_S_no9_ni1_tElSSeq_1_Int__vTrue_inst0_O_0_0;
wire [7:0] Partition_S_no9_ni1_tElSSeq_1_Int__vTrue_inst0_O_1_0;
wire [7:0] Partition_S_no9_ni1_tElSSeq_1_Int__vTrue_inst0_O_2_0;
wire [7:0] Partition_S_no9_ni1_tElSSeq_1_Int__vTrue_inst0_O_3_0;
wire [7:0] Partition_S_no9_ni1_tElSSeq_1_Int__vTrue_inst0_O_4_0;
wire [7:0] Partition_S_no9_ni1_tElSSeq_1_Int__vTrue_inst0_O_5_0;
wire [7:0] Partition_S_no9_ni1_tElSSeq_1_Int__vTrue_inst0_O_6_0;
wire [7:0] Partition_S_no9_ni1_tElSSeq_1_Int__vTrue_inst0_O_7_0;
wire [7:0] Partition_S_no9_ni1_tElSSeq_1_Int__vTrue_inst0_O_8_0;
wire Partition_S_no9_ni1_tElSSeq_1_Int__vTrue_inst0_valid_down;
wire [7:0] Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_0_0_0;
wire [7:0] Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_0_1_0;
wire [7:0] Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_0_2_0;
wire [7:0] Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_1_0_0;
wire [7:0] Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_1_1_0;
wire [7:0] Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_1_2_0;
wire [7:0] Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_2_0_0;
wire [7:0] Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_2_1_0;
wire [7:0] Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_2_2_0;
wire [7:0] Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_3_0_0;
wire [7:0] Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_3_1_0;
wire [7:0] Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_3_2_0;
wire [7:0] Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_4_0_0;
wire [7:0] Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_4_1_0;
wire [7:0] Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_4_2_0;
wire [7:0] Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_5_0_0;
wire [7:0] Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_5_1_0;
wire [7:0] Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_5_2_0;
wire [7:0] Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_6_0_0;
wire [7:0] Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_6_1_0;
wire [7:0] Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_6_2_0;
wire [7:0] Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_7_0_0;
wire [7:0] Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_7_1_0;
wire [7:0] Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_7_2_0;
wire [7:0] Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_8_0_0;
wire [7:0] Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_8_1_0;
wire [7:0] Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_8_2_0;
wire Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_valid_down;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_0_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_10_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_11_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_12_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_13_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_14_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_15_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_16_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_17_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_18_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_19_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_1_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_20_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_21_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_22_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_23_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_24_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_25_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_26_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_2_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_3_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_4_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_5_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_6_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_7_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_8_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_9_0;
wire Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_valid_down;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_0_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_10_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_11_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_12_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_13_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_14_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_15_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_16_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_17_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_18_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_19_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_1_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_20_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_21_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_22_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_23_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_24_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_25_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_26_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_2_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_3_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_4_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_5_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_6_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_7_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_8_0;
wire [7:0] Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_9_0;
wire Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_valid_down;
wire [7:0] Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_0_0;
wire [7:0] Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_1_0;
wire [7:0] Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_2_0;
wire [7:0] Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_3_0;
wire [7:0] Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_4_0;
wire [7:0] Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_5_0;
wire [7:0] Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_6_0;
wire [7:0] Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_7_0;
wire [7:0] Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_8_0;
wire Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst0_valid_down;
wire [7:0] Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_0_0;
wire [7:0] Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_1_0;
wire [7:0] Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_2_0;
wire [7:0] Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_3_0;
wire [7:0] Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_4_0;
wire [7:0] Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_5_0;
wire [7:0] Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_6_0;
wire [7:0] Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_7_0;
wire [7:0] Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_8_0;
wire Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst1_valid_down;
wire and_inst0_out;
wire and_inst1_out;
wire and_inst2_out;
wire and_inst3_out;
FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0(.CLK(CLK), .I_0_0(I_0_0), .I_10_0(I_10_0), .I_11_0(I_11_0), .I_12_0(I_12_0), .I_13_0(I_13_0), .I_14_0(I_14_0), .I_15_0(I_15_0), .I_16_0(I_16_0), .I_17_0(I_17_0), .I_18_0(I_18_0), .I_19_0(I_19_0), .I_1_0(I_1_0), .I_20_0(I_20_0), .I_21_0(I_21_0), .I_22_0(I_22_0), .I_23_0(I_23_0), .I_24_0(I_24_0), .I_25_0(I_25_0), .I_26_0(I_26_0), .I_2_0(I_2_0), .I_3_0(I_3_0), .I_4_0(I_4_0), .I_5_0(I_5_0), .I_6_0(I_6_0), .I_7_0(I_7_0), .I_8_0(I_8_0), .I_9_0(I_9_0), .O_0_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0_0), .O_10_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_10_0), .O_11_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_11_0), .O_12_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_12_0), .O_13_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_13_0), .O_14_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_14_0), .O_15_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_15_0), .O_16_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_16_0), .O_17_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_17_0), .O_18_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_18_0), .O_19_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_19_0), .O_1_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_1_0), .O_20_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_20_0), .O_21_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_21_0), .O_22_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_22_0), .O_23_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_23_0), .O_24_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_24_0), .O_25_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_25_0), .O_26_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_26_0), .O_2_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_2_0), .O_3_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_3_0), .O_4_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_4_0), .O_5_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_5_0), .O_6_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_6_0), .O_7_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_7_0), .O_8_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_8_0), .O_9_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_9_0), .valid_down(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down), .valid_up(valid_up));
FIFO_tSSeq_3_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue FIFO_tSSeq_3_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0(.CLK(CLK), .I_0_0(Partition_S_no3_ni1_tElSSeq_1_Int__vTrue_inst0_O_0_0), .I_1_0(Partition_S_no3_ni1_tElSSeq_1_Int__vTrue_inst0_O_1_0), .I_2_0(Partition_S_no3_ni1_tElSSeq_1_Int__vTrue_inst0_O_2_0), .O_0_0(FIFO_tSSeq_3_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0_0), .O_1_0(FIFO_tSSeq_3_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_1_0), .O_2_0(FIFO_tSSeq_3_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_2_0), .valid_down(FIFO_tSSeq_3_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down), .valid_up(Partition_S_no3_ni1_tElSSeq_1_Int__vTrue_inst0_valid_down));
FIFO_tSSeq_3_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue FIFO_tSSeq_3_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1(.CLK(CLK), .I_0_0(FIFO_tSSeq_3_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0_0), .I_1_0(FIFO_tSSeq_3_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_1_0), .I_2_0(FIFO_tSSeq_3_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_2_0), .O_0_0(FIFO_tSSeq_3_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_0_0), .O_1_0(FIFO_tSSeq_3_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_1_0), .O_2_0(FIFO_tSSeq_3_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_2_0), .valid_down(FIFO_tSSeq_3_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_valid_down), .valid_up(FIFO_tSSeq_3_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down));
FIFO_tSSeq_3_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue FIFO_tSSeq_3_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2(.CLK(CLK), .I_0_0(FIFO_tSSeq_3_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_0_0), .I_1_0(FIFO_tSSeq_3_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_1_0), .I_2_0(FIFO_tSSeq_3_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_2_0), .O_0_0(FIFO_tSSeq_3_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_0_0), .O_1_0(FIFO_tSSeq_3_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_1_0), .O_2_0(FIFO_tSSeq_3_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_2_0), .valid_down(FIFO_tSSeq_3_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_valid_down), .valid_up(FIFO_tSSeq_3_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_valid_down));
NativeMapParallel_n27 NativeMapParallel_n27_inst0(.I0_0_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_0_0), .I0_10_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_10_0), .I0_11_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_11_0), .I0_12_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_12_0), .I0_13_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_13_0), .I0_14_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_14_0), .I0_15_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_15_0), .I0_16_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_16_0), .I0_17_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_17_0), .I0_18_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_18_0), .I0_19_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_19_0), .I0_1_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_1_0), .I0_20_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_20_0), .I0_21_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_21_0), .I0_22_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_22_0), .I0_23_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_23_0), .I0_24_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_24_0), .I0_25_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_25_0), .I0_26_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_26_0), .I0_2_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_2_0), .I0_3_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_3_0), .I0_4_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_4_0), .I0_5_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_5_0), .I0_6_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_6_0), .I0_7_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_7_0), .I0_8_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_8_0), .I0_9_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_9_0), .I1_0_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_0_0), .I1_10_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_10_0), .I1_11_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_11_0), .I1_12_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_12_0), .I1_13_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_13_0), .I1_14_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_14_0), .I1_15_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_15_0), .I1_16_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_16_0), .I1_17_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_17_0), .I1_18_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_18_0), .I1_19_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_19_0), .I1_1_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_1_0), .I1_20_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_20_0), .I1_21_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_21_0), .I1_22_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_22_0), .I1_23_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_23_0), .I1_24_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_24_0), .I1_25_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_25_0), .I1_26_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_26_0), .I1_2_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_2_0), .I1_3_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_3_0), .I1_4_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_4_0), .I1_5_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_5_0), .I1_6_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_6_0), .I1_7_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_7_0), .I1_8_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_8_0), .I1_9_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_9_0), .O_0_0_0(NativeMapParallel_n27_inst0_O_0_0_0), .O_0_0_1(NativeMapParallel_n27_inst0_O_0_0_1), .O_10_0_0(NativeMapParallel_n27_inst0_O_10_0_0), .O_10_0_1(NativeMapParallel_n27_inst0_O_10_0_1), .O_11_0_0(NativeMapParallel_n27_inst0_O_11_0_0), .O_11_0_1(NativeMapParallel_n27_inst0_O_11_0_1), .O_12_0_0(NativeMapParallel_n27_inst0_O_12_0_0), .O_12_0_1(NativeMapParallel_n27_inst0_O_12_0_1), .O_13_0_0(NativeMapParallel_n27_inst0_O_13_0_0), .O_13_0_1(NativeMapParallel_n27_inst0_O_13_0_1), .O_14_0_0(NativeMapParallel_n27_inst0_O_14_0_0), .O_14_0_1(NativeMapParallel_n27_inst0_O_14_0_1), .O_15_0_0(NativeMapParallel_n27_inst0_O_15_0_0), .O_15_0_1(NativeMapParallel_n27_inst0_O_15_0_1), .O_16_0_0(NativeMapParallel_n27_inst0_O_16_0_0), .O_16_0_1(NativeMapParallel_n27_inst0_O_16_0_1), .O_17_0_0(NativeMapParallel_n27_inst0_O_17_0_0), .O_17_0_1(NativeMapParallel_n27_inst0_O_17_0_1), .O_18_0_0(NativeMapParallel_n27_inst0_O_18_0_0), .O_18_0_1(NativeMapParallel_n27_inst0_O_18_0_1), .O_19_0_0(NativeMapParallel_n27_inst0_O_19_0_0), .O_19_0_1(NativeMapParallel_n27_inst0_O_19_0_1), .O_1_0_0(NativeMapParallel_n27_inst0_O_1_0_0), .O_1_0_1(NativeMapParallel_n27_inst0_O_1_0_1), .O_20_0_0(NativeMapParallel_n27_inst0_O_20_0_0), .O_20_0_1(NativeMapParallel_n27_inst0_O_20_0_1), .O_21_0_0(NativeMapParallel_n27_inst0_O_21_0_0), .O_21_0_1(NativeMapParallel_n27_inst0_O_21_0_1), .O_22_0_0(NativeMapParallel_n27_inst0_O_22_0_0), .O_22_0_1(NativeMapParallel_n27_inst0_O_22_0_1), .O_23_0_0(NativeMapParallel_n27_inst0_O_23_0_0), .O_23_0_1(NativeMapParallel_n27_inst0_O_23_0_1), .O_24_0_0(NativeMapParallel_n27_inst0_O_24_0_0), .O_24_0_1(NativeMapParallel_n27_inst0_O_24_0_1), .O_25_0_0(NativeMapParallel_n27_inst0_O_25_0_0), .O_25_0_1(NativeMapParallel_n27_inst0_O_25_0_1), .O_26_0_0(NativeMapParallel_n27_inst0_O_26_0_0), .O_26_0_1(NativeMapParallel_n27_inst0_O_26_0_1), .O_2_0_0(NativeMapParallel_n27_inst0_O_2_0_0), .O_2_0_1(NativeMapParallel_n27_inst0_O_2_0_1), .O_3_0_0(NativeMapParallel_n27_inst0_O_3_0_0), .O_3_0_1(NativeMapParallel_n27_inst0_O_3_0_1), .O_4_0_0(NativeMapParallel_n27_inst0_O_4_0_0), .O_4_0_1(NativeMapParallel_n27_inst0_O_4_0_1), .O_5_0_0(NativeMapParallel_n27_inst0_O_5_0_0), .O_5_0_1(NativeMapParallel_n27_inst0_O_5_0_1), .O_6_0_0(NativeMapParallel_n27_inst0_O_6_0_0), .O_6_0_1(NativeMapParallel_n27_inst0_O_6_0_1), .O_7_0_0(NativeMapParallel_n27_inst0_O_7_0_0), .O_7_0_1(NativeMapParallel_n27_inst0_O_7_0_1), .O_8_0_0(NativeMapParallel_n27_inst0_O_8_0_0), .O_8_0_1(NativeMapParallel_n27_inst0_O_8_0_1), .O_9_0_0(NativeMapParallel_n27_inst0_O_9_0_0), .O_9_0_1(NativeMapParallel_n27_inst0_O_9_0_1), .valid_down(NativeMapParallel_n27_inst0_valid_down), .valid_up(and_inst0_out));
NativeMapParallel_n27_unq1 NativeMapParallel_n27_inst1(.I0_0_0_0(NativeMapParallel_n27_inst0_O_0_0_0), .I0_0_0_1(NativeMapParallel_n27_inst0_O_0_0_1), .I0_10_0_0(NativeMapParallel_n27_inst0_O_10_0_0), .I0_10_0_1(NativeMapParallel_n27_inst0_O_10_0_1), .I0_11_0_0(NativeMapParallel_n27_inst0_O_11_0_0), .I0_11_0_1(NativeMapParallel_n27_inst0_O_11_0_1), .I0_12_0_0(NativeMapParallel_n27_inst0_O_12_0_0), .I0_12_0_1(NativeMapParallel_n27_inst0_O_12_0_1), .I0_13_0_0(NativeMapParallel_n27_inst0_O_13_0_0), .I0_13_0_1(NativeMapParallel_n27_inst0_O_13_0_1), .I0_14_0_0(NativeMapParallel_n27_inst0_O_14_0_0), .I0_14_0_1(NativeMapParallel_n27_inst0_O_14_0_1), .I0_15_0_0(NativeMapParallel_n27_inst0_O_15_0_0), .I0_15_0_1(NativeMapParallel_n27_inst0_O_15_0_1), .I0_16_0_0(NativeMapParallel_n27_inst0_O_16_0_0), .I0_16_0_1(NativeMapParallel_n27_inst0_O_16_0_1), .I0_17_0_0(NativeMapParallel_n27_inst0_O_17_0_0), .I0_17_0_1(NativeMapParallel_n27_inst0_O_17_0_1), .I0_18_0_0(NativeMapParallel_n27_inst0_O_18_0_0), .I0_18_0_1(NativeMapParallel_n27_inst0_O_18_0_1), .I0_19_0_0(NativeMapParallel_n27_inst0_O_19_0_0), .I0_19_0_1(NativeMapParallel_n27_inst0_O_19_0_1), .I0_1_0_0(NativeMapParallel_n27_inst0_O_1_0_0), .I0_1_0_1(NativeMapParallel_n27_inst0_O_1_0_1), .I0_20_0_0(NativeMapParallel_n27_inst0_O_20_0_0), .I0_20_0_1(NativeMapParallel_n27_inst0_O_20_0_1), .I0_21_0_0(NativeMapParallel_n27_inst0_O_21_0_0), .I0_21_0_1(NativeMapParallel_n27_inst0_O_21_0_1), .I0_22_0_0(NativeMapParallel_n27_inst0_O_22_0_0), .I0_22_0_1(NativeMapParallel_n27_inst0_O_22_0_1), .I0_23_0_0(NativeMapParallel_n27_inst0_O_23_0_0), .I0_23_0_1(NativeMapParallel_n27_inst0_O_23_0_1), .I0_24_0_0(NativeMapParallel_n27_inst0_O_24_0_0), .I0_24_0_1(NativeMapParallel_n27_inst0_O_24_0_1), .I0_25_0_0(NativeMapParallel_n27_inst0_O_25_0_0), .I0_25_0_1(NativeMapParallel_n27_inst0_O_25_0_1), .I0_26_0_0(NativeMapParallel_n27_inst0_O_26_0_0), .I0_26_0_1(NativeMapParallel_n27_inst0_O_26_0_1), .I0_2_0_0(NativeMapParallel_n27_inst0_O_2_0_0), .I0_2_0_1(NativeMapParallel_n27_inst0_O_2_0_1), .I0_3_0_0(NativeMapParallel_n27_inst0_O_3_0_0), .I0_3_0_1(NativeMapParallel_n27_inst0_O_3_0_1), .I0_4_0_0(NativeMapParallel_n27_inst0_O_4_0_0), .I0_4_0_1(NativeMapParallel_n27_inst0_O_4_0_1), .I0_5_0_0(NativeMapParallel_n27_inst0_O_5_0_0), .I0_5_0_1(NativeMapParallel_n27_inst0_O_5_0_1), .I0_6_0_0(NativeMapParallel_n27_inst0_O_6_0_0), .I0_6_0_1(NativeMapParallel_n27_inst0_O_6_0_1), .I0_7_0_0(NativeMapParallel_n27_inst0_O_7_0_0), .I0_7_0_1(NativeMapParallel_n27_inst0_O_7_0_1), .I0_8_0_0(NativeMapParallel_n27_inst0_O_8_0_0), .I0_8_0_1(NativeMapParallel_n27_inst0_O_8_0_1), .I0_9_0_0(NativeMapParallel_n27_inst0_O_9_0_0), .I0_9_0_1(NativeMapParallel_n27_inst0_O_9_0_1), .I1_0_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0_0), .I1_10_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_10_0), .I1_11_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_11_0), .I1_12_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_12_0), .I1_13_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_13_0), .I1_14_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_14_0), .I1_15_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_15_0), .I1_16_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_16_0), .I1_17_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_17_0), .I1_18_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_18_0), .I1_19_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_19_0), .I1_1_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_1_0), .I1_20_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_20_0), .I1_21_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_21_0), .I1_22_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_22_0), .I1_23_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_23_0), .I1_24_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_24_0), .I1_25_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_25_0), .I1_26_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_26_0), .I1_2_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_2_0), .I1_3_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_3_0), .I1_4_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_4_0), .I1_5_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_5_0), .I1_6_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_6_0), .I1_7_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_7_0), .I1_8_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_8_0), .I1_9_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_9_0), .O_0_0_0(NativeMapParallel_n27_inst1_O_0_0_0), .O_0_0_1(NativeMapParallel_n27_inst1_O_0_0_1), .O_0_0_2(NativeMapParallel_n27_inst1_O_0_0_2), .O_10_0_0(NativeMapParallel_n27_inst1_O_10_0_0), .O_10_0_1(NativeMapParallel_n27_inst1_O_10_0_1), .O_10_0_2(NativeMapParallel_n27_inst1_O_10_0_2), .O_11_0_0(NativeMapParallel_n27_inst1_O_11_0_0), .O_11_0_1(NativeMapParallel_n27_inst1_O_11_0_1), .O_11_0_2(NativeMapParallel_n27_inst1_O_11_0_2), .O_12_0_0(NativeMapParallel_n27_inst1_O_12_0_0), .O_12_0_1(NativeMapParallel_n27_inst1_O_12_0_1), .O_12_0_2(NativeMapParallel_n27_inst1_O_12_0_2), .O_13_0_0(NativeMapParallel_n27_inst1_O_13_0_0), .O_13_0_1(NativeMapParallel_n27_inst1_O_13_0_1), .O_13_0_2(NativeMapParallel_n27_inst1_O_13_0_2), .O_14_0_0(NativeMapParallel_n27_inst1_O_14_0_0), .O_14_0_1(NativeMapParallel_n27_inst1_O_14_0_1), .O_14_0_2(NativeMapParallel_n27_inst1_O_14_0_2), .O_15_0_0(NativeMapParallel_n27_inst1_O_15_0_0), .O_15_0_1(NativeMapParallel_n27_inst1_O_15_0_1), .O_15_0_2(NativeMapParallel_n27_inst1_O_15_0_2), .O_16_0_0(NativeMapParallel_n27_inst1_O_16_0_0), .O_16_0_1(NativeMapParallel_n27_inst1_O_16_0_1), .O_16_0_2(NativeMapParallel_n27_inst1_O_16_0_2), .O_17_0_0(NativeMapParallel_n27_inst1_O_17_0_0), .O_17_0_1(NativeMapParallel_n27_inst1_O_17_0_1), .O_17_0_2(NativeMapParallel_n27_inst1_O_17_0_2), .O_18_0_0(NativeMapParallel_n27_inst1_O_18_0_0), .O_18_0_1(NativeMapParallel_n27_inst1_O_18_0_1), .O_18_0_2(NativeMapParallel_n27_inst1_O_18_0_2), .O_19_0_0(NativeMapParallel_n27_inst1_O_19_0_0), .O_19_0_1(NativeMapParallel_n27_inst1_O_19_0_1), .O_19_0_2(NativeMapParallel_n27_inst1_O_19_0_2), .O_1_0_0(NativeMapParallel_n27_inst1_O_1_0_0), .O_1_0_1(NativeMapParallel_n27_inst1_O_1_0_1), .O_1_0_2(NativeMapParallel_n27_inst1_O_1_0_2), .O_20_0_0(NativeMapParallel_n27_inst1_O_20_0_0), .O_20_0_1(NativeMapParallel_n27_inst1_O_20_0_1), .O_20_0_2(NativeMapParallel_n27_inst1_O_20_0_2), .O_21_0_0(NativeMapParallel_n27_inst1_O_21_0_0), .O_21_0_1(NativeMapParallel_n27_inst1_O_21_0_1), .O_21_0_2(NativeMapParallel_n27_inst1_O_21_0_2), .O_22_0_0(NativeMapParallel_n27_inst1_O_22_0_0), .O_22_0_1(NativeMapParallel_n27_inst1_O_22_0_1), .O_22_0_2(NativeMapParallel_n27_inst1_O_22_0_2), .O_23_0_0(NativeMapParallel_n27_inst1_O_23_0_0), .O_23_0_1(NativeMapParallel_n27_inst1_O_23_0_1), .O_23_0_2(NativeMapParallel_n27_inst1_O_23_0_2), .O_24_0_0(NativeMapParallel_n27_inst1_O_24_0_0), .O_24_0_1(NativeMapParallel_n27_inst1_O_24_0_1), .O_24_0_2(NativeMapParallel_n27_inst1_O_24_0_2), .O_25_0_0(NativeMapParallel_n27_inst1_O_25_0_0), .O_25_0_1(NativeMapParallel_n27_inst1_O_25_0_1), .O_25_0_2(NativeMapParallel_n27_inst1_O_25_0_2), .O_26_0_0(NativeMapParallel_n27_inst1_O_26_0_0), .O_26_0_1(NativeMapParallel_n27_inst1_O_26_0_1), .O_26_0_2(NativeMapParallel_n27_inst1_O_26_0_2), .O_2_0_0(NativeMapParallel_n27_inst1_O_2_0_0), .O_2_0_1(NativeMapParallel_n27_inst1_O_2_0_1), .O_2_0_2(NativeMapParallel_n27_inst1_O_2_0_2), .O_3_0_0(NativeMapParallel_n27_inst1_O_3_0_0), .O_3_0_1(NativeMapParallel_n27_inst1_O_3_0_1), .O_3_0_2(NativeMapParallel_n27_inst1_O_3_0_2), .O_4_0_0(NativeMapParallel_n27_inst1_O_4_0_0), .O_4_0_1(NativeMapParallel_n27_inst1_O_4_0_1), .O_4_0_2(NativeMapParallel_n27_inst1_O_4_0_2), .O_5_0_0(NativeMapParallel_n27_inst1_O_5_0_0), .O_5_0_1(NativeMapParallel_n27_inst1_O_5_0_1), .O_5_0_2(NativeMapParallel_n27_inst1_O_5_0_2), .O_6_0_0(NativeMapParallel_n27_inst1_O_6_0_0), .O_6_0_1(NativeMapParallel_n27_inst1_O_6_0_1), .O_6_0_2(NativeMapParallel_n27_inst1_O_6_0_2), .O_7_0_0(NativeMapParallel_n27_inst1_O_7_0_0), .O_7_0_1(NativeMapParallel_n27_inst1_O_7_0_1), .O_7_0_2(NativeMapParallel_n27_inst1_O_7_0_2), .O_8_0_0(NativeMapParallel_n27_inst1_O_8_0_0), .O_8_0_1(NativeMapParallel_n27_inst1_O_8_0_1), .O_8_0_2(NativeMapParallel_n27_inst1_O_8_0_2), .O_9_0_0(NativeMapParallel_n27_inst1_O_9_0_0), .O_9_0_1(NativeMapParallel_n27_inst1_O_9_0_1), .O_9_0_2(NativeMapParallel_n27_inst1_O_9_0_2), .valid_down(NativeMapParallel_n27_inst1_valid_down), .valid_up(and_inst1_out));
NativeMapParallel_n27_unq2 NativeMapParallel_n27_inst2(.I_0_0_0(NativeMapParallel_n27_inst1_O_0_0_0), .I_0_0_1(NativeMapParallel_n27_inst1_O_0_0_1), .I_0_0_2(NativeMapParallel_n27_inst1_O_0_0_2), .I_10_0_0(NativeMapParallel_n27_inst1_O_10_0_0), .I_10_0_1(NativeMapParallel_n27_inst1_O_10_0_1), .I_10_0_2(NativeMapParallel_n27_inst1_O_10_0_2), .I_11_0_0(NativeMapParallel_n27_inst1_O_11_0_0), .I_11_0_1(NativeMapParallel_n27_inst1_O_11_0_1), .I_11_0_2(NativeMapParallel_n27_inst1_O_11_0_2), .I_12_0_0(NativeMapParallel_n27_inst1_O_12_0_0), .I_12_0_1(NativeMapParallel_n27_inst1_O_12_0_1), .I_12_0_2(NativeMapParallel_n27_inst1_O_12_0_2), .I_13_0_0(NativeMapParallel_n27_inst1_O_13_0_0), .I_13_0_1(NativeMapParallel_n27_inst1_O_13_0_1), .I_13_0_2(NativeMapParallel_n27_inst1_O_13_0_2), .I_14_0_0(NativeMapParallel_n27_inst1_O_14_0_0), .I_14_0_1(NativeMapParallel_n27_inst1_O_14_0_1), .I_14_0_2(NativeMapParallel_n27_inst1_O_14_0_2), .I_15_0_0(NativeMapParallel_n27_inst1_O_15_0_0), .I_15_0_1(NativeMapParallel_n27_inst1_O_15_0_1), .I_15_0_2(NativeMapParallel_n27_inst1_O_15_0_2), .I_16_0_0(NativeMapParallel_n27_inst1_O_16_0_0), .I_16_0_1(NativeMapParallel_n27_inst1_O_16_0_1), .I_16_0_2(NativeMapParallel_n27_inst1_O_16_0_2), .I_17_0_0(NativeMapParallel_n27_inst1_O_17_0_0), .I_17_0_1(NativeMapParallel_n27_inst1_O_17_0_1), .I_17_0_2(NativeMapParallel_n27_inst1_O_17_0_2), .I_18_0_0(NativeMapParallel_n27_inst1_O_18_0_0), .I_18_0_1(NativeMapParallel_n27_inst1_O_18_0_1), .I_18_0_2(NativeMapParallel_n27_inst1_O_18_0_2), .I_19_0_0(NativeMapParallel_n27_inst1_O_19_0_0), .I_19_0_1(NativeMapParallel_n27_inst1_O_19_0_1), .I_19_0_2(NativeMapParallel_n27_inst1_O_19_0_2), .I_1_0_0(NativeMapParallel_n27_inst1_O_1_0_0), .I_1_0_1(NativeMapParallel_n27_inst1_O_1_0_1), .I_1_0_2(NativeMapParallel_n27_inst1_O_1_0_2), .I_20_0_0(NativeMapParallel_n27_inst1_O_20_0_0), .I_20_0_1(NativeMapParallel_n27_inst1_O_20_0_1), .I_20_0_2(NativeMapParallel_n27_inst1_O_20_0_2), .I_21_0_0(NativeMapParallel_n27_inst1_O_21_0_0), .I_21_0_1(NativeMapParallel_n27_inst1_O_21_0_1), .I_21_0_2(NativeMapParallel_n27_inst1_O_21_0_2), .I_22_0_0(NativeMapParallel_n27_inst1_O_22_0_0), .I_22_0_1(NativeMapParallel_n27_inst1_O_22_0_1), .I_22_0_2(NativeMapParallel_n27_inst1_O_22_0_2), .I_23_0_0(NativeMapParallel_n27_inst1_O_23_0_0), .I_23_0_1(NativeMapParallel_n27_inst1_O_23_0_1), .I_23_0_2(NativeMapParallel_n27_inst1_O_23_0_2), .I_24_0_0(NativeMapParallel_n27_inst1_O_24_0_0), .I_24_0_1(NativeMapParallel_n27_inst1_O_24_0_1), .I_24_0_2(NativeMapParallel_n27_inst1_O_24_0_2), .I_25_0_0(NativeMapParallel_n27_inst1_O_25_0_0), .I_25_0_1(NativeMapParallel_n27_inst1_O_25_0_1), .I_25_0_2(NativeMapParallel_n27_inst1_O_25_0_2), .I_26_0_0(NativeMapParallel_n27_inst1_O_26_0_0), .I_26_0_1(NativeMapParallel_n27_inst1_O_26_0_1), .I_26_0_2(NativeMapParallel_n27_inst1_O_26_0_2), .I_2_0_0(NativeMapParallel_n27_inst1_O_2_0_0), .I_2_0_1(NativeMapParallel_n27_inst1_O_2_0_1), .I_2_0_2(NativeMapParallel_n27_inst1_O_2_0_2), .I_3_0_0(NativeMapParallel_n27_inst1_O_3_0_0), .I_3_0_1(NativeMapParallel_n27_inst1_O_3_0_1), .I_3_0_2(NativeMapParallel_n27_inst1_O_3_0_2), .I_4_0_0(NativeMapParallel_n27_inst1_O_4_0_0), .I_4_0_1(NativeMapParallel_n27_inst1_O_4_0_1), .I_4_0_2(NativeMapParallel_n27_inst1_O_4_0_2), .I_5_0_0(NativeMapParallel_n27_inst1_O_5_0_0), .I_5_0_1(NativeMapParallel_n27_inst1_O_5_0_1), .I_5_0_2(NativeMapParallel_n27_inst1_O_5_0_2), .I_6_0_0(NativeMapParallel_n27_inst1_O_6_0_0), .I_6_0_1(NativeMapParallel_n27_inst1_O_6_0_1), .I_6_0_2(NativeMapParallel_n27_inst1_O_6_0_2), .I_7_0_0(NativeMapParallel_n27_inst1_O_7_0_0), .I_7_0_1(NativeMapParallel_n27_inst1_O_7_0_1), .I_7_0_2(NativeMapParallel_n27_inst1_O_7_0_2), .I_8_0_0(NativeMapParallel_n27_inst1_O_8_0_0), .I_8_0_1(NativeMapParallel_n27_inst1_O_8_0_1), .I_8_0_2(NativeMapParallel_n27_inst1_O_8_0_2), .I_9_0_0(NativeMapParallel_n27_inst1_O_9_0_0), .I_9_0_1(NativeMapParallel_n27_inst1_O_9_0_1), .I_9_0_2(NativeMapParallel_n27_inst1_O_9_0_2), .O_0_0(NativeMapParallel_n27_inst2_O_0_0), .O_0_1(NativeMapParallel_n27_inst2_O_0_1), .O_0_2(NativeMapParallel_n27_inst2_O_0_2), .O_10_0(NativeMapParallel_n27_inst2_O_10_0), .O_10_1(NativeMapParallel_n27_inst2_O_10_1), .O_10_2(NativeMapParallel_n27_inst2_O_10_2), .O_11_0(NativeMapParallel_n27_inst2_O_11_0), .O_11_1(NativeMapParallel_n27_inst2_O_11_1), .O_11_2(NativeMapParallel_n27_inst2_O_11_2), .O_12_0(NativeMapParallel_n27_inst2_O_12_0), .O_12_1(NativeMapParallel_n27_inst2_O_12_1), .O_12_2(NativeMapParallel_n27_inst2_O_12_2), .O_13_0(NativeMapParallel_n27_inst2_O_13_0), .O_13_1(NativeMapParallel_n27_inst2_O_13_1), .O_13_2(NativeMapParallel_n27_inst2_O_13_2), .O_14_0(NativeMapParallel_n27_inst2_O_14_0), .O_14_1(NativeMapParallel_n27_inst2_O_14_1), .O_14_2(NativeMapParallel_n27_inst2_O_14_2), .O_15_0(NativeMapParallel_n27_inst2_O_15_0), .O_15_1(NativeMapParallel_n27_inst2_O_15_1), .O_15_2(NativeMapParallel_n27_inst2_O_15_2), .O_16_0(NativeMapParallel_n27_inst2_O_16_0), .O_16_1(NativeMapParallel_n27_inst2_O_16_1), .O_16_2(NativeMapParallel_n27_inst2_O_16_2), .O_17_0(NativeMapParallel_n27_inst2_O_17_0), .O_17_1(NativeMapParallel_n27_inst2_O_17_1), .O_17_2(NativeMapParallel_n27_inst2_O_17_2), .O_18_0(NativeMapParallel_n27_inst2_O_18_0), .O_18_1(NativeMapParallel_n27_inst2_O_18_1), .O_18_2(NativeMapParallel_n27_inst2_O_18_2), .O_19_0(NativeMapParallel_n27_inst2_O_19_0), .O_19_1(NativeMapParallel_n27_inst2_O_19_1), .O_19_2(NativeMapParallel_n27_inst2_O_19_2), .O_1_0(NativeMapParallel_n27_inst2_O_1_0), .O_1_1(NativeMapParallel_n27_inst2_O_1_1), .O_1_2(NativeMapParallel_n27_inst2_O_1_2), .O_20_0(NativeMapParallel_n27_inst2_O_20_0), .O_20_1(NativeMapParallel_n27_inst2_O_20_1), .O_20_2(NativeMapParallel_n27_inst2_O_20_2), .O_21_0(NativeMapParallel_n27_inst2_O_21_0), .O_21_1(NativeMapParallel_n27_inst2_O_21_1), .O_21_2(NativeMapParallel_n27_inst2_O_21_2), .O_22_0(NativeMapParallel_n27_inst2_O_22_0), .O_22_1(NativeMapParallel_n27_inst2_O_22_1), .O_22_2(NativeMapParallel_n27_inst2_O_22_2), .O_23_0(NativeMapParallel_n27_inst2_O_23_0), .O_23_1(NativeMapParallel_n27_inst2_O_23_1), .O_23_2(NativeMapParallel_n27_inst2_O_23_2), .O_24_0(NativeMapParallel_n27_inst2_O_24_0), .O_24_1(NativeMapParallel_n27_inst2_O_24_1), .O_24_2(NativeMapParallel_n27_inst2_O_24_2), .O_25_0(NativeMapParallel_n27_inst2_O_25_0), .O_25_1(NativeMapParallel_n27_inst2_O_25_1), .O_25_2(NativeMapParallel_n27_inst2_O_25_2), .O_26_0(NativeMapParallel_n27_inst2_O_26_0), .O_26_1(NativeMapParallel_n27_inst2_O_26_1), .O_26_2(NativeMapParallel_n27_inst2_O_26_2), .O_2_0(NativeMapParallel_n27_inst2_O_2_0), .O_2_1(NativeMapParallel_n27_inst2_O_2_1), .O_2_2(NativeMapParallel_n27_inst2_O_2_2), .O_3_0(NativeMapParallel_n27_inst2_O_3_0), .O_3_1(NativeMapParallel_n27_inst2_O_3_1), .O_3_2(NativeMapParallel_n27_inst2_O_3_2), .O_4_0(NativeMapParallel_n27_inst2_O_4_0), .O_4_1(NativeMapParallel_n27_inst2_O_4_1), .O_4_2(NativeMapParallel_n27_inst2_O_4_2), .O_5_0(NativeMapParallel_n27_inst2_O_5_0), .O_5_1(NativeMapParallel_n27_inst2_O_5_1), .O_5_2(NativeMapParallel_n27_inst2_O_5_2), .O_6_0(NativeMapParallel_n27_inst2_O_6_0), .O_6_1(NativeMapParallel_n27_inst2_O_6_1), .O_6_2(NativeMapParallel_n27_inst2_O_6_2), .O_7_0(NativeMapParallel_n27_inst2_O_7_0), .O_7_1(NativeMapParallel_n27_inst2_O_7_1), .O_7_2(NativeMapParallel_n27_inst2_O_7_2), .O_8_0(NativeMapParallel_n27_inst2_O_8_0), .O_8_1(NativeMapParallel_n27_inst2_O_8_1), .O_8_2(NativeMapParallel_n27_inst2_O_8_2), .O_9_0(NativeMapParallel_n27_inst2_O_9_0), .O_9_1(NativeMapParallel_n27_inst2_O_9_1), .O_9_2(NativeMapParallel_n27_inst2_O_9_2), .valid_down(NativeMapParallel_n27_inst2_valid_down), .valid_up(NativeMapParallel_n27_inst1_valid_down));
NativeMapParallel_n27_unq3 NativeMapParallel_n27_inst3(.CLK(CLK), .I_0_0(NativeMapParallel_n27_inst2_O_0_0), .I_0_1(NativeMapParallel_n27_inst2_O_0_1), .I_0_2(NativeMapParallel_n27_inst2_O_0_2), .I_10_0(NativeMapParallel_n27_inst2_O_10_0), .I_10_1(NativeMapParallel_n27_inst2_O_10_1), .I_10_2(NativeMapParallel_n27_inst2_O_10_2), .I_11_0(NativeMapParallel_n27_inst2_O_11_0), .I_11_1(NativeMapParallel_n27_inst2_O_11_1), .I_11_2(NativeMapParallel_n27_inst2_O_11_2), .I_12_0(NativeMapParallel_n27_inst2_O_12_0), .I_12_1(NativeMapParallel_n27_inst2_O_12_1), .I_12_2(NativeMapParallel_n27_inst2_O_12_2), .I_13_0(NativeMapParallel_n27_inst2_O_13_0), .I_13_1(NativeMapParallel_n27_inst2_O_13_1), .I_13_2(NativeMapParallel_n27_inst2_O_13_2), .I_14_0(NativeMapParallel_n27_inst2_O_14_0), .I_14_1(NativeMapParallel_n27_inst2_O_14_1), .I_14_2(NativeMapParallel_n27_inst2_O_14_2), .I_15_0(NativeMapParallel_n27_inst2_O_15_0), .I_15_1(NativeMapParallel_n27_inst2_O_15_1), .I_15_2(NativeMapParallel_n27_inst2_O_15_2), .I_16_0(NativeMapParallel_n27_inst2_O_16_0), .I_16_1(NativeMapParallel_n27_inst2_O_16_1), .I_16_2(NativeMapParallel_n27_inst2_O_16_2), .I_17_0(NativeMapParallel_n27_inst2_O_17_0), .I_17_1(NativeMapParallel_n27_inst2_O_17_1), .I_17_2(NativeMapParallel_n27_inst2_O_17_2), .I_18_0(NativeMapParallel_n27_inst2_O_18_0), .I_18_1(NativeMapParallel_n27_inst2_O_18_1), .I_18_2(NativeMapParallel_n27_inst2_O_18_2), .I_19_0(NativeMapParallel_n27_inst2_O_19_0), .I_19_1(NativeMapParallel_n27_inst2_O_19_1), .I_19_2(NativeMapParallel_n27_inst2_O_19_2), .I_1_0(NativeMapParallel_n27_inst2_O_1_0), .I_1_1(NativeMapParallel_n27_inst2_O_1_1), .I_1_2(NativeMapParallel_n27_inst2_O_1_2), .I_20_0(NativeMapParallel_n27_inst2_O_20_0), .I_20_1(NativeMapParallel_n27_inst2_O_20_1), .I_20_2(NativeMapParallel_n27_inst2_O_20_2), .I_21_0(NativeMapParallel_n27_inst2_O_21_0), .I_21_1(NativeMapParallel_n27_inst2_O_21_1), .I_21_2(NativeMapParallel_n27_inst2_O_21_2), .I_22_0(NativeMapParallel_n27_inst2_O_22_0), .I_22_1(NativeMapParallel_n27_inst2_O_22_1), .I_22_2(NativeMapParallel_n27_inst2_O_22_2), .I_23_0(NativeMapParallel_n27_inst2_O_23_0), .I_23_1(NativeMapParallel_n27_inst2_O_23_1), .I_23_2(NativeMapParallel_n27_inst2_O_23_2), .I_24_0(NativeMapParallel_n27_inst2_O_24_0), .I_24_1(NativeMapParallel_n27_inst2_O_24_1), .I_24_2(NativeMapParallel_n27_inst2_O_24_2), .I_25_0(NativeMapParallel_n27_inst2_O_25_0), .I_25_1(NativeMapParallel_n27_inst2_O_25_1), .I_25_2(NativeMapParallel_n27_inst2_O_25_2), .I_26_0(NativeMapParallel_n27_inst2_O_26_0), .I_26_1(NativeMapParallel_n27_inst2_O_26_1), .I_26_2(NativeMapParallel_n27_inst2_O_26_2), .I_2_0(NativeMapParallel_n27_inst2_O_2_0), .I_2_1(NativeMapParallel_n27_inst2_O_2_1), .I_2_2(NativeMapParallel_n27_inst2_O_2_2), .I_3_0(NativeMapParallel_n27_inst2_O_3_0), .I_3_1(NativeMapParallel_n27_inst2_O_3_1), .I_3_2(NativeMapParallel_n27_inst2_O_3_2), .I_4_0(NativeMapParallel_n27_inst2_O_4_0), .I_4_1(NativeMapParallel_n27_inst2_O_4_1), .I_4_2(NativeMapParallel_n27_inst2_O_4_2), .I_5_0(NativeMapParallel_n27_inst2_O_5_0), .I_5_1(NativeMapParallel_n27_inst2_O_5_1), .I_5_2(NativeMapParallel_n27_inst2_O_5_2), .I_6_0(NativeMapParallel_n27_inst2_O_6_0), .I_6_1(NativeMapParallel_n27_inst2_O_6_1), .I_6_2(NativeMapParallel_n27_inst2_O_6_2), .I_7_0(NativeMapParallel_n27_inst2_O_7_0), .I_7_1(NativeMapParallel_n27_inst2_O_7_1), .I_7_2(NativeMapParallel_n27_inst2_O_7_2), .I_8_0(NativeMapParallel_n27_inst2_O_8_0), .I_8_1(NativeMapParallel_n27_inst2_O_8_1), .I_8_2(NativeMapParallel_n27_inst2_O_8_2), .I_9_0(NativeMapParallel_n27_inst2_O_9_0), .I_9_1(NativeMapParallel_n27_inst2_O_9_1), .I_9_2(NativeMapParallel_n27_inst2_O_9_2), .O_0_0(NativeMapParallel_n27_inst3_O_0_0), .O_10_0(NativeMapParallel_n27_inst3_O_10_0), .O_11_0(NativeMapParallel_n27_inst3_O_11_0), .O_12_0(NativeMapParallel_n27_inst3_O_12_0), .O_13_0(NativeMapParallel_n27_inst3_O_13_0), .O_14_0(NativeMapParallel_n27_inst3_O_14_0), .O_15_0(NativeMapParallel_n27_inst3_O_15_0), .O_16_0(NativeMapParallel_n27_inst3_O_16_0), .O_17_0(NativeMapParallel_n27_inst3_O_17_0), .O_18_0(NativeMapParallel_n27_inst3_O_18_0), .O_19_0(NativeMapParallel_n27_inst3_O_19_0), .O_1_0(NativeMapParallel_n27_inst3_O_1_0), .O_20_0(NativeMapParallel_n27_inst3_O_20_0), .O_21_0(NativeMapParallel_n27_inst3_O_21_0), .O_22_0(NativeMapParallel_n27_inst3_O_22_0), .O_23_0(NativeMapParallel_n27_inst3_O_23_0), .O_24_0(NativeMapParallel_n27_inst3_O_24_0), .O_25_0(NativeMapParallel_n27_inst3_O_25_0), .O_26_0(NativeMapParallel_n27_inst3_O_26_0), .O_2_0(NativeMapParallel_n27_inst3_O_2_0), .O_3_0(NativeMapParallel_n27_inst3_O_3_0), .O_4_0(NativeMapParallel_n27_inst3_O_4_0), .O_5_0(NativeMapParallel_n27_inst3_O_5_0), .O_6_0(NativeMapParallel_n27_inst3_O_6_0), .O_7_0(NativeMapParallel_n27_inst3_O_7_0), .O_8_0(NativeMapParallel_n27_inst3_O_8_0), .O_9_0(NativeMapParallel_n27_inst3_O_9_0), .valid_down(NativeMapParallel_n27_inst3_valid_down), .valid_up(NativeMapParallel_n27_inst2_valid_down));
NativeMapParallel_n3_unq2 NativeMapParallel_n3_inst0(.CLK(CLK), .I_0_0_0(Partition_S_no3_ni3_tElSSeq_1_Int__vTrue_inst0_O_0_0_0), .I_0_1_0(Partition_S_no3_ni3_tElSSeq_1_Int__vTrue_inst0_O_0_1_0), .I_0_2_0(Partition_S_no3_ni3_tElSSeq_1_Int__vTrue_inst0_O_0_2_0), .I_1_0_0(Partition_S_no3_ni3_tElSSeq_1_Int__vTrue_inst0_O_1_0_0), .I_1_1_0(Partition_S_no3_ni3_tElSSeq_1_Int__vTrue_inst0_O_1_1_0), .I_1_2_0(Partition_S_no3_ni3_tElSSeq_1_Int__vTrue_inst0_O_1_2_0), .I_2_0_0(Partition_S_no3_ni3_tElSSeq_1_Int__vTrue_inst0_O_2_0_0), .I_2_1_0(Partition_S_no3_ni3_tElSSeq_1_Int__vTrue_inst0_O_2_1_0), .I_2_2_0(Partition_S_no3_ni3_tElSSeq_1_Int__vTrue_inst0_O_2_2_0), .O_0_0_0(NativeMapParallel_n3_inst0_O_0_0_0), .O_1_0_0(NativeMapParallel_n3_inst0_O_1_0_0), .O_2_0_0(NativeMapParallel_n3_inst0_O_2_0_0), .valid_down(NativeMapParallel_n3_inst0_valid_down), .valid_up(Partition_S_no3_ni3_tElSSeq_1_Int__vTrue_inst0_valid_down));
NativeMapParallel_n9 NativeMapParallel_n9_inst0(.CLK(CLK), .I_0_0_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_0_0_0), .I_0_1_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_0_1_0), .I_0_2_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_0_2_0), .I_1_0_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_1_0_0), .I_1_1_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_1_1_0), .I_1_2_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_1_2_0), .I_2_0_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_2_0_0), .I_2_1_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_2_1_0), .I_2_2_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_2_2_0), .I_3_0_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_3_0_0), .I_3_1_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_3_1_0), .I_3_2_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_3_2_0), .I_4_0_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_4_0_0), .I_4_1_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_4_1_0), .I_4_2_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_4_2_0), .I_5_0_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_5_0_0), .I_5_1_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_5_1_0), .I_5_2_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_5_2_0), .I_6_0_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_6_0_0), .I_6_1_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_6_1_0), .I_6_2_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_6_2_0), .I_7_0_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_7_0_0), .I_7_1_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_7_1_0), .I_7_2_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_7_2_0), .I_8_0_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_8_0_0), .I_8_1_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_8_1_0), .I_8_2_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_8_2_0), .O_0_0_0(NativeMapParallel_n9_inst0_O_0_0_0), .O_1_0_0(NativeMapParallel_n9_inst0_O_1_0_0), .O_2_0_0(NativeMapParallel_n9_inst0_O_2_0_0), .O_3_0_0(NativeMapParallel_n9_inst0_O_3_0_0), .O_4_0_0(NativeMapParallel_n9_inst0_O_4_0_0), .O_5_0_0(NativeMapParallel_n9_inst0_O_5_0_0), .O_6_0_0(NativeMapParallel_n9_inst0_O_6_0_0), .O_7_0_0(NativeMapParallel_n9_inst0_O_7_0_0), .O_8_0_0(NativeMapParallel_n9_inst0_O_8_0_0), .valid_down(NativeMapParallel_n9_inst0_valid_down), .valid_up(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_valid_down));
NativeMapParallel_n9_unq1 NativeMapParallel_n9_inst1(.I0_0_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_0_0), .I0_1_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_1_0), .I0_2_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_2_0), .I0_3_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_3_0), .I0_4_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_4_0), .I0_5_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_5_0), .I0_6_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_6_0), .I0_7_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_7_0), .I0_8_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_8_0), .I1_0_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_0_0), .I1_1_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_1_0), .I1_2_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_2_0), .I1_3_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_3_0), .I1_4_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_4_0), .I1_5_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_5_0), .I1_6_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_6_0), .I1_7_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_7_0), .I1_8_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_8_0), .O_0_0_0(NativeMapParallel_n9_inst1_O_0_0_0), .O_0_0_1(NativeMapParallel_n9_inst1_O_0_0_1), .O_1_0_0(NativeMapParallel_n9_inst1_O_1_0_0), .O_1_0_1(NativeMapParallel_n9_inst1_O_1_0_1), .O_2_0_0(NativeMapParallel_n9_inst1_O_2_0_0), .O_2_0_1(NativeMapParallel_n9_inst1_O_2_0_1), .O_3_0_0(NativeMapParallel_n9_inst1_O_3_0_0), .O_3_0_1(NativeMapParallel_n9_inst1_O_3_0_1), .O_4_0_0(NativeMapParallel_n9_inst1_O_4_0_0), .O_4_0_1(NativeMapParallel_n9_inst1_O_4_0_1), .O_5_0_0(NativeMapParallel_n9_inst1_O_5_0_0), .O_5_0_1(NativeMapParallel_n9_inst1_O_5_0_1), .O_6_0_0(NativeMapParallel_n9_inst1_O_6_0_0), .O_6_0_1(NativeMapParallel_n9_inst1_O_6_0_1), .O_7_0_0(NativeMapParallel_n9_inst1_O_7_0_0), .O_7_0_1(NativeMapParallel_n9_inst1_O_7_0_1), .O_8_0_0(NativeMapParallel_n9_inst1_O_8_0_0), .O_8_0_1(NativeMapParallel_n9_inst1_O_8_0_1), .valid_down(NativeMapParallel_n9_inst1_valid_down), .valid_up(and_inst2_out));
NativeMapParallel_n9_unq2 NativeMapParallel_n9_inst2(.I0_0_0_0(NativeMapParallel_n9_inst1_O_0_0_0), .I0_0_0_1(NativeMapParallel_n9_inst1_O_0_0_1), .I0_1_0_0(NativeMapParallel_n9_inst1_O_1_0_0), .I0_1_0_1(NativeMapParallel_n9_inst1_O_1_0_1), .I0_2_0_0(NativeMapParallel_n9_inst1_O_2_0_0), .I0_2_0_1(NativeMapParallel_n9_inst1_O_2_0_1), .I0_3_0_0(NativeMapParallel_n9_inst1_O_3_0_0), .I0_3_0_1(NativeMapParallel_n9_inst1_O_3_0_1), .I0_4_0_0(NativeMapParallel_n9_inst1_O_4_0_0), .I0_4_0_1(NativeMapParallel_n9_inst1_O_4_0_1), .I0_5_0_0(NativeMapParallel_n9_inst1_O_5_0_0), .I0_5_0_1(NativeMapParallel_n9_inst1_O_5_0_1), .I0_6_0_0(NativeMapParallel_n9_inst1_O_6_0_0), .I0_6_0_1(NativeMapParallel_n9_inst1_O_6_0_1), .I0_7_0_0(NativeMapParallel_n9_inst1_O_7_0_0), .I0_7_0_1(NativeMapParallel_n9_inst1_O_7_0_1), .I0_8_0_0(NativeMapParallel_n9_inst1_O_8_0_0), .I0_8_0_1(NativeMapParallel_n9_inst1_O_8_0_1), .I1_0_0(Partition_S_no9_ni1_tElSSeq_1_Int__vTrue_inst0_O_0_0), .I1_1_0(Partition_S_no9_ni1_tElSSeq_1_Int__vTrue_inst0_O_1_0), .I1_2_0(Partition_S_no9_ni1_tElSSeq_1_Int__vTrue_inst0_O_2_0), .I1_3_0(Partition_S_no9_ni1_tElSSeq_1_Int__vTrue_inst0_O_3_0), .I1_4_0(Partition_S_no9_ni1_tElSSeq_1_Int__vTrue_inst0_O_4_0), .I1_5_0(Partition_S_no9_ni1_tElSSeq_1_Int__vTrue_inst0_O_5_0), .I1_6_0(Partition_S_no9_ni1_tElSSeq_1_Int__vTrue_inst0_O_6_0), .I1_7_0(Partition_S_no9_ni1_tElSSeq_1_Int__vTrue_inst0_O_7_0), .I1_8_0(Partition_S_no9_ni1_tElSSeq_1_Int__vTrue_inst0_O_8_0), .O_0_0_0(NativeMapParallel_n9_inst2_O_0_0_0), .O_0_0_1(NativeMapParallel_n9_inst2_O_0_0_1), .O_0_0_2(NativeMapParallel_n9_inst2_O_0_0_2), .O_1_0_0(NativeMapParallel_n9_inst2_O_1_0_0), .O_1_0_1(NativeMapParallel_n9_inst2_O_1_0_1), .O_1_0_2(NativeMapParallel_n9_inst2_O_1_0_2), .O_2_0_0(NativeMapParallel_n9_inst2_O_2_0_0), .O_2_0_1(NativeMapParallel_n9_inst2_O_2_0_1), .O_2_0_2(NativeMapParallel_n9_inst2_O_2_0_2), .O_3_0_0(NativeMapParallel_n9_inst2_O_3_0_0), .O_3_0_1(NativeMapParallel_n9_inst2_O_3_0_1), .O_3_0_2(NativeMapParallel_n9_inst2_O_3_0_2), .O_4_0_0(NativeMapParallel_n9_inst2_O_4_0_0), .O_4_0_1(NativeMapParallel_n9_inst2_O_4_0_1), .O_4_0_2(NativeMapParallel_n9_inst2_O_4_0_2), .O_5_0_0(NativeMapParallel_n9_inst2_O_5_0_0), .O_5_0_1(NativeMapParallel_n9_inst2_O_5_0_1), .O_5_0_2(NativeMapParallel_n9_inst2_O_5_0_2), .O_6_0_0(NativeMapParallel_n9_inst2_O_6_0_0), .O_6_0_1(NativeMapParallel_n9_inst2_O_6_0_1), .O_6_0_2(NativeMapParallel_n9_inst2_O_6_0_2), .O_7_0_0(NativeMapParallel_n9_inst2_O_7_0_0), .O_7_0_1(NativeMapParallel_n9_inst2_O_7_0_1), .O_7_0_2(NativeMapParallel_n9_inst2_O_7_0_2), .O_8_0_0(NativeMapParallel_n9_inst2_O_8_0_0), .O_8_0_1(NativeMapParallel_n9_inst2_O_8_0_1), .O_8_0_2(NativeMapParallel_n9_inst2_O_8_0_2), .valid_down(NativeMapParallel_n9_inst2_valid_down), .valid_up(and_inst3_out));
NativeMapParallel_n9_unq3 NativeMapParallel_n9_inst3(.I_0_0_0(NativeMapParallel_n9_inst2_O_0_0_0), .I_0_0_1(NativeMapParallel_n9_inst2_O_0_0_1), .I_0_0_2(NativeMapParallel_n9_inst2_O_0_0_2), .I_1_0_0(NativeMapParallel_n9_inst2_O_1_0_0), .I_1_0_1(NativeMapParallel_n9_inst2_O_1_0_1), .I_1_0_2(NativeMapParallel_n9_inst2_O_1_0_2), .I_2_0_0(NativeMapParallel_n9_inst2_O_2_0_0), .I_2_0_1(NativeMapParallel_n9_inst2_O_2_0_1), .I_2_0_2(NativeMapParallel_n9_inst2_O_2_0_2), .I_3_0_0(NativeMapParallel_n9_inst2_O_3_0_0), .I_3_0_1(NativeMapParallel_n9_inst2_O_3_0_1), .I_3_0_2(NativeMapParallel_n9_inst2_O_3_0_2), .I_4_0_0(NativeMapParallel_n9_inst2_O_4_0_0), .I_4_0_1(NativeMapParallel_n9_inst2_O_4_0_1), .I_4_0_2(NativeMapParallel_n9_inst2_O_4_0_2), .I_5_0_0(NativeMapParallel_n9_inst2_O_5_0_0), .I_5_0_1(NativeMapParallel_n9_inst2_O_5_0_1), .I_5_0_2(NativeMapParallel_n9_inst2_O_5_0_2), .I_6_0_0(NativeMapParallel_n9_inst2_O_6_0_0), .I_6_0_1(NativeMapParallel_n9_inst2_O_6_0_1), .I_6_0_2(NativeMapParallel_n9_inst2_O_6_0_2), .I_7_0_0(NativeMapParallel_n9_inst2_O_7_0_0), .I_7_0_1(NativeMapParallel_n9_inst2_O_7_0_1), .I_7_0_2(NativeMapParallel_n9_inst2_O_7_0_2), .I_8_0_0(NativeMapParallel_n9_inst2_O_8_0_0), .I_8_0_1(NativeMapParallel_n9_inst2_O_8_0_1), .I_8_0_2(NativeMapParallel_n9_inst2_O_8_0_2), .O_0_0(NativeMapParallel_n9_inst3_O_0_0), .O_0_1(NativeMapParallel_n9_inst3_O_0_1), .O_0_2(NativeMapParallel_n9_inst3_O_0_2), .O_1_0(NativeMapParallel_n9_inst3_O_1_0), .O_1_1(NativeMapParallel_n9_inst3_O_1_1), .O_1_2(NativeMapParallel_n9_inst3_O_1_2), .O_2_0(NativeMapParallel_n9_inst3_O_2_0), .O_2_1(NativeMapParallel_n9_inst3_O_2_1), .O_2_2(NativeMapParallel_n9_inst3_O_2_2), .O_3_0(NativeMapParallel_n9_inst3_O_3_0), .O_3_1(NativeMapParallel_n9_inst3_O_3_1), .O_3_2(NativeMapParallel_n9_inst3_O_3_2), .O_4_0(NativeMapParallel_n9_inst3_O_4_0), .O_4_1(NativeMapParallel_n9_inst3_O_4_1), .O_4_2(NativeMapParallel_n9_inst3_O_4_2), .O_5_0(NativeMapParallel_n9_inst3_O_5_0), .O_5_1(NativeMapParallel_n9_inst3_O_5_1), .O_5_2(NativeMapParallel_n9_inst3_O_5_2), .O_6_0(NativeMapParallel_n9_inst3_O_6_0), .O_6_1(NativeMapParallel_n9_inst3_O_6_1), .O_6_2(NativeMapParallel_n9_inst3_O_6_2), .O_7_0(NativeMapParallel_n9_inst3_O_7_0), .O_7_1(NativeMapParallel_n9_inst3_O_7_1), .O_7_2(NativeMapParallel_n9_inst3_O_7_2), .O_8_0(NativeMapParallel_n9_inst3_O_8_0), .O_8_1(NativeMapParallel_n9_inst3_O_8_1), .O_8_2(NativeMapParallel_n9_inst3_O_8_2), .valid_down(NativeMapParallel_n9_inst3_valid_down), .valid_up(NativeMapParallel_n9_inst2_valid_down));
NativeMapParallel_n9_unq4 NativeMapParallel_n9_inst4(.CLK(CLK), .I_0_0(NativeMapParallel_n9_inst3_O_0_0), .I_0_1(NativeMapParallel_n9_inst3_O_0_1), .I_0_2(NativeMapParallel_n9_inst3_O_0_2), .I_1_0(NativeMapParallel_n9_inst3_O_1_0), .I_1_1(NativeMapParallel_n9_inst3_O_1_1), .I_1_2(NativeMapParallel_n9_inst3_O_1_2), .I_2_0(NativeMapParallel_n9_inst3_O_2_0), .I_2_1(NativeMapParallel_n9_inst3_O_2_1), .I_2_2(NativeMapParallel_n9_inst3_O_2_2), .I_3_0(NativeMapParallel_n9_inst3_O_3_0), .I_3_1(NativeMapParallel_n9_inst3_O_3_1), .I_3_2(NativeMapParallel_n9_inst3_O_3_2), .I_4_0(NativeMapParallel_n9_inst3_O_4_0), .I_4_1(NativeMapParallel_n9_inst3_O_4_1), .I_4_2(NativeMapParallel_n9_inst3_O_4_2), .I_5_0(NativeMapParallel_n9_inst3_O_5_0), .I_5_1(NativeMapParallel_n9_inst3_O_5_1), .I_5_2(NativeMapParallel_n9_inst3_O_5_2), .I_6_0(NativeMapParallel_n9_inst3_O_6_0), .I_6_1(NativeMapParallel_n9_inst3_O_6_1), .I_6_2(NativeMapParallel_n9_inst3_O_6_2), .I_7_0(NativeMapParallel_n9_inst3_O_7_0), .I_7_1(NativeMapParallel_n9_inst3_O_7_1), .I_7_2(NativeMapParallel_n9_inst3_O_7_2), .I_8_0(NativeMapParallel_n9_inst3_O_8_0), .I_8_1(NativeMapParallel_n9_inst3_O_8_1), .I_8_2(NativeMapParallel_n9_inst3_O_8_2), .O_0_0(NativeMapParallel_n9_inst4_O_0_0), .O_1_0(NativeMapParallel_n9_inst4_O_1_0), .O_2_0(NativeMapParallel_n9_inst4_O_2_0), .O_3_0(NativeMapParallel_n9_inst4_O_3_0), .O_4_0(NativeMapParallel_n9_inst4_O_4_0), .O_5_0(NativeMapParallel_n9_inst4_O_5_0), .O_6_0(NativeMapParallel_n9_inst4_O_6_0), .O_7_0(NativeMapParallel_n9_inst4_O_7_0), .O_8_0(NativeMapParallel_n9_inst4_O_8_0), .valid_down(NativeMapParallel_n9_inst4_valid_down), .valid_up(NativeMapParallel_n9_inst3_valid_down));
Partition_S_no3_ni1_tElSSeq_1_Int__vTrue Partition_S_no3_ni1_tElSSeq_1_Int__vTrue_inst0(.CLK(CLK), .I_0_0_0(NativeMapParallel_n3_inst0_O_0_0_0), .I_1_0_0(NativeMapParallel_n3_inst0_O_1_0_0), .I_2_0_0(NativeMapParallel_n3_inst0_O_2_0_0), .O_0_0(Partition_S_no3_ni1_tElSSeq_1_Int__vTrue_inst0_O_0_0), .O_1_0(Partition_S_no3_ni1_tElSSeq_1_Int__vTrue_inst0_O_1_0), .O_2_0(Partition_S_no3_ni1_tElSSeq_1_Int__vTrue_inst0_O_2_0), .valid_down(Partition_S_no3_ni1_tElSSeq_1_Int__vTrue_inst0_valid_down), .valid_up(NativeMapParallel_n3_inst0_valid_down));
Partition_S_no3_ni3_tElSSeq_1_Int__vTrue Partition_S_no3_ni3_tElSSeq_1_Int__vTrue_inst0(.CLK(CLK), .I_0_0(NativeMapParallel_n9_inst4_O_0_0), .I_1_0(NativeMapParallel_n9_inst4_O_1_0), .I_2_0(NativeMapParallel_n9_inst4_O_2_0), .I_3_0(NativeMapParallel_n9_inst4_O_3_0), .I_4_0(NativeMapParallel_n9_inst4_O_4_0), .I_5_0(NativeMapParallel_n9_inst4_O_5_0), .I_6_0(NativeMapParallel_n9_inst4_O_6_0), .I_7_0(NativeMapParallel_n9_inst4_O_7_0), .I_8_0(NativeMapParallel_n9_inst4_O_8_0), .O_0_0_0(Partition_S_no3_ni3_tElSSeq_1_Int__vTrue_inst0_O_0_0_0), .O_0_1_0(Partition_S_no3_ni3_tElSSeq_1_Int__vTrue_inst0_O_0_1_0), .O_0_2_0(Partition_S_no3_ni3_tElSSeq_1_Int__vTrue_inst0_O_0_2_0), .O_1_0_0(Partition_S_no3_ni3_tElSSeq_1_Int__vTrue_inst0_O_1_0_0), .O_1_1_0(Partition_S_no3_ni3_tElSSeq_1_Int__vTrue_inst0_O_1_1_0), .O_1_2_0(Partition_S_no3_ni3_tElSSeq_1_Int__vTrue_inst0_O_1_2_0), .O_2_0_0(Partition_S_no3_ni3_tElSSeq_1_Int__vTrue_inst0_O_2_0_0), .O_2_1_0(Partition_S_no3_ni3_tElSSeq_1_Int__vTrue_inst0_O_2_1_0), .O_2_2_0(Partition_S_no3_ni3_tElSSeq_1_Int__vTrue_inst0_O_2_2_0), .valid_down(Partition_S_no3_ni3_tElSSeq_1_Int__vTrue_inst0_valid_down), .valid_up(NativeMapParallel_n9_inst4_valid_down));
Partition_S_no9_ni1_tElSSeq_1_Int__vTrue Partition_S_no9_ni1_tElSSeq_1_Int__vTrue_inst0(.CLK(CLK), .I_0_0_0(NativeMapParallel_n9_inst0_O_0_0_0), .I_1_0_0(NativeMapParallel_n9_inst0_O_1_0_0), .I_2_0_0(NativeMapParallel_n9_inst0_O_2_0_0), .I_3_0_0(NativeMapParallel_n9_inst0_O_3_0_0), .I_4_0_0(NativeMapParallel_n9_inst0_O_4_0_0), .I_5_0_0(NativeMapParallel_n9_inst0_O_5_0_0), .I_6_0_0(NativeMapParallel_n9_inst0_O_6_0_0), .I_7_0_0(NativeMapParallel_n9_inst0_O_7_0_0), .I_8_0_0(NativeMapParallel_n9_inst0_O_8_0_0), .O_0_0(Partition_S_no9_ni1_tElSSeq_1_Int__vTrue_inst0_O_0_0), .O_1_0(Partition_S_no9_ni1_tElSSeq_1_Int__vTrue_inst0_O_1_0), .O_2_0(Partition_S_no9_ni1_tElSSeq_1_Int__vTrue_inst0_O_2_0), .O_3_0(Partition_S_no9_ni1_tElSSeq_1_Int__vTrue_inst0_O_3_0), .O_4_0(Partition_S_no9_ni1_tElSSeq_1_Int__vTrue_inst0_O_4_0), .O_5_0(Partition_S_no9_ni1_tElSSeq_1_Int__vTrue_inst0_O_5_0), .O_6_0(Partition_S_no9_ni1_tElSSeq_1_Int__vTrue_inst0_O_6_0), .O_7_0(Partition_S_no9_ni1_tElSSeq_1_Int__vTrue_inst0_O_7_0), .O_8_0(Partition_S_no9_ni1_tElSSeq_1_Int__vTrue_inst0_O_8_0), .valid_down(Partition_S_no9_ni1_tElSSeq_1_Int__vTrue_inst0_valid_down), .valid_up(NativeMapParallel_n9_inst0_valid_down));
Partition_S_no9_ni3_tElSSeq_1_Int__vTrue Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0(.CLK(CLK), .I_0_0(NativeMapParallel_n27_inst3_O_0_0), .I_10_0(NativeMapParallel_n27_inst3_O_10_0), .I_11_0(NativeMapParallel_n27_inst3_O_11_0), .I_12_0(NativeMapParallel_n27_inst3_O_12_0), .I_13_0(NativeMapParallel_n27_inst3_O_13_0), .I_14_0(NativeMapParallel_n27_inst3_O_14_0), .I_15_0(NativeMapParallel_n27_inst3_O_15_0), .I_16_0(NativeMapParallel_n27_inst3_O_16_0), .I_17_0(NativeMapParallel_n27_inst3_O_17_0), .I_18_0(NativeMapParallel_n27_inst3_O_18_0), .I_19_0(NativeMapParallel_n27_inst3_O_19_0), .I_1_0(NativeMapParallel_n27_inst3_O_1_0), .I_20_0(NativeMapParallel_n27_inst3_O_20_0), .I_21_0(NativeMapParallel_n27_inst3_O_21_0), .I_22_0(NativeMapParallel_n27_inst3_O_22_0), .I_23_0(NativeMapParallel_n27_inst3_O_23_0), .I_24_0(NativeMapParallel_n27_inst3_O_24_0), .I_25_0(NativeMapParallel_n27_inst3_O_25_0), .I_26_0(NativeMapParallel_n27_inst3_O_26_0), .I_2_0(NativeMapParallel_n27_inst3_O_2_0), .I_3_0(NativeMapParallel_n27_inst3_O_3_0), .I_4_0(NativeMapParallel_n27_inst3_O_4_0), .I_5_0(NativeMapParallel_n27_inst3_O_5_0), .I_6_0(NativeMapParallel_n27_inst3_O_6_0), .I_7_0(NativeMapParallel_n27_inst3_O_7_0), .I_8_0(NativeMapParallel_n27_inst3_O_8_0), .I_9_0(NativeMapParallel_n27_inst3_O_9_0), .O_0_0_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_0_0_0), .O_0_1_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_0_1_0), .O_0_2_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_0_2_0), .O_1_0_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_1_0_0), .O_1_1_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_1_1_0), .O_1_2_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_1_2_0), .O_2_0_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_2_0_0), .O_2_1_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_2_1_0), .O_2_2_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_2_2_0), .O_3_0_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_3_0_0), .O_3_1_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_3_1_0), .O_3_2_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_3_2_0), .O_4_0_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_4_0_0), .O_4_1_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_4_1_0), .O_4_2_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_4_2_0), .O_5_0_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_5_0_0), .O_5_1_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_5_1_0), .O_5_2_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_5_2_0), .O_6_0_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_6_0_0), .O_6_1_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_6_1_0), .O_6_2_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_6_2_0), .O_7_0_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_7_0_0), .O_7_1_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_7_1_0), .O_7_2_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_7_2_0), .O_8_0_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_8_0_0), .O_8_1_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_8_1_0), .O_8_2_0(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_O_8_2_0), .valid_down(Partition_S_no9_ni3_tElSSeq_1_Int__vTrue_inst0_valid_down), .valid_up(NativeMapParallel_n27_inst3_valid_down));
Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0(.CLK(CLK), .I_0_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0_0), .I_10_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_10_0), .I_11_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_11_0), .I_12_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_12_0), .I_13_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_13_0), .I_14_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_14_0), .I_15_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_15_0), .I_16_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_16_0), .I_17_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_17_0), .I_18_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_18_0), .I_19_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_19_0), .I_1_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_1_0), .I_20_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_20_0), .I_21_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_21_0), .I_22_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_22_0), .I_23_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_23_0), .I_24_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_24_0), .I_25_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_25_0), .I_26_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_26_0), .I_2_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_2_0), .I_3_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_3_0), .I_4_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_4_0), .I_5_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_5_0), .I_6_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_6_0), .I_7_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_7_0), .I_8_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_8_0), .I_9_0(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_9_0), .O_0_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_0_0), .O_10_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_10_0), .O_11_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_11_0), .O_12_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_12_0), .O_13_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_13_0), .O_14_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_14_0), .O_15_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_15_0), .O_16_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_16_0), .O_17_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_17_0), .O_18_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_18_0), .O_19_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_19_0), .O_1_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_1_0), .O_20_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_20_0), .O_21_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_21_0), .O_22_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_22_0), .O_23_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_23_0), .O_24_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_24_0), .O_25_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_25_0), .O_26_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_26_0), .O_2_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_2_0), .O_3_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_3_0), .O_4_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_4_0), .O_5_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_5_0), .O_6_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_6_0), .O_7_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_7_0), .O_8_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_8_0), .O_9_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_9_0), .valid_down(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_valid_down), .valid_up(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down));
Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1(.CLK(CLK), .I_0_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_0_0), .I_10_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_10_0), .I_11_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_11_0), .I_12_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_12_0), .I_13_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_13_0), .I_14_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_14_0), .I_15_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_15_0), .I_16_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_16_0), .I_17_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_17_0), .I_18_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_18_0), .I_19_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_19_0), .I_1_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_1_0), .I_20_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_20_0), .I_21_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_21_0), .I_22_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_22_0), .I_23_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_23_0), .I_24_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_24_0), .I_25_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_25_0), .I_26_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_26_0), .I_2_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_2_0), .I_3_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_3_0), .I_4_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_4_0), .I_5_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_5_0), .I_6_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_6_0), .I_7_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_7_0), .I_8_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_8_0), .I_9_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_9_0), .O_0_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_0_0), .O_10_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_10_0), .O_11_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_11_0), .O_12_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_12_0), .O_13_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_13_0), .O_14_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_14_0), .O_15_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_15_0), .O_16_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_16_0), .O_17_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_17_0), .O_18_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_18_0), .O_19_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_19_0), .O_1_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_1_0), .O_20_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_20_0), .O_21_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_21_0), .O_22_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_22_0), .O_23_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_23_0), .O_24_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_24_0), .O_25_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_25_0), .O_26_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_26_0), .O_2_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_2_0), .O_3_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_3_0), .O_4_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_4_0), .O_5_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_5_0), .O_6_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_6_0), .O_7_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_7_0), .O_8_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_8_0), .O_9_0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_9_0), .valid_down(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_valid_down), .valid_up(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_valid_down));
Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst0(.CLK(CLK), .I_0_0(Partition_S_no9_ni1_tElSSeq_1_Int__vTrue_inst0_O_0_0), .I_1_0(Partition_S_no9_ni1_tElSSeq_1_Int__vTrue_inst0_O_1_0), .I_2_0(Partition_S_no9_ni1_tElSSeq_1_Int__vTrue_inst0_O_2_0), .I_3_0(Partition_S_no9_ni1_tElSSeq_1_Int__vTrue_inst0_O_3_0), .I_4_0(Partition_S_no9_ni1_tElSSeq_1_Int__vTrue_inst0_O_4_0), .I_5_0(Partition_S_no9_ni1_tElSSeq_1_Int__vTrue_inst0_O_5_0), .I_6_0(Partition_S_no9_ni1_tElSSeq_1_Int__vTrue_inst0_O_6_0), .I_7_0(Partition_S_no9_ni1_tElSSeq_1_Int__vTrue_inst0_O_7_0), .I_8_0(Partition_S_no9_ni1_tElSSeq_1_Int__vTrue_inst0_O_8_0), .O_0_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_0_0), .O_1_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_1_0), .O_2_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_2_0), .O_3_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_3_0), .O_4_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_4_0), .O_5_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_5_0), .O_6_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_6_0), .O_7_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_7_0), .O_8_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_8_0), .valid_down(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst0_valid_down), .valid_up(Partition_S_no9_ni1_tElSSeq_1_Int__vTrue_inst0_valid_down));
Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst1(.CLK(CLK), .I_0_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_0_0), .I_1_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_1_0), .I_2_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_2_0), .I_3_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_3_0), .I_4_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_4_0), .I_5_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_5_0), .I_6_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_6_0), .I_7_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_7_0), .I_8_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst0_O_8_0), .O_0_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_0_0), .O_1_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_1_0), .O_2_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_2_0), .O_3_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_3_0), .O_4_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_4_0), .O_5_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_5_0), .O_6_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_6_0), .O_7_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_7_0), .O_8_0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst1_O_8_0), .valid_down(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst1_valid_down), .valid_up(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst0_valid_down));
corebit_and and_inst0(.in0(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst1_valid_down), .in1(Shift_S_n27_amt1_tElSSeq_1_Int__hasValidTrue_inst0_valid_down), .out(and_inst0_out));
corebit_and and_inst1(.in0(NativeMapParallel_n27_inst0_valid_down), .in1(FIFO_tSSeq_27_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down), .out(and_inst1_out));
corebit_and and_inst2(.in0(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst1_valid_down), .in1(Shift_S_n9_amt1_tElSSeq_1_Int__hasValidTrue_inst0_valid_down), .out(and_inst2_out));
corebit_and and_inst3(.in0(NativeMapParallel_n9_inst1_valid_down), .in1(Partition_S_no9_ni1_tElSSeq_1_Int__vTrue_inst0_valid_down), .out(and_inst3_out));
assign O_0_0 = FIFO_tSSeq_3_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_0_0;
assign O_1_0 = FIFO_tSSeq_3_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_1_0;
assign O_2_0 = FIFO_tSSeq_3_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_2_0;
assign valid_down = FIFO_tSSeq_3_SSeq_1_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_valid_down;
endmodule

