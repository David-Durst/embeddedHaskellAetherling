// Latency = 4
module top(
  input CLK/*verilator public*/, 
  input [7:0] I/*verilator public*/, 
  output [7:0] O/*verilator public*/, 
  output valid_down/*verilator public*/, 
  input valid_up/*verilator public*/
);
  wire dontcare;
  x35_inr_Foreach_SAMPLER_BOX_kernelx35_inr_Foreach_SAMPLER_BOX_concrete1 sampler_box ( // @[m_x55_ctr_0.scala 26:17:@1721.4]
    .clock(CLK), // @[:@1296.4]
    .reset('b0), // @[:@1297.4]
    .io_in_x21_TREADY(dontcare), // @[:@1298.4]
    .io_in_x21_TDATA(I), // @[:@1298.4]
    .io_in_x21_TID(8'h0),
    .io_in_x21_TDEST(8'h0),
    .io_in_x22_TVALID(valid_down), // @[:@1298.4]
    .io_in_x22_TDATA(O), // @[:@1298.4]
    .io_sigsIn_datapathEn(valid_up), // @[:@1298.4]
    .io_sigsIn_cchainOutputs_0_oobs_0('b0), // @[:@1298.4]
    .io_rr('b1) // @[:@1298.4]
  );

endmodule

module RetimeShiftRegister
#(
    parameter WIDTH = 1,
    parameter STAGES = 1)
(
    input clock,
    input reset,
    input flow,
    input [WIDTH-1:0] init,
    input [WIDTH-1:0] in,
    output reg [WIDTH-1:0] out
);
  integer i;
  reg [WIDTH-1:0] sr[STAGES:0]; // Create 'STAGES' number of register, each 'WIDTH' bits wide

   /* synopsys dc_tcl_script_begin
    set_ungroup [current_design] true
    set_flatten true -effort high -phase true -design [current_design]
    set_dont_retime [current_design] false
    set_optimize_registers true -design [current_design]
    */
  always @(posedge clock) begin
    if (reset) begin
      for(i=0; i<STAGES; i=i+1) begin
        sr[i] <= init;
      end
    end else begin
      if (flow) begin 
        sr[0] <= in;
        for(i=1; i<STAGES; i=i+1) begin
          sr[i] <= sr[i-1];
        end
      end
    end
  end

  always @(*) begin
    out = sr[STAGES-1];
  end
endmodule

module FF( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  output [31:0] io_rPort_0_output_0, // @[:@6.4]
  input  [31:0] io_wPort_0_data_0, // @[:@6.4]
  input         io_wPort_0_reset, // @[:@6.4]
  input         io_wPort_0_en_0 // @[:@6.4]
);
  reg [31:0] ff; // @[MemPrimitives.scala 173:19:@21.4]
  reg [31:0] _RAND_0;
  wire [31:0] _T_68; // @[MemPrimitives.scala 177:32:@23.4]
  wire [31:0] _T_69; // @[MemPrimitives.scala 177:12:@24.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 177:32:@23.4]
  assign _T_69 = io_wPort_0_reset ? 32'h0 : _T_68; // @[MemPrimitives.scala 177:12:@24.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 178:34:@26.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 32'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 32'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SRFF( // @[:@28.2]
  input   clock, // @[:@29.4]
  input   reset, // @[:@30.4]
  input   io_input_set, // @[:@31.4]
  input   io_input_reset, // @[:@31.4]
  input   io_input_asyn_reset, // @[:@31.4]
  output  io_output // @[:@31.4]
);
  reg  _T_15; // @[SRFF.scala 20:21:@33.4]
  reg [31:0] _RAND_0;
  wire  _T_19; // @[SRFF.scala 21:74:@34.4]
  wire  _T_20; // @[SRFF.scala 21:48:@35.4]
  wire  _T_21; // @[SRFF.scala 21:14:@36.4]
  assign _T_19 = io_input_reset ? 1'h0 : _T_15; // @[SRFF.scala 21:74:@34.4]
  assign _T_20 = io_input_set ? 1'h1 : _T_19; // @[SRFF.scala 21:48:@35.4]
  assign _T_21 = io_input_asyn_reset ? 1'h0 : _T_20; // @[SRFF.scala 21:14:@36.4]
  assign io_output = io_input_asyn_reset ? 1'h0 : _T_15; // @[SRFF.scala 22:15:@39.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_15 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_15 <= 1'h0;
    end else begin
      if (io_input_asyn_reset) begin
        _T_15 <= 1'h0;
      end else begin
        if (io_input_set) begin
          _T_15 <= 1'h1;
        end else begin
          if (io_input_reset) begin
            _T_15 <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module SingleCounter( // @[:@41.2]
  input   clock, // @[:@42.4]
  input   reset, // @[:@43.4]
  input   io_input_reset, // @[:@44.4]
  output  io_output_done // @[:@44.4]
);
  wire  bases_0_clock; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_reset; // @[Counter.scala 253:53:@57.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 253:53:@57.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 253:53:@57.4]
  wire  SRFF_clock; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_set; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_output; // @[Counter.scala 255:22:@73.4]
  wire [31:0] _T_48; // @[Counter.scala 279:52:@101.4]
  wire [32:0] _T_50; // @[Counter.scala 283:33:@102.4]
  wire [31:0] _T_51; // @[Counter.scala 283:33:@103.4]
  wire [31:0] _T_52; // @[Counter.scala 283:33:@104.4]
  wire  _T_57; // @[Counter.scala 285:18:@106.4]
  wire [31:0] _T_68; // @[Counter.scala 291:115:@114.4]
  wire [31:0] _T_71; // @[Counter.scala 291:152:@117.4]
  wire [31:0] _T_72; // @[Counter.scala 291:74:@118.4]
  FF bases_0 ( // @[Counter.scala 253:53:@57.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 255:22:@73.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 279:52:@101.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@102.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@103.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 283:33:@104.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh4); // @[Counter.scala 285:18:@106.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 291:115:@114.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 291:152:@117.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 291:74:@118.4]
  assign io_output_done = $signed(_T_52) >= $signed(32'sh4); // @[Counter.scala 325:20:@127.4]
  assign bases_0_clock = clock; // @[:@58.4]
  assign bases_0_reset = reset; // @[:@59.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 291:31:@120.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 273:27:@99.4]
  assign bases_0_io_wPort_0_en_0 = 1'h1; // @[Counter.scala 276:29:@100.4]
  assign SRFF_clock = clock; // @[:@74.4]
  assign SRFF_reset = reset; // @[:@75.4]
  assign SRFF_io_input_set = io_input_reset == 1'h0; // @[Counter.scala 256:23:@78.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 257:25:@80.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 258:30:@81.4]
endmodule
module RetimeWrapper( // @[:@144.2]
  input   clock, // @[:@145.4]
  input   reset, // @[:@146.4]
  input   io_flow, // @[:@147.4]
  input   io_in, // @[:@147.4]
  output  io_out // @[:@147.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@149.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@149.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@162.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@161.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@160.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@159.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@158.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@156.4]
endmodule
module RootController_sm( // @[:@312.2]
  input   clock, // @[:@313.4]
  input   reset, // @[:@314.4]
  input   io_enable, // @[:@315.4]
  output  io_done, // @[:@315.4]
  input   io_rst, // @[:@315.4]
  input   io_ctrDone, // @[:@315.4]
  output  io_ctrInc, // @[:@315.4]
  input   io_doneIn_0, // @[:@315.4]
  output  io_enableOut_0, // @[:@315.4]
  output  io_childAck_0 // @[:@315.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@318.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@321.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@338.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@433.4]
  wire  finished; // @[Controllers.scala 81:26:@324.4]
  wire  synchronize; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  wire  _T_122; // @[Controllers.scala 128:33:@371.4]
  wire  _T_124; // @[Controllers.scala 128:54:@372.4]
  wire  _T_125; // @[Controllers.scala 128:52:@373.4]
  wire  _T_126; // @[Controllers.scala 128:66:@374.4]
  wire  _T_128; // @[Controllers.scala 128:98:@376.4]
  wire  _T_129; // @[Controllers.scala 128:96:@377.4]
  wire  _T_131; // @[Controllers.scala 128:123:@378.4]
  wire  _T_133; // @[Controllers.scala 129:48:@381.4]
  wire  _T_138; // @[Controllers.scala 130:52:@386.4]
  wire  _T_139; // @[Controllers.scala 130:50:@387.4]
  wire  _T_147; // @[Controllers.scala 130:129:@393.4]
  wire  _T_150; // @[Controllers.scala 131:45:@396.4]
  wire  _T_154; // @[Controllers.scala 213:68:@402.4]
  wire  _T_156; // @[Controllers.scala 213:90:@404.4]
  wire  _T_158; // @[Controllers.scala 213:132:@406.4]
  wire  _T_159; // @[Controllers.scala 213:130:@407.4]
  wire  _T_160; // @[Controllers.scala 213:156:@408.4]
  reg  _T_166; // @[package.scala 48:56:@412.4]
  reg [31:0] _RAND_0;
  reg  _T_180; // @[package.scala 48:56:@430.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@318.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@321.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@338.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@357.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@416.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@433.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  assign finished = done_0_io_output | io_done; // @[Controllers.scala 81:26:@324.4]
  assign synchronize = RetimeWrapper_io_out; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  assign _T_122 = done_0_io_output == 1'h0; // @[Controllers.scala 128:33:@371.4]
  assign _T_124 = io_ctrDone == 1'h0; // @[Controllers.scala 128:54:@372.4]
  assign _T_125 = _T_122 & _T_124; // @[Controllers.scala 128:52:@373.4]
  assign _T_126 = _T_125 & io_enable; // @[Controllers.scala 128:66:@374.4]
  assign _T_128 = ~ iterDone_0_io_output; // @[Controllers.scala 128:98:@376.4]
  assign _T_129 = _T_126 & _T_128; // @[Controllers.scala 128:96:@377.4]
  assign _T_131 = io_doneIn_0 == 1'h0; // @[Controllers.scala 128:123:@378.4]
  assign _T_133 = io_doneIn_0 | io_rst; // @[Controllers.scala 129:48:@381.4]
  assign _T_138 = synchronize == 1'h0; // @[Controllers.scala 130:52:@386.4]
  assign _T_139 = io_doneIn_0 & _T_138; // @[Controllers.scala 130:50:@387.4]
  assign _T_147 = finished == 1'h0; // @[Controllers.scala 130:129:@393.4]
  assign _T_150 = io_rst == 1'h0; // @[Controllers.scala 131:45:@396.4]
  assign _T_154 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@402.4]
  assign _T_156 = _T_154 & _T_128; // @[Controllers.scala 213:90:@404.4]
  assign _T_158 = ~ done_0_io_output; // @[Controllers.scala 213:132:@406.4]
  assign _T_159 = _T_156 & _T_158; // @[Controllers.scala 213:130:@407.4]
  assign _T_160 = ~ io_ctrDone; // @[Controllers.scala 213:156:@408.4]
  assign io_done = RetimeWrapper_2_io_out; // @[Controllers.scala 245:13:@440.4]
  assign io_ctrInc = io_doneIn_0; // @[Controllers.scala 122:17:@356.4]
  assign io_enableOut_0 = _T_159 & _T_160; // @[Controllers.scala 213:55:@410.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@401.4]
  assign active_0_clock = clock; // @[:@319.4]
  assign active_0_reset = reset; // @[:@320.4]
  assign active_0_io_input_set = _T_129 & _T_131; // @[Controllers.scala 128:30:@380.4]
  assign active_0_io_input_reset = _T_133 | done_0_io_output; // @[Controllers.scala 129:32:@385.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@326.4]
  assign done_0_clock = clock; // @[:@322.4]
  assign done_0_reset = reset; // @[:@323.4]
  assign done_0_io_input_set = io_ctrDone & _T_150; // @[Controllers.scala 131:28:@399.4]
  assign done_0_io_input_reset = io_rst | done_0_io_output; // @[Controllers.scala 86:33:@336.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@327.4]
  assign iterDone_0_clock = clock; // @[:@339.4]
  assign iterDone_0_reset = reset; // @[:@340.4]
  assign iterDone_0_io_input_set = _T_139 & _T_147; // @[Controllers.scala 130:32:@395.4]
  assign iterDone_0_io_input_reset = synchronize | io_rst; // @[Controllers.scala 92:37:@350.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@341.4]
  assign RetimeWrapper_clock = clock; // @[:@358.4]
  assign RetimeWrapper_reset = reset; // @[:@359.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@361.4]
  assign RetimeWrapper_io_in = io_doneIn_0; // @[package.scala 94:16:@360.4]
  assign RetimeWrapper_1_clock = clock; // @[:@417.4]
  assign RetimeWrapper_1_reset = reset; // @[:@418.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@420.4]
  assign RetimeWrapper_1_io_in = done_0_io_output & _T_166; // @[package.scala 94:16:@419.4]
  assign RetimeWrapper_2_clock = clock; // @[:@434.4]
  assign RetimeWrapper_2_reset = reset; // @[:@435.4]
  assign RetimeWrapper_2_io_flow = io_enable; // @[package.scala 95:18:@437.4]
  assign RetimeWrapper_2_io_in = done_0_io_output & _T_180; // @[package.scala 94:16:@436.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_166 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_180 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_166 <= 1'h0;
    end else begin
      _T_166 <= _T_122;
    end
    if (reset) begin
      _T_180 <= 1'h0;
    end else begin
      _T_180 <= _T_122;
    end
  end
endmodule
module SingleCounter_1( // @[:@515.2]
  input   clock, // @[:@516.4]
  input   reset, // @[:@517.4]
  input   io_input_reset, // @[:@518.4]
  input   io_input_enable // @[:@518.4]
);
  wire  bases_0_clock; // @[Counter.scala 253:53:@531.4]
  wire  bases_0_reset; // @[Counter.scala 253:53:@531.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 253:53:@531.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 253:53:@531.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 253:53:@531.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 253:53:@531.4]
  wire [31:0] _T_36; // @[Counter.scala 339:61:@550.4]
  wire [32:0] _T_38; // @[Counter.scala 339:68:@551.4]
  wire [31:0] _T_39; // @[Counter.scala 339:68:@552.4]
  wire [31:0] _T_40; // @[Counter.scala 339:68:@553.4]
  FF bases_0 ( // @[Counter.scala 253:53:@531.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  assign _T_36 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 339:61:@550.4]
  assign _T_38 = $signed(_T_36) + $signed(32'sh1); // @[Counter.scala 339:68:@551.4]
  assign _T_39 = $signed(_T_36) + $signed(32'sh1); // @[Counter.scala 339:68:@552.4]
  assign _T_40 = $signed(_T_39); // @[Counter.scala 339:68:@553.4]
  assign bases_0_clock = clock; // @[:@532.4]
  assign bases_0_reset = reset; // @[:@533.4]
  assign bases_0_io_wPort_0_data_0 = $unsigned(_T_40); // @[Counter.scala 339:31:@555.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 337:27:@548.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 338:29:@549.4]
endmodule
module x24_ctrchain( // @[:@562.2]
  input   clock, // @[:@563.4]
  input   reset, // @[:@564.4]
  input   io_input_reset, // @[:@565.4]
  input   io_input_enable, // @[:@565.4]
  output  io_output_oobs_0 // @[:@565.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 505:46:@567.4]
  wire  ctrs_0_reset; // @[Counter.scala 505:46:@567.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 505:46:@567.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 505:46:@567.4]
  reg  doneLatch; // @[Counter.scala 542:26:@588.4]
  reg [31:0] _RAND_0;
  wire  _T_55; // @[Counter.scala 543:19:@590.4]
  SingleCounter_1 ctrs_0 ( // @[Counter.scala 505:46:@567.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable)
  );
  assign _T_55 = io_input_reset ? 1'h0 : doneLatch; // @[Counter.scala 543:19:@590.4]
  assign io_output_oobs_0 = doneLatch; // @[Counter.scala 550:30:@594.4]
  assign ctrs_0_clock = clock; // @[:@568.4]
  assign ctrs_0_reset = reset; // @[:@569.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 512:24:@573.4]
  assign ctrs_0_io_input_enable = io_input_enable; // @[Counter.scala 516:33:@574.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  doneLatch = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end
    end
  end
endmodule
module RetimeWrapper_5( // @[:@634.2]
  input   clock, // @[:@635.4]
  input   reset, // @[:@636.4]
  input   io_in, // @[:@637.4]
  output  io_out // @[:@637.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@639.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@639.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@639.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@639.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@639.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@639.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(5)) sr ( // @[RetimeShiftRegister.scala 15:20:@639.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@652.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@651.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@650.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@649.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@648.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@646.4]
endmodule
module RetimeWrapper_9( // @[:@762.2]
  input   clock, // @[:@763.4]
  input   reset, // @[:@764.4]
  input   io_in, // @[:@765.4]
  output  io_out // @[:@765.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@767.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@767.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@767.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@767.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@767.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@767.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(4)) sr ( // @[RetimeShiftRegister.scala 15:20:@767.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@780.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@779.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@778.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@777.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@776.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@774.4]
endmodule
module x35_inr_Foreach_SAMPLER_BOX_sm( // @[:@782.2]
  input   clock, // @[:@783.4]
  input   reset, // @[:@784.4]
  input   io_enable, // @[:@785.4]
  output  io_done, // @[:@785.4]
  input   io_ctrDone, // @[:@785.4]
  output  io_datapathEn, // @[:@785.4]
  output  io_ctrInc, // @[:@785.4]
  output  io_ctrRst, // @[:@785.4]
  input   io_parentAck // @[:@785.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@787.4]
  wire  active_reset; // @[Controllers.scala 261:22:@787.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@787.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@787.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@787.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@787.4]
  wire  done_clock; // @[Controllers.scala 262:20:@790.4]
  wire  done_reset; // @[Controllers.scala 262:20:@790.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@790.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@790.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@790.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@790.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@824.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@824.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@824.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@824.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@846.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@846.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@846.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@846.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@858.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@858.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@858.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@858.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@858.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@866.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@866.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@866.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@866.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@866.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@882.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@882.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@882.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@882.4]
  wire  _T_80; // @[Controllers.scala 264:48:@795.4]
  wire  _T_81; // @[Controllers.scala 264:46:@796.4]
  wire  _T_82; // @[Controllers.scala 264:62:@797.4]
  wire  _T_100; // @[package.scala 100:49:@815.4]
  reg  _T_103; // @[package.scala 48:56:@816.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@829.4 package.scala 96:25:@830.4]
  wire  _T_110; // @[package.scala 100:49:@831.4]
  reg  _T_113; // @[package.scala 48:56:@832.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@834.4]
  wire  _T_118; // @[Controllers.scala 283:41:@839.4]
  wire  _T_124; // @[package.scala 96:25:@851.4 package.scala 96:25:@852.4]
  wire  _T_126; // @[package.scala 100:49:@853.4]
  reg  _T_129; // @[package.scala 48:56:@854.4]
  reg [31:0] _RAND_2;
  wire  _T_150; // @[package.scala 100:49:@878.4]
  reg  _T_153; // @[package.scala 48:56:@879.4]
  reg [31:0] _RAND_3;
  SRFF active ( // @[Controllers.scala 261:22:@787.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@790.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_5 RetimeWrapper ( // @[package.scala 93:22:@824.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_5 RetimeWrapper_1 ( // @[package.scala 93:22:@846.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@858.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@866.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_9 RetimeWrapper_4 ( // @[package.scala 93:22:@882.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@795.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@796.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@797.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@815.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@829.4 package.scala 96:25:@830.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@831.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@834.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@839.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@851.4 package.scala 96:25:@852.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@853.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@878.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@857.4]
  assign io_datapathEn = _T_118 & io_enable; // @[Controllers.scala 283:21:@842.4]
  assign io_ctrInc = active_io_output & io_enable; // @[Controllers.scala 284:17:@845.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@837.4]
  assign active_clock = clock; // @[:@788.4]
  assign active_reset = reset; // @[:@789.4]
  assign active_io_input_set = _T_81 & _T_82; // @[Controllers.scala 264:23:@800.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@804.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@805.4]
  assign done_clock = clock; // @[:@791.4]
  assign done_reset = reset; // @[:@792.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@820.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@813.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@814.4]
  assign RetimeWrapper_clock = clock; // @[:@825.4]
  assign RetimeWrapper_reset = reset; // @[:@826.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@827.4]
  assign RetimeWrapper_1_clock = clock; // @[:@847.4]
  assign RetimeWrapper_1_reset = reset; // @[:@848.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@849.4]
  assign RetimeWrapper_2_clock = clock; // @[:@859.4]
  assign RetimeWrapper_2_reset = reset; // @[:@860.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@862.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@861.4]
  assign RetimeWrapper_3_clock = clock; // @[:@867.4]
  assign RetimeWrapper_3_reset = reset; // @[:@868.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@870.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@869.4]
  assign RetimeWrapper_4_clock = clock; // @[:@883.4]
  assign RetimeWrapper_4_reset = reset; // @[:@884.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@885.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_153 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module RetimeWrapper_13( // @[:@1048.2]
  input        clock, // @[:@1049.4]
  input        reset, // @[:@1050.4]
  input  [7:0] io_in, // @[:@1051.4]
  output [7:0] io_out // @[:@1051.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@1053.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@1053.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@1053.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@1053.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@1053.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@1053.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@1053.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@1066.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@1065.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@1064.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@1063.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@1062.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@1060.4]
endmodule
module SimBlackBoxesfix2fixBox_1( // @[:@1068.2]
  input  [7:0] io_a, // @[:@1071.4]
  output [8:0] io_b // @[:@1071.4]
);
  wire  _T_20; // @[implicits.scala 69:16:@1078.4]
  assign _T_20 = io_a[7]; // @[implicits.scala 69:16:@1078.4]
  assign io_b = {_T_20,io_a}; // @[SimBlackBoxes.scala 99:40:@1083.4]
endmodule
module __1( // @[:@1085.2]
  input  [7:0] io_b, // @[:@1088.4]
  output [8:0] io_result // @[:@1088.4]
);
  wire [7:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@1093.4]
  wire [8:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@1093.4]
  SimBlackBoxesfix2fixBox_1 SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@1093.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@1106.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@1101.4]
endmodule
module RetimeWrapper_14( // @[:@1160.2]
  input        clock, // @[:@1161.4]
  input        reset, // @[:@1162.4]
  input  [7:0] io_in, // @[:@1163.4]
  output [7:0] io_out // @[:@1163.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@1165.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@1165.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@1165.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@1165.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@1165.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@1165.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@1165.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@1178.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@1177.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@1176.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@1175.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@1174.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@1172.4]
endmodule
module fix2fixBox( // @[:@1180.2]
  input        clock, // @[:@1181.4]
  input        reset, // @[:@1182.4]
  input  [8:0] io_a, // @[:@1183.4]
  output [7:0] io_b // @[:@1183.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@1193.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@1193.4]
  wire [7:0] RetimeWrapper_io_in; // @[package.scala 93:22:@1193.4]
  wire [7:0] RetimeWrapper_io_out; // @[package.scala 93:22:@1193.4]
  RetimeWrapper_14 RetimeWrapper ( // @[package.scala 93:22:@1193.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@1200.4]
  assign RetimeWrapper_clock = clock; // @[:@1194.4]
  assign RetimeWrapper_reset = reset; // @[:@1195.4]
  assign RetimeWrapper_io_in = io_a[7:0]; // @[package.scala 94:16:@1196.4]
endmodule
module x31_sum( // @[:@1202.2]
  input        clock, // @[:@1203.4]
  input        reset, // @[:@1204.4]
  input  [7:0] io_a, // @[:@1205.4]
  output [7:0] io_result // @[:@1205.4]
);
  wire [7:0] __io_b; // @[Math.scala 709:24:@1213.4]
  wire [8:0] __io_result; // @[Math.scala 709:24:@1213.4]
  wire [7:0] __1_io_b; // @[Math.scala 709:24:@1220.4]
  wire [8:0] __1_io_result; // @[Math.scala 709:24:@1220.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@1238.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@1238.4]
  wire [8:0] fix2fixBox_io_a; // @[Math.scala 141:30:@1238.4]
  wire [7:0] fix2fixBox_io_b; // @[Math.scala 141:30:@1238.4]
  wire [8:0] a_upcast_number; // @[Math.scala 712:22:@1218.4 Math.scala 713:14:@1219.4]
  wire [8:0] b_upcast_number; // @[Math.scala 712:22:@1225.4 Math.scala 713:14:@1226.4]
  wire [9:0] _T_21; // @[Math.scala 136:37:@1227.4]
  __1 _ ( // @[Math.scala 709:24:@1213.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __1 __1 ( // @[Math.scala 709:24:@1220.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox fix2fixBox ( // @[Math.scala 141:30:@1238.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@1218.4 Math.scala 713:14:@1219.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@1225.4 Math.scala 713:14:@1226.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@1227.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@1246.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@1216.4]
  assign __1_io_b = 8'h5; // @[Math.scala 710:17:@1223.4]
  assign fix2fixBox_clock = clock; // @[:@1239.4]
  assign fix2fixBox_reset = reset; // @[:@1240.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@1241.4]
endmodule
module x35_inr_Foreach_SAMPLER_BOX_kernelx35_inr_Foreach_SAMPLER_BOX_concrete1( // @[:@1344.2]
  input          clock, // @[:@1345.4]
  input          reset, // @[:@1346.4]
  output         io_in_x21_TREADY, // @[:@1347.4]
  input  [255:0] io_in_x21_TDATA, // @[:@1347.4]
  input  [7:0]   io_in_x21_TID, // @[:@1347.4]
  input  [7:0]   io_in_x21_TDEST, // @[:@1347.4]
  output         io_in_x22_TVALID, // @[:@1347.4]
  output [255:0] io_in_x22_TDATA, // @[:@1347.4]
  input          io_sigsIn_datapathEn, // @[:@1347.4]
  input          io_sigsIn_cchainOutputs_0_oobs_0, // @[:@1347.4]
  input          io_rr // @[:@1347.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@1381.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@1381.4]
  wire [7:0] RetimeWrapper_io_in; // @[package.scala 93:22:@1381.4]
  wire [7:0] RetimeWrapper_io_out; // @[package.scala 93:22:@1381.4]
  wire  x31_sum_1_clock; // @[Math.scala 150:24:@1399.4]
  wire  x31_sum_1_reset; // @[Math.scala 150:24:@1399.4]
  wire [7:0] x31_sum_1_io_a; // @[Math.scala 150:24:@1399.4]
  wire [7:0] x31_sum_1_io_result; // @[Math.scala 150:24:@1399.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@1409.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@1409.4]
  wire [7:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@1409.4]
  wire [7:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@1409.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@1422.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@1422.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@1422.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@1422.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@1431.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@1431.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@1431.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@1431.4]
  wire  b26; // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 61:17:@1369.4]
  wire  _T_186; // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 63:24:@1371.4]
  wire  _T_189; // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 65:62:@1375.4]
  wire  _T_190; // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 65:49:@1376.4]
  wire  _T_192; // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 65:86:@1377.4]
  wire  _T_234; // @[package.scala 96:25:@1436.4 package.scala 96:25:@1437.4]
  wire  _T_236; // @[implicits.scala 55:10:@1438.4]
  wire  x38_b26_D4; // @[package.scala 96:25:@1427.4 package.scala 96:25:@1428.4]
  RetimeWrapper_13 RetimeWrapper ( // @[package.scala 93:22:@1381.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x31_sum x31_sum_1 ( // @[Math.scala 150:24:@1399.4]
    .clock(x31_sum_1_clock),
    .reset(x31_sum_1_reset),
    .io_a(x31_sum_1_io_a),
    .io_result(x31_sum_1_io_result)
  );
  RetimeWrapper_14 RetimeWrapper_1 ( // @[package.scala 93:22:@1409.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_9 RetimeWrapper_2 ( // @[package.scala 93:22:@1422.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_9 RetimeWrapper_3 ( // @[package.scala 93:22:@1431.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  assign b26 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 61:17:@1369.4]
  assign _T_186 = b26 & io_sigsIn_datapathEn; // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 63:24:@1371.4]
  assign _T_189 = 8'h0 == 8'h0; // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 65:62:@1375.4]
  assign _T_190 = _T_186 & _T_189; // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 65:49:@1376.4]
  assign _T_192 = io_in_x21_TDEST == 8'h0; // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 65:86:@1377.4]
  assign _T_234 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@1436.4 package.scala 96:25:@1437.4]
  assign _T_236 = io_rr ? _T_234 : 1'h0; // @[implicits.scala 55:10:@1438.4]
  assign x38_b26_D4 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@1427.4 package.scala 96:25:@1428.4]
  assign io_in_x21_TREADY = _T_190 & _T_192; // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 63:17:@1372.4 sm_x35_inr_Foreach_SAMPLER_BOX.scala 65:17:@1379.4]
  assign io_in_x22_TVALID = _T_236 & x38_b26_D4; // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 83:17:@1441.4]
  assign io_in_x22_TDATA = {{248'd0}, RetimeWrapper_1_io_out}; // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 84:19:@1442.4]
  assign RetimeWrapper_clock = clock; // @[:@1382.4]
  assign RetimeWrapper_reset = reset; // @[:@1383.4]
  assign RetimeWrapper_io_in = io_in_x21_TDATA[7:0]; // @[package.scala 94:16:@1384.4]
  assign x31_sum_1_clock = clock; // @[:@1400.4]
  assign x31_sum_1_reset = reset; // @[:@1401.4]
  assign x31_sum_1_io_a = RetimeWrapper_io_out; // @[Math.scala 151:17:@1402.4]
  assign RetimeWrapper_1_clock = clock; // @[:@1410.4]
  assign RetimeWrapper_1_reset = reset; // @[:@1411.4]
  assign RetimeWrapper_1_io_in = x31_sum_1_io_result; // @[package.scala 94:16:@1412.4]
  assign RetimeWrapper_2_clock = clock; // @[:@1423.4]
  assign RetimeWrapper_2_reset = reset; // @[:@1424.4]
  assign RetimeWrapper_2_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@1425.4]
  assign RetimeWrapper_3_clock = clock; // @[:@1432.4]
  assign RetimeWrapper_3_reset = reset; // @[:@1433.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@1434.4]
endmodule
module RootController_kernelRootController_concrete1( // @[:@1452.2]
  input          clock, // @[:@1453.4]
  input          reset, // @[:@1454.4]
  output         io_in_x21_TREADY, // @[:@1455.4]
  input  [255:0] io_in_x21_TDATA, // @[:@1455.4]
  input  [7:0]   io_in_x21_TID, // @[:@1455.4]
  input  [7:0]   io_in_x21_TDEST, // @[:@1455.4]
  output         io_in_x22_TVALID, // @[:@1455.4]
  output [255:0] io_in_x22_TDATA, // @[:@1455.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@1455.4]
  input          io_sigsIn_smChildAcks_0, // @[:@1455.4]
  output         io_sigsOut_smDoneIn_0, // @[:@1455.4]
  input          io_rr // @[:@1455.4]
);
  wire  x24_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@1465.4]
  wire  x24_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@1465.4]
  wire  x24_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@1465.4]
  wire  x24_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@1465.4]
  wire  x24_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@1465.4]
  wire  x35_inr_Foreach_SAMPLER_BOX_sm_clock; // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 32:18:@1517.4]
  wire  x35_inr_Foreach_SAMPLER_BOX_sm_reset; // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 32:18:@1517.4]
  wire  x35_inr_Foreach_SAMPLER_BOX_sm_io_enable; // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 32:18:@1517.4]
  wire  x35_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 32:18:@1517.4]
  wire  x35_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 32:18:@1517.4]
  wire  x35_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 32:18:@1517.4]
  wire  x35_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 32:18:@1517.4]
  wire  x35_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 32:18:@1517.4]
  wire  x35_inr_Foreach_SAMPLER_BOX_sm_io_parentAck; // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 32:18:@1517.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@1545.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@1545.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@1545.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@1545.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@1545.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@1585.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@1585.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@1585.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@1585.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@1585.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@1593.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@1593.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@1593.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@1593.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@1593.4]
  wire  x35_inr_Foreach_SAMPLER_BOX_kernelx35_inr_Foreach_SAMPLER_BOX_concrete1_clock; // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 92:24:@1624.4]
  wire  x35_inr_Foreach_SAMPLER_BOX_kernelx35_inr_Foreach_SAMPLER_BOX_concrete1_reset; // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 92:24:@1624.4]
  wire  x35_inr_Foreach_SAMPLER_BOX_kernelx35_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x21_TREADY; // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 92:24:@1624.4]
  wire [255:0] x35_inr_Foreach_SAMPLER_BOX_kernelx35_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x21_TDATA; // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 92:24:@1624.4]
  wire [7:0] x35_inr_Foreach_SAMPLER_BOX_kernelx35_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x21_TID; // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 92:24:@1624.4]
  wire [7:0] x35_inr_Foreach_SAMPLER_BOX_kernelx35_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x21_TDEST; // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 92:24:@1624.4]
  wire  x35_inr_Foreach_SAMPLER_BOX_kernelx35_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x22_TVALID; // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 92:24:@1624.4]
  wire [255:0] x35_inr_Foreach_SAMPLER_BOX_kernelx35_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x22_TDATA; // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 92:24:@1624.4]
  wire  x35_inr_Foreach_SAMPLER_BOX_kernelx35_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn; // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 92:24:@1624.4]
  wire  x35_inr_Foreach_SAMPLER_BOX_kernelx35_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 92:24:@1624.4]
  wire  x35_inr_Foreach_SAMPLER_BOX_kernelx35_inr_Foreach_SAMPLER_BOX_concrete1_io_rr; // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 92:24:@1624.4]
  wire  _T_233; // @[package.scala 96:25:@1550.4 package.scala 96:25:@1551.4]
  wire  _T_248; // @[package.scala 96:25:@1590.4 package.scala 96:25:@1591.4]
  wire  _T_254; // @[package.scala 96:25:@1598.4 package.scala 96:25:@1599.4]
  wire  _T_257; // @[SpatialBlocks.scala 110:93:@1601.4]
  wire  _T_259; // @[SpatialBlocks.scala 128:36:@1610.4]
  wire  _T_260; // @[SpatialBlocks.scala 128:78:@1611.4]
  x24_ctrchain x24_ctrchain ( // @[SpatialBlocks.scala 37:22:@1465.4]
    .clock(x24_ctrchain_clock),
    .reset(x24_ctrchain_reset),
    .io_input_reset(x24_ctrchain_io_input_reset),
    .io_input_enable(x24_ctrchain_io_input_enable),
    .io_output_oobs_0(x24_ctrchain_io_output_oobs_0)
  );
  x35_inr_Foreach_SAMPLER_BOX_sm x35_inr_Foreach_SAMPLER_BOX_sm ( // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 32:18:@1517.4]
    .clock(x35_inr_Foreach_SAMPLER_BOX_sm_clock),
    .reset(x35_inr_Foreach_SAMPLER_BOX_sm_reset),
    .io_enable(x35_inr_Foreach_SAMPLER_BOX_sm_io_enable),
    .io_done(x35_inr_Foreach_SAMPLER_BOX_sm_io_done),
    .io_ctrDone(x35_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone),
    .io_datapathEn(x35_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn),
    .io_ctrInc(x35_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc),
    .io_ctrRst(x35_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst),
    .io_parentAck(x35_inr_Foreach_SAMPLER_BOX_sm_io_parentAck)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@1545.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@1585.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@1593.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x35_inr_Foreach_SAMPLER_BOX_kernelx35_inr_Foreach_SAMPLER_BOX_concrete1 x35_inr_Foreach_SAMPLER_BOX_kernelx35_inr_Foreach_SAMPLER_BOX_concrete1 ( // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 92:24:@1624.4]
    .clock(x35_inr_Foreach_SAMPLER_BOX_kernelx35_inr_Foreach_SAMPLER_BOX_concrete1_clock),
    .reset(x35_inr_Foreach_SAMPLER_BOX_kernelx35_inr_Foreach_SAMPLER_BOX_concrete1_reset),
    .io_in_x21_TREADY(x35_inr_Foreach_SAMPLER_BOX_kernelx35_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x21_TREADY),
    .io_in_x21_TDATA(x35_inr_Foreach_SAMPLER_BOX_kernelx35_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x21_TDATA),
    .io_in_x21_TID(x35_inr_Foreach_SAMPLER_BOX_kernelx35_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x21_TID),
    .io_in_x21_TDEST(x35_inr_Foreach_SAMPLER_BOX_kernelx35_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x21_TDEST),
    .io_in_x22_TVALID(x35_inr_Foreach_SAMPLER_BOX_kernelx35_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x22_TVALID),
    .io_in_x22_TDATA(x35_inr_Foreach_SAMPLER_BOX_kernelx35_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x22_TDATA),
    .io_sigsIn_datapathEn(x35_inr_Foreach_SAMPLER_BOX_kernelx35_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_cchainOutputs_0_oobs_0(x35_inr_Foreach_SAMPLER_BOX_kernelx35_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_rr(x35_inr_Foreach_SAMPLER_BOX_kernelx35_inr_Foreach_SAMPLER_BOX_concrete1_io_rr)
  );
  assign _T_233 = RetimeWrapper_io_out; // @[package.scala 96:25:@1550.4 package.scala 96:25:@1551.4]
  assign _T_248 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@1590.4 package.scala 96:25:@1591.4]
  assign _T_254 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@1598.4 package.scala 96:25:@1599.4]
  assign _T_257 = ~ _T_254; // @[SpatialBlocks.scala 110:93:@1601.4]
  assign _T_259 = x35_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[SpatialBlocks.scala 128:36:@1610.4]
  assign _T_260 = ~ x35_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[SpatialBlocks.scala 128:78:@1611.4]
  assign io_in_x21_TREADY = x35_inr_Foreach_SAMPLER_BOX_kernelx35_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x21_TREADY; // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 48:22:@1679.4]
  assign io_in_x22_TVALID = x35_inr_Foreach_SAMPLER_BOX_kernelx35_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x22_TVALID; // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 49:22:@1689.4]
  assign io_in_x22_TDATA = x35_inr_Foreach_SAMPLER_BOX_kernelx35_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x22_TDATA; // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 49:22:@1687.4]
  assign io_sigsOut_smDoneIn_0 = x35_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[SpatialBlocks.scala 127:53:@1608.4]
  assign x24_ctrchain_clock = clock; // @[:@1466.4]
  assign x24_ctrchain_reset = reset; // @[:@1467.4]
  assign x24_ctrchain_io_input_reset = x35_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[SpatialBlocks.scala 130:103:@1623.4]
  assign x24_ctrchain_io_input_enable = x35_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[SpatialBlocks.scala 104:75:@1578.4 SpatialBlocks.scala 130:45:@1622.4]
  assign x35_inr_Foreach_SAMPLER_BOX_sm_clock = clock; // @[:@1518.4]
  assign x35_inr_Foreach_SAMPLER_BOX_sm_reset = reset; // @[:@1519.4]
  assign x35_inr_Foreach_SAMPLER_BOX_sm_io_enable = _T_248 & _T_257; // @[SpatialBlocks.scala 112:18:@1605.4]
  assign x35_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone = io_rr ? _T_233 : 1'h0; // @[sm_RootController.scala 65:49:@1553.4]
  assign x35_inr_Foreach_SAMPLER_BOX_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 114:21:@1607.4]
  assign RetimeWrapper_clock = clock; // @[:@1546.4]
  assign RetimeWrapper_reset = reset; // @[:@1547.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@1549.4]
  assign RetimeWrapper_io_in = 1'h0; // @[package.scala 94:16:@1548.4]
  assign RetimeWrapper_1_clock = clock; // @[:@1586.4]
  assign RetimeWrapper_1_reset = reset; // @[:@1587.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@1589.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@1588.4]
  assign RetimeWrapper_2_clock = clock; // @[:@1594.4]
  assign RetimeWrapper_2_reset = reset; // @[:@1595.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@1597.4]
  assign RetimeWrapper_2_io_in = x35_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[package.scala 94:16:@1596.4]
  assign x35_inr_Foreach_SAMPLER_BOX_kernelx35_inr_Foreach_SAMPLER_BOX_concrete1_clock = clock; // @[:@1625.4]
  assign x35_inr_Foreach_SAMPLER_BOX_kernelx35_inr_Foreach_SAMPLER_BOX_concrete1_reset = reset; // @[:@1626.4]
  assign x35_inr_Foreach_SAMPLER_BOX_kernelx35_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x21_TDATA = io_in_x21_TDATA; // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 48:22:@1678.4]
  assign x35_inr_Foreach_SAMPLER_BOX_kernelx35_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x21_TID = io_in_x21_TID; // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 48:22:@1674.4]
  assign x35_inr_Foreach_SAMPLER_BOX_kernelx35_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x21_TDEST = io_in_x21_TDEST; // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 48:22:@1673.4]
  assign x35_inr_Foreach_SAMPLER_BOX_kernelx35_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn = _T_259 & _T_260; // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 96:22:@1702.4]
  assign x35_inr_Foreach_SAMPLER_BOX_kernelx35_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x24_ctrchain_io_output_oobs_0; // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 96:22:@1694.4]
  assign x35_inr_Foreach_SAMPLER_BOX_kernelx35_inr_Foreach_SAMPLER_BOX_concrete1_io_rr = io_rr; // @[sm_x35_inr_Foreach_SAMPLER_BOX.scala 95:18:@1690.4]
endmodule
module AccelUnit( // @[:@1717.2]
  input          clock, // @[:@1718.4]
  input          reset, // @[:@1719.4]
  input          io_enable, // @[:@1720.4]
  output         io_done, // @[:@1720.4]
  input          io_reset, // @[:@1720.4]
  input          io_memStreams_loads_0_cmd_ready, // @[:@1720.4]
  output         io_memStreams_loads_0_cmd_valid, // @[:@1720.4]
  output [63:0]  io_memStreams_loads_0_cmd_bits_addr, // @[:@1720.4]
  output [31:0]  io_memStreams_loads_0_cmd_bits_size, // @[:@1720.4]
  output         io_memStreams_loads_0_data_ready, // @[:@1720.4]
  input          io_memStreams_loads_0_data_valid, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_0, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_1, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_2, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_3, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_4, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_5, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_6, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_7, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_8, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_9, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_10, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_11, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_12, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_13, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_14, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_15, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_16, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_17, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_18, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_19, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_20, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_21, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_22, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_23, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_24, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_25, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_26, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_27, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_28, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_29, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_30, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_31, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_32, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_33, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_34, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_35, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_36, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_37, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_38, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_39, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_40, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_41, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_42, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_43, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_44, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_45, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_46, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_47, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_48, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_49, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_50, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_51, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_52, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_53, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_54, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_55, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_56, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_57, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_58, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_59, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_60, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_61, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_62, // @[:@1720.4]
  input  [7:0]   io_memStreams_loads_0_data_bits_rdata_63, // @[:@1720.4]
  input          io_memStreams_stores_0_cmd_ready, // @[:@1720.4]
  output         io_memStreams_stores_0_cmd_valid, // @[:@1720.4]
  output [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@1720.4]
  output [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@1720.4]
  input          io_memStreams_stores_0_data_ready, // @[:@1720.4]
  output         io_memStreams_stores_0_data_valid, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_0, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_1, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_2, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_3, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_4, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_5, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_6, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_7, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_8, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_9, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_10, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_11, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_12, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_13, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_14, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_15, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_16, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_17, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_18, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_19, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_20, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_21, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_22, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_23, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_24, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_25, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_26, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_27, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_28, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_29, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_30, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_31, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_32, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_33, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_34, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_35, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_36, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_37, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_38, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_39, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_40, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_41, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_42, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_43, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_44, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_45, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_46, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_47, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_48, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_49, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_50, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_51, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_52, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_53, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_54, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_55, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_56, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_57, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_58, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_59, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_60, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_61, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_62, // @[:@1720.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_63, // @[:@1720.4]
  output [63:0]  io_memStreams_stores_0_data_bits_wstrb, // @[:@1720.4]
  output         io_memStreams_stores_0_wresp_ready, // @[:@1720.4]
  input          io_memStreams_stores_0_wresp_valid, // @[:@1720.4]
  input          io_memStreams_stores_0_wresp_bits, // @[:@1720.4]
  input          io_memStreams_gathers_0_cmd_ready, // @[:@1720.4]
  output         io_memStreams_gathers_0_cmd_valid, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_0, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_1, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_2, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_3, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_4, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_5, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_6, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_7, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_8, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_9, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_10, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_11, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_12, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_13, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_14, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_15, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_16, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_17, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_18, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_19, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_20, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_21, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_22, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_23, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_24, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_25, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_26, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_27, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_28, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_29, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_30, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_31, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_32, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_33, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_34, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_35, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_36, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_37, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_38, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_39, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_40, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_41, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_42, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_43, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_44, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_45, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_46, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_47, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_48, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_49, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_50, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_51, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_52, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_53, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_54, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_55, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_56, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_57, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_58, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_59, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_60, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_61, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_62, // @[:@1720.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_63, // @[:@1720.4]
  output         io_memStreams_gathers_0_data_ready, // @[:@1720.4]
  input          io_memStreams_gathers_0_data_valid, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_0, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_1, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_2, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_3, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_4, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_5, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_6, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_7, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_8, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_9, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_10, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_11, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_12, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_13, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_14, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_15, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_16, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_17, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_18, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_19, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_20, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_21, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_22, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_23, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_24, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_25, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_26, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_27, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_28, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_29, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_30, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_31, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_32, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_33, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_34, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_35, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_36, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_37, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_38, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_39, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_40, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_41, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_42, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_43, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_44, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_45, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_46, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_47, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_48, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_49, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_50, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_51, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_52, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_53, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_54, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_55, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_56, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_57, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_58, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_59, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_60, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_61, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_62, // @[:@1720.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_63, // @[:@1720.4]
  input          io_memStreams_scatters_0_cmd_ready, // @[:@1720.4]
  output         io_memStreams_scatters_0_cmd_valid, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_0, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_1, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_2, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_3, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_4, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_5, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_6, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_7, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_8, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_9, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_10, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_11, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_12, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_13, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_14, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_15, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_16, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_17, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_18, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_19, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_20, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_21, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_22, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_23, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_24, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_25, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_26, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_27, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_28, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_29, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_30, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_31, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_32, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_33, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_34, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_35, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_36, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_37, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_38, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_39, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_40, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_41, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_42, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_43, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_44, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_45, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_46, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_47, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_48, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_49, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_50, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_51, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_52, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_53, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_54, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_55, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_56, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_57, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_58, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_59, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_60, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_61, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_62, // @[:@1720.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_63, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_0, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_1, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_2, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_3, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_4, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_5, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_6, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_7, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_8, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_9, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_10, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_11, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_12, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_13, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_14, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_15, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_16, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_17, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_18, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_19, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_20, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_21, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_22, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_23, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_24, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_25, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_26, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_27, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_28, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_29, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_30, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_31, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_32, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_33, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_34, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_35, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_36, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_37, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_38, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_39, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_40, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_41, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_42, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_43, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_44, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_45, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_46, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_47, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_48, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_49, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_50, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_51, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_52, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_53, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_54, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_55, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_56, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_57, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_58, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_59, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_60, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_61, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_62, // @[:@1720.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_63, // @[:@1720.4]
  output         io_memStreams_scatters_0_wresp_ready, // @[:@1720.4]
  input          io_memStreams_scatters_0_wresp_valid, // @[:@1720.4]
  input          io_memStreams_scatters_0_wresp_bits, // @[:@1720.4]
  input          io_axiStreamsIn_0_TVALID, // @[:@1720.4]
  output         io_axiStreamsIn_0_TREADY, // @[:@1720.4]
  input  [255:0] io_axiStreamsIn_0_TDATA, // @[:@1720.4]
  input  [31:0]  io_axiStreamsIn_0_TSTRB, // @[:@1720.4]
  input  [31:0]  io_axiStreamsIn_0_TKEEP, // @[:@1720.4]
  input          io_axiStreamsIn_0_TLAST, // @[:@1720.4]
  input  [7:0]   io_axiStreamsIn_0_TID, // @[:@1720.4]
  input  [7:0]   io_axiStreamsIn_0_TDEST, // @[:@1720.4]
  input  [31:0]  io_axiStreamsIn_0_TUSER, // @[:@1720.4]
  output         io_axiStreamsOut_0_TVALID, // @[:@1720.4]
  input          io_axiStreamsOut_0_TREADY, // @[:@1720.4]
  output [255:0] io_axiStreamsOut_0_TDATA, // @[:@1720.4]
  output [31:0]  io_axiStreamsOut_0_TSTRB, // @[:@1720.4]
  output [31:0]  io_axiStreamsOut_0_TKEEP, // @[:@1720.4]
  output         io_axiStreamsOut_0_TLAST, // @[:@1720.4]
  output [7:0]   io_axiStreamsOut_0_TID, // @[:@1720.4]
  output [7:0]   io_axiStreamsOut_0_TDEST, // @[:@1720.4]
  output [31:0]  io_axiStreamsOut_0_TUSER, // @[:@1720.4]
  output         io_heap_0_req_valid, // @[:@1720.4]
  output         io_heap_0_req_bits_allocDealloc, // @[:@1720.4]
  output [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@1720.4]
  input          io_heap_0_resp_valid, // @[:@1720.4]
  input          io_heap_0_resp_bits_allocDealloc, // @[:@1720.4]
  input  [63:0]  io_heap_0_resp_bits_sizeAddr, // @[:@1720.4]
  input  [63:0]  io_argIns_0, // @[:@1720.4]
  input          io_argOuts_0_port_ready, // @[:@1720.4]
  output         io_argOuts_0_port_valid, // @[:@1720.4]
  output [63:0]  io_argOuts_0_port_bits, // @[:@1720.4]
  input  [63:0]  io_argOuts_0_echo // @[:@1720.4]
);
  wire  SingleCounter_clock; // @[Main.scala 29:32:@2166.4]
  wire  SingleCounter_reset; // @[Main.scala 29:32:@2166.4]
  wire  SingleCounter_io_input_reset; // @[Main.scala 29:32:@2166.4]
  wire  SingleCounter_io_output_done; // @[Main.scala 29:32:@2166.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@2184.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@2184.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@2184.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@2184.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@2184.4]
  wire  SRFF_clock; // @[Main.scala 33:28:@2193.4]
  wire  SRFF_reset; // @[Main.scala 33:28:@2193.4]
  wire  SRFF_io_input_set; // @[Main.scala 33:28:@2193.4]
  wire  SRFF_io_input_reset; // @[Main.scala 33:28:@2193.4]
  wire  SRFF_io_input_asyn_reset; // @[Main.scala 33:28:@2193.4]
  wire  SRFF_io_output; // @[Main.scala 33:28:@2193.4]
  wire  RootController_sm_clock; // @[sm_RootController.scala 32:18:@2231.4]
  wire  RootController_sm_reset; // @[sm_RootController.scala 32:18:@2231.4]
  wire  RootController_sm_io_enable; // @[sm_RootController.scala 32:18:@2231.4]
  wire  RootController_sm_io_done; // @[sm_RootController.scala 32:18:@2231.4]
  wire  RootController_sm_io_rst; // @[sm_RootController.scala 32:18:@2231.4]
  wire  RootController_sm_io_ctrDone; // @[sm_RootController.scala 32:18:@2231.4]
  wire  RootController_sm_io_ctrInc; // @[sm_RootController.scala 32:18:@2231.4]
  wire  RootController_sm_io_doneIn_0; // @[sm_RootController.scala 32:18:@2231.4]
  wire  RootController_sm_io_enableOut_0; // @[sm_RootController.scala 32:18:@2231.4]
  wire  RootController_sm_io_childAck_0; // @[sm_RootController.scala 32:18:@2231.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@2263.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@2263.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@2263.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@2263.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@2263.4]
  wire  RootController_kernelRootController_concrete1_clock; // @[sm_RootController.scala 74:24:@2322.4]
  wire  RootController_kernelRootController_concrete1_reset; // @[sm_RootController.scala 74:24:@2322.4]
  wire  RootController_kernelRootController_concrete1_io_in_x21_TREADY; // @[sm_RootController.scala 74:24:@2322.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x21_TDATA; // @[sm_RootController.scala 74:24:@2322.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x21_TID; // @[sm_RootController.scala 74:24:@2322.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x21_TDEST; // @[sm_RootController.scala 74:24:@2322.4]
  wire  RootController_kernelRootController_concrete1_io_in_x22_TVALID; // @[sm_RootController.scala 74:24:@2322.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x22_TDATA; // @[sm_RootController.scala 74:24:@2322.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_RootController.scala 74:24:@2322.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0; // @[sm_RootController.scala 74:24:@2322.4]
  wire  RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[sm_RootController.scala 74:24:@2322.4]
  wire  RootController_kernelRootController_concrete1_io_rr; // @[sm_RootController.scala 74:24:@2322.4]
  wire  _T_785; // @[package.scala 96:25:@2189.4 package.scala 96:25:@2190.4]
  wire  _T_850; // @[Main.scala 35:50:@2259.4]
  wire  _T_851; // @[Main.scala 35:59:@2260.4]
  wire  _T_863; // @[package.scala 100:49:@2280.4]
  reg  _T_866; // @[package.scala 48:56:@2281.4]
  reg [31:0] _RAND_0;
  SingleCounter SingleCounter ( // @[Main.scala 29:32:@2166.4]
    .clock(SingleCounter_clock),
    .reset(SingleCounter_reset),
    .io_input_reset(SingleCounter_io_input_reset),
    .io_output_done(SingleCounter_io_output_done)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@2184.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  SRFF SRFF ( // @[Main.scala 33:28:@2193.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  RootController_sm RootController_sm ( // @[sm_RootController.scala 32:18:@2231.4]
    .clock(RootController_sm_clock),
    .reset(RootController_sm_reset),
    .io_enable(RootController_sm_io_enable),
    .io_done(RootController_sm_io_done),
    .io_rst(RootController_sm_io_rst),
    .io_ctrDone(RootController_sm_io_ctrDone),
    .io_ctrInc(RootController_sm_io_ctrInc),
    .io_doneIn_0(RootController_sm_io_doneIn_0),
    .io_enableOut_0(RootController_sm_io_enableOut_0),
    .io_childAck_0(RootController_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@2263.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RootController_kernelRootController_concrete1 RootController_kernelRootController_concrete1 ( // @[sm_RootController.scala 74:24:@2322.4]
    .clock(RootController_kernelRootController_concrete1_clock),
    .reset(RootController_kernelRootController_concrete1_reset),
    .io_in_x21_TREADY(RootController_kernelRootController_concrete1_io_in_x21_TREADY),
    .io_in_x21_TDATA(RootController_kernelRootController_concrete1_io_in_x21_TDATA),
    .io_in_x21_TID(RootController_kernelRootController_concrete1_io_in_x21_TID),
    .io_in_x21_TDEST(RootController_kernelRootController_concrete1_io_in_x21_TDEST),
    .io_in_x22_TVALID(RootController_kernelRootController_concrete1_io_in_x22_TVALID),
    .io_in_x22_TDATA(RootController_kernelRootController_concrete1_io_in_x22_TDATA),
    .io_sigsIn_smEnableOuts_0(RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(RootController_kernelRootController_concrete1_io_rr)
  );
  assign _T_785 = RetimeWrapper_io_out; // @[package.scala 96:25:@2189.4 package.scala 96:25:@2190.4]
  assign _T_850 = io_enable & _T_785; // @[Main.scala 35:50:@2259.4]
  assign _T_851 = ~ SRFF_io_output; // @[Main.scala 35:59:@2260.4]
  assign _T_863 = RootController_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@2280.4]
  assign io_done = SRFF_io_output; // @[Main.scala 42:23:@2279.4]
  assign io_memStreams_loads_0_cmd_valid = 1'h0;
  assign io_memStreams_loads_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_loads_0_cmd_bits_size = 32'h0;
  assign io_memStreams_loads_0_data_ready = 1'h0;
  assign io_memStreams_stores_0_cmd_valid = 1'h0;
  assign io_memStreams_stores_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_stores_0_cmd_bits_size = 32'h0;
  assign io_memStreams_stores_0_data_valid = 1'h0;
  assign io_memStreams_stores_0_data_bits_wdata_0 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_1 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_2 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_3 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_4 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_5 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_6 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_7 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_8 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_9 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_10 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_11 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_12 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_13 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_14 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_15 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_16 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_17 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_18 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_19 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_20 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_21 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_22 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_23 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_24 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_25 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_26 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_27 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_28 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_29 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_30 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_31 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_32 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_33 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_34 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_35 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_36 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_37 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_38 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_39 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_40 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_41 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_42 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_43 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_44 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_45 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_46 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_47 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_48 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_49 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_50 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_51 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_52 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_53 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_54 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_55 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_56 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_57 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_58 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_59 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_60 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_61 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_62 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wdata_63 = 8'h0;
  assign io_memStreams_stores_0_data_bits_wstrb = 64'h0;
  assign io_memStreams_stores_0_wresp_ready = 1'h0;
  assign io_memStreams_gathers_0_cmd_valid = 1'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_0 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_1 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_2 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_3 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_4 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_5 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_6 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_7 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_8 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_9 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_10 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_11 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_12 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_13 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_14 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_15 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_16 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_17 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_18 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_19 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_20 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_21 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_22 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_23 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_24 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_25 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_26 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_27 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_28 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_29 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_30 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_31 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_32 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_33 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_34 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_35 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_36 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_37 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_38 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_39 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_40 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_41 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_42 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_43 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_44 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_45 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_46 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_47 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_48 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_49 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_50 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_51 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_52 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_53 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_54 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_55 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_56 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_57 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_58 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_59 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_60 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_61 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_62 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_63 = 64'h0;
  assign io_memStreams_gathers_0_data_ready = 1'h0;
  assign io_memStreams_scatters_0_cmd_valid = 1'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_0 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_1 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_2 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_3 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_4 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_5 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_6 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_7 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_8 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_9 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_10 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_11 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_12 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_13 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_14 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_15 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_16 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_17 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_18 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_19 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_20 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_21 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_22 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_23 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_24 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_25 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_26 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_27 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_28 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_29 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_30 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_31 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_32 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_33 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_34 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_35 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_36 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_37 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_38 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_39 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_40 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_41 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_42 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_43 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_44 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_45 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_46 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_47 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_48 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_49 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_50 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_51 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_52 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_53 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_54 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_55 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_56 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_57 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_58 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_59 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_60 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_61 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_62 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_63 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_0 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_1 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_2 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_3 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_4 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_5 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_6 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_7 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_8 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_9 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_10 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_11 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_12 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_13 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_14 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_15 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_16 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_17 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_18 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_19 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_20 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_21 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_22 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_23 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_24 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_25 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_26 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_27 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_28 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_29 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_30 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_31 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_32 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_33 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_34 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_35 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_36 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_37 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_38 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_39 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_40 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_41 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_42 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_43 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_44 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_45 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_46 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_47 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_48 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_49 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_50 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_51 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_52 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_53 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_54 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_55 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_56 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_57 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_58 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_59 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_60 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_61 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_62 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_63 = 8'h0;
  assign io_memStreams_scatters_0_wresp_ready = 1'h0;
  assign io_axiStreamsIn_0_TREADY = RootController_kernelRootController_concrete1_io_in_x21_TREADY; // @[sm_RootController.scala 48:22:@2377.4]
  assign io_axiStreamsOut_0_TVALID = RootController_kernelRootController_concrete1_io_in_x22_TVALID; // @[sm_RootController.scala 49:22:@2387.4]
  assign io_axiStreamsOut_0_TDATA = RootController_kernelRootController_concrete1_io_in_x22_TDATA; // @[sm_RootController.scala 49:22:@2385.4]
  assign io_axiStreamsOut_0_TSTRB = 32'hffffffff; // @[sm_RootController.scala 49:22:@2384.4]
  assign io_axiStreamsOut_0_TKEEP = 32'hffffffff; // @[sm_RootController.scala 49:22:@2383.4]
  assign io_axiStreamsOut_0_TLAST = 1'h0; // @[sm_RootController.scala 49:22:@2382.4]
  assign io_axiStreamsOut_0_TID = 8'h0; // @[sm_RootController.scala 49:22:@2381.4]
  assign io_axiStreamsOut_0_TDEST = 8'h0; // @[sm_RootController.scala 49:22:@2380.4]
  assign io_axiStreamsOut_0_TUSER = 32'h4; // @[sm_RootController.scala 49:22:@2379.4]
  assign io_heap_0_req_valid = 1'h0;
  assign io_heap_0_req_bits_allocDealloc = 1'h0;
  assign io_heap_0_req_bits_sizeAddr = 64'h0;
  assign io_argOuts_0_port_valid = 1'h0;
  assign io_argOuts_0_port_bits = 64'h0;
  assign SingleCounter_clock = clock; // @[:@2167.4]
  assign SingleCounter_reset = reset; // @[:@2168.4]
  assign SingleCounter_io_input_reset = reset; // @[Main.scala 30:79:@2182.4]
  assign RetimeWrapper_clock = clock; // @[:@2185.4]
  assign RetimeWrapper_reset = reset; // @[:@2186.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@2188.4]
  assign RetimeWrapper_io_in = SingleCounter_io_output_done; // @[package.scala 94:16:@2187.4]
  assign SRFF_clock = clock; // @[:@2194.4]
  assign SRFF_reset = reset; // @[:@2195.4]
  assign SRFF_io_input_set = RootController_sm_io_done; // @[Main.scala 51:29:@2414.4]
  assign SRFF_io_input_reset = RetimeWrapper_1_io_out; // @[Main.scala 40:31:@2277.4]
  assign SRFF_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[Main.scala 41:36:@2278.4]
  assign RootController_sm_clock = clock; // @[:@2232.4]
  assign RootController_sm_reset = reset; // @[:@2233.4]
  assign RootController_sm_io_enable = _T_850 & _T_851; // @[Main.scala 39:33:@2276.4 SpatialBlocks.scala 112:18:@2310.4]
  assign RootController_sm_io_rst = RetimeWrapper_1_io_out; // @[SpatialBlocks.scala 106:15:@2304.4]
  assign RootController_sm_io_ctrDone = RootController_sm_io_ctrInc & _T_866; // @[Main.scala 43:34:@2284.4]
  assign RootController_sm_io_doneIn_0 = RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 102:67:@2301.4]
  assign RetimeWrapper_1_clock = clock; // @[:@2264.4]
  assign RetimeWrapper_1_reset = reset; // @[:@2265.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@2267.4]
  assign RetimeWrapper_1_io_in = reset | io_reset; // @[package.scala 94:16:@2266.4]
  assign RootController_kernelRootController_concrete1_clock = clock; // @[:@2323.4]
  assign RootController_kernelRootController_concrete1_reset = reset; // @[:@2324.4]
  assign RootController_kernelRootController_concrete1_io_in_x21_TDATA = io_axiStreamsIn_0_TDATA; // @[sm_RootController.scala 48:22:@2376.4]
  assign RootController_kernelRootController_concrete1_io_in_x21_TID = io_axiStreamsIn_0_TID; // @[sm_RootController.scala 48:22:@2372.4]
  assign RootController_kernelRootController_concrete1_io_in_x21_TDEST = io_axiStreamsIn_0_TDEST; // @[sm_RootController.scala 48:22:@2371.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0 = RootController_sm_io_enableOut_0; // @[sm_RootController.scala 78:22:@2396.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0 = RootController_sm_io_childAck_0; // @[sm_RootController.scala 78:22:@2394.4]
  assign RootController_kernelRootController_concrete1_io_rr = RetimeWrapper_io_out; // @[sm_RootController.scala 77:18:@2388.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_866 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_866 <= 1'h0;
    end else begin
      _T_866 <= _T_863;
    end
  end
endmodule
module DRAMHeap( // @[:@3705.2]
  input         io_accel_0_req_valid, // @[:@3708.4]
  input         io_accel_0_req_bits_allocDealloc, // @[:@3708.4]
  input  [63:0] io_accel_0_req_bits_sizeAddr, // @[:@3708.4]
  output        io_accel_0_resp_valid, // @[:@3708.4]
  output        io_accel_0_resp_bits_allocDealloc, // @[:@3708.4]
  output [63:0] io_accel_0_resp_bits_sizeAddr, // @[:@3708.4]
  output        io_host_0_req_valid, // @[:@3708.4]
  output        io_host_0_req_bits_allocDealloc, // @[:@3708.4]
  output [63:0] io_host_0_req_bits_sizeAddr, // @[:@3708.4]
  input         io_host_0_resp_valid, // @[:@3708.4]
  input         io_host_0_resp_bits_allocDealloc, // @[:@3708.4]
  input  [63:0] io_host_0_resp_bits_sizeAddr // @[:@3708.4]
);
  assign io_accel_0_resp_valid = io_host_0_resp_valid; // @[DRAMHeap.scala 24:18:@3715.4]
  assign io_accel_0_resp_bits_allocDealloc = io_host_0_resp_bits_allocDealloc; // @[DRAMHeap.scala 25:17:@3717.4]
  assign io_accel_0_resp_bits_sizeAddr = io_host_0_resp_bits_sizeAddr; // @[DRAMHeap.scala 25:17:@3716.4]
  assign io_host_0_req_valid = io_accel_0_req_valid; // @[DRAMHeap.scala 21:18:@3712.4]
  assign io_host_0_req_bits_allocDealloc = io_accel_0_req_bits_allocDealloc; // @[DRAMHeap.scala 21:18:@3711.4]
  assign io_host_0_req_bits_sizeAddr = io_accel_0_req_bits_sizeAddr; // @[DRAMHeap.scala 21:18:@3710.4]
endmodule
module RetimeWrapper_18( // @[:@3731.2]
  input         clock, // @[:@3732.4]
  input         reset, // @[:@3733.4]
  input         io_flow, // @[:@3734.4]
  input  [63:0] io_in, // @[:@3734.4]
  output [63:0] io_out // @[:@3734.4]
);
  wire [63:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@3736.4]
  wire [63:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@3736.4]
  wire [63:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@3736.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3736.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3736.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3736.4]
  RetimeShiftRegister #(.WIDTH(64), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@3736.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3749.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3748.4]
  assign sr_init = 64'h0; // @[RetimeShiftRegister.scala 19:16:@3747.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3746.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3745.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3743.4]
endmodule
module FringeFF( // @[:@3751.2]
  input         clock, // @[:@3752.4]
  input         reset, // @[:@3753.4]
  input  [63:0] io_in, // @[:@3754.4]
  input         io_reset, // @[:@3754.4]
  output [63:0] io_out, // @[:@3754.4]
  input         io_enable // @[:@3754.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3757.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3757.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3757.4]
  wire [63:0] RetimeWrapper_io_in; // @[package.scala 93:22:@3757.4]
  wire [63:0] RetimeWrapper_io_out; // @[package.scala 93:22:@3757.4]
  wire [63:0] _T_18; // @[package.scala 96:25:@3762.4 package.scala 96:25:@3763.4]
  wire [63:0] _GEN_0; // @[FringeFF.scala 21:27:@3768.6]
  RetimeWrapper_18 RetimeWrapper ( // @[package.scala 93:22:@3757.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@3762.4 package.scala 96:25:@3763.4]
  assign _GEN_0 = io_reset ? 64'h0 : _T_18; // @[FringeFF.scala 21:27:@3768.6]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@3774.4]
  assign RetimeWrapper_clock = clock; // @[:@3758.4]
  assign RetimeWrapper_reset = reset; // @[:@3759.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@3761.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _GEN_0; // @[package.scala 94:16:@3760.4]
endmodule
module MuxN( // @[:@32390.2]
  input  [63:0] io_ins_0, // @[:@32393.4]
  input  [63:0] io_ins_1, // @[:@32393.4]
  input  [63:0] io_ins_2, // @[:@32393.4]
  input  [63:0] io_ins_3, // @[:@32393.4]
  input  [63:0] io_ins_4, // @[:@32393.4]
  input  [63:0] io_ins_5, // @[:@32393.4]
  input  [63:0] io_ins_6, // @[:@32393.4]
  input  [63:0] io_ins_7, // @[:@32393.4]
  input  [63:0] io_ins_8, // @[:@32393.4]
  input  [63:0] io_ins_9, // @[:@32393.4]
  input  [63:0] io_ins_10, // @[:@32393.4]
  input  [63:0] io_ins_11, // @[:@32393.4]
  input  [63:0] io_ins_12, // @[:@32393.4]
  input  [63:0] io_ins_13, // @[:@32393.4]
  input  [63:0] io_ins_14, // @[:@32393.4]
  input  [63:0] io_ins_15, // @[:@32393.4]
  input  [63:0] io_ins_16, // @[:@32393.4]
  input  [63:0] io_ins_17, // @[:@32393.4]
  input  [63:0] io_ins_18, // @[:@32393.4]
  input  [63:0] io_ins_19, // @[:@32393.4]
  input  [63:0] io_ins_20, // @[:@32393.4]
  input  [63:0] io_ins_21, // @[:@32393.4]
  input  [63:0] io_ins_22, // @[:@32393.4]
  input  [63:0] io_ins_23, // @[:@32393.4]
  input  [63:0] io_ins_24, // @[:@32393.4]
  input  [63:0] io_ins_25, // @[:@32393.4]
  input  [63:0] io_ins_26, // @[:@32393.4]
  input  [63:0] io_ins_27, // @[:@32393.4]
  input  [63:0] io_ins_28, // @[:@32393.4]
  input  [63:0] io_ins_29, // @[:@32393.4]
  input  [63:0] io_ins_30, // @[:@32393.4]
  input  [63:0] io_ins_31, // @[:@32393.4]
  input  [63:0] io_ins_32, // @[:@32393.4]
  input  [63:0] io_ins_33, // @[:@32393.4]
  input  [63:0] io_ins_34, // @[:@32393.4]
  input  [63:0] io_ins_35, // @[:@32393.4]
  input  [63:0] io_ins_36, // @[:@32393.4]
  input  [63:0] io_ins_37, // @[:@32393.4]
  input  [63:0] io_ins_38, // @[:@32393.4]
  input  [63:0] io_ins_39, // @[:@32393.4]
  input  [63:0] io_ins_40, // @[:@32393.4]
  input  [63:0] io_ins_41, // @[:@32393.4]
  input  [63:0] io_ins_42, // @[:@32393.4]
  input  [63:0] io_ins_43, // @[:@32393.4]
  input  [63:0] io_ins_44, // @[:@32393.4]
  input  [63:0] io_ins_45, // @[:@32393.4]
  input  [63:0] io_ins_46, // @[:@32393.4]
  input  [63:0] io_ins_47, // @[:@32393.4]
  input  [63:0] io_ins_48, // @[:@32393.4]
  input  [63:0] io_ins_49, // @[:@32393.4]
  input  [63:0] io_ins_50, // @[:@32393.4]
  input  [63:0] io_ins_51, // @[:@32393.4]
  input  [63:0] io_ins_52, // @[:@32393.4]
  input  [63:0] io_ins_53, // @[:@32393.4]
  input  [63:0] io_ins_54, // @[:@32393.4]
  input  [63:0] io_ins_55, // @[:@32393.4]
  input  [63:0] io_ins_56, // @[:@32393.4]
  input  [63:0] io_ins_57, // @[:@32393.4]
  input  [63:0] io_ins_58, // @[:@32393.4]
  input  [63:0] io_ins_59, // @[:@32393.4]
  input  [63:0] io_ins_60, // @[:@32393.4]
  input  [63:0] io_ins_61, // @[:@32393.4]
  input  [63:0] io_ins_62, // @[:@32393.4]
  input  [63:0] io_ins_63, // @[:@32393.4]
  input  [63:0] io_ins_64, // @[:@32393.4]
  input  [63:0] io_ins_65, // @[:@32393.4]
  input  [63:0] io_ins_66, // @[:@32393.4]
  input  [63:0] io_ins_67, // @[:@32393.4]
  input  [63:0] io_ins_68, // @[:@32393.4]
  input  [63:0] io_ins_69, // @[:@32393.4]
  input  [63:0] io_ins_70, // @[:@32393.4]
  input  [63:0] io_ins_71, // @[:@32393.4]
  input  [63:0] io_ins_72, // @[:@32393.4]
  input  [63:0] io_ins_73, // @[:@32393.4]
  input  [63:0] io_ins_74, // @[:@32393.4]
  input  [63:0] io_ins_75, // @[:@32393.4]
  input  [63:0] io_ins_76, // @[:@32393.4]
  input  [63:0] io_ins_77, // @[:@32393.4]
  input  [63:0] io_ins_78, // @[:@32393.4]
  input  [63:0] io_ins_79, // @[:@32393.4]
  input  [63:0] io_ins_80, // @[:@32393.4]
  input  [63:0] io_ins_81, // @[:@32393.4]
  input  [63:0] io_ins_82, // @[:@32393.4]
  input  [63:0] io_ins_83, // @[:@32393.4]
  input  [63:0] io_ins_84, // @[:@32393.4]
  input  [63:0] io_ins_85, // @[:@32393.4]
  input  [63:0] io_ins_86, // @[:@32393.4]
  input  [63:0] io_ins_87, // @[:@32393.4]
  input  [63:0] io_ins_88, // @[:@32393.4]
  input  [63:0] io_ins_89, // @[:@32393.4]
  input  [63:0] io_ins_90, // @[:@32393.4]
  input  [63:0] io_ins_91, // @[:@32393.4]
  input  [63:0] io_ins_92, // @[:@32393.4]
  input  [63:0] io_ins_93, // @[:@32393.4]
  input  [63:0] io_ins_94, // @[:@32393.4]
  input  [63:0] io_ins_95, // @[:@32393.4]
  input  [63:0] io_ins_96, // @[:@32393.4]
  input  [63:0] io_ins_97, // @[:@32393.4]
  input  [63:0] io_ins_98, // @[:@32393.4]
  input  [63:0] io_ins_99, // @[:@32393.4]
  input  [63:0] io_ins_100, // @[:@32393.4]
  input  [63:0] io_ins_101, // @[:@32393.4]
  input  [63:0] io_ins_102, // @[:@32393.4]
  input  [63:0] io_ins_103, // @[:@32393.4]
  input  [63:0] io_ins_104, // @[:@32393.4]
  input  [63:0] io_ins_105, // @[:@32393.4]
  input  [63:0] io_ins_106, // @[:@32393.4]
  input  [63:0] io_ins_107, // @[:@32393.4]
  input  [63:0] io_ins_108, // @[:@32393.4]
  input  [63:0] io_ins_109, // @[:@32393.4]
  input  [63:0] io_ins_110, // @[:@32393.4]
  input  [63:0] io_ins_111, // @[:@32393.4]
  input  [63:0] io_ins_112, // @[:@32393.4]
  input  [63:0] io_ins_113, // @[:@32393.4]
  input  [63:0] io_ins_114, // @[:@32393.4]
  input  [63:0] io_ins_115, // @[:@32393.4]
  input  [63:0] io_ins_116, // @[:@32393.4]
  input  [63:0] io_ins_117, // @[:@32393.4]
  input  [63:0] io_ins_118, // @[:@32393.4]
  input  [63:0] io_ins_119, // @[:@32393.4]
  input  [63:0] io_ins_120, // @[:@32393.4]
  input  [63:0] io_ins_121, // @[:@32393.4]
  input  [63:0] io_ins_122, // @[:@32393.4]
  input  [63:0] io_ins_123, // @[:@32393.4]
  input  [63:0] io_ins_124, // @[:@32393.4]
  input  [63:0] io_ins_125, // @[:@32393.4]
  input  [63:0] io_ins_126, // @[:@32393.4]
  input  [63:0] io_ins_127, // @[:@32393.4]
  input  [63:0] io_ins_128, // @[:@32393.4]
  input  [63:0] io_ins_129, // @[:@32393.4]
  input  [63:0] io_ins_130, // @[:@32393.4]
  input  [63:0] io_ins_131, // @[:@32393.4]
  input  [63:0] io_ins_132, // @[:@32393.4]
  input  [63:0] io_ins_133, // @[:@32393.4]
  input  [63:0] io_ins_134, // @[:@32393.4]
  input  [63:0] io_ins_135, // @[:@32393.4]
  input  [63:0] io_ins_136, // @[:@32393.4]
  input  [63:0] io_ins_137, // @[:@32393.4]
  input  [63:0] io_ins_138, // @[:@32393.4]
  input  [63:0] io_ins_139, // @[:@32393.4]
  input  [63:0] io_ins_140, // @[:@32393.4]
  input  [63:0] io_ins_141, // @[:@32393.4]
  input  [63:0] io_ins_142, // @[:@32393.4]
  input  [63:0] io_ins_143, // @[:@32393.4]
  input  [63:0] io_ins_144, // @[:@32393.4]
  input  [63:0] io_ins_145, // @[:@32393.4]
  input  [63:0] io_ins_146, // @[:@32393.4]
  input  [63:0] io_ins_147, // @[:@32393.4]
  input  [63:0] io_ins_148, // @[:@32393.4]
  input  [63:0] io_ins_149, // @[:@32393.4]
  input  [63:0] io_ins_150, // @[:@32393.4]
  input  [63:0] io_ins_151, // @[:@32393.4]
  input  [63:0] io_ins_152, // @[:@32393.4]
  input  [63:0] io_ins_153, // @[:@32393.4]
  input  [63:0] io_ins_154, // @[:@32393.4]
  input  [63:0] io_ins_155, // @[:@32393.4]
  input  [63:0] io_ins_156, // @[:@32393.4]
  input  [63:0] io_ins_157, // @[:@32393.4]
  input  [63:0] io_ins_158, // @[:@32393.4]
  input  [63:0] io_ins_159, // @[:@32393.4]
  input  [63:0] io_ins_160, // @[:@32393.4]
  input  [63:0] io_ins_161, // @[:@32393.4]
  input  [63:0] io_ins_162, // @[:@32393.4]
  input  [63:0] io_ins_163, // @[:@32393.4]
  input  [63:0] io_ins_164, // @[:@32393.4]
  input  [63:0] io_ins_165, // @[:@32393.4]
  input  [63:0] io_ins_166, // @[:@32393.4]
  input  [63:0] io_ins_167, // @[:@32393.4]
  input  [63:0] io_ins_168, // @[:@32393.4]
  input  [63:0] io_ins_169, // @[:@32393.4]
  input  [63:0] io_ins_170, // @[:@32393.4]
  input  [63:0] io_ins_171, // @[:@32393.4]
  input  [63:0] io_ins_172, // @[:@32393.4]
  input  [63:0] io_ins_173, // @[:@32393.4]
  input  [63:0] io_ins_174, // @[:@32393.4]
  input  [63:0] io_ins_175, // @[:@32393.4]
  input  [63:0] io_ins_176, // @[:@32393.4]
  input  [63:0] io_ins_177, // @[:@32393.4]
  input  [63:0] io_ins_178, // @[:@32393.4]
  input  [63:0] io_ins_179, // @[:@32393.4]
  input  [63:0] io_ins_180, // @[:@32393.4]
  input  [63:0] io_ins_181, // @[:@32393.4]
  input  [63:0] io_ins_182, // @[:@32393.4]
  input  [63:0] io_ins_183, // @[:@32393.4]
  input  [63:0] io_ins_184, // @[:@32393.4]
  input  [63:0] io_ins_185, // @[:@32393.4]
  input  [63:0] io_ins_186, // @[:@32393.4]
  input  [63:0] io_ins_187, // @[:@32393.4]
  input  [63:0] io_ins_188, // @[:@32393.4]
  input  [63:0] io_ins_189, // @[:@32393.4]
  input  [63:0] io_ins_190, // @[:@32393.4]
  input  [63:0] io_ins_191, // @[:@32393.4]
  input  [63:0] io_ins_192, // @[:@32393.4]
  input  [63:0] io_ins_193, // @[:@32393.4]
  input  [63:0] io_ins_194, // @[:@32393.4]
  input  [63:0] io_ins_195, // @[:@32393.4]
  input  [63:0] io_ins_196, // @[:@32393.4]
  input  [63:0] io_ins_197, // @[:@32393.4]
  input  [63:0] io_ins_198, // @[:@32393.4]
  input  [63:0] io_ins_199, // @[:@32393.4]
  input  [63:0] io_ins_200, // @[:@32393.4]
  input  [63:0] io_ins_201, // @[:@32393.4]
  input  [63:0] io_ins_202, // @[:@32393.4]
  input  [63:0] io_ins_203, // @[:@32393.4]
  input  [63:0] io_ins_204, // @[:@32393.4]
  input  [63:0] io_ins_205, // @[:@32393.4]
  input  [63:0] io_ins_206, // @[:@32393.4]
  input  [63:0] io_ins_207, // @[:@32393.4]
  input  [63:0] io_ins_208, // @[:@32393.4]
  input  [63:0] io_ins_209, // @[:@32393.4]
  input  [63:0] io_ins_210, // @[:@32393.4]
  input  [63:0] io_ins_211, // @[:@32393.4]
  input  [63:0] io_ins_212, // @[:@32393.4]
  input  [63:0] io_ins_213, // @[:@32393.4]
  input  [63:0] io_ins_214, // @[:@32393.4]
  input  [63:0] io_ins_215, // @[:@32393.4]
  input  [63:0] io_ins_216, // @[:@32393.4]
  input  [63:0] io_ins_217, // @[:@32393.4]
  input  [63:0] io_ins_218, // @[:@32393.4]
  input  [63:0] io_ins_219, // @[:@32393.4]
  input  [63:0] io_ins_220, // @[:@32393.4]
  input  [63:0] io_ins_221, // @[:@32393.4]
  input  [63:0] io_ins_222, // @[:@32393.4]
  input  [63:0] io_ins_223, // @[:@32393.4]
  input  [63:0] io_ins_224, // @[:@32393.4]
  input  [63:0] io_ins_225, // @[:@32393.4]
  input  [63:0] io_ins_226, // @[:@32393.4]
  input  [63:0] io_ins_227, // @[:@32393.4]
  input  [63:0] io_ins_228, // @[:@32393.4]
  input  [63:0] io_ins_229, // @[:@32393.4]
  input  [63:0] io_ins_230, // @[:@32393.4]
  input  [63:0] io_ins_231, // @[:@32393.4]
  input  [63:0] io_ins_232, // @[:@32393.4]
  input  [63:0] io_ins_233, // @[:@32393.4]
  input  [63:0] io_ins_234, // @[:@32393.4]
  input  [63:0] io_ins_235, // @[:@32393.4]
  input  [63:0] io_ins_236, // @[:@32393.4]
  input  [63:0] io_ins_237, // @[:@32393.4]
  input  [63:0] io_ins_238, // @[:@32393.4]
  input  [63:0] io_ins_239, // @[:@32393.4]
  input  [63:0] io_ins_240, // @[:@32393.4]
  input  [63:0] io_ins_241, // @[:@32393.4]
  input  [63:0] io_ins_242, // @[:@32393.4]
  input  [63:0] io_ins_243, // @[:@32393.4]
  input  [63:0] io_ins_244, // @[:@32393.4]
  input  [63:0] io_ins_245, // @[:@32393.4]
  input  [63:0] io_ins_246, // @[:@32393.4]
  input  [63:0] io_ins_247, // @[:@32393.4]
  input  [63:0] io_ins_248, // @[:@32393.4]
  input  [63:0] io_ins_249, // @[:@32393.4]
  input  [63:0] io_ins_250, // @[:@32393.4]
  input  [63:0] io_ins_251, // @[:@32393.4]
  input  [63:0] io_ins_252, // @[:@32393.4]
  input  [63:0] io_ins_253, // @[:@32393.4]
  input  [63:0] io_ins_254, // @[:@32393.4]
  input  [63:0] io_ins_255, // @[:@32393.4]
  input  [63:0] io_ins_256, // @[:@32393.4]
  input  [63:0] io_ins_257, // @[:@32393.4]
  input  [63:0] io_ins_258, // @[:@32393.4]
  input  [63:0] io_ins_259, // @[:@32393.4]
  input  [63:0] io_ins_260, // @[:@32393.4]
  input  [63:0] io_ins_261, // @[:@32393.4]
  input  [63:0] io_ins_262, // @[:@32393.4]
  input  [63:0] io_ins_263, // @[:@32393.4]
  input  [63:0] io_ins_264, // @[:@32393.4]
  input  [63:0] io_ins_265, // @[:@32393.4]
  input  [63:0] io_ins_266, // @[:@32393.4]
  input  [63:0] io_ins_267, // @[:@32393.4]
  input  [63:0] io_ins_268, // @[:@32393.4]
  input  [63:0] io_ins_269, // @[:@32393.4]
  input  [63:0] io_ins_270, // @[:@32393.4]
  input  [63:0] io_ins_271, // @[:@32393.4]
  input  [63:0] io_ins_272, // @[:@32393.4]
  input  [63:0] io_ins_273, // @[:@32393.4]
  input  [63:0] io_ins_274, // @[:@32393.4]
  input  [63:0] io_ins_275, // @[:@32393.4]
  input  [63:0] io_ins_276, // @[:@32393.4]
  input  [63:0] io_ins_277, // @[:@32393.4]
  input  [63:0] io_ins_278, // @[:@32393.4]
  input  [63:0] io_ins_279, // @[:@32393.4]
  input  [63:0] io_ins_280, // @[:@32393.4]
  input  [63:0] io_ins_281, // @[:@32393.4]
  input  [63:0] io_ins_282, // @[:@32393.4]
  input  [63:0] io_ins_283, // @[:@32393.4]
  input  [63:0] io_ins_284, // @[:@32393.4]
  input  [63:0] io_ins_285, // @[:@32393.4]
  input  [63:0] io_ins_286, // @[:@32393.4]
  input  [63:0] io_ins_287, // @[:@32393.4]
  input  [63:0] io_ins_288, // @[:@32393.4]
  input  [63:0] io_ins_289, // @[:@32393.4]
  input  [63:0] io_ins_290, // @[:@32393.4]
  input  [63:0] io_ins_291, // @[:@32393.4]
  input  [63:0] io_ins_292, // @[:@32393.4]
  input  [63:0] io_ins_293, // @[:@32393.4]
  input  [63:0] io_ins_294, // @[:@32393.4]
  input  [63:0] io_ins_295, // @[:@32393.4]
  input  [63:0] io_ins_296, // @[:@32393.4]
  input  [63:0] io_ins_297, // @[:@32393.4]
  input  [63:0] io_ins_298, // @[:@32393.4]
  input  [63:0] io_ins_299, // @[:@32393.4]
  input  [63:0] io_ins_300, // @[:@32393.4]
  input  [63:0] io_ins_301, // @[:@32393.4]
  input  [63:0] io_ins_302, // @[:@32393.4]
  input  [63:0] io_ins_303, // @[:@32393.4]
  input  [63:0] io_ins_304, // @[:@32393.4]
  input  [63:0] io_ins_305, // @[:@32393.4]
  input  [63:0] io_ins_306, // @[:@32393.4]
  input  [63:0] io_ins_307, // @[:@32393.4]
  input  [63:0] io_ins_308, // @[:@32393.4]
  input  [63:0] io_ins_309, // @[:@32393.4]
  input  [63:0] io_ins_310, // @[:@32393.4]
  input  [63:0] io_ins_311, // @[:@32393.4]
  input  [63:0] io_ins_312, // @[:@32393.4]
  input  [63:0] io_ins_313, // @[:@32393.4]
  input  [63:0] io_ins_314, // @[:@32393.4]
  input  [63:0] io_ins_315, // @[:@32393.4]
  input  [63:0] io_ins_316, // @[:@32393.4]
  input  [63:0] io_ins_317, // @[:@32393.4]
  input  [63:0] io_ins_318, // @[:@32393.4]
  input  [63:0] io_ins_319, // @[:@32393.4]
  input  [63:0] io_ins_320, // @[:@32393.4]
  input  [63:0] io_ins_321, // @[:@32393.4]
  input  [63:0] io_ins_322, // @[:@32393.4]
  input  [63:0] io_ins_323, // @[:@32393.4]
  input  [63:0] io_ins_324, // @[:@32393.4]
  input  [63:0] io_ins_325, // @[:@32393.4]
  input  [63:0] io_ins_326, // @[:@32393.4]
  input  [63:0] io_ins_327, // @[:@32393.4]
  input  [63:0] io_ins_328, // @[:@32393.4]
  input  [63:0] io_ins_329, // @[:@32393.4]
  input  [63:0] io_ins_330, // @[:@32393.4]
  input  [63:0] io_ins_331, // @[:@32393.4]
  input  [63:0] io_ins_332, // @[:@32393.4]
  input  [63:0] io_ins_333, // @[:@32393.4]
  input  [63:0] io_ins_334, // @[:@32393.4]
  input  [63:0] io_ins_335, // @[:@32393.4]
  input  [63:0] io_ins_336, // @[:@32393.4]
  input  [63:0] io_ins_337, // @[:@32393.4]
  input  [63:0] io_ins_338, // @[:@32393.4]
  input  [63:0] io_ins_339, // @[:@32393.4]
  input  [63:0] io_ins_340, // @[:@32393.4]
  input  [63:0] io_ins_341, // @[:@32393.4]
  input  [63:0] io_ins_342, // @[:@32393.4]
  input  [63:0] io_ins_343, // @[:@32393.4]
  input  [63:0] io_ins_344, // @[:@32393.4]
  input  [63:0] io_ins_345, // @[:@32393.4]
  input  [63:0] io_ins_346, // @[:@32393.4]
  input  [63:0] io_ins_347, // @[:@32393.4]
  input  [63:0] io_ins_348, // @[:@32393.4]
  input  [63:0] io_ins_349, // @[:@32393.4]
  input  [63:0] io_ins_350, // @[:@32393.4]
  input  [63:0] io_ins_351, // @[:@32393.4]
  input  [63:0] io_ins_352, // @[:@32393.4]
  input  [63:0] io_ins_353, // @[:@32393.4]
  input  [63:0] io_ins_354, // @[:@32393.4]
  input  [63:0] io_ins_355, // @[:@32393.4]
  input  [63:0] io_ins_356, // @[:@32393.4]
  input  [63:0] io_ins_357, // @[:@32393.4]
  input  [63:0] io_ins_358, // @[:@32393.4]
  input  [63:0] io_ins_359, // @[:@32393.4]
  input  [63:0] io_ins_360, // @[:@32393.4]
  input  [63:0] io_ins_361, // @[:@32393.4]
  input  [63:0] io_ins_362, // @[:@32393.4]
  input  [63:0] io_ins_363, // @[:@32393.4]
  input  [63:0] io_ins_364, // @[:@32393.4]
  input  [63:0] io_ins_365, // @[:@32393.4]
  input  [63:0] io_ins_366, // @[:@32393.4]
  input  [63:0] io_ins_367, // @[:@32393.4]
  input  [63:0] io_ins_368, // @[:@32393.4]
  input  [63:0] io_ins_369, // @[:@32393.4]
  input  [63:0] io_ins_370, // @[:@32393.4]
  input  [63:0] io_ins_371, // @[:@32393.4]
  input  [63:0] io_ins_372, // @[:@32393.4]
  input  [63:0] io_ins_373, // @[:@32393.4]
  input  [63:0] io_ins_374, // @[:@32393.4]
  input  [63:0] io_ins_375, // @[:@32393.4]
  input  [63:0] io_ins_376, // @[:@32393.4]
  input  [63:0] io_ins_377, // @[:@32393.4]
  input  [63:0] io_ins_378, // @[:@32393.4]
  input  [63:0] io_ins_379, // @[:@32393.4]
  input  [63:0] io_ins_380, // @[:@32393.4]
  input  [63:0] io_ins_381, // @[:@32393.4]
  input  [63:0] io_ins_382, // @[:@32393.4]
  input  [63:0] io_ins_383, // @[:@32393.4]
  input  [63:0] io_ins_384, // @[:@32393.4]
  input  [63:0] io_ins_385, // @[:@32393.4]
  input  [63:0] io_ins_386, // @[:@32393.4]
  input  [63:0] io_ins_387, // @[:@32393.4]
  input  [63:0] io_ins_388, // @[:@32393.4]
  input  [63:0] io_ins_389, // @[:@32393.4]
  input  [63:0] io_ins_390, // @[:@32393.4]
  input  [63:0] io_ins_391, // @[:@32393.4]
  input  [63:0] io_ins_392, // @[:@32393.4]
  input  [63:0] io_ins_393, // @[:@32393.4]
  input  [63:0] io_ins_394, // @[:@32393.4]
  input  [63:0] io_ins_395, // @[:@32393.4]
  input  [63:0] io_ins_396, // @[:@32393.4]
  input  [63:0] io_ins_397, // @[:@32393.4]
  input  [63:0] io_ins_398, // @[:@32393.4]
  input  [63:0] io_ins_399, // @[:@32393.4]
  input  [63:0] io_ins_400, // @[:@32393.4]
  input  [63:0] io_ins_401, // @[:@32393.4]
  input  [63:0] io_ins_402, // @[:@32393.4]
  input  [63:0] io_ins_403, // @[:@32393.4]
  input  [63:0] io_ins_404, // @[:@32393.4]
  input  [63:0] io_ins_405, // @[:@32393.4]
  input  [63:0] io_ins_406, // @[:@32393.4]
  input  [63:0] io_ins_407, // @[:@32393.4]
  input  [63:0] io_ins_408, // @[:@32393.4]
  input  [63:0] io_ins_409, // @[:@32393.4]
  input  [63:0] io_ins_410, // @[:@32393.4]
  input  [63:0] io_ins_411, // @[:@32393.4]
  input  [63:0] io_ins_412, // @[:@32393.4]
  input  [63:0] io_ins_413, // @[:@32393.4]
  input  [63:0] io_ins_414, // @[:@32393.4]
  input  [63:0] io_ins_415, // @[:@32393.4]
  input  [63:0] io_ins_416, // @[:@32393.4]
  input  [63:0] io_ins_417, // @[:@32393.4]
  input  [63:0] io_ins_418, // @[:@32393.4]
  input  [63:0] io_ins_419, // @[:@32393.4]
  input  [63:0] io_ins_420, // @[:@32393.4]
  input  [63:0] io_ins_421, // @[:@32393.4]
  input  [63:0] io_ins_422, // @[:@32393.4]
  input  [63:0] io_ins_423, // @[:@32393.4]
  input  [63:0] io_ins_424, // @[:@32393.4]
  input  [63:0] io_ins_425, // @[:@32393.4]
  input  [63:0] io_ins_426, // @[:@32393.4]
  input  [63:0] io_ins_427, // @[:@32393.4]
  input  [63:0] io_ins_428, // @[:@32393.4]
  input  [63:0] io_ins_429, // @[:@32393.4]
  input  [63:0] io_ins_430, // @[:@32393.4]
  input  [63:0] io_ins_431, // @[:@32393.4]
  input  [63:0] io_ins_432, // @[:@32393.4]
  input  [63:0] io_ins_433, // @[:@32393.4]
  input  [63:0] io_ins_434, // @[:@32393.4]
  input  [63:0] io_ins_435, // @[:@32393.4]
  input  [63:0] io_ins_436, // @[:@32393.4]
  input  [63:0] io_ins_437, // @[:@32393.4]
  input  [63:0] io_ins_438, // @[:@32393.4]
  input  [63:0] io_ins_439, // @[:@32393.4]
  input  [63:0] io_ins_440, // @[:@32393.4]
  input  [63:0] io_ins_441, // @[:@32393.4]
  input  [63:0] io_ins_442, // @[:@32393.4]
  input  [63:0] io_ins_443, // @[:@32393.4]
  input  [63:0] io_ins_444, // @[:@32393.4]
  input  [63:0] io_ins_445, // @[:@32393.4]
  input  [63:0] io_ins_446, // @[:@32393.4]
  input  [63:0] io_ins_447, // @[:@32393.4]
  input  [63:0] io_ins_448, // @[:@32393.4]
  input  [63:0] io_ins_449, // @[:@32393.4]
  input  [63:0] io_ins_450, // @[:@32393.4]
  input  [63:0] io_ins_451, // @[:@32393.4]
  input  [63:0] io_ins_452, // @[:@32393.4]
  input  [63:0] io_ins_453, // @[:@32393.4]
  input  [63:0] io_ins_454, // @[:@32393.4]
  input  [63:0] io_ins_455, // @[:@32393.4]
  input  [63:0] io_ins_456, // @[:@32393.4]
  input  [63:0] io_ins_457, // @[:@32393.4]
  input  [63:0] io_ins_458, // @[:@32393.4]
  input  [63:0] io_ins_459, // @[:@32393.4]
  input  [63:0] io_ins_460, // @[:@32393.4]
  input  [63:0] io_ins_461, // @[:@32393.4]
  input  [63:0] io_ins_462, // @[:@32393.4]
  input  [63:0] io_ins_463, // @[:@32393.4]
  input  [63:0] io_ins_464, // @[:@32393.4]
  input  [63:0] io_ins_465, // @[:@32393.4]
  input  [63:0] io_ins_466, // @[:@32393.4]
  input  [63:0] io_ins_467, // @[:@32393.4]
  input  [63:0] io_ins_468, // @[:@32393.4]
  input  [63:0] io_ins_469, // @[:@32393.4]
  input  [63:0] io_ins_470, // @[:@32393.4]
  input  [63:0] io_ins_471, // @[:@32393.4]
  input  [63:0] io_ins_472, // @[:@32393.4]
  input  [63:0] io_ins_473, // @[:@32393.4]
  input  [63:0] io_ins_474, // @[:@32393.4]
  input  [63:0] io_ins_475, // @[:@32393.4]
  input  [63:0] io_ins_476, // @[:@32393.4]
  input  [63:0] io_ins_477, // @[:@32393.4]
  input  [63:0] io_ins_478, // @[:@32393.4]
  input  [63:0] io_ins_479, // @[:@32393.4]
  input  [63:0] io_ins_480, // @[:@32393.4]
  input  [63:0] io_ins_481, // @[:@32393.4]
  input  [63:0] io_ins_482, // @[:@32393.4]
  input  [63:0] io_ins_483, // @[:@32393.4]
  input  [63:0] io_ins_484, // @[:@32393.4]
  input  [63:0] io_ins_485, // @[:@32393.4]
  input  [63:0] io_ins_486, // @[:@32393.4]
  input  [63:0] io_ins_487, // @[:@32393.4]
  input  [63:0] io_ins_488, // @[:@32393.4]
  input  [63:0] io_ins_489, // @[:@32393.4]
  input  [63:0] io_ins_490, // @[:@32393.4]
  input  [63:0] io_ins_491, // @[:@32393.4]
  input  [63:0] io_ins_492, // @[:@32393.4]
  input  [63:0] io_ins_493, // @[:@32393.4]
  input  [63:0] io_ins_494, // @[:@32393.4]
  input  [63:0] io_ins_495, // @[:@32393.4]
  input  [63:0] io_ins_496, // @[:@32393.4]
  input  [63:0] io_ins_497, // @[:@32393.4]
  input  [63:0] io_ins_498, // @[:@32393.4]
  input  [63:0] io_ins_499, // @[:@32393.4]
  input  [63:0] io_ins_500, // @[:@32393.4]
  input  [63:0] io_ins_501, // @[:@32393.4]
  input  [63:0] io_ins_502, // @[:@32393.4]
  input  [8:0]  io_sel, // @[:@32393.4]
  output [63:0] io_out // @[:@32393.4]
);
  wire [63:0] _GEN_1; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_2; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_3; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_4; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_5; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_6; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_7; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_8; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_9; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_10; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_11; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_12; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_13; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_14; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_15; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_16; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_17; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_18; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_19; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_20; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_21; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_22; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_23; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_24; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_25; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_26; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_27; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_28; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_29; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_30; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_31; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_32; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_33; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_34; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_35; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_36; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_37; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_38; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_39; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_40; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_41; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_42; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_43; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_44; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_45; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_46; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_47; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_48; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_49; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_50; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_51; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_52; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_53; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_54; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_55; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_56; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_57; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_58; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_59; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_60; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_61; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_62; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_63; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_64; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_65; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_66; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_67; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_68; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_69; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_70; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_71; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_72; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_73; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_74; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_75; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_76; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_77; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_78; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_79; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_80; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_81; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_82; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_83; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_84; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_85; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_86; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_87; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_88; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_89; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_90; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_91; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_92; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_93; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_94; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_95; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_96; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_97; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_98; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_99; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_100; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_101; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_102; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_103; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_104; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_105; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_106; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_107; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_108; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_109; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_110; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_111; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_112; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_113; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_114; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_115; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_116; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_117; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_118; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_119; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_120; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_121; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_122; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_123; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_124; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_125; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_126; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_127; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_128; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_129; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_130; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_131; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_132; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_133; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_134; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_135; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_136; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_137; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_138; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_139; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_140; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_141; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_142; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_143; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_144; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_145; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_146; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_147; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_148; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_149; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_150; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_151; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_152; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_153; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_154; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_155; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_156; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_157; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_158; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_159; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_160; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_161; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_162; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_163; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_164; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_165; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_166; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_167; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_168; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_169; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_170; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_171; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_172; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_173; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_174; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_175; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_176; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_177; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_178; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_179; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_180; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_181; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_182; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_183; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_184; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_185; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_186; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_187; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_188; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_189; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_190; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_191; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_192; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_193; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_194; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_195; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_196; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_197; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_198; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_199; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_200; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_201; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_202; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_203; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_204; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_205; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_206; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_207; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_208; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_209; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_210; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_211; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_212; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_213; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_214; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_215; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_216; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_217; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_218; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_219; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_220; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_221; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_222; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_223; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_224; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_225; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_226; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_227; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_228; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_229; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_230; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_231; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_232; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_233; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_234; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_235; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_236; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_237; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_238; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_239; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_240; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_241; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_242; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_243; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_244; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_245; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_246; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_247; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_248; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_249; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_250; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_251; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_252; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_253; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_254; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_255; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_256; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_257; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_258; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_259; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_260; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_261; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_262; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_263; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_264; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_265; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_266; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_267; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_268; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_269; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_270; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_271; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_272; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_273; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_274; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_275; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_276; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_277; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_278; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_279; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_280; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_281; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_282; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_283; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_284; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_285; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_286; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_287; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_288; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_289; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_290; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_291; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_292; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_293; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_294; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_295; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_296; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_297; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_298; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_299; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_300; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_301; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_302; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_303; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_304; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_305; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_306; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_307; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_308; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_309; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_310; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_311; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_312; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_313; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_314; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_315; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_316; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_317; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_318; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_319; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_320; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_321; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_322; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_323; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_324; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_325; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_326; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_327; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_328; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_329; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_330; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_331; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_332; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_333; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_334; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_335; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_336; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_337; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_338; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_339; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_340; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_341; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_342; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_343; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_344; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_345; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_346; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_347; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_348; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_349; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_350; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_351; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_352; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_353; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_354; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_355; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_356; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_357; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_358; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_359; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_360; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_361; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_362; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_363; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_364; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_365; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_366; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_367; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_368; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_369; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_370; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_371; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_372; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_373; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_374; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_375; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_376; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_377; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_378; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_379; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_380; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_381; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_382; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_383; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_384; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_385; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_386; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_387; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_388; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_389; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_390; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_391; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_392; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_393; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_394; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_395; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_396; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_397; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_398; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_399; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_400; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_401; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_402; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_403; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_404; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_405; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_406; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_407; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_408; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_409; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_410; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_411; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_412; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_413; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_414; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_415; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_416; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_417; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_418; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_419; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_420; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_421; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_422; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_423; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_424; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_425; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_426; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_427; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_428; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_429; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_430; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_431; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_432; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_433; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_434; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_435; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_436; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_437; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_438; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_439; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_440; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_441; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_442; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_443; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_444; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_445; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_446; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_447; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_448; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_449; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_450; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_451; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_452; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_453; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_454; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_455; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_456; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_457; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_458; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_459; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_460; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_461; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_462; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_463; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_464; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_465; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_466; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_467; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_468; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_469; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_470; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_471; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_472; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_473; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_474; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_475; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_476; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_477; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_478; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_479; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_480; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_481; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_482; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_483; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_484; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_485; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_486; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_487; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_488; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_489; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_490; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_491; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_492; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_493; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_494; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_495; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_496; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_497; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_498; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_499; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_500; // @[MuxN.scala 16:10:@32395.4]
  wire [63:0] _GEN_501; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_1 = 9'h1 == io_sel ? io_ins_1 : io_ins_0; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_2 = 9'h2 == io_sel ? io_ins_2 : _GEN_1; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_3 = 9'h3 == io_sel ? io_ins_3 : _GEN_2; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_4 = 9'h4 == io_sel ? io_ins_4 : _GEN_3; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_5 = 9'h5 == io_sel ? io_ins_5 : _GEN_4; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_6 = 9'h6 == io_sel ? io_ins_6 : _GEN_5; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_7 = 9'h7 == io_sel ? io_ins_7 : _GEN_6; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_8 = 9'h8 == io_sel ? io_ins_8 : _GEN_7; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_9 = 9'h9 == io_sel ? io_ins_9 : _GEN_8; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_10 = 9'ha == io_sel ? io_ins_10 : _GEN_9; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_11 = 9'hb == io_sel ? io_ins_11 : _GEN_10; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_12 = 9'hc == io_sel ? io_ins_12 : _GEN_11; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_13 = 9'hd == io_sel ? io_ins_13 : _GEN_12; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_14 = 9'he == io_sel ? io_ins_14 : _GEN_13; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_15 = 9'hf == io_sel ? io_ins_15 : _GEN_14; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_16 = 9'h10 == io_sel ? io_ins_16 : _GEN_15; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_17 = 9'h11 == io_sel ? io_ins_17 : _GEN_16; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_18 = 9'h12 == io_sel ? io_ins_18 : _GEN_17; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_19 = 9'h13 == io_sel ? io_ins_19 : _GEN_18; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_20 = 9'h14 == io_sel ? io_ins_20 : _GEN_19; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_21 = 9'h15 == io_sel ? io_ins_21 : _GEN_20; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_22 = 9'h16 == io_sel ? io_ins_22 : _GEN_21; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_23 = 9'h17 == io_sel ? io_ins_23 : _GEN_22; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_24 = 9'h18 == io_sel ? io_ins_24 : _GEN_23; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_25 = 9'h19 == io_sel ? io_ins_25 : _GEN_24; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_26 = 9'h1a == io_sel ? io_ins_26 : _GEN_25; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_27 = 9'h1b == io_sel ? io_ins_27 : _GEN_26; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_28 = 9'h1c == io_sel ? io_ins_28 : _GEN_27; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_29 = 9'h1d == io_sel ? io_ins_29 : _GEN_28; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_30 = 9'h1e == io_sel ? io_ins_30 : _GEN_29; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_31 = 9'h1f == io_sel ? io_ins_31 : _GEN_30; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_32 = 9'h20 == io_sel ? io_ins_32 : _GEN_31; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_33 = 9'h21 == io_sel ? io_ins_33 : _GEN_32; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_34 = 9'h22 == io_sel ? io_ins_34 : _GEN_33; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_35 = 9'h23 == io_sel ? io_ins_35 : _GEN_34; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_36 = 9'h24 == io_sel ? io_ins_36 : _GEN_35; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_37 = 9'h25 == io_sel ? io_ins_37 : _GEN_36; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_38 = 9'h26 == io_sel ? io_ins_38 : _GEN_37; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_39 = 9'h27 == io_sel ? io_ins_39 : _GEN_38; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_40 = 9'h28 == io_sel ? io_ins_40 : _GEN_39; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_41 = 9'h29 == io_sel ? io_ins_41 : _GEN_40; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_42 = 9'h2a == io_sel ? io_ins_42 : _GEN_41; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_43 = 9'h2b == io_sel ? io_ins_43 : _GEN_42; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_44 = 9'h2c == io_sel ? io_ins_44 : _GEN_43; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_45 = 9'h2d == io_sel ? io_ins_45 : _GEN_44; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_46 = 9'h2e == io_sel ? io_ins_46 : _GEN_45; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_47 = 9'h2f == io_sel ? io_ins_47 : _GEN_46; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_48 = 9'h30 == io_sel ? io_ins_48 : _GEN_47; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_49 = 9'h31 == io_sel ? io_ins_49 : _GEN_48; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_50 = 9'h32 == io_sel ? io_ins_50 : _GEN_49; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_51 = 9'h33 == io_sel ? io_ins_51 : _GEN_50; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_52 = 9'h34 == io_sel ? io_ins_52 : _GEN_51; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_53 = 9'h35 == io_sel ? io_ins_53 : _GEN_52; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_54 = 9'h36 == io_sel ? io_ins_54 : _GEN_53; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_55 = 9'h37 == io_sel ? io_ins_55 : _GEN_54; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_56 = 9'h38 == io_sel ? io_ins_56 : _GEN_55; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_57 = 9'h39 == io_sel ? io_ins_57 : _GEN_56; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_58 = 9'h3a == io_sel ? io_ins_58 : _GEN_57; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_59 = 9'h3b == io_sel ? io_ins_59 : _GEN_58; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_60 = 9'h3c == io_sel ? io_ins_60 : _GEN_59; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_61 = 9'h3d == io_sel ? io_ins_61 : _GEN_60; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_62 = 9'h3e == io_sel ? io_ins_62 : _GEN_61; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_63 = 9'h3f == io_sel ? io_ins_63 : _GEN_62; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_64 = 9'h40 == io_sel ? io_ins_64 : _GEN_63; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_65 = 9'h41 == io_sel ? io_ins_65 : _GEN_64; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_66 = 9'h42 == io_sel ? io_ins_66 : _GEN_65; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_67 = 9'h43 == io_sel ? io_ins_67 : _GEN_66; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_68 = 9'h44 == io_sel ? io_ins_68 : _GEN_67; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_69 = 9'h45 == io_sel ? io_ins_69 : _GEN_68; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_70 = 9'h46 == io_sel ? io_ins_70 : _GEN_69; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_71 = 9'h47 == io_sel ? io_ins_71 : _GEN_70; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_72 = 9'h48 == io_sel ? io_ins_72 : _GEN_71; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_73 = 9'h49 == io_sel ? io_ins_73 : _GEN_72; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_74 = 9'h4a == io_sel ? io_ins_74 : _GEN_73; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_75 = 9'h4b == io_sel ? io_ins_75 : _GEN_74; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_76 = 9'h4c == io_sel ? io_ins_76 : _GEN_75; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_77 = 9'h4d == io_sel ? io_ins_77 : _GEN_76; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_78 = 9'h4e == io_sel ? io_ins_78 : _GEN_77; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_79 = 9'h4f == io_sel ? io_ins_79 : _GEN_78; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_80 = 9'h50 == io_sel ? io_ins_80 : _GEN_79; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_81 = 9'h51 == io_sel ? io_ins_81 : _GEN_80; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_82 = 9'h52 == io_sel ? io_ins_82 : _GEN_81; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_83 = 9'h53 == io_sel ? io_ins_83 : _GEN_82; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_84 = 9'h54 == io_sel ? io_ins_84 : _GEN_83; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_85 = 9'h55 == io_sel ? io_ins_85 : _GEN_84; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_86 = 9'h56 == io_sel ? io_ins_86 : _GEN_85; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_87 = 9'h57 == io_sel ? io_ins_87 : _GEN_86; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_88 = 9'h58 == io_sel ? io_ins_88 : _GEN_87; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_89 = 9'h59 == io_sel ? io_ins_89 : _GEN_88; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_90 = 9'h5a == io_sel ? io_ins_90 : _GEN_89; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_91 = 9'h5b == io_sel ? io_ins_91 : _GEN_90; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_92 = 9'h5c == io_sel ? io_ins_92 : _GEN_91; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_93 = 9'h5d == io_sel ? io_ins_93 : _GEN_92; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_94 = 9'h5e == io_sel ? io_ins_94 : _GEN_93; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_95 = 9'h5f == io_sel ? io_ins_95 : _GEN_94; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_96 = 9'h60 == io_sel ? io_ins_96 : _GEN_95; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_97 = 9'h61 == io_sel ? io_ins_97 : _GEN_96; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_98 = 9'h62 == io_sel ? io_ins_98 : _GEN_97; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_99 = 9'h63 == io_sel ? io_ins_99 : _GEN_98; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_100 = 9'h64 == io_sel ? io_ins_100 : _GEN_99; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_101 = 9'h65 == io_sel ? io_ins_101 : _GEN_100; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_102 = 9'h66 == io_sel ? io_ins_102 : _GEN_101; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_103 = 9'h67 == io_sel ? io_ins_103 : _GEN_102; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_104 = 9'h68 == io_sel ? io_ins_104 : _GEN_103; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_105 = 9'h69 == io_sel ? io_ins_105 : _GEN_104; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_106 = 9'h6a == io_sel ? io_ins_106 : _GEN_105; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_107 = 9'h6b == io_sel ? io_ins_107 : _GEN_106; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_108 = 9'h6c == io_sel ? io_ins_108 : _GEN_107; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_109 = 9'h6d == io_sel ? io_ins_109 : _GEN_108; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_110 = 9'h6e == io_sel ? io_ins_110 : _GEN_109; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_111 = 9'h6f == io_sel ? io_ins_111 : _GEN_110; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_112 = 9'h70 == io_sel ? io_ins_112 : _GEN_111; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_113 = 9'h71 == io_sel ? io_ins_113 : _GEN_112; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_114 = 9'h72 == io_sel ? io_ins_114 : _GEN_113; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_115 = 9'h73 == io_sel ? io_ins_115 : _GEN_114; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_116 = 9'h74 == io_sel ? io_ins_116 : _GEN_115; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_117 = 9'h75 == io_sel ? io_ins_117 : _GEN_116; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_118 = 9'h76 == io_sel ? io_ins_118 : _GEN_117; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_119 = 9'h77 == io_sel ? io_ins_119 : _GEN_118; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_120 = 9'h78 == io_sel ? io_ins_120 : _GEN_119; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_121 = 9'h79 == io_sel ? io_ins_121 : _GEN_120; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_122 = 9'h7a == io_sel ? io_ins_122 : _GEN_121; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_123 = 9'h7b == io_sel ? io_ins_123 : _GEN_122; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_124 = 9'h7c == io_sel ? io_ins_124 : _GEN_123; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_125 = 9'h7d == io_sel ? io_ins_125 : _GEN_124; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_126 = 9'h7e == io_sel ? io_ins_126 : _GEN_125; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_127 = 9'h7f == io_sel ? io_ins_127 : _GEN_126; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_128 = 9'h80 == io_sel ? io_ins_128 : _GEN_127; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_129 = 9'h81 == io_sel ? io_ins_129 : _GEN_128; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_130 = 9'h82 == io_sel ? io_ins_130 : _GEN_129; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_131 = 9'h83 == io_sel ? io_ins_131 : _GEN_130; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_132 = 9'h84 == io_sel ? io_ins_132 : _GEN_131; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_133 = 9'h85 == io_sel ? io_ins_133 : _GEN_132; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_134 = 9'h86 == io_sel ? io_ins_134 : _GEN_133; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_135 = 9'h87 == io_sel ? io_ins_135 : _GEN_134; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_136 = 9'h88 == io_sel ? io_ins_136 : _GEN_135; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_137 = 9'h89 == io_sel ? io_ins_137 : _GEN_136; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_138 = 9'h8a == io_sel ? io_ins_138 : _GEN_137; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_139 = 9'h8b == io_sel ? io_ins_139 : _GEN_138; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_140 = 9'h8c == io_sel ? io_ins_140 : _GEN_139; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_141 = 9'h8d == io_sel ? io_ins_141 : _GEN_140; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_142 = 9'h8e == io_sel ? io_ins_142 : _GEN_141; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_143 = 9'h8f == io_sel ? io_ins_143 : _GEN_142; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_144 = 9'h90 == io_sel ? io_ins_144 : _GEN_143; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_145 = 9'h91 == io_sel ? io_ins_145 : _GEN_144; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_146 = 9'h92 == io_sel ? io_ins_146 : _GEN_145; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_147 = 9'h93 == io_sel ? io_ins_147 : _GEN_146; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_148 = 9'h94 == io_sel ? io_ins_148 : _GEN_147; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_149 = 9'h95 == io_sel ? io_ins_149 : _GEN_148; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_150 = 9'h96 == io_sel ? io_ins_150 : _GEN_149; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_151 = 9'h97 == io_sel ? io_ins_151 : _GEN_150; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_152 = 9'h98 == io_sel ? io_ins_152 : _GEN_151; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_153 = 9'h99 == io_sel ? io_ins_153 : _GEN_152; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_154 = 9'h9a == io_sel ? io_ins_154 : _GEN_153; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_155 = 9'h9b == io_sel ? io_ins_155 : _GEN_154; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_156 = 9'h9c == io_sel ? io_ins_156 : _GEN_155; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_157 = 9'h9d == io_sel ? io_ins_157 : _GEN_156; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_158 = 9'h9e == io_sel ? io_ins_158 : _GEN_157; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_159 = 9'h9f == io_sel ? io_ins_159 : _GEN_158; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_160 = 9'ha0 == io_sel ? io_ins_160 : _GEN_159; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_161 = 9'ha1 == io_sel ? io_ins_161 : _GEN_160; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_162 = 9'ha2 == io_sel ? io_ins_162 : _GEN_161; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_163 = 9'ha3 == io_sel ? io_ins_163 : _GEN_162; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_164 = 9'ha4 == io_sel ? io_ins_164 : _GEN_163; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_165 = 9'ha5 == io_sel ? io_ins_165 : _GEN_164; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_166 = 9'ha6 == io_sel ? io_ins_166 : _GEN_165; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_167 = 9'ha7 == io_sel ? io_ins_167 : _GEN_166; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_168 = 9'ha8 == io_sel ? io_ins_168 : _GEN_167; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_169 = 9'ha9 == io_sel ? io_ins_169 : _GEN_168; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_170 = 9'haa == io_sel ? io_ins_170 : _GEN_169; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_171 = 9'hab == io_sel ? io_ins_171 : _GEN_170; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_172 = 9'hac == io_sel ? io_ins_172 : _GEN_171; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_173 = 9'had == io_sel ? io_ins_173 : _GEN_172; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_174 = 9'hae == io_sel ? io_ins_174 : _GEN_173; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_175 = 9'haf == io_sel ? io_ins_175 : _GEN_174; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_176 = 9'hb0 == io_sel ? io_ins_176 : _GEN_175; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_177 = 9'hb1 == io_sel ? io_ins_177 : _GEN_176; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_178 = 9'hb2 == io_sel ? io_ins_178 : _GEN_177; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_179 = 9'hb3 == io_sel ? io_ins_179 : _GEN_178; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_180 = 9'hb4 == io_sel ? io_ins_180 : _GEN_179; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_181 = 9'hb5 == io_sel ? io_ins_181 : _GEN_180; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_182 = 9'hb6 == io_sel ? io_ins_182 : _GEN_181; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_183 = 9'hb7 == io_sel ? io_ins_183 : _GEN_182; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_184 = 9'hb8 == io_sel ? io_ins_184 : _GEN_183; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_185 = 9'hb9 == io_sel ? io_ins_185 : _GEN_184; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_186 = 9'hba == io_sel ? io_ins_186 : _GEN_185; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_187 = 9'hbb == io_sel ? io_ins_187 : _GEN_186; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_188 = 9'hbc == io_sel ? io_ins_188 : _GEN_187; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_189 = 9'hbd == io_sel ? io_ins_189 : _GEN_188; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_190 = 9'hbe == io_sel ? io_ins_190 : _GEN_189; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_191 = 9'hbf == io_sel ? io_ins_191 : _GEN_190; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_192 = 9'hc0 == io_sel ? io_ins_192 : _GEN_191; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_193 = 9'hc1 == io_sel ? io_ins_193 : _GEN_192; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_194 = 9'hc2 == io_sel ? io_ins_194 : _GEN_193; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_195 = 9'hc3 == io_sel ? io_ins_195 : _GEN_194; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_196 = 9'hc4 == io_sel ? io_ins_196 : _GEN_195; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_197 = 9'hc5 == io_sel ? io_ins_197 : _GEN_196; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_198 = 9'hc6 == io_sel ? io_ins_198 : _GEN_197; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_199 = 9'hc7 == io_sel ? io_ins_199 : _GEN_198; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_200 = 9'hc8 == io_sel ? io_ins_200 : _GEN_199; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_201 = 9'hc9 == io_sel ? io_ins_201 : _GEN_200; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_202 = 9'hca == io_sel ? io_ins_202 : _GEN_201; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_203 = 9'hcb == io_sel ? io_ins_203 : _GEN_202; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_204 = 9'hcc == io_sel ? io_ins_204 : _GEN_203; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_205 = 9'hcd == io_sel ? io_ins_205 : _GEN_204; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_206 = 9'hce == io_sel ? io_ins_206 : _GEN_205; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_207 = 9'hcf == io_sel ? io_ins_207 : _GEN_206; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_208 = 9'hd0 == io_sel ? io_ins_208 : _GEN_207; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_209 = 9'hd1 == io_sel ? io_ins_209 : _GEN_208; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_210 = 9'hd2 == io_sel ? io_ins_210 : _GEN_209; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_211 = 9'hd3 == io_sel ? io_ins_211 : _GEN_210; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_212 = 9'hd4 == io_sel ? io_ins_212 : _GEN_211; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_213 = 9'hd5 == io_sel ? io_ins_213 : _GEN_212; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_214 = 9'hd6 == io_sel ? io_ins_214 : _GEN_213; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_215 = 9'hd7 == io_sel ? io_ins_215 : _GEN_214; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_216 = 9'hd8 == io_sel ? io_ins_216 : _GEN_215; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_217 = 9'hd9 == io_sel ? io_ins_217 : _GEN_216; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_218 = 9'hda == io_sel ? io_ins_218 : _GEN_217; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_219 = 9'hdb == io_sel ? io_ins_219 : _GEN_218; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_220 = 9'hdc == io_sel ? io_ins_220 : _GEN_219; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_221 = 9'hdd == io_sel ? io_ins_221 : _GEN_220; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_222 = 9'hde == io_sel ? io_ins_222 : _GEN_221; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_223 = 9'hdf == io_sel ? io_ins_223 : _GEN_222; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_224 = 9'he0 == io_sel ? io_ins_224 : _GEN_223; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_225 = 9'he1 == io_sel ? io_ins_225 : _GEN_224; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_226 = 9'he2 == io_sel ? io_ins_226 : _GEN_225; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_227 = 9'he3 == io_sel ? io_ins_227 : _GEN_226; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_228 = 9'he4 == io_sel ? io_ins_228 : _GEN_227; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_229 = 9'he5 == io_sel ? io_ins_229 : _GEN_228; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_230 = 9'he6 == io_sel ? io_ins_230 : _GEN_229; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_231 = 9'he7 == io_sel ? io_ins_231 : _GEN_230; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_232 = 9'he8 == io_sel ? io_ins_232 : _GEN_231; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_233 = 9'he9 == io_sel ? io_ins_233 : _GEN_232; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_234 = 9'hea == io_sel ? io_ins_234 : _GEN_233; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_235 = 9'heb == io_sel ? io_ins_235 : _GEN_234; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_236 = 9'hec == io_sel ? io_ins_236 : _GEN_235; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_237 = 9'hed == io_sel ? io_ins_237 : _GEN_236; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_238 = 9'hee == io_sel ? io_ins_238 : _GEN_237; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_239 = 9'hef == io_sel ? io_ins_239 : _GEN_238; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_240 = 9'hf0 == io_sel ? io_ins_240 : _GEN_239; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_241 = 9'hf1 == io_sel ? io_ins_241 : _GEN_240; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_242 = 9'hf2 == io_sel ? io_ins_242 : _GEN_241; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_243 = 9'hf3 == io_sel ? io_ins_243 : _GEN_242; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_244 = 9'hf4 == io_sel ? io_ins_244 : _GEN_243; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_245 = 9'hf5 == io_sel ? io_ins_245 : _GEN_244; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_246 = 9'hf6 == io_sel ? io_ins_246 : _GEN_245; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_247 = 9'hf7 == io_sel ? io_ins_247 : _GEN_246; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_248 = 9'hf8 == io_sel ? io_ins_248 : _GEN_247; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_249 = 9'hf9 == io_sel ? io_ins_249 : _GEN_248; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_250 = 9'hfa == io_sel ? io_ins_250 : _GEN_249; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_251 = 9'hfb == io_sel ? io_ins_251 : _GEN_250; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_252 = 9'hfc == io_sel ? io_ins_252 : _GEN_251; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_253 = 9'hfd == io_sel ? io_ins_253 : _GEN_252; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_254 = 9'hfe == io_sel ? io_ins_254 : _GEN_253; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_255 = 9'hff == io_sel ? io_ins_255 : _GEN_254; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_256 = 9'h100 == io_sel ? io_ins_256 : _GEN_255; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_257 = 9'h101 == io_sel ? io_ins_257 : _GEN_256; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_258 = 9'h102 == io_sel ? io_ins_258 : _GEN_257; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_259 = 9'h103 == io_sel ? io_ins_259 : _GEN_258; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_260 = 9'h104 == io_sel ? io_ins_260 : _GEN_259; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_261 = 9'h105 == io_sel ? io_ins_261 : _GEN_260; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_262 = 9'h106 == io_sel ? io_ins_262 : _GEN_261; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_263 = 9'h107 == io_sel ? io_ins_263 : _GEN_262; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_264 = 9'h108 == io_sel ? io_ins_264 : _GEN_263; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_265 = 9'h109 == io_sel ? io_ins_265 : _GEN_264; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_266 = 9'h10a == io_sel ? io_ins_266 : _GEN_265; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_267 = 9'h10b == io_sel ? io_ins_267 : _GEN_266; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_268 = 9'h10c == io_sel ? io_ins_268 : _GEN_267; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_269 = 9'h10d == io_sel ? io_ins_269 : _GEN_268; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_270 = 9'h10e == io_sel ? io_ins_270 : _GEN_269; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_271 = 9'h10f == io_sel ? io_ins_271 : _GEN_270; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_272 = 9'h110 == io_sel ? io_ins_272 : _GEN_271; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_273 = 9'h111 == io_sel ? io_ins_273 : _GEN_272; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_274 = 9'h112 == io_sel ? io_ins_274 : _GEN_273; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_275 = 9'h113 == io_sel ? io_ins_275 : _GEN_274; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_276 = 9'h114 == io_sel ? io_ins_276 : _GEN_275; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_277 = 9'h115 == io_sel ? io_ins_277 : _GEN_276; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_278 = 9'h116 == io_sel ? io_ins_278 : _GEN_277; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_279 = 9'h117 == io_sel ? io_ins_279 : _GEN_278; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_280 = 9'h118 == io_sel ? io_ins_280 : _GEN_279; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_281 = 9'h119 == io_sel ? io_ins_281 : _GEN_280; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_282 = 9'h11a == io_sel ? io_ins_282 : _GEN_281; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_283 = 9'h11b == io_sel ? io_ins_283 : _GEN_282; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_284 = 9'h11c == io_sel ? io_ins_284 : _GEN_283; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_285 = 9'h11d == io_sel ? io_ins_285 : _GEN_284; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_286 = 9'h11e == io_sel ? io_ins_286 : _GEN_285; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_287 = 9'h11f == io_sel ? io_ins_287 : _GEN_286; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_288 = 9'h120 == io_sel ? io_ins_288 : _GEN_287; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_289 = 9'h121 == io_sel ? io_ins_289 : _GEN_288; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_290 = 9'h122 == io_sel ? io_ins_290 : _GEN_289; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_291 = 9'h123 == io_sel ? io_ins_291 : _GEN_290; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_292 = 9'h124 == io_sel ? io_ins_292 : _GEN_291; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_293 = 9'h125 == io_sel ? io_ins_293 : _GEN_292; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_294 = 9'h126 == io_sel ? io_ins_294 : _GEN_293; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_295 = 9'h127 == io_sel ? io_ins_295 : _GEN_294; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_296 = 9'h128 == io_sel ? io_ins_296 : _GEN_295; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_297 = 9'h129 == io_sel ? io_ins_297 : _GEN_296; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_298 = 9'h12a == io_sel ? io_ins_298 : _GEN_297; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_299 = 9'h12b == io_sel ? io_ins_299 : _GEN_298; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_300 = 9'h12c == io_sel ? io_ins_300 : _GEN_299; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_301 = 9'h12d == io_sel ? io_ins_301 : _GEN_300; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_302 = 9'h12e == io_sel ? io_ins_302 : _GEN_301; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_303 = 9'h12f == io_sel ? io_ins_303 : _GEN_302; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_304 = 9'h130 == io_sel ? io_ins_304 : _GEN_303; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_305 = 9'h131 == io_sel ? io_ins_305 : _GEN_304; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_306 = 9'h132 == io_sel ? io_ins_306 : _GEN_305; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_307 = 9'h133 == io_sel ? io_ins_307 : _GEN_306; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_308 = 9'h134 == io_sel ? io_ins_308 : _GEN_307; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_309 = 9'h135 == io_sel ? io_ins_309 : _GEN_308; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_310 = 9'h136 == io_sel ? io_ins_310 : _GEN_309; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_311 = 9'h137 == io_sel ? io_ins_311 : _GEN_310; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_312 = 9'h138 == io_sel ? io_ins_312 : _GEN_311; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_313 = 9'h139 == io_sel ? io_ins_313 : _GEN_312; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_314 = 9'h13a == io_sel ? io_ins_314 : _GEN_313; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_315 = 9'h13b == io_sel ? io_ins_315 : _GEN_314; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_316 = 9'h13c == io_sel ? io_ins_316 : _GEN_315; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_317 = 9'h13d == io_sel ? io_ins_317 : _GEN_316; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_318 = 9'h13e == io_sel ? io_ins_318 : _GEN_317; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_319 = 9'h13f == io_sel ? io_ins_319 : _GEN_318; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_320 = 9'h140 == io_sel ? io_ins_320 : _GEN_319; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_321 = 9'h141 == io_sel ? io_ins_321 : _GEN_320; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_322 = 9'h142 == io_sel ? io_ins_322 : _GEN_321; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_323 = 9'h143 == io_sel ? io_ins_323 : _GEN_322; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_324 = 9'h144 == io_sel ? io_ins_324 : _GEN_323; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_325 = 9'h145 == io_sel ? io_ins_325 : _GEN_324; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_326 = 9'h146 == io_sel ? io_ins_326 : _GEN_325; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_327 = 9'h147 == io_sel ? io_ins_327 : _GEN_326; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_328 = 9'h148 == io_sel ? io_ins_328 : _GEN_327; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_329 = 9'h149 == io_sel ? io_ins_329 : _GEN_328; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_330 = 9'h14a == io_sel ? io_ins_330 : _GEN_329; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_331 = 9'h14b == io_sel ? io_ins_331 : _GEN_330; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_332 = 9'h14c == io_sel ? io_ins_332 : _GEN_331; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_333 = 9'h14d == io_sel ? io_ins_333 : _GEN_332; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_334 = 9'h14e == io_sel ? io_ins_334 : _GEN_333; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_335 = 9'h14f == io_sel ? io_ins_335 : _GEN_334; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_336 = 9'h150 == io_sel ? io_ins_336 : _GEN_335; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_337 = 9'h151 == io_sel ? io_ins_337 : _GEN_336; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_338 = 9'h152 == io_sel ? io_ins_338 : _GEN_337; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_339 = 9'h153 == io_sel ? io_ins_339 : _GEN_338; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_340 = 9'h154 == io_sel ? io_ins_340 : _GEN_339; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_341 = 9'h155 == io_sel ? io_ins_341 : _GEN_340; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_342 = 9'h156 == io_sel ? io_ins_342 : _GEN_341; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_343 = 9'h157 == io_sel ? io_ins_343 : _GEN_342; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_344 = 9'h158 == io_sel ? io_ins_344 : _GEN_343; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_345 = 9'h159 == io_sel ? io_ins_345 : _GEN_344; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_346 = 9'h15a == io_sel ? io_ins_346 : _GEN_345; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_347 = 9'h15b == io_sel ? io_ins_347 : _GEN_346; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_348 = 9'h15c == io_sel ? io_ins_348 : _GEN_347; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_349 = 9'h15d == io_sel ? io_ins_349 : _GEN_348; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_350 = 9'h15e == io_sel ? io_ins_350 : _GEN_349; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_351 = 9'h15f == io_sel ? io_ins_351 : _GEN_350; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_352 = 9'h160 == io_sel ? io_ins_352 : _GEN_351; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_353 = 9'h161 == io_sel ? io_ins_353 : _GEN_352; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_354 = 9'h162 == io_sel ? io_ins_354 : _GEN_353; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_355 = 9'h163 == io_sel ? io_ins_355 : _GEN_354; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_356 = 9'h164 == io_sel ? io_ins_356 : _GEN_355; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_357 = 9'h165 == io_sel ? io_ins_357 : _GEN_356; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_358 = 9'h166 == io_sel ? io_ins_358 : _GEN_357; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_359 = 9'h167 == io_sel ? io_ins_359 : _GEN_358; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_360 = 9'h168 == io_sel ? io_ins_360 : _GEN_359; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_361 = 9'h169 == io_sel ? io_ins_361 : _GEN_360; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_362 = 9'h16a == io_sel ? io_ins_362 : _GEN_361; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_363 = 9'h16b == io_sel ? io_ins_363 : _GEN_362; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_364 = 9'h16c == io_sel ? io_ins_364 : _GEN_363; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_365 = 9'h16d == io_sel ? io_ins_365 : _GEN_364; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_366 = 9'h16e == io_sel ? io_ins_366 : _GEN_365; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_367 = 9'h16f == io_sel ? io_ins_367 : _GEN_366; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_368 = 9'h170 == io_sel ? io_ins_368 : _GEN_367; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_369 = 9'h171 == io_sel ? io_ins_369 : _GEN_368; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_370 = 9'h172 == io_sel ? io_ins_370 : _GEN_369; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_371 = 9'h173 == io_sel ? io_ins_371 : _GEN_370; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_372 = 9'h174 == io_sel ? io_ins_372 : _GEN_371; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_373 = 9'h175 == io_sel ? io_ins_373 : _GEN_372; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_374 = 9'h176 == io_sel ? io_ins_374 : _GEN_373; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_375 = 9'h177 == io_sel ? io_ins_375 : _GEN_374; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_376 = 9'h178 == io_sel ? io_ins_376 : _GEN_375; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_377 = 9'h179 == io_sel ? io_ins_377 : _GEN_376; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_378 = 9'h17a == io_sel ? io_ins_378 : _GEN_377; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_379 = 9'h17b == io_sel ? io_ins_379 : _GEN_378; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_380 = 9'h17c == io_sel ? io_ins_380 : _GEN_379; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_381 = 9'h17d == io_sel ? io_ins_381 : _GEN_380; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_382 = 9'h17e == io_sel ? io_ins_382 : _GEN_381; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_383 = 9'h17f == io_sel ? io_ins_383 : _GEN_382; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_384 = 9'h180 == io_sel ? io_ins_384 : _GEN_383; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_385 = 9'h181 == io_sel ? io_ins_385 : _GEN_384; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_386 = 9'h182 == io_sel ? io_ins_386 : _GEN_385; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_387 = 9'h183 == io_sel ? io_ins_387 : _GEN_386; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_388 = 9'h184 == io_sel ? io_ins_388 : _GEN_387; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_389 = 9'h185 == io_sel ? io_ins_389 : _GEN_388; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_390 = 9'h186 == io_sel ? io_ins_390 : _GEN_389; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_391 = 9'h187 == io_sel ? io_ins_391 : _GEN_390; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_392 = 9'h188 == io_sel ? io_ins_392 : _GEN_391; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_393 = 9'h189 == io_sel ? io_ins_393 : _GEN_392; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_394 = 9'h18a == io_sel ? io_ins_394 : _GEN_393; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_395 = 9'h18b == io_sel ? io_ins_395 : _GEN_394; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_396 = 9'h18c == io_sel ? io_ins_396 : _GEN_395; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_397 = 9'h18d == io_sel ? io_ins_397 : _GEN_396; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_398 = 9'h18e == io_sel ? io_ins_398 : _GEN_397; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_399 = 9'h18f == io_sel ? io_ins_399 : _GEN_398; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_400 = 9'h190 == io_sel ? io_ins_400 : _GEN_399; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_401 = 9'h191 == io_sel ? io_ins_401 : _GEN_400; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_402 = 9'h192 == io_sel ? io_ins_402 : _GEN_401; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_403 = 9'h193 == io_sel ? io_ins_403 : _GEN_402; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_404 = 9'h194 == io_sel ? io_ins_404 : _GEN_403; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_405 = 9'h195 == io_sel ? io_ins_405 : _GEN_404; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_406 = 9'h196 == io_sel ? io_ins_406 : _GEN_405; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_407 = 9'h197 == io_sel ? io_ins_407 : _GEN_406; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_408 = 9'h198 == io_sel ? io_ins_408 : _GEN_407; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_409 = 9'h199 == io_sel ? io_ins_409 : _GEN_408; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_410 = 9'h19a == io_sel ? io_ins_410 : _GEN_409; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_411 = 9'h19b == io_sel ? io_ins_411 : _GEN_410; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_412 = 9'h19c == io_sel ? io_ins_412 : _GEN_411; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_413 = 9'h19d == io_sel ? io_ins_413 : _GEN_412; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_414 = 9'h19e == io_sel ? io_ins_414 : _GEN_413; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_415 = 9'h19f == io_sel ? io_ins_415 : _GEN_414; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_416 = 9'h1a0 == io_sel ? io_ins_416 : _GEN_415; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_417 = 9'h1a1 == io_sel ? io_ins_417 : _GEN_416; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_418 = 9'h1a2 == io_sel ? io_ins_418 : _GEN_417; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_419 = 9'h1a3 == io_sel ? io_ins_419 : _GEN_418; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_420 = 9'h1a4 == io_sel ? io_ins_420 : _GEN_419; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_421 = 9'h1a5 == io_sel ? io_ins_421 : _GEN_420; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_422 = 9'h1a6 == io_sel ? io_ins_422 : _GEN_421; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_423 = 9'h1a7 == io_sel ? io_ins_423 : _GEN_422; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_424 = 9'h1a8 == io_sel ? io_ins_424 : _GEN_423; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_425 = 9'h1a9 == io_sel ? io_ins_425 : _GEN_424; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_426 = 9'h1aa == io_sel ? io_ins_426 : _GEN_425; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_427 = 9'h1ab == io_sel ? io_ins_427 : _GEN_426; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_428 = 9'h1ac == io_sel ? io_ins_428 : _GEN_427; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_429 = 9'h1ad == io_sel ? io_ins_429 : _GEN_428; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_430 = 9'h1ae == io_sel ? io_ins_430 : _GEN_429; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_431 = 9'h1af == io_sel ? io_ins_431 : _GEN_430; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_432 = 9'h1b0 == io_sel ? io_ins_432 : _GEN_431; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_433 = 9'h1b1 == io_sel ? io_ins_433 : _GEN_432; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_434 = 9'h1b2 == io_sel ? io_ins_434 : _GEN_433; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_435 = 9'h1b3 == io_sel ? io_ins_435 : _GEN_434; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_436 = 9'h1b4 == io_sel ? io_ins_436 : _GEN_435; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_437 = 9'h1b5 == io_sel ? io_ins_437 : _GEN_436; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_438 = 9'h1b6 == io_sel ? io_ins_438 : _GEN_437; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_439 = 9'h1b7 == io_sel ? io_ins_439 : _GEN_438; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_440 = 9'h1b8 == io_sel ? io_ins_440 : _GEN_439; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_441 = 9'h1b9 == io_sel ? io_ins_441 : _GEN_440; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_442 = 9'h1ba == io_sel ? io_ins_442 : _GEN_441; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_443 = 9'h1bb == io_sel ? io_ins_443 : _GEN_442; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_444 = 9'h1bc == io_sel ? io_ins_444 : _GEN_443; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_445 = 9'h1bd == io_sel ? io_ins_445 : _GEN_444; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_446 = 9'h1be == io_sel ? io_ins_446 : _GEN_445; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_447 = 9'h1bf == io_sel ? io_ins_447 : _GEN_446; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_448 = 9'h1c0 == io_sel ? io_ins_448 : _GEN_447; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_449 = 9'h1c1 == io_sel ? io_ins_449 : _GEN_448; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_450 = 9'h1c2 == io_sel ? io_ins_450 : _GEN_449; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_451 = 9'h1c3 == io_sel ? io_ins_451 : _GEN_450; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_452 = 9'h1c4 == io_sel ? io_ins_452 : _GEN_451; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_453 = 9'h1c5 == io_sel ? io_ins_453 : _GEN_452; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_454 = 9'h1c6 == io_sel ? io_ins_454 : _GEN_453; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_455 = 9'h1c7 == io_sel ? io_ins_455 : _GEN_454; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_456 = 9'h1c8 == io_sel ? io_ins_456 : _GEN_455; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_457 = 9'h1c9 == io_sel ? io_ins_457 : _GEN_456; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_458 = 9'h1ca == io_sel ? io_ins_458 : _GEN_457; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_459 = 9'h1cb == io_sel ? io_ins_459 : _GEN_458; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_460 = 9'h1cc == io_sel ? io_ins_460 : _GEN_459; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_461 = 9'h1cd == io_sel ? io_ins_461 : _GEN_460; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_462 = 9'h1ce == io_sel ? io_ins_462 : _GEN_461; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_463 = 9'h1cf == io_sel ? io_ins_463 : _GEN_462; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_464 = 9'h1d0 == io_sel ? io_ins_464 : _GEN_463; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_465 = 9'h1d1 == io_sel ? io_ins_465 : _GEN_464; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_466 = 9'h1d2 == io_sel ? io_ins_466 : _GEN_465; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_467 = 9'h1d3 == io_sel ? io_ins_467 : _GEN_466; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_468 = 9'h1d4 == io_sel ? io_ins_468 : _GEN_467; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_469 = 9'h1d5 == io_sel ? io_ins_469 : _GEN_468; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_470 = 9'h1d6 == io_sel ? io_ins_470 : _GEN_469; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_471 = 9'h1d7 == io_sel ? io_ins_471 : _GEN_470; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_472 = 9'h1d8 == io_sel ? io_ins_472 : _GEN_471; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_473 = 9'h1d9 == io_sel ? io_ins_473 : _GEN_472; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_474 = 9'h1da == io_sel ? io_ins_474 : _GEN_473; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_475 = 9'h1db == io_sel ? io_ins_475 : _GEN_474; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_476 = 9'h1dc == io_sel ? io_ins_476 : _GEN_475; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_477 = 9'h1dd == io_sel ? io_ins_477 : _GEN_476; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_478 = 9'h1de == io_sel ? io_ins_478 : _GEN_477; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_479 = 9'h1df == io_sel ? io_ins_479 : _GEN_478; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_480 = 9'h1e0 == io_sel ? io_ins_480 : _GEN_479; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_481 = 9'h1e1 == io_sel ? io_ins_481 : _GEN_480; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_482 = 9'h1e2 == io_sel ? io_ins_482 : _GEN_481; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_483 = 9'h1e3 == io_sel ? io_ins_483 : _GEN_482; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_484 = 9'h1e4 == io_sel ? io_ins_484 : _GEN_483; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_485 = 9'h1e5 == io_sel ? io_ins_485 : _GEN_484; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_486 = 9'h1e6 == io_sel ? io_ins_486 : _GEN_485; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_487 = 9'h1e7 == io_sel ? io_ins_487 : _GEN_486; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_488 = 9'h1e8 == io_sel ? io_ins_488 : _GEN_487; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_489 = 9'h1e9 == io_sel ? io_ins_489 : _GEN_488; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_490 = 9'h1ea == io_sel ? io_ins_490 : _GEN_489; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_491 = 9'h1eb == io_sel ? io_ins_491 : _GEN_490; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_492 = 9'h1ec == io_sel ? io_ins_492 : _GEN_491; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_493 = 9'h1ed == io_sel ? io_ins_493 : _GEN_492; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_494 = 9'h1ee == io_sel ? io_ins_494 : _GEN_493; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_495 = 9'h1ef == io_sel ? io_ins_495 : _GEN_494; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_496 = 9'h1f0 == io_sel ? io_ins_496 : _GEN_495; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_497 = 9'h1f1 == io_sel ? io_ins_497 : _GEN_496; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_498 = 9'h1f2 == io_sel ? io_ins_498 : _GEN_497; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_499 = 9'h1f3 == io_sel ? io_ins_499 : _GEN_498; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_500 = 9'h1f4 == io_sel ? io_ins_500 : _GEN_499; // @[MuxN.scala 16:10:@32395.4]
  assign _GEN_501 = 9'h1f5 == io_sel ? io_ins_501 : _GEN_500; // @[MuxN.scala 16:10:@32395.4]
  assign io_out = 9'h1f6 == io_sel ? io_ins_502 : _GEN_501; // @[MuxN.scala 16:10:@32395.4]
endmodule
module RegFile( // @[:@32397.2]
  input         clock, // @[:@32398.4]
  input         reset, // @[:@32399.4]
  input  [9:0]  io_raddr, // @[:@32400.4]
  input         io_wen, // @[:@32400.4]
  input  [9:0]  io_waddr, // @[:@32400.4]
  input  [63:0] io_wdata, // @[:@32400.4]
  output [63:0] io_rdata, // @[:@32400.4]
  input         io_reset, // @[:@32400.4]
  output [63:0] io_argIns_0, // @[:@32400.4]
  output [63:0] io_argIns_1, // @[:@32400.4]
  output [63:0] io_argIns_2, // @[:@32400.4]
  input         io_argOuts_0_valid, // @[:@32400.4]
  input  [63:0] io_argOuts_0_bits, // @[:@32400.4]
  input         io_argOuts_1_valid, // @[:@32400.4]
  input  [63:0] io_argOuts_1_bits, // @[:@32400.4]
  output [63:0] io_argEchos_1 // @[:@32400.4]
);
  wire  regs_0_clock; // @[RegFile.scala 66:20:@34410.4]
  wire  regs_0_reset; // @[RegFile.scala 66:20:@34410.4]
  wire [63:0] regs_0_io_in; // @[RegFile.scala 66:20:@34410.4]
  wire  regs_0_io_reset; // @[RegFile.scala 66:20:@34410.4]
  wire [63:0] regs_0_io_out; // @[RegFile.scala 66:20:@34410.4]
  wire  regs_0_io_enable; // @[RegFile.scala 66:20:@34410.4]
  wire  regs_1_clock; // @[RegFile.scala 66:20:@34422.4]
  wire  regs_1_reset; // @[RegFile.scala 66:20:@34422.4]
  wire [63:0] regs_1_io_in; // @[RegFile.scala 66:20:@34422.4]
  wire  regs_1_io_reset; // @[RegFile.scala 66:20:@34422.4]
  wire [63:0] regs_1_io_out; // @[RegFile.scala 66:20:@34422.4]
  wire  regs_1_io_enable; // @[RegFile.scala 66:20:@34422.4]
  wire  regs_2_clock; // @[RegFile.scala 66:20:@34441.4]
  wire  regs_2_reset; // @[RegFile.scala 66:20:@34441.4]
  wire [63:0] regs_2_io_in; // @[RegFile.scala 66:20:@34441.4]
  wire  regs_2_io_reset; // @[RegFile.scala 66:20:@34441.4]
  wire [63:0] regs_2_io_out; // @[RegFile.scala 66:20:@34441.4]
  wire  regs_2_io_enable; // @[RegFile.scala 66:20:@34441.4]
  wire  regs_3_clock; // @[RegFile.scala 66:20:@34453.4]
  wire  regs_3_reset; // @[RegFile.scala 66:20:@34453.4]
  wire [63:0] regs_3_io_in; // @[RegFile.scala 66:20:@34453.4]
  wire  regs_3_io_reset; // @[RegFile.scala 66:20:@34453.4]
  wire [63:0] regs_3_io_out; // @[RegFile.scala 66:20:@34453.4]
  wire  regs_3_io_enable; // @[RegFile.scala 66:20:@34453.4]
  wire  regs_4_clock; // @[RegFile.scala 66:20:@34467.4]
  wire  regs_4_reset; // @[RegFile.scala 66:20:@34467.4]
  wire [63:0] regs_4_io_in; // @[RegFile.scala 66:20:@34467.4]
  wire  regs_4_io_reset; // @[RegFile.scala 66:20:@34467.4]
  wire [63:0] regs_4_io_out; // @[RegFile.scala 66:20:@34467.4]
  wire  regs_4_io_enable; // @[RegFile.scala 66:20:@34467.4]
  wire  regs_5_clock; // @[RegFile.scala 66:20:@34481.4]
  wire  regs_5_reset; // @[RegFile.scala 66:20:@34481.4]
  wire [63:0] regs_5_io_in; // @[RegFile.scala 66:20:@34481.4]
  wire  regs_5_io_reset; // @[RegFile.scala 66:20:@34481.4]
  wire [63:0] regs_5_io_out; // @[RegFile.scala 66:20:@34481.4]
  wire  regs_5_io_enable; // @[RegFile.scala 66:20:@34481.4]
  wire  regs_6_clock; // @[RegFile.scala 66:20:@34495.4]
  wire  regs_6_reset; // @[RegFile.scala 66:20:@34495.4]
  wire [63:0] regs_6_io_in; // @[RegFile.scala 66:20:@34495.4]
  wire  regs_6_io_reset; // @[RegFile.scala 66:20:@34495.4]
  wire [63:0] regs_6_io_out; // @[RegFile.scala 66:20:@34495.4]
  wire  regs_6_io_enable; // @[RegFile.scala 66:20:@34495.4]
  wire  regs_7_clock; // @[RegFile.scala 66:20:@34509.4]
  wire  regs_7_reset; // @[RegFile.scala 66:20:@34509.4]
  wire [63:0] regs_7_io_in; // @[RegFile.scala 66:20:@34509.4]
  wire  regs_7_io_reset; // @[RegFile.scala 66:20:@34509.4]
  wire [63:0] regs_7_io_out; // @[RegFile.scala 66:20:@34509.4]
  wire  regs_7_io_enable; // @[RegFile.scala 66:20:@34509.4]
  wire  regs_8_clock; // @[RegFile.scala 66:20:@34523.4]
  wire  regs_8_reset; // @[RegFile.scala 66:20:@34523.4]
  wire [63:0] regs_8_io_in; // @[RegFile.scala 66:20:@34523.4]
  wire  regs_8_io_reset; // @[RegFile.scala 66:20:@34523.4]
  wire [63:0] regs_8_io_out; // @[RegFile.scala 66:20:@34523.4]
  wire  regs_8_io_enable; // @[RegFile.scala 66:20:@34523.4]
  wire  regs_9_clock; // @[RegFile.scala 66:20:@34537.4]
  wire  regs_9_reset; // @[RegFile.scala 66:20:@34537.4]
  wire [63:0] regs_9_io_in; // @[RegFile.scala 66:20:@34537.4]
  wire  regs_9_io_reset; // @[RegFile.scala 66:20:@34537.4]
  wire [63:0] regs_9_io_out; // @[RegFile.scala 66:20:@34537.4]
  wire  regs_9_io_enable; // @[RegFile.scala 66:20:@34537.4]
  wire  regs_10_clock; // @[RegFile.scala 66:20:@34551.4]
  wire  regs_10_reset; // @[RegFile.scala 66:20:@34551.4]
  wire [63:0] regs_10_io_in; // @[RegFile.scala 66:20:@34551.4]
  wire  regs_10_io_reset; // @[RegFile.scala 66:20:@34551.4]
  wire [63:0] regs_10_io_out; // @[RegFile.scala 66:20:@34551.4]
  wire  regs_10_io_enable; // @[RegFile.scala 66:20:@34551.4]
  wire  regs_11_clock; // @[RegFile.scala 66:20:@34565.4]
  wire  regs_11_reset; // @[RegFile.scala 66:20:@34565.4]
  wire [63:0] regs_11_io_in; // @[RegFile.scala 66:20:@34565.4]
  wire  regs_11_io_reset; // @[RegFile.scala 66:20:@34565.4]
  wire [63:0] regs_11_io_out; // @[RegFile.scala 66:20:@34565.4]
  wire  regs_11_io_enable; // @[RegFile.scala 66:20:@34565.4]
  wire  regs_12_clock; // @[RegFile.scala 66:20:@34579.4]
  wire  regs_12_reset; // @[RegFile.scala 66:20:@34579.4]
  wire [63:0] regs_12_io_in; // @[RegFile.scala 66:20:@34579.4]
  wire  regs_12_io_reset; // @[RegFile.scala 66:20:@34579.4]
  wire [63:0] regs_12_io_out; // @[RegFile.scala 66:20:@34579.4]
  wire  regs_12_io_enable; // @[RegFile.scala 66:20:@34579.4]
  wire  regs_13_clock; // @[RegFile.scala 66:20:@34593.4]
  wire  regs_13_reset; // @[RegFile.scala 66:20:@34593.4]
  wire [63:0] regs_13_io_in; // @[RegFile.scala 66:20:@34593.4]
  wire  regs_13_io_reset; // @[RegFile.scala 66:20:@34593.4]
  wire [63:0] regs_13_io_out; // @[RegFile.scala 66:20:@34593.4]
  wire  regs_13_io_enable; // @[RegFile.scala 66:20:@34593.4]
  wire  regs_14_clock; // @[RegFile.scala 66:20:@34607.4]
  wire  regs_14_reset; // @[RegFile.scala 66:20:@34607.4]
  wire [63:0] regs_14_io_in; // @[RegFile.scala 66:20:@34607.4]
  wire  regs_14_io_reset; // @[RegFile.scala 66:20:@34607.4]
  wire [63:0] regs_14_io_out; // @[RegFile.scala 66:20:@34607.4]
  wire  regs_14_io_enable; // @[RegFile.scala 66:20:@34607.4]
  wire  regs_15_clock; // @[RegFile.scala 66:20:@34621.4]
  wire  regs_15_reset; // @[RegFile.scala 66:20:@34621.4]
  wire [63:0] regs_15_io_in; // @[RegFile.scala 66:20:@34621.4]
  wire  regs_15_io_reset; // @[RegFile.scala 66:20:@34621.4]
  wire [63:0] regs_15_io_out; // @[RegFile.scala 66:20:@34621.4]
  wire  regs_15_io_enable; // @[RegFile.scala 66:20:@34621.4]
  wire  regs_16_clock; // @[RegFile.scala 66:20:@34635.4]
  wire  regs_16_reset; // @[RegFile.scala 66:20:@34635.4]
  wire [63:0] regs_16_io_in; // @[RegFile.scala 66:20:@34635.4]
  wire  regs_16_io_reset; // @[RegFile.scala 66:20:@34635.4]
  wire [63:0] regs_16_io_out; // @[RegFile.scala 66:20:@34635.4]
  wire  regs_16_io_enable; // @[RegFile.scala 66:20:@34635.4]
  wire  regs_17_clock; // @[RegFile.scala 66:20:@34649.4]
  wire  regs_17_reset; // @[RegFile.scala 66:20:@34649.4]
  wire [63:0] regs_17_io_in; // @[RegFile.scala 66:20:@34649.4]
  wire  regs_17_io_reset; // @[RegFile.scala 66:20:@34649.4]
  wire [63:0] regs_17_io_out; // @[RegFile.scala 66:20:@34649.4]
  wire  regs_17_io_enable; // @[RegFile.scala 66:20:@34649.4]
  wire  regs_18_clock; // @[RegFile.scala 66:20:@34663.4]
  wire  regs_18_reset; // @[RegFile.scala 66:20:@34663.4]
  wire [63:0] regs_18_io_in; // @[RegFile.scala 66:20:@34663.4]
  wire  regs_18_io_reset; // @[RegFile.scala 66:20:@34663.4]
  wire [63:0] regs_18_io_out; // @[RegFile.scala 66:20:@34663.4]
  wire  regs_18_io_enable; // @[RegFile.scala 66:20:@34663.4]
  wire  regs_19_clock; // @[RegFile.scala 66:20:@34677.4]
  wire  regs_19_reset; // @[RegFile.scala 66:20:@34677.4]
  wire [63:0] regs_19_io_in; // @[RegFile.scala 66:20:@34677.4]
  wire  regs_19_io_reset; // @[RegFile.scala 66:20:@34677.4]
  wire [63:0] regs_19_io_out; // @[RegFile.scala 66:20:@34677.4]
  wire  regs_19_io_enable; // @[RegFile.scala 66:20:@34677.4]
  wire  regs_20_clock; // @[RegFile.scala 66:20:@34691.4]
  wire  regs_20_reset; // @[RegFile.scala 66:20:@34691.4]
  wire [63:0] regs_20_io_in; // @[RegFile.scala 66:20:@34691.4]
  wire  regs_20_io_reset; // @[RegFile.scala 66:20:@34691.4]
  wire [63:0] regs_20_io_out; // @[RegFile.scala 66:20:@34691.4]
  wire  regs_20_io_enable; // @[RegFile.scala 66:20:@34691.4]
  wire  regs_21_clock; // @[RegFile.scala 66:20:@34705.4]
  wire  regs_21_reset; // @[RegFile.scala 66:20:@34705.4]
  wire [63:0] regs_21_io_in; // @[RegFile.scala 66:20:@34705.4]
  wire  regs_21_io_reset; // @[RegFile.scala 66:20:@34705.4]
  wire [63:0] regs_21_io_out; // @[RegFile.scala 66:20:@34705.4]
  wire  regs_21_io_enable; // @[RegFile.scala 66:20:@34705.4]
  wire  regs_22_clock; // @[RegFile.scala 66:20:@34719.4]
  wire  regs_22_reset; // @[RegFile.scala 66:20:@34719.4]
  wire [63:0] regs_22_io_in; // @[RegFile.scala 66:20:@34719.4]
  wire  regs_22_io_reset; // @[RegFile.scala 66:20:@34719.4]
  wire [63:0] regs_22_io_out; // @[RegFile.scala 66:20:@34719.4]
  wire  regs_22_io_enable; // @[RegFile.scala 66:20:@34719.4]
  wire  regs_23_clock; // @[RegFile.scala 66:20:@34733.4]
  wire  regs_23_reset; // @[RegFile.scala 66:20:@34733.4]
  wire [63:0] regs_23_io_in; // @[RegFile.scala 66:20:@34733.4]
  wire  regs_23_io_reset; // @[RegFile.scala 66:20:@34733.4]
  wire [63:0] regs_23_io_out; // @[RegFile.scala 66:20:@34733.4]
  wire  regs_23_io_enable; // @[RegFile.scala 66:20:@34733.4]
  wire  regs_24_clock; // @[RegFile.scala 66:20:@34747.4]
  wire  regs_24_reset; // @[RegFile.scala 66:20:@34747.4]
  wire [63:0] regs_24_io_in; // @[RegFile.scala 66:20:@34747.4]
  wire  regs_24_io_reset; // @[RegFile.scala 66:20:@34747.4]
  wire [63:0] regs_24_io_out; // @[RegFile.scala 66:20:@34747.4]
  wire  regs_24_io_enable; // @[RegFile.scala 66:20:@34747.4]
  wire  regs_25_clock; // @[RegFile.scala 66:20:@34761.4]
  wire  regs_25_reset; // @[RegFile.scala 66:20:@34761.4]
  wire [63:0] regs_25_io_in; // @[RegFile.scala 66:20:@34761.4]
  wire  regs_25_io_reset; // @[RegFile.scala 66:20:@34761.4]
  wire [63:0] regs_25_io_out; // @[RegFile.scala 66:20:@34761.4]
  wire  regs_25_io_enable; // @[RegFile.scala 66:20:@34761.4]
  wire  regs_26_clock; // @[RegFile.scala 66:20:@34775.4]
  wire  regs_26_reset; // @[RegFile.scala 66:20:@34775.4]
  wire [63:0] regs_26_io_in; // @[RegFile.scala 66:20:@34775.4]
  wire  regs_26_io_reset; // @[RegFile.scala 66:20:@34775.4]
  wire [63:0] regs_26_io_out; // @[RegFile.scala 66:20:@34775.4]
  wire  regs_26_io_enable; // @[RegFile.scala 66:20:@34775.4]
  wire  regs_27_clock; // @[RegFile.scala 66:20:@34789.4]
  wire  regs_27_reset; // @[RegFile.scala 66:20:@34789.4]
  wire [63:0] regs_27_io_in; // @[RegFile.scala 66:20:@34789.4]
  wire  regs_27_io_reset; // @[RegFile.scala 66:20:@34789.4]
  wire [63:0] regs_27_io_out; // @[RegFile.scala 66:20:@34789.4]
  wire  regs_27_io_enable; // @[RegFile.scala 66:20:@34789.4]
  wire  regs_28_clock; // @[RegFile.scala 66:20:@34803.4]
  wire  regs_28_reset; // @[RegFile.scala 66:20:@34803.4]
  wire [63:0] regs_28_io_in; // @[RegFile.scala 66:20:@34803.4]
  wire  regs_28_io_reset; // @[RegFile.scala 66:20:@34803.4]
  wire [63:0] regs_28_io_out; // @[RegFile.scala 66:20:@34803.4]
  wire  regs_28_io_enable; // @[RegFile.scala 66:20:@34803.4]
  wire  regs_29_clock; // @[RegFile.scala 66:20:@34817.4]
  wire  regs_29_reset; // @[RegFile.scala 66:20:@34817.4]
  wire [63:0] regs_29_io_in; // @[RegFile.scala 66:20:@34817.4]
  wire  regs_29_io_reset; // @[RegFile.scala 66:20:@34817.4]
  wire [63:0] regs_29_io_out; // @[RegFile.scala 66:20:@34817.4]
  wire  regs_29_io_enable; // @[RegFile.scala 66:20:@34817.4]
  wire  regs_30_clock; // @[RegFile.scala 66:20:@34831.4]
  wire  regs_30_reset; // @[RegFile.scala 66:20:@34831.4]
  wire [63:0] regs_30_io_in; // @[RegFile.scala 66:20:@34831.4]
  wire  regs_30_io_reset; // @[RegFile.scala 66:20:@34831.4]
  wire [63:0] regs_30_io_out; // @[RegFile.scala 66:20:@34831.4]
  wire  regs_30_io_enable; // @[RegFile.scala 66:20:@34831.4]
  wire  regs_31_clock; // @[RegFile.scala 66:20:@34845.4]
  wire  regs_31_reset; // @[RegFile.scala 66:20:@34845.4]
  wire [63:0] regs_31_io_in; // @[RegFile.scala 66:20:@34845.4]
  wire  regs_31_io_reset; // @[RegFile.scala 66:20:@34845.4]
  wire [63:0] regs_31_io_out; // @[RegFile.scala 66:20:@34845.4]
  wire  regs_31_io_enable; // @[RegFile.scala 66:20:@34845.4]
  wire  regs_32_clock; // @[RegFile.scala 66:20:@34859.4]
  wire  regs_32_reset; // @[RegFile.scala 66:20:@34859.4]
  wire [63:0] regs_32_io_in; // @[RegFile.scala 66:20:@34859.4]
  wire  regs_32_io_reset; // @[RegFile.scala 66:20:@34859.4]
  wire [63:0] regs_32_io_out; // @[RegFile.scala 66:20:@34859.4]
  wire  regs_32_io_enable; // @[RegFile.scala 66:20:@34859.4]
  wire  regs_33_clock; // @[RegFile.scala 66:20:@34873.4]
  wire  regs_33_reset; // @[RegFile.scala 66:20:@34873.4]
  wire [63:0] regs_33_io_in; // @[RegFile.scala 66:20:@34873.4]
  wire  regs_33_io_reset; // @[RegFile.scala 66:20:@34873.4]
  wire [63:0] regs_33_io_out; // @[RegFile.scala 66:20:@34873.4]
  wire  regs_33_io_enable; // @[RegFile.scala 66:20:@34873.4]
  wire  regs_34_clock; // @[RegFile.scala 66:20:@34887.4]
  wire  regs_34_reset; // @[RegFile.scala 66:20:@34887.4]
  wire [63:0] regs_34_io_in; // @[RegFile.scala 66:20:@34887.4]
  wire  regs_34_io_reset; // @[RegFile.scala 66:20:@34887.4]
  wire [63:0] regs_34_io_out; // @[RegFile.scala 66:20:@34887.4]
  wire  regs_34_io_enable; // @[RegFile.scala 66:20:@34887.4]
  wire  regs_35_clock; // @[RegFile.scala 66:20:@34901.4]
  wire  regs_35_reset; // @[RegFile.scala 66:20:@34901.4]
  wire [63:0] regs_35_io_in; // @[RegFile.scala 66:20:@34901.4]
  wire  regs_35_io_reset; // @[RegFile.scala 66:20:@34901.4]
  wire [63:0] regs_35_io_out; // @[RegFile.scala 66:20:@34901.4]
  wire  regs_35_io_enable; // @[RegFile.scala 66:20:@34901.4]
  wire  regs_36_clock; // @[RegFile.scala 66:20:@34915.4]
  wire  regs_36_reset; // @[RegFile.scala 66:20:@34915.4]
  wire [63:0] regs_36_io_in; // @[RegFile.scala 66:20:@34915.4]
  wire  regs_36_io_reset; // @[RegFile.scala 66:20:@34915.4]
  wire [63:0] regs_36_io_out; // @[RegFile.scala 66:20:@34915.4]
  wire  regs_36_io_enable; // @[RegFile.scala 66:20:@34915.4]
  wire  regs_37_clock; // @[RegFile.scala 66:20:@34929.4]
  wire  regs_37_reset; // @[RegFile.scala 66:20:@34929.4]
  wire [63:0] regs_37_io_in; // @[RegFile.scala 66:20:@34929.4]
  wire  regs_37_io_reset; // @[RegFile.scala 66:20:@34929.4]
  wire [63:0] regs_37_io_out; // @[RegFile.scala 66:20:@34929.4]
  wire  regs_37_io_enable; // @[RegFile.scala 66:20:@34929.4]
  wire  regs_38_clock; // @[RegFile.scala 66:20:@34943.4]
  wire  regs_38_reset; // @[RegFile.scala 66:20:@34943.4]
  wire [63:0] regs_38_io_in; // @[RegFile.scala 66:20:@34943.4]
  wire  regs_38_io_reset; // @[RegFile.scala 66:20:@34943.4]
  wire [63:0] regs_38_io_out; // @[RegFile.scala 66:20:@34943.4]
  wire  regs_38_io_enable; // @[RegFile.scala 66:20:@34943.4]
  wire  regs_39_clock; // @[RegFile.scala 66:20:@34957.4]
  wire  regs_39_reset; // @[RegFile.scala 66:20:@34957.4]
  wire [63:0] regs_39_io_in; // @[RegFile.scala 66:20:@34957.4]
  wire  regs_39_io_reset; // @[RegFile.scala 66:20:@34957.4]
  wire [63:0] regs_39_io_out; // @[RegFile.scala 66:20:@34957.4]
  wire  regs_39_io_enable; // @[RegFile.scala 66:20:@34957.4]
  wire  regs_40_clock; // @[RegFile.scala 66:20:@34971.4]
  wire  regs_40_reset; // @[RegFile.scala 66:20:@34971.4]
  wire [63:0] regs_40_io_in; // @[RegFile.scala 66:20:@34971.4]
  wire  regs_40_io_reset; // @[RegFile.scala 66:20:@34971.4]
  wire [63:0] regs_40_io_out; // @[RegFile.scala 66:20:@34971.4]
  wire  regs_40_io_enable; // @[RegFile.scala 66:20:@34971.4]
  wire  regs_41_clock; // @[RegFile.scala 66:20:@34985.4]
  wire  regs_41_reset; // @[RegFile.scala 66:20:@34985.4]
  wire [63:0] regs_41_io_in; // @[RegFile.scala 66:20:@34985.4]
  wire  regs_41_io_reset; // @[RegFile.scala 66:20:@34985.4]
  wire [63:0] regs_41_io_out; // @[RegFile.scala 66:20:@34985.4]
  wire  regs_41_io_enable; // @[RegFile.scala 66:20:@34985.4]
  wire  regs_42_clock; // @[RegFile.scala 66:20:@34999.4]
  wire  regs_42_reset; // @[RegFile.scala 66:20:@34999.4]
  wire [63:0] regs_42_io_in; // @[RegFile.scala 66:20:@34999.4]
  wire  regs_42_io_reset; // @[RegFile.scala 66:20:@34999.4]
  wire [63:0] regs_42_io_out; // @[RegFile.scala 66:20:@34999.4]
  wire  regs_42_io_enable; // @[RegFile.scala 66:20:@34999.4]
  wire  regs_43_clock; // @[RegFile.scala 66:20:@35013.4]
  wire  regs_43_reset; // @[RegFile.scala 66:20:@35013.4]
  wire [63:0] regs_43_io_in; // @[RegFile.scala 66:20:@35013.4]
  wire  regs_43_io_reset; // @[RegFile.scala 66:20:@35013.4]
  wire [63:0] regs_43_io_out; // @[RegFile.scala 66:20:@35013.4]
  wire  regs_43_io_enable; // @[RegFile.scala 66:20:@35013.4]
  wire  regs_44_clock; // @[RegFile.scala 66:20:@35027.4]
  wire  regs_44_reset; // @[RegFile.scala 66:20:@35027.4]
  wire [63:0] regs_44_io_in; // @[RegFile.scala 66:20:@35027.4]
  wire  regs_44_io_reset; // @[RegFile.scala 66:20:@35027.4]
  wire [63:0] regs_44_io_out; // @[RegFile.scala 66:20:@35027.4]
  wire  regs_44_io_enable; // @[RegFile.scala 66:20:@35027.4]
  wire  regs_45_clock; // @[RegFile.scala 66:20:@35041.4]
  wire  regs_45_reset; // @[RegFile.scala 66:20:@35041.4]
  wire [63:0] regs_45_io_in; // @[RegFile.scala 66:20:@35041.4]
  wire  regs_45_io_reset; // @[RegFile.scala 66:20:@35041.4]
  wire [63:0] regs_45_io_out; // @[RegFile.scala 66:20:@35041.4]
  wire  regs_45_io_enable; // @[RegFile.scala 66:20:@35041.4]
  wire  regs_46_clock; // @[RegFile.scala 66:20:@35055.4]
  wire  regs_46_reset; // @[RegFile.scala 66:20:@35055.4]
  wire [63:0] regs_46_io_in; // @[RegFile.scala 66:20:@35055.4]
  wire  regs_46_io_reset; // @[RegFile.scala 66:20:@35055.4]
  wire [63:0] regs_46_io_out; // @[RegFile.scala 66:20:@35055.4]
  wire  regs_46_io_enable; // @[RegFile.scala 66:20:@35055.4]
  wire  regs_47_clock; // @[RegFile.scala 66:20:@35069.4]
  wire  regs_47_reset; // @[RegFile.scala 66:20:@35069.4]
  wire [63:0] regs_47_io_in; // @[RegFile.scala 66:20:@35069.4]
  wire  regs_47_io_reset; // @[RegFile.scala 66:20:@35069.4]
  wire [63:0] regs_47_io_out; // @[RegFile.scala 66:20:@35069.4]
  wire  regs_47_io_enable; // @[RegFile.scala 66:20:@35069.4]
  wire  regs_48_clock; // @[RegFile.scala 66:20:@35083.4]
  wire  regs_48_reset; // @[RegFile.scala 66:20:@35083.4]
  wire [63:0] regs_48_io_in; // @[RegFile.scala 66:20:@35083.4]
  wire  regs_48_io_reset; // @[RegFile.scala 66:20:@35083.4]
  wire [63:0] regs_48_io_out; // @[RegFile.scala 66:20:@35083.4]
  wire  regs_48_io_enable; // @[RegFile.scala 66:20:@35083.4]
  wire  regs_49_clock; // @[RegFile.scala 66:20:@35097.4]
  wire  regs_49_reset; // @[RegFile.scala 66:20:@35097.4]
  wire [63:0] regs_49_io_in; // @[RegFile.scala 66:20:@35097.4]
  wire  regs_49_io_reset; // @[RegFile.scala 66:20:@35097.4]
  wire [63:0] regs_49_io_out; // @[RegFile.scala 66:20:@35097.4]
  wire  regs_49_io_enable; // @[RegFile.scala 66:20:@35097.4]
  wire  regs_50_clock; // @[RegFile.scala 66:20:@35111.4]
  wire  regs_50_reset; // @[RegFile.scala 66:20:@35111.4]
  wire [63:0] regs_50_io_in; // @[RegFile.scala 66:20:@35111.4]
  wire  regs_50_io_reset; // @[RegFile.scala 66:20:@35111.4]
  wire [63:0] regs_50_io_out; // @[RegFile.scala 66:20:@35111.4]
  wire  regs_50_io_enable; // @[RegFile.scala 66:20:@35111.4]
  wire  regs_51_clock; // @[RegFile.scala 66:20:@35125.4]
  wire  regs_51_reset; // @[RegFile.scala 66:20:@35125.4]
  wire [63:0] regs_51_io_in; // @[RegFile.scala 66:20:@35125.4]
  wire  regs_51_io_reset; // @[RegFile.scala 66:20:@35125.4]
  wire [63:0] regs_51_io_out; // @[RegFile.scala 66:20:@35125.4]
  wire  regs_51_io_enable; // @[RegFile.scala 66:20:@35125.4]
  wire  regs_52_clock; // @[RegFile.scala 66:20:@35139.4]
  wire  regs_52_reset; // @[RegFile.scala 66:20:@35139.4]
  wire [63:0] regs_52_io_in; // @[RegFile.scala 66:20:@35139.4]
  wire  regs_52_io_reset; // @[RegFile.scala 66:20:@35139.4]
  wire [63:0] regs_52_io_out; // @[RegFile.scala 66:20:@35139.4]
  wire  regs_52_io_enable; // @[RegFile.scala 66:20:@35139.4]
  wire  regs_53_clock; // @[RegFile.scala 66:20:@35153.4]
  wire  regs_53_reset; // @[RegFile.scala 66:20:@35153.4]
  wire [63:0] regs_53_io_in; // @[RegFile.scala 66:20:@35153.4]
  wire  regs_53_io_reset; // @[RegFile.scala 66:20:@35153.4]
  wire [63:0] regs_53_io_out; // @[RegFile.scala 66:20:@35153.4]
  wire  regs_53_io_enable; // @[RegFile.scala 66:20:@35153.4]
  wire  regs_54_clock; // @[RegFile.scala 66:20:@35167.4]
  wire  regs_54_reset; // @[RegFile.scala 66:20:@35167.4]
  wire [63:0] regs_54_io_in; // @[RegFile.scala 66:20:@35167.4]
  wire  regs_54_io_reset; // @[RegFile.scala 66:20:@35167.4]
  wire [63:0] regs_54_io_out; // @[RegFile.scala 66:20:@35167.4]
  wire  regs_54_io_enable; // @[RegFile.scala 66:20:@35167.4]
  wire  regs_55_clock; // @[RegFile.scala 66:20:@35181.4]
  wire  regs_55_reset; // @[RegFile.scala 66:20:@35181.4]
  wire [63:0] regs_55_io_in; // @[RegFile.scala 66:20:@35181.4]
  wire  regs_55_io_reset; // @[RegFile.scala 66:20:@35181.4]
  wire [63:0] regs_55_io_out; // @[RegFile.scala 66:20:@35181.4]
  wire  regs_55_io_enable; // @[RegFile.scala 66:20:@35181.4]
  wire  regs_56_clock; // @[RegFile.scala 66:20:@35195.4]
  wire  regs_56_reset; // @[RegFile.scala 66:20:@35195.4]
  wire [63:0] regs_56_io_in; // @[RegFile.scala 66:20:@35195.4]
  wire  regs_56_io_reset; // @[RegFile.scala 66:20:@35195.4]
  wire [63:0] regs_56_io_out; // @[RegFile.scala 66:20:@35195.4]
  wire  regs_56_io_enable; // @[RegFile.scala 66:20:@35195.4]
  wire  regs_57_clock; // @[RegFile.scala 66:20:@35209.4]
  wire  regs_57_reset; // @[RegFile.scala 66:20:@35209.4]
  wire [63:0] regs_57_io_in; // @[RegFile.scala 66:20:@35209.4]
  wire  regs_57_io_reset; // @[RegFile.scala 66:20:@35209.4]
  wire [63:0] regs_57_io_out; // @[RegFile.scala 66:20:@35209.4]
  wire  regs_57_io_enable; // @[RegFile.scala 66:20:@35209.4]
  wire  regs_58_clock; // @[RegFile.scala 66:20:@35223.4]
  wire  regs_58_reset; // @[RegFile.scala 66:20:@35223.4]
  wire [63:0] regs_58_io_in; // @[RegFile.scala 66:20:@35223.4]
  wire  regs_58_io_reset; // @[RegFile.scala 66:20:@35223.4]
  wire [63:0] regs_58_io_out; // @[RegFile.scala 66:20:@35223.4]
  wire  regs_58_io_enable; // @[RegFile.scala 66:20:@35223.4]
  wire  regs_59_clock; // @[RegFile.scala 66:20:@35237.4]
  wire  regs_59_reset; // @[RegFile.scala 66:20:@35237.4]
  wire [63:0] regs_59_io_in; // @[RegFile.scala 66:20:@35237.4]
  wire  regs_59_io_reset; // @[RegFile.scala 66:20:@35237.4]
  wire [63:0] regs_59_io_out; // @[RegFile.scala 66:20:@35237.4]
  wire  regs_59_io_enable; // @[RegFile.scala 66:20:@35237.4]
  wire  regs_60_clock; // @[RegFile.scala 66:20:@35251.4]
  wire  regs_60_reset; // @[RegFile.scala 66:20:@35251.4]
  wire [63:0] regs_60_io_in; // @[RegFile.scala 66:20:@35251.4]
  wire  regs_60_io_reset; // @[RegFile.scala 66:20:@35251.4]
  wire [63:0] regs_60_io_out; // @[RegFile.scala 66:20:@35251.4]
  wire  regs_60_io_enable; // @[RegFile.scala 66:20:@35251.4]
  wire  regs_61_clock; // @[RegFile.scala 66:20:@35265.4]
  wire  regs_61_reset; // @[RegFile.scala 66:20:@35265.4]
  wire [63:0] regs_61_io_in; // @[RegFile.scala 66:20:@35265.4]
  wire  regs_61_io_reset; // @[RegFile.scala 66:20:@35265.4]
  wire [63:0] regs_61_io_out; // @[RegFile.scala 66:20:@35265.4]
  wire  regs_61_io_enable; // @[RegFile.scala 66:20:@35265.4]
  wire  regs_62_clock; // @[RegFile.scala 66:20:@35279.4]
  wire  regs_62_reset; // @[RegFile.scala 66:20:@35279.4]
  wire [63:0] regs_62_io_in; // @[RegFile.scala 66:20:@35279.4]
  wire  regs_62_io_reset; // @[RegFile.scala 66:20:@35279.4]
  wire [63:0] regs_62_io_out; // @[RegFile.scala 66:20:@35279.4]
  wire  regs_62_io_enable; // @[RegFile.scala 66:20:@35279.4]
  wire  regs_63_clock; // @[RegFile.scala 66:20:@35293.4]
  wire  regs_63_reset; // @[RegFile.scala 66:20:@35293.4]
  wire [63:0] regs_63_io_in; // @[RegFile.scala 66:20:@35293.4]
  wire  regs_63_io_reset; // @[RegFile.scala 66:20:@35293.4]
  wire [63:0] regs_63_io_out; // @[RegFile.scala 66:20:@35293.4]
  wire  regs_63_io_enable; // @[RegFile.scala 66:20:@35293.4]
  wire  regs_64_clock; // @[RegFile.scala 66:20:@35307.4]
  wire  regs_64_reset; // @[RegFile.scala 66:20:@35307.4]
  wire [63:0] regs_64_io_in; // @[RegFile.scala 66:20:@35307.4]
  wire  regs_64_io_reset; // @[RegFile.scala 66:20:@35307.4]
  wire [63:0] regs_64_io_out; // @[RegFile.scala 66:20:@35307.4]
  wire  regs_64_io_enable; // @[RegFile.scala 66:20:@35307.4]
  wire  regs_65_clock; // @[RegFile.scala 66:20:@35321.4]
  wire  regs_65_reset; // @[RegFile.scala 66:20:@35321.4]
  wire [63:0] regs_65_io_in; // @[RegFile.scala 66:20:@35321.4]
  wire  regs_65_io_reset; // @[RegFile.scala 66:20:@35321.4]
  wire [63:0] regs_65_io_out; // @[RegFile.scala 66:20:@35321.4]
  wire  regs_65_io_enable; // @[RegFile.scala 66:20:@35321.4]
  wire  regs_66_clock; // @[RegFile.scala 66:20:@35335.4]
  wire  regs_66_reset; // @[RegFile.scala 66:20:@35335.4]
  wire [63:0] regs_66_io_in; // @[RegFile.scala 66:20:@35335.4]
  wire  regs_66_io_reset; // @[RegFile.scala 66:20:@35335.4]
  wire [63:0] regs_66_io_out; // @[RegFile.scala 66:20:@35335.4]
  wire  regs_66_io_enable; // @[RegFile.scala 66:20:@35335.4]
  wire  regs_67_clock; // @[RegFile.scala 66:20:@35349.4]
  wire  regs_67_reset; // @[RegFile.scala 66:20:@35349.4]
  wire [63:0] regs_67_io_in; // @[RegFile.scala 66:20:@35349.4]
  wire  regs_67_io_reset; // @[RegFile.scala 66:20:@35349.4]
  wire [63:0] regs_67_io_out; // @[RegFile.scala 66:20:@35349.4]
  wire  regs_67_io_enable; // @[RegFile.scala 66:20:@35349.4]
  wire  regs_68_clock; // @[RegFile.scala 66:20:@35363.4]
  wire  regs_68_reset; // @[RegFile.scala 66:20:@35363.4]
  wire [63:0] regs_68_io_in; // @[RegFile.scala 66:20:@35363.4]
  wire  regs_68_io_reset; // @[RegFile.scala 66:20:@35363.4]
  wire [63:0] regs_68_io_out; // @[RegFile.scala 66:20:@35363.4]
  wire  regs_68_io_enable; // @[RegFile.scala 66:20:@35363.4]
  wire  regs_69_clock; // @[RegFile.scala 66:20:@35377.4]
  wire  regs_69_reset; // @[RegFile.scala 66:20:@35377.4]
  wire [63:0] regs_69_io_in; // @[RegFile.scala 66:20:@35377.4]
  wire  regs_69_io_reset; // @[RegFile.scala 66:20:@35377.4]
  wire [63:0] regs_69_io_out; // @[RegFile.scala 66:20:@35377.4]
  wire  regs_69_io_enable; // @[RegFile.scala 66:20:@35377.4]
  wire  regs_70_clock; // @[RegFile.scala 66:20:@35391.4]
  wire  regs_70_reset; // @[RegFile.scala 66:20:@35391.4]
  wire [63:0] regs_70_io_in; // @[RegFile.scala 66:20:@35391.4]
  wire  regs_70_io_reset; // @[RegFile.scala 66:20:@35391.4]
  wire [63:0] regs_70_io_out; // @[RegFile.scala 66:20:@35391.4]
  wire  regs_70_io_enable; // @[RegFile.scala 66:20:@35391.4]
  wire  regs_71_clock; // @[RegFile.scala 66:20:@35405.4]
  wire  regs_71_reset; // @[RegFile.scala 66:20:@35405.4]
  wire [63:0] regs_71_io_in; // @[RegFile.scala 66:20:@35405.4]
  wire  regs_71_io_reset; // @[RegFile.scala 66:20:@35405.4]
  wire [63:0] regs_71_io_out; // @[RegFile.scala 66:20:@35405.4]
  wire  regs_71_io_enable; // @[RegFile.scala 66:20:@35405.4]
  wire  regs_72_clock; // @[RegFile.scala 66:20:@35419.4]
  wire  regs_72_reset; // @[RegFile.scala 66:20:@35419.4]
  wire [63:0] regs_72_io_in; // @[RegFile.scala 66:20:@35419.4]
  wire  regs_72_io_reset; // @[RegFile.scala 66:20:@35419.4]
  wire [63:0] regs_72_io_out; // @[RegFile.scala 66:20:@35419.4]
  wire  regs_72_io_enable; // @[RegFile.scala 66:20:@35419.4]
  wire  regs_73_clock; // @[RegFile.scala 66:20:@35433.4]
  wire  regs_73_reset; // @[RegFile.scala 66:20:@35433.4]
  wire [63:0] regs_73_io_in; // @[RegFile.scala 66:20:@35433.4]
  wire  regs_73_io_reset; // @[RegFile.scala 66:20:@35433.4]
  wire [63:0] regs_73_io_out; // @[RegFile.scala 66:20:@35433.4]
  wire  regs_73_io_enable; // @[RegFile.scala 66:20:@35433.4]
  wire  regs_74_clock; // @[RegFile.scala 66:20:@35447.4]
  wire  regs_74_reset; // @[RegFile.scala 66:20:@35447.4]
  wire [63:0] regs_74_io_in; // @[RegFile.scala 66:20:@35447.4]
  wire  regs_74_io_reset; // @[RegFile.scala 66:20:@35447.4]
  wire [63:0] regs_74_io_out; // @[RegFile.scala 66:20:@35447.4]
  wire  regs_74_io_enable; // @[RegFile.scala 66:20:@35447.4]
  wire  regs_75_clock; // @[RegFile.scala 66:20:@35461.4]
  wire  regs_75_reset; // @[RegFile.scala 66:20:@35461.4]
  wire [63:0] regs_75_io_in; // @[RegFile.scala 66:20:@35461.4]
  wire  regs_75_io_reset; // @[RegFile.scala 66:20:@35461.4]
  wire [63:0] regs_75_io_out; // @[RegFile.scala 66:20:@35461.4]
  wire  regs_75_io_enable; // @[RegFile.scala 66:20:@35461.4]
  wire  regs_76_clock; // @[RegFile.scala 66:20:@35475.4]
  wire  regs_76_reset; // @[RegFile.scala 66:20:@35475.4]
  wire [63:0] regs_76_io_in; // @[RegFile.scala 66:20:@35475.4]
  wire  regs_76_io_reset; // @[RegFile.scala 66:20:@35475.4]
  wire [63:0] regs_76_io_out; // @[RegFile.scala 66:20:@35475.4]
  wire  regs_76_io_enable; // @[RegFile.scala 66:20:@35475.4]
  wire  regs_77_clock; // @[RegFile.scala 66:20:@35489.4]
  wire  regs_77_reset; // @[RegFile.scala 66:20:@35489.4]
  wire [63:0] regs_77_io_in; // @[RegFile.scala 66:20:@35489.4]
  wire  regs_77_io_reset; // @[RegFile.scala 66:20:@35489.4]
  wire [63:0] regs_77_io_out; // @[RegFile.scala 66:20:@35489.4]
  wire  regs_77_io_enable; // @[RegFile.scala 66:20:@35489.4]
  wire  regs_78_clock; // @[RegFile.scala 66:20:@35503.4]
  wire  regs_78_reset; // @[RegFile.scala 66:20:@35503.4]
  wire [63:0] regs_78_io_in; // @[RegFile.scala 66:20:@35503.4]
  wire  regs_78_io_reset; // @[RegFile.scala 66:20:@35503.4]
  wire [63:0] regs_78_io_out; // @[RegFile.scala 66:20:@35503.4]
  wire  regs_78_io_enable; // @[RegFile.scala 66:20:@35503.4]
  wire  regs_79_clock; // @[RegFile.scala 66:20:@35517.4]
  wire  regs_79_reset; // @[RegFile.scala 66:20:@35517.4]
  wire [63:0] regs_79_io_in; // @[RegFile.scala 66:20:@35517.4]
  wire  regs_79_io_reset; // @[RegFile.scala 66:20:@35517.4]
  wire [63:0] regs_79_io_out; // @[RegFile.scala 66:20:@35517.4]
  wire  regs_79_io_enable; // @[RegFile.scala 66:20:@35517.4]
  wire  regs_80_clock; // @[RegFile.scala 66:20:@35531.4]
  wire  regs_80_reset; // @[RegFile.scala 66:20:@35531.4]
  wire [63:0] regs_80_io_in; // @[RegFile.scala 66:20:@35531.4]
  wire  regs_80_io_reset; // @[RegFile.scala 66:20:@35531.4]
  wire [63:0] regs_80_io_out; // @[RegFile.scala 66:20:@35531.4]
  wire  regs_80_io_enable; // @[RegFile.scala 66:20:@35531.4]
  wire  regs_81_clock; // @[RegFile.scala 66:20:@35545.4]
  wire  regs_81_reset; // @[RegFile.scala 66:20:@35545.4]
  wire [63:0] regs_81_io_in; // @[RegFile.scala 66:20:@35545.4]
  wire  regs_81_io_reset; // @[RegFile.scala 66:20:@35545.4]
  wire [63:0] regs_81_io_out; // @[RegFile.scala 66:20:@35545.4]
  wire  regs_81_io_enable; // @[RegFile.scala 66:20:@35545.4]
  wire  regs_82_clock; // @[RegFile.scala 66:20:@35559.4]
  wire  regs_82_reset; // @[RegFile.scala 66:20:@35559.4]
  wire [63:0] regs_82_io_in; // @[RegFile.scala 66:20:@35559.4]
  wire  regs_82_io_reset; // @[RegFile.scala 66:20:@35559.4]
  wire [63:0] regs_82_io_out; // @[RegFile.scala 66:20:@35559.4]
  wire  regs_82_io_enable; // @[RegFile.scala 66:20:@35559.4]
  wire  regs_83_clock; // @[RegFile.scala 66:20:@35573.4]
  wire  regs_83_reset; // @[RegFile.scala 66:20:@35573.4]
  wire [63:0] regs_83_io_in; // @[RegFile.scala 66:20:@35573.4]
  wire  regs_83_io_reset; // @[RegFile.scala 66:20:@35573.4]
  wire [63:0] regs_83_io_out; // @[RegFile.scala 66:20:@35573.4]
  wire  regs_83_io_enable; // @[RegFile.scala 66:20:@35573.4]
  wire  regs_84_clock; // @[RegFile.scala 66:20:@35587.4]
  wire  regs_84_reset; // @[RegFile.scala 66:20:@35587.4]
  wire [63:0] regs_84_io_in; // @[RegFile.scala 66:20:@35587.4]
  wire  regs_84_io_reset; // @[RegFile.scala 66:20:@35587.4]
  wire [63:0] regs_84_io_out; // @[RegFile.scala 66:20:@35587.4]
  wire  regs_84_io_enable; // @[RegFile.scala 66:20:@35587.4]
  wire  regs_85_clock; // @[RegFile.scala 66:20:@35601.4]
  wire  regs_85_reset; // @[RegFile.scala 66:20:@35601.4]
  wire [63:0] regs_85_io_in; // @[RegFile.scala 66:20:@35601.4]
  wire  regs_85_io_reset; // @[RegFile.scala 66:20:@35601.4]
  wire [63:0] regs_85_io_out; // @[RegFile.scala 66:20:@35601.4]
  wire  regs_85_io_enable; // @[RegFile.scala 66:20:@35601.4]
  wire  regs_86_clock; // @[RegFile.scala 66:20:@35615.4]
  wire  regs_86_reset; // @[RegFile.scala 66:20:@35615.4]
  wire [63:0] regs_86_io_in; // @[RegFile.scala 66:20:@35615.4]
  wire  regs_86_io_reset; // @[RegFile.scala 66:20:@35615.4]
  wire [63:0] regs_86_io_out; // @[RegFile.scala 66:20:@35615.4]
  wire  regs_86_io_enable; // @[RegFile.scala 66:20:@35615.4]
  wire  regs_87_clock; // @[RegFile.scala 66:20:@35629.4]
  wire  regs_87_reset; // @[RegFile.scala 66:20:@35629.4]
  wire [63:0] regs_87_io_in; // @[RegFile.scala 66:20:@35629.4]
  wire  regs_87_io_reset; // @[RegFile.scala 66:20:@35629.4]
  wire [63:0] regs_87_io_out; // @[RegFile.scala 66:20:@35629.4]
  wire  regs_87_io_enable; // @[RegFile.scala 66:20:@35629.4]
  wire  regs_88_clock; // @[RegFile.scala 66:20:@35643.4]
  wire  regs_88_reset; // @[RegFile.scala 66:20:@35643.4]
  wire [63:0] regs_88_io_in; // @[RegFile.scala 66:20:@35643.4]
  wire  regs_88_io_reset; // @[RegFile.scala 66:20:@35643.4]
  wire [63:0] regs_88_io_out; // @[RegFile.scala 66:20:@35643.4]
  wire  regs_88_io_enable; // @[RegFile.scala 66:20:@35643.4]
  wire  regs_89_clock; // @[RegFile.scala 66:20:@35657.4]
  wire  regs_89_reset; // @[RegFile.scala 66:20:@35657.4]
  wire [63:0] regs_89_io_in; // @[RegFile.scala 66:20:@35657.4]
  wire  regs_89_io_reset; // @[RegFile.scala 66:20:@35657.4]
  wire [63:0] regs_89_io_out; // @[RegFile.scala 66:20:@35657.4]
  wire  regs_89_io_enable; // @[RegFile.scala 66:20:@35657.4]
  wire  regs_90_clock; // @[RegFile.scala 66:20:@35671.4]
  wire  regs_90_reset; // @[RegFile.scala 66:20:@35671.4]
  wire [63:0] regs_90_io_in; // @[RegFile.scala 66:20:@35671.4]
  wire  regs_90_io_reset; // @[RegFile.scala 66:20:@35671.4]
  wire [63:0] regs_90_io_out; // @[RegFile.scala 66:20:@35671.4]
  wire  regs_90_io_enable; // @[RegFile.scala 66:20:@35671.4]
  wire  regs_91_clock; // @[RegFile.scala 66:20:@35685.4]
  wire  regs_91_reset; // @[RegFile.scala 66:20:@35685.4]
  wire [63:0] regs_91_io_in; // @[RegFile.scala 66:20:@35685.4]
  wire  regs_91_io_reset; // @[RegFile.scala 66:20:@35685.4]
  wire [63:0] regs_91_io_out; // @[RegFile.scala 66:20:@35685.4]
  wire  regs_91_io_enable; // @[RegFile.scala 66:20:@35685.4]
  wire  regs_92_clock; // @[RegFile.scala 66:20:@35699.4]
  wire  regs_92_reset; // @[RegFile.scala 66:20:@35699.4]
  wire [63:0] regs_92_io_in; // @[RegFile.scala 66:20:@35699.4]
  wire  regs_92_io_reset; // @[RegFile.scala 66:20:@35699.4]
  wire [63:0] regs_92_io_out; // @[RegFile.scala 66:20:@35699.4]
  wire  regs_92_io_enable; // @[RegFile.scala 66:20:@35699.4]
  wire  regs_93_clock; // @[RegFile.scala 66:20:@35713.4]
  wire  regs_93_reset; // @[RegFile.scala 66:20:@35713.4]
  wire [63:0] regs_93_io_in; // @[RegFile.scala 66:20:@35713.4]
  wire  regs_93_io_reset; // @[RegFile.scala 66:20:@35713.4]
  wire [63:0] regs_93_io_out; // @[RegFile.scala 66:20:@35713.4]
  wire  regs_93_io_enable; // @[RegFile.scala 66:20:@35713.4]
  wire  regs_94_clock; // @[RegFile.scala 66:20:@35727.4]
  wire  regs_94_reset; // @[RegFile.scala 66:20:@35727.4]
  wire [63:0] regs_94_io_in; // @[RegFile.scala 66:20:@35727.4]
  wire  regs_94_io_reset; // @[RegFile.scala 66:20:@35727.4]
  wire [63:0] regs_94_io_out; // @[RegFile.scala 66:20:@35727.4]
  wire  regs_94_io_enable; // @[RegFile.scala 66:20:@35727.4]
  wire  regs_95_clock; // @[RegFile.scala 66:20:@35741.4]
  wire  regs_95_reset; // @[RegFile.scala 66:20:@35741.4]
  wire [63:0] regs_95_io_in; // @[RegFile.scala 66:20:@35741.4]
  wire  regs_95_io_reset; // @[RegFile.scala 66:20:@35741.4]
  wire [63:0] regs_95_io_out; // @[RegFile.scala 66:20:@35741.4]
  wire  regs_95_io_enable; // @[RegFile.scala 66:20:@35741.4]
  wire  regs_96_clock; // @[RegFile.scala 66:20:@35755.4]
  wire  regs_96_reset; // @[RegFile.scala 66:20:@35755.4]
  wire [63:0] regs_96_io_in; // @[RegFile.scala 66:20:@35755.4]
  wire  regs_96_io_reset; // @[RegFile.scala 66:20:@35755.4]
  wire [63:0] regs_96_io_out; // @[RegFile.scala 66:20:@35755.4]
  wire  regs_96_io_enable; // @[RegFile.scala 66:20:@35755.4]
  wire  regs_97_clock; // @[RegFile.scala 66:20:@35769.4]
  wire  regs_97_reset; // @[RegFile.scala 66:20:@35769.4]
  wire [63:0] regs_97_io_in; // @[RegFile.scala 66:20:@35769.4]
  wire  regs_97_io_reset; // @[RegFile.scala 66:20:@35769.4]
  wire [63:0] regs_97_io_out; // @[RegFile.scala 66:20:@35769.4]
  wire  regs_97_io_enable; // @[RegFile.scala 66:20:@35769.4]
  wire  regs_98_clock; // @[RegFile.scala 66:20:@35783.4]
  wire  regs_98_reset; // @[RegFile.scala 66:20:@35783.4]
  wire [63:0] regs_98_io_in; // @[RegFile.scala 66:20:@35783.4]
  wire  regs_98_io_reset; // @[RegFile.scala 66:20:@35783.4]
  wire [63:0] regs_98_io_out; // @[RegFile.scala 66:20:@35783.4]
  wire  regs_98_io_enable; // @[RegFile.scala 66:20:@35783.4]
  wire  regs_99_clock; // @[RegFile.scala 66:20:@35797.4]
  wire  regs_99_reset; // @[RegFile.scala 66:20:@35797.4]
  wire [63:0] regs_99_io_in; // @[RegFile.scala 66:20:@35797.4]
  wire  regs_99_io_reset; // @[RegFile.scala 66:20:@35797.4]
  wire [63:0] regs_99_io_out; // @[RegFile.scala 66:20:@35797.4]
  wire  regs_99_io_enable; // @[RegFile.scala 66:20:@35797.4]
  wire  regs_100_clock; // @[RegFile.scala 66:20:@35811.4]
  wire  regs_100_reset; // @[RegFile.scala 66:20:@35811.4]
  wire [63:0] regs_100_io_in; // @[RegFile.scala 66:20:@35811.4]
  wire  regs_100_io_reset; // @[RegFile.scala 66:20:@35811.4]
  wire [63:0] regs_100_io_out; // @[RegFile.scala 66:20:@35811.4]
  wire  regs_100_io_enable; // @[RegFile.scala 66:20:@35811.4]
  wire  regs_101_clock; // @[RegFile.scala 66:20:@35825.4]
  wire  regs_101_reset; // @[RegFile.scala 66:20:@35825.4]
  wire [63:0] regs_101_io_in; // @[RegFile.scala 66:20:@35825.4]
  wire  regs_101_io_reset; // @[RegFile.scala 66:20:@35825.4]
  wire [63:0] regs_101_io_out; // @[RegFile.scala 66:20:@35825.4]
  wire  regs_101_io_enable; // @[RegFile.scala 66:20:@35825.4]
  wire  regs_102_clock; // @[RegFile.scala 66:20:@35839.4]
  wire  regs_102_reset; // @[RegFile.scala 66:20:@35839.4]
  wire [63:0] regs_102_io_in; // @[RegFile.scala 66:20:@35839.4]
  wire  regs_102_io_reset; // @[RegFile.scala 66:20:@35839.4]
  wire [63:0] regs_102_io_out; // @[RegFile.scala 66:20:@35839.4]
  wire  regs_102_io_enable; // @[RegFile.scala 66:20:@35839.4]
  wire  regs_103_clock; // @[RegFile.scala 66:20:@35853.4]
  wire  regs_103_reset; // @[RegFile.scala 66:20:@35853.4]
  wire [63:0] regs_103_io_in; // @[RegFile.scala 66:20:@35853.4]
  wire  regs_103_io_reset; // @[RegFile.scala 66:20:@35853.4]
  wire [63:0] regs_103_io_out; // @[RegFile.scala 66:20:@35853.4]
  wire  regs_103_io_enable; // @[RegFile.scala 66:20:@35853.4]
  wire  regs_104_clock; // @[RegFile.scala 66:20:@35867.4]
  wire  regs_104_reset; // @[RegFile.scala 66:20:@35867.4]
  wire [63:0] regs_104_io_in; // @[RegFile.scala 66:20:@35867.4]
  wire  regs_104_io_reset; // @[RegFile.scala 66:20:@35867.4]
  wire [63:0] regs_104_io_out; // @[RegFile.scala 66:20:@35867.4]
  wire  regs_104_io_enable; // @[RegFile.scala 66:20:@35867.4]
  wire  regs_105_clock; // @[RegFile.scala 66:20:@35881.4]
  wire  regs_105_reset; // @[RegFile.scala 66:20:@35881.4]
  wire [63:0] regs_105_io_in; // @[RegFile.scala 66:20:@35881.4]
  wire  regs_105_io_reset; // @[RegFile.scala 66:20:@35881.4]
  wire [63:0] regs_105_io_out; // @[RegFile.scala 66:20:@35881.4]
  wire  regs_105_io_enable; // @[RegFile.scala 66:20:@35881.4]
  wire  regs_106_clock; // @[RegFile.scala 66:20:@35895.4]
  wire  regs_106_reset; // @[RegFile.scala 66:20:@35895.4]
  wire [63:0] regs_106_io_in; // @[RegFile.scala 66:20:@35895.4]
  wire  regs_106_io_reset; // @[RegFile.scala 66:20:@35895.4]
  wire [63:0] regs_106_io_out; // @[RegFile.scala 66:20:@35895.4]
  wire  regs_106_io_enable; // @[RegFile.scala 66:20:@35895.4]
  wire  regs_107_clock; // @[RegFile.scala 66:20:@35909.4]
  wire  regs_107_reset; // @[RegFile.scala 66:20:@35909.4]
  wire [63:0] regs_107_io_in; // @[RegFile.scala 66:20:@35909.4]
  wire  regs_107_io_reset; // @[RegFile.scala 66:20:@35909.4]
  wire [63:0] regs_107_io_out; // @[RegFile.scala 66:20:@35909.4]
  wire  regs_107_io_enable; // @[RegFile.scala 66:20:@35909.4]
  wire  regs_108_clock; // @[RegFile.scala 66:20:@35923.4]
  wire  regs_108_reset; // @[RegFile.scala 66:20:@35923.4]
  wire [63:0] regs_108_io_in; // @[RegFile.scala 66:20:@35923.4]
  wire  regs_108_io_reset; // @[RegFile.scala 66:20:@35923.4]
  wire [63:0] regs_108_io_out; // @[RegFile.scala 66:20:@35923.4]
  wire  regs_108_io_enable; // @[RegFile.scala 66:20:@35923.4]
  wire  regs_109_clock; // @[RegFile.scala 66:20:@35937.4]
  wire  regs_109_reset; // @[RegFile.scala 66:20:@35937.4]
  wire [63:0] regs_109_io_in; // @[RegFile.scala 66:20:@35937.4]
  wire  regs_109_io_reset; // @[RegFile.scala 66:20:@35937.4]
  wire [63:0] regs_109_io_out; // @[RegFile.scala 66:20:@35937.4]
  wire  regs_109_io_enable; // @[RegFile.scala 66:20:@35937.4]
  wire  regs_110_clock; // @[RegFile.scala 66:20:@35951.4]
  wire  regs_110_reset; // @[RegFile.scala 66:20:@35951.4]
  wire [63:0] regs_110_io_in; // @[RegFile.scala 66:20:@35951.4]
  wire  regs_110_io_reset; // @[RegFile.scala 66:20:@35951.4]
  wire [63:0] regs_110_io_out; // @[RegFile.scala 66:20:@35951.4]
  wire  regs_110_io_enable; // @[RegFile.scala 66:20:@35951.4]
  wire  regs_111_clock; // @[RegFile.scala 66:20:@35965.4]
  wire  regs_111_reset; // @[RegFile.scala 66:20:@35965.4]
  wire [63:0] regs_111_io_in; // @[RegFile.scala 66:20:@35965.4]
  wire  regs_111_io_reset; // @[RegFile.scala 66:20:@35965.4]
  wire [63:0] regs_111_io_out; // @[RegFile.scala 66:20:@35965.4]
  wire  regs_111_io_enable; // @[RegFile.scala 66:20:@35965.4]
  wire  regs_112_clock; // @[RegFile.scala 66:20:@35979.4]
  wire  regs_112_reset; // @[RegFile.scala 66:20:@35979.4]
  wire [63:0] regs_112_io_in; // @[RegFile.scala 66:20:@35979.4]
  wire  regs_112_io_reset; // @[RegFile.scala 66:20:@35979.4]
  wire [63:0] regs_112_io_out; // @[RegFile.scala 66:20:@35979.4]
  wire  regs_112_io_enable; // @[RegFile.scala 66:20:@35979.4]
  wire  regs_113_clock; // @[RegFile.scala 66:20:@35993.4]
  wire  regs_113_reset; // @[RegFile.scala 66:20:@35993.4]
  wire [63:0] regs_113_io_in; // @[RegFile.scala 66:20:@35993.4]
  wire  regs_113_io_reset; // @[RegFile.scala 66:20:@35993.4]
  wire [63:0] regs_113_io_out; // @[RegFile.scala 66:20:@35993.4]
  wire  regs_113_io_enable; // @[RegFile.scala 66:20:@35993.4]
  wire  regs_114_clock; // @[RegFile.scala 66:20:@36007.4]
  wire  regs_114_reset; // @[RegFile.scala 66:20:@36007.4]
  wire [63:0] regs_114_io_in; // @[RegFile.scala 66:20:@36007.4]
  wire  regs_114_io_reset; // @[RegFile.scala 66:20:@36007.4]
  wire [63:0] regs_114_io_out; // @[RegFile.scala 66:20:@36007.4]
  wire  regs_114_io_enable; // @[RegFile.scala 66:20:@36007.4]
  wire  regs_115_clock; // @[RegFile.scala 66:20:@36021.4]
  wire  regs_115_reset; // @[RegFile.scala 66:20:@36021.4]
  wire [63:0] regs_115_io_in; // @[RegFile.scala 66:20:@36021.4]
  wire  regs_115_io_reset; // @[RegFile.scala 66:20:@36021.4]
  wire [63:0] regs_115_io_out; // @[RegFile.scala 66:20:@36021.4]
  wire  regs_115_io_enable; // @[RegFile.scala 66:20:@36021.4]
  wire  regs_116_clock; // @[RegFile.scala 66:20:@36035.4]
  wire  regs_116_reset; // @[RegFile.scala 66:20:@36035.4]
  wire [63:0] regs_116_io_in; // @[RegFile.scala 66:20:@36035.4]
  wire  regs_116_io_reset; // @[RegFile.scala 66:20:@36035.4]
  wire [63:0] regs_116_io_out; // @[RegFile.scala 66:20:@36035.4]
  wire  regs_116_io_enable; // @[RegFile.scala 66:20:@36035.4]
  wire  regs_117_clock; // @[RegFile.scala 66:20:@36049.4]
  wire  regs_117_reset; // @[RegFile.scala 66:20:@36049.4]
  wire [63:0] regs_117_io_in; // @[RegFile.scala 66:20:@36049.4]
  wire  regs_117_io_reset; // @[RegFile.scala 66:20:@36049.4]
  wire [63:0] regs_117_io_out; // @[RegFile.scala 66:20:@36049.4]
  wire  regs_117_io_enable; // @[RegFile.scala 66:20:@36049.4]
  wire  regs_118_clock; // @[RegFile.scala 66:20:@36063.4]
  wire  regs_118_reset; // @[RegFile.scala 66:20:@36063.4]
  wire [63:0] regs_118_io_in; // @[RegFile.scala 66:20:@36063.4]
  wire  regs_118_io_reset; // @[RegFile.scala 66:20:@36063.4]
  wire [63:0] regs_118_io_out; // @[RegFile.scala 66:20:@36063.4]
  wire  regs_118_io_enable; // @[RegFile.scala 66:20:@36063.4]
  wire  regs_119_clock; // @[RegFile.scala 66:20:@36077.4]
  wire  regs_119_reset; // @[RegFile.scala 66:20:@36077.4]
  wire [63:0] regs_119_io_in; // @[RegFile.scala 66:20:@36077.4]
  wire  regs_119_io_reset; // @[RegFile.scala 66:20:@36077.4]
  wire [63:0] regs_119_io_out; // @[RegFile.scala 66:20:@36077.4]
  wire  regs_119_io_enable; // @[RegFile.scala 66:20:@36077.4]
  wire  regs_120_clock; // @[RegFile.scala 66:20:@36091.4]
  wire  regs_120_reset; // @[RegFile.scala 66:20:@36091.4]
  wire [63:0] regs_120_io_in; // @[RegFile.scala 66:20:@36091.4]
  wire  regs_120_io_reset; // @[RegFile.scala 66:20:@36091.4]
  wire [63:0] regs_120_io_out; // @[RegFile.scala 66:20:@36091.4]
  wire  regs_120_io_enable; // @[RegFile.scala 66:20:@36091.4]
  wire  regs_121_clock; // @[RegFile.scala 66:20:@36105.4]
  wire  regs_121_reset; // @[RegFile.scala 66:20:@36105.4]
  wire [63:0] regs_121_io_in; // @[RegFile.scala 66:20:@36105.4]
  wire  regs_121_io_reset; // @[RegFile.scala 66:20:@36105.4]
  wire [63:0] regs_121_io_out; // @[RegFile.scala 66:20:@36105.4]
  wire  regs_121_io_enable; // @[RegFile.scala 66:20:@36105.4]
  wire  regs_122_clock; // @[RegFile.scala 66:20:@36119.4]
  wire  regs_122_reset; // @[RegFile.scala 66:20:@36119.4]
  wire [63:0] regs_122_io_in; // @[RegFile.scala 66:20:@36119.4]
  wire  regs_122_io_reset; // @[RegFile.scala 66:20:@36119.4]
  wire [63:0] regs_122_io_out; // @[RegFile.scala 66:20:@36119.4]
  wire  regs_122_io_enable; // @[RegFile.scala 66:20:@36119.4]
  wire  regs_123_clock; // @[RegFile.scala 66:20:@36133.4]
  wire  regs_123_reset; // @[RegFile.scala 66:20:@36133.4]
  wire [63:0] regs_123_io_in; // @[RegFile.scala 66:20:@36133.4]
  wire  regs_123_io_reset; // @[RegFile.scala 66:20:@36133.4]
  wire [63:0] regs_123_io_out; // @[RegFile.scala 66:20:@36133.4]
  wire  regs_123_io_enable; // @[RegFile.scala 66:20:@36133.4]
  wire  regs_124_clock; // @[RegFile.scala 66:20:@36147.4]
  wire  regs_124_reset; // @[RegFile.scala 66:20:@36147.4]
  wire [63:0] regs_124_io_in; // @[RegFile.scala 66:20:@36147.4]
  wire  regs_124_io_reset; // @[RegFile.scala 66:20:@36147.4]
  wire [63:0] regs_124_io_out; // @[RegFile.scala 66:20:@36147.4]
  wire  regs_124_io_enable; // @[RegFile.scala 66:20:@36147.4]
  wire  regs_125_clock; // @[RegFile.scala 66:20:@36161.4]
  wire  regs_125_reset; // @[RegFile.scala 66:20:@36161.4]
  wire [63:0] regs_125_io_in; // @[RegFile.scala 66:20:@36161.4]
  wire  regs_125_io_reset; // @[RegFile.scala 66:20:@36161.4]
  wire [63:0] regs_125_io_out; // @[RegFile.scala 66:20:@36161.4]
  wire  regs_125_io_enable; // @[RegFile.scala 66:20:@36161.4]
  wire  regs_126_clock; // @[RegFile.scala 66:20:@36175.4]
  wire  regs_126_reset; // @[RegFile.scala 66:20:@36175.4]
  wire [63:0] regs_126_io_in; // @[RegFile.scala 66:20:@36175.4]
  wire  regs_126_io_reset; // @[RegFile.scala 66:20:@36175.4]
  wire [63:0] regs_126_io_out; // @[RegFile.scala 66:20:@36175.4]
  wire  regs_126_io_enable; // @[RegFile.scala 66:20:@36175.4]
  wire  regs_127_clock; // @[RegFile.scala 66:20:@36189.4]
  wire  regs_127_reset; // @[RegFile.scala 66:20:@36189.4]
  wire [63:0] regs_127_io_in; // @[RegFile.scala 66:20:@36189.4]
  wire  regs_127_io_reset; // @[RegFile.scala 66:20:@36189.4]
  wire [63:0] regs_127_io_out; // @[RegFile.scala 66:20:@36189.4]
  wire  regs_127_io_enable; // @[RegFile.scala 66:20:@36189.4]
  wire  regs_128_clock; // @[RegFile.scala 66:20:@36203.4]
  wire  regs_128_reset; // @[RegFile.scala 66:20:@36203.4]
  wire [63:0] regs_128_io_in; // @[RegFile.scala 66:20:@36203.4]
  wire  regs_128_io_reset; // @[RegFile.scala 66:20:@36203.4]
  wire [63:0] regs_128_io_out; // @[RegFile.scala 66:20:@36203.4]
  wire  regs_128_io_enable; // @[RegFile.scala 66:20:@36203.4]
  wire  regs_129_clock; // @[RegFile.scala 66:20:@36217.4]
  wire  regs_129_reset; // @[RegFile.scala 66:20:@36217.4]
  wire [63:0] regs_129_io_in; // @[RegFile.scala 66:20:@36217.4]
  wire  regs_129_io_reset; // @[RegFile.scala 66:20:@36217.4]
  wire [63:0] regs_129_io_out; // @[RegFile.scala 66:20:@36217.4]
  wire  regs_129_io_enable; // @[RegFile.scala 66:20:@36217.4]
  wire  regs_130_clock; // @[RegFile.scala 66:20:@36231.4]
  wire  regs_130_reset; // @[RegFile.scala 66:20:@36231.4]
  wire [63:0] regs_130_io_in; // @[RegFile.scala 66:20:@36231.4]
  wire  regs_130_io_reset; // @[RegFile.scala 66:20:@36231.4]
  wire [63:0] regs_130_io_out; // @[RegFile.scala 66:20:@36231.4]
  wire  regs_130_io_enable; // @[RegFile.scala 66:20:@36231.4]
  wire  regs_131_clock; // @[RegFile.scala 66:20:@36245.4]
  wire  regs_131_reset; // @[RegFile.scala 66:20:@36245.4]
  wire [63:0] regs_131_io_in; // @[RegFile.scala 66:20:@36245.4]
  wire  regs_131_io_reset; // @[RegFile.scala 66:20:@36245.4]
  wire [63:0] regs_131_io_out; // @[RegFile.scala 66:20:@36245.4]
  wire  regs_131_io_enable; // @[RegFile.scala 66:20:@36245.4]
  wire  regs_132_clock; // @[RegFile.scala 66:20:@36259.4]
  wire  regs_132_reset; // @[RegFile.scala 66:20:@36259.4]
  wire [63:0] regs_132_io_in; // @[RegFile.scala 66:20:@36259.4]
  wire  regs_132_io_reset; // @[RegFile.scala 66:20:@36259.4]
  wire [63:0] regs_132_io_out; // @[RegFile.scala 66:20:@36259.4]
  wire  regs_132_io_enable; // @[RegFile.scala 66:20:@36259.4]
  wire  regs_133_clock; // @[RegFile.scala 66:20:@36273.4]
  wire  regs_133_reset; // @[RegFile.scala 66:20:@36273.4]
  wire [63:0] regs_133_io_in; // @[RegFile.scala 66:20:@36273.4]
  wire  regs_133_io_reset; // @[RegFile.scala 66:20:@36273.4]
  wire [63:0] regs_133_io_out; // @[RegFile.scala 66:20:@36273.4]
  wire  regs_133_io_enable; // @[RegFile.scala 66:20:@36273.4]
  wire  regs_134_clock; // @[RegFile.scala 66:20:@36287.4]
  wire  regs_134_reset; // @[RegFile.scala 66:20:@36287.4]
  wire [63:0] regs_134_io_in; // @[RegFile.scala 66:20:@36287.4]
  wire  regs_134_io_reset; // @[RegFile.scala 66:20:@36287.4]
  wire [63:0] regs_134_io_out; // @[RegFile.scala 66:20:@36287.4]
  wire  regs_134_io_enable; // @[RegFile.scala 66:20:@36287.4]
  wire  regs_135_clock; // @[RegFile.scala 66:20:@36301.4]
  wire  regs_135_reset; // @[RegFile.scala 66:20:@36301.4]
  wire [63:0] regs_135_io_in; // @[RegFile.scala 66:20:@36301.4]
  wire  regs_135_io_reset; // @[RegFile.scala 66:20:@36301.4]
  wire [63:0] regs_135_io_out; // @[RegFile.scala 66:20:@36301.4]
  wire  regs_135_io_enable; // @[RegFile.scala 66:20:@36301.4]
  wire  regs_136_clock; // @[RegFile.scala 66:20:@36315.4]
  wire  regs_136_reset; // @[RegFile.scala 66:20:@36315.4]
  wire [63:0] regs_136_io_in; // @[RegFile.scala 66:20:@36315.4]
  wire  regs_136_io_reset; // @[RegFile.scala 66:20:@36315.4]
  wire [63:0] regs_136_io_out; // @[RegFile.scala 66:20:@36315.4]
  wire  regs_136_io_enable; // @[RegFile.scala 66:20:@36315.4]
  wire  regs_137_clock; // @[RegFile.scala 66:20:@36329.4]
  wire  regs_137_reset; // @[RegFile.scala 66:20:@36329.4]
  wire [63:0] regs_137_io_in; // @[RegFile.scala 66:20:@36329.4]
  wire  regs_137_io_reset; // @[RegFile.scala 66:20:@36329.4]
  wire [63:0] regs_137_io_out; // @[RegFile.scala 66:20:@36329.4]
  wire  regs_137_io_enable; // @[RegFile.scala 66:20:@36329.4]
  wire  regs_138_clock; // @[RegFile.scala 66:20:@36343.4]
  wire  regs_138_reset; // @[RegFile.scala 66:20:@36343.4]
  wire [63:0] regs_138_io_in; // @[RegFile.scala 66:20:@36343.4]
  wire  regs_138_io_reset; // @[RegFile.scala 66:20:@36343.4]
  wire [63:0] regs_138_io_out; // @[RegFile.scala 66:20:@36343.4]
  wire  regs_138_io_enable; // @[RegFile.scala 66:20:@36343.4]
  wire  regs_139_clock; // @[RegFile.scala 66:20:@36357.4]
  wire  regs_139_reset; // @[RegFile.scala 66:20:@36357.4]
  wire [63:0] regs_139_io_in; // @[RegFile.scala 66:20:@36357.4]
  wire  regs_139_io_reset; // @[RegFile.scala 66:20:@36357.4]
  wire [63:0] regs_139_io_out; // @[RegFile.scala 66:20:@36357.4]
  wire  regs_139_io_enable; // @[RegFile.scala 66:20:@36357.4]
  wire  regs_140_clock; // @[RegFile.scala 66:20:@36371.4]
  wire  regs_140_reset; // @[RegFile.scala 66:20:@36371.4]
  wire [63:0] regs_140_io_in; // @[RegFile.scala 66:20:@36371.4]
  wire  regs_140_io_reset; // @[RegFile.scala 66:20:@36371.4]
  wire [63:0] regs_140_io_out; // @[RegFile.scala 66:20:@36371.4]
  wire  regs_140_io_enable; // @[RegFile.scala 66:20:@36371.4]
  wire  regs_141_clock; // @[RegFile.scala 66:20:@36385.4]
  wire  regs_141_reset; // @[RegFile.scala 66:20:@36385.4]
  wire [63:0] regs_141_io_in; // @[RegFile.scala 66:20:@36385.4]
  wire  regs_141_io_reset; // @[RegFile.scala 66:20:@36385.4]
  wire [63:0] regs_141_io_out; // @[RegFile.scala 66:20:@36385.4]
  wire  regs_141_io_enable; // @[RegFile.scala 66:20:@36385.4]
  wire  regs_142_clock; // @[RegFile.scala 66:20:@36399.4]
  wire  regs_142_reset; // @[RegFile.scala 66:20:@36399.4]
  wire [63:0] regs_142_io_in; // @[RegFile.scala 66:20:@36399.4]
  wire  regs_142_io_reset; // @[RegFile.scala 66:20:@36399.4]
  wire [63:0] regs_142_io_out; // @[RegFile.scala 66:20:@36399.4]
  wire  regs_142_io_enable; // @[RegFile.scala 66:20:@36399.4]
  wire  regs_143_clock; // @[RegFile.scala 66:20:@36413.4]
  wire  regs_143_reset; // @[RegFile.scala 66:20:@36413.4]
  wire [63:0] regs_143_io_in; // @[RegFile.scala 66:20:@36413.4]
  wire  regs_143_io_reset; // @[RegFile.scala 66:20:@36413.4]
  wire [63:0] regs_143_io_out; // @[RegFile.scala 66:20:@36413.4]
  wire  regs_143_io_enable; // @[RegFile.scala 66:20:@36413.4]
  wire  regs_144_clock; // @[RegFile.scala 66:20:@36427.4]
  wire  regs_144_reset; // @[RegFile.scala 66:20:@36427.4]
  wire [63:0] regs_144_io_in; // @[RegFile.scala 66:20:@36427.4]
  wire  regs_144_io_reset; // @[RegFile.scala 66:20:@36427.4]
  wire [63:0] regs_144_io_out; // @[RegFile.scala 66:20:@36427.4]
  wire  regs_144_io_enable; // @[RegFile.scala 66:20:@36427.4]
  wire  regs_145_clock; // @[RegFile.scala 66:20:@36441.4]
  wire  regs_145_reset; // @[RegFile.scala 66:20:@36441.4]
  wire [63:0] regs_145_io_in; // @[RegFile.scala 66:20:@36441.4]
  wire  regs_145_io_reset; // @[RegFile.scala 66:20:@36441.4]
  wire [63:0] regs_145_io_out; // @[RegFile.scala 66:20:@36441.4]
  wire  regs_145_io_enable; // @[RegFile.scala 66:20:@36441.4]
  wire  regs_146_clock; // @[RegFile.scala 66:20:@36455.4]
  wire  regs_146_reset; // @[RegFile.scala 66:20:@36455.4]
  wire [63:0] regs_146_io_in; // @[RegFile.scala 66:20:@36455.4]
  wire  regs_146_io_reset; // @[RegFile.scala 66:20:@36455.4]
  wire [63:0] regs_146_io_out; // @[RegFile.scala 66:20:@36455.4]
  wire  regs_146_io_enable; // @[RegFile.scala 66:20:@36455.4]
  wire  regs_147_clock; // @[RegFile.scala 66:20:@36469.4]
  wire  regs_147_reset; // @[RegFile.scala 66:20:@36469.4]
  wire [63:0] regs_147_io_in; // @[RegFile.scala 66:20:@36469.4]
  wire  regs_147_io_reset; // @[RegFile.scala 66:20:@36469.4]
  wire [63:0] regs_147_io_out; // @[RegFile.scala 66:20:@36469.4]
  wire  regs_147_io_enable; // @[RegFile.scala 66:20:@36469.4]
  wire  regs_148_clock; // @[RegFile.scala 66:20:@36483.4]
  wire  regs_148_reset; // @[RegFile.scala 66:20:@36483.4]
  wire [63:0] regs_148_io_in; // @[RegFile.scala 66:20:@36483.4]
  wire  regs_148_io_reset; // @[RegFile.scala 66:20:@36483.4]
  wire [63:0] regs_148_io_out; // @[RegFile.scala 66:20:@36483.4]
  wire  regs_148_io_enable; // @[RegFile.scala 66:20:@36483.4]
  wire  regs_149_clock; // @[RegFile.scala 66:20:@36497.4]
  wire  regs_149_reset; // @[RegFile.scala 66:20:@36497.4]
  wire [63:0] regs_149_io_in; // @[RegFile.scala 66:20:@36497.4]
  wire  regs_149_io_reset; // @[RegFile.scala 66:20:@36497.4]
  wire [63:0] regs_149_io_out; // @[RegFile.scala 66:20:@36497.4]
  wire  regs_149_io_enable; // @[RegFile.scala 66:20:@36497.4]
  wire  regs_150_clock; // @[RegFile.scala 66:20:@36511.4]
  wire  regs_150_reset; // @[RegFile.scala 66:20:@36511.4]
  wire [63:0] regs_150_io_in; // @[RegFile.scala 66:20:@36511.4]
  wire  regs_150_io_reset; // @[RegFile.scala 66:20:@36511.4]
  wire [63:0] regs_150_io_out; // @[RegFile.scala 66:20:@36511.4]
  wire  regs_150_io_enable; // @[RegFile.scala 66:20:@36511.4]
  wire  regs_151_clock; // @[RegFile.scala 66:20:@36525.4]
  wire  regs_151_reset; // @[RegFile.scala 66:20:@36525.4]
  wire [63:0] regs_151_io_in; // @[RegFile.scala 66:20:@36525.4]
  wire  regs_151_io_reset; // @[RegFile.scala 66:20:@36525.4]
  wire [63:0] regs_151_io_out; // @[RegFile.scala 66:20:@36525.4]
  wire  regs_151_io_enable; // @[RegFile.scala 66:20:@36525.4]
  wire  regs_152_clock; // @[RegFile.scala 66:20:@36539.4]
  wire  regs_152_reset; // @[RegFile.scala 66:20:@36539.4]
  wire [63:0] regs_152_io_in; // @[RegFile.scala 66:20:@36539.4]
  wire  regs_152_io_reset; // @[RegFile.scala 66:20:@36539.4]
  wire [63:0] regs_152_io_out; // @[RegFile.scala 66:20:@36539.4]
  wire  regs_152_io_enable; // @[RegFile.scala 66:20:@36539.4]
  wire  regs_153_clock; // @[RegFile.scala 66:20:@36553.4]
  wire  regs_153_reset; // @[RegFile.scala 66:20:@36553.4]
  wire [63:0] regs_153_io_in; // @[RegFile.scala 66:20:@36553.4]
  wire  regs_153_io_reset; // @[RegFile.scala 66:20:@36553.4]
  wire [63:0] regs_153_io_out; // @[RegFile.scala 66:20:@36553.4]
  wire  regs_153_io_enable; // @[RegFile.scala 66:20:@36553.4]
  wire  regs_154_clock; // @[RegFile.scala 66:20:@36567.4]
  wire  regs_154_reset; // @[RegFile.scala 66:20:@36567.4]
  wire [63:0] regs_154_io_in; // @[RegFile.scala 66:20:@36567.4]
  wire  regs_154_io_reset; // @[RegFile.scala 66:20:@36567.4]
  wire [63:0] regs_154_io_out; // @[RegFile.scala 66:20:@36567.4]
  wire  regs_154_io_enable; // @[RegFile.scala 66:20:@36567.4]
  wire  regs_155_clock; // @[RegFile.scala 66:20:@36581.4]
  wire  regs_155_reset; // @[RegFile.scala 66:20:@36581.4]
  wire [63:0] regs_155_io_in; // @[RegFile.scala 66:20:@36581.4]
  wire  regs_155_io_reset; // @[RegFile.scala 66:20:@36581.4]
  wire [63:0] regs_155_io_out; // @[RegFile.scala 66:20:@36581.4]
  wire  regs_155_io_enable; // @[RegFile.scala 66:20:@36581.4]
  wire  regs_156_clock; // @[RegFile.scala 66:20:@36595.4]
  wire  regs_156_reset; // @[RegFile.scala 66:20:@36595.4]
  wire [63:0] regs_156_io_in; // @[RegFile.scala 66:20:@36595.4]
  wire  regs_156_io_reset; // @[RegFile.scala 66:20:@36595.4]
  wire [63:0] regs_156_io_out; // @[RegFile.scala 66:20:@36595.4]
  wire  regs_156_io_enable; // @[RegFile.scala 66:20:@36595.4]
  wire  regs_157_clock; // @[RegFile.scala 66:20:@36609.4]
  wire  regs_157_reset; // @[RegFile.scala 66:20:@36609.4]
  wire [63:0] regs_157_io_in; // @[RegFile.scala 66:20:@36609.4]
  wire  regs_157_io_reset; // @[RegFile.scala 66:20:@36609.4]
  wire [63:0] regs_157_io_out; // @[RegFile.scala 66:20:@36609.4]
  wire  regs_157_io_enable; // @[RegFile.scala 66:20:@36609.4]
  wire  regs_158_clock; // @[RegFile.scala 66:20:@36623.4]
  wire  regs_158_reset; // @[RegFile.scala 66:20:@36623.4]
  wire [63:0] regs_158_io_in; // @[RegFile.scala 66:20:@36623.4]
  wire  regs_158_io_reset; // @[RegFile.scala 66:20:@36623.4]
  wire [63:0] regs_158_io_out; // @[RegFile.scala 66:20:@36623.4]
  wire  regs_158_io_enable; // @[RegFile.scala 66:20:@36623.4]
  wire  regs_159_clock; // @[RegFile.scala 66:20:@36637.4]
  wire  regs_159_reset; // @[RegFile.scala 66:20:@36637.4]
  wire [63:0] regs_159_io_in; // @[RegFile.scala 66:20:@36637.4]
  wire  regs_159_io_reset; // @[RegFile.scala 66:20:@36637.4]
  wire [63:0] regs_159_io_out; // @[RegFile.scala 66:20:@36637.4]
  wire  regs_159_io_enable; // @[RegFile.scala 66:20:@36637.4]
  wire  regs_160_clock; // @[RegFile.scala 66:20:@36651.4]
  wire  regs_160_reset; // @[RegFile.scala 66:20:@36651.4]
  wire [63:0] regs_160_io_in; // @[RegFile.scala 66:20:@36651.4]
  wire  regs_160_io_reset; // @[RegFile.scala 66:20:@36651.4]
  wire [63:0] regs_160_io_out; // @[RegFile.scala 66:20:@36651.4]
  wire  regs_160_io_enable; // @[RegFile.scala 66:20:@36651.4]
  wire  regs_161_clock; // @[RegFile.scala 66:20:@36665.4]
  wire  regs_161_reset; // @[RegFile.scala 66:20:@36665.4]
  wire [63:0] regs_161_io_in; // @[RegFile.scala 66:20:@36665.4]
  wire  regs_161_io_reset; // @[RegFile.scala 66:20:@36665.4]
  wire [63:0] regs_161_io_out; // @[RegFile.scala 66:20:@36665.4]
  wire  regs_161_io_enable; // @[RegFile.scala 66:20:@36665.4]
  wire  regs_162_clock; // @[RegFile.scala 66:20:@36679.4]
  wire  regs_162_reset; // @[RegFile.scala 66:20:@36679.4]
  wire [63:0] regs_162_io_in; // @[RegFile.scala 66:20:@36679.4]
  wire  regs_162_io_reset; // @[RegFile.scala 66:20:@36679.4]
  wire [63:0] regs_162_io_out; // @[RegFile.scala 66:20:@36679.4]
  wire  regs_162_io_enable; // @[RegFile.scala 66:20:@36679.4]
  wire  regs_163_clock; // @[RegFile.scala 66:20:@36693.4]
  wire  regs_163_reset; // @[RegFile.scala 66:20:@36693.4]
  wire [63:0] regs_163_io_in; // @[RegFile.scala 66:20:@36693.4]
  wire  regs_163_io_reset; // @[RegFile.scala 66:20:@36693.4]
  wire [63:0] regs_163_io_out; // @[RegFile.scala 66:20:@36693.4]
  wire  regs_163_io_enable; // @[RegFile.scala 66:20:@36693.4]
  wire  regs_164_clock; // @[RegFile.scala 66:20:@36707.4]
  wire  regs_164_reset; // @[RegFile.scala 66:20:@36707.4]
  wire [63:0] regs_164_io_in; // @[RegFile.scala 66:20:@36707.4]
  wire  regs_164_io_reset; // @[RegFile.scala 66:20:@36707.4]
  wire [63:0] regs_164_io_out; // @[RegFile.scala 66:20:@36707.4]
  wire  regs_164_io_enable; // @[RegFile.scala 66:20:@36707.4]
  wire  regs_165_clock; // @[RegFile.scala 66:20:@36721.4]
  wire  regs_165_reset; // @[RegFile.scala 66:20:@36721.4]
  wire [63:0] regs_165_io_in; // @[RegFile.scala 66:20:@36721.4]
  wire  regs_165_io_reset; // @[RegFile.scala 66:20:@36721.4]
  wire [63:0] regs_165_io_out; // @[RegFile.scala 66:20:@36721.4]
  wire  regs_165_io_enable; // @[RegFile.scala 66:20:@36721.4]
  wire  regs_166_clock; // @[RegFile.scala 66:20:@36735.4]
  wire  regs_166_reset; // @[RegFile.scala 66:20:@36735.4]
  wire [63:0] regs_166_io_in; // @[RegFile.scala 66:20:@36735.4]
  wire  regs_166_io_reset; // @[RegFile.scala 66:20:@36735.4]
  wire [63:0] regs_166_io_out; // @[RegFile.scala 66:20:@36735.4]
  wire  regs_166_io_enable; // @[RegFile.scala 66:20:@36735.4]
  wire  regs_167_clock; // @[RegFile.scala 66:20:@36749.4]
  wire  regs_167_reset; // @[RegFile.scala 66:20:@36749.4]
  wire [63:0] regs_167_io_in; // @[RegFile.scala 66:20:@36749.4]
  wire  regs_167_io_reset; // @[RegFile.scala 66:20:@36749.4]
  wire [63:0] regs_167_io_out; // @[RegFile.scala 66:20:@36749.4]
  wire  regs_167_io_enable; // @[RegFile.scala 66:20:@36749.4]
  wire  regs_168_clock; // @[RegFile.scala 66:20:@36763.4]
  wire  regs_168_reset; // @[RegFile.scala 66:20:@36763.4]
  wire [63:0] regs_168_io_in; // @[RegFile.scala 66:20:@36763.4]
  wire  regs_168_io_reset; // @[RegFile.scala 66:20:@36763.4]
  wire [63:0] regs_168_io_out; // @[RegFile.scala 66:20:@36763.4]
  wire  regs_168_io_enable; // @[RegFile.scala 66:20:@36763.4]
  wire  regs_169_clock; // @[RegFile.scala 66:20:@36777.4]
  wire  regs_169_reset; // @[RegFile.scala 66:20:@36777.4]
  wire [63:0] regs_169_io_in; // @[RegFile.scala 66:20:@36777.4]
  wire  regs_169_io_reset; // @[RegFile.scala 66:20:@36777.4]
  wire [63:0] regs_169_io_out; // @[RegFile.scala 66:20:@36777.4]
  wire  regs_169_io_enable; // @[RegFile.scala 66:20:@36777.4]
  wire  regs_170_clock; // @[RegFile.scala 66:20:@36791.4]
  wire  regs_170_reset; // @[RegFile.scala 66:20:@36791.4]
  wire [63:0] regs_170_io_in; // @[RegFile.scala 66:20:@36791.4]
  wire  regs_170_io_reset; // @[RegFile.scala 66:20:@36791.4]
  wire [63:0] regs_170_io_out; // @[RegFile.scala 66:20:@36791.4]
  wire  regs_170_io_enable; // @[RegFile.scala 66:20:@36791.4]
  wire  regs_171_clock; // @[RegFile.scala 66:20:@36805.4]
  wire  regs_171_reset; // @[RegFile.scala 66:20:@36805.4]
  wire [63:0] regs_171_io_in; // @[RegFile.scala 66:20:@36805.4]
  wire  regs_171_io_reset; // @[RegFile.scala 66:20:@36805.4]
  wire [63:0] regs_171_io_out; // @[RegFile.scala 66:20:@36805.4]
  wire  regs_171_io_enable; // @[RegFile.scala 66:20:@36805.4]
  wire  regs_172_clock; // @[RegFile.scala 66:20:@36819.4]
  wire  regs_172_reset; // @[RegFile.scala 66:20:@36819.4]
  wire [63:0] regs_172_io_in; // @[RegFile.scala 66:20:@36819.4]
  wire  regs_172_io_reset; // @[RegFile.scala 66:20:@36819.4]
  wire [63:0] regs_172_io_out; // @[RegFile.scala 66:20:@36819.4]
  wire  regs_172_io_enable; // @[RegFile.scala 66:20:@36819.4]
  wire  regs_173_clock; // @[RegFile.scala 66:20:@36833.4]
  wire  regs_173_reset; // @[RegFile.scala 66:20:@36833.4]
  wire [63:0] regs_173_io_in; // @[RegFile.scala 66:20:@36833.4]
  wire  regs_173_io_reset; // @[RegFile.scala 66:20:@36833.4]
  wire [63:0] regs_173_io_out; // @[RegFile.scala 66:20:@36833.4]
  wire  regs_173_io_enable; // @[RegFile.scala 66:20:@36833.4]
  wire  regs_174_clock; // @[RegFile.scala 66:20:@36847.4]
  wire  regs_174_reset; // @[RegFile.scala 66:20:@36847.4]
  wire [63:0] regs_174_io_in; // @[RegFile.scala 66:20:@36847.4]
  wire  regs_174_io_reset; // @[RegFile.scala 66:20:@36847.4]
  wire [63:0] regs_174_io_out; // @[RegFile.scala 66:20:@36847.4]
  wire  regs_174_io_enable; // @[RegFile.scala 66:20:@36847.4]
  wire  regs_175_clock; // @[RegFile.scala 66:20:@36861.4]
  wire  regs_175_reset; // @[RegFile.scala 66:20:@36861.4]
  wire [63:0] regs_175_io_in; // @[RegFile.scala 66:20:@36861.4]
  wire  regs_175_io_reset; // @[RegFile.scala 66:20:@36861.4]
  wire [63:0] regs_175_io_out; // @[RegFile.scala 66:20:@36861.4]
  wire  regs_175_io_enable; // @[RegFile.scala 66:20:@36861.4]
  wire  regs_176_clock; // @[RegFile.scala 66:20:@36875.4]
  wire  regs_176_reset; // @[RegFile.scala 66:20:@36875.4]
  wire [63:0] regs_176_io_in; // @[RegFile.scala 66:20:@36875.4]
  wire  regs_176_io_reset; // @[RegFile.scala 66:20:@36875.4]
  wire [63:0] regs_176_io_out; // @[RegFile.scala 66:20:@36875.4]
  wire  regs_176_io_enable; // @[RegFile.scala 66:20:@36875.4]
  wire  regs_177_clock; // @[RegFile.scala 66:20:@36889.4]
  wire  regs_177_reset; // @[RegFile.scala 66:20:@36889.4]
  wire [63:0] regs_177_io_in; // @[RegFile.scala 66:20:@36889.4]
  wire  regs_177_io_reset; // @[RegFile.scala 66:20:@36889.4]
  wire [63:0] regs_177_io_out; // @[RegFile.scala 66:20:@36889.4]
  wire  regs_177_io_enable; // @[RegFile.scala 66:20:@36889.4]
  wire  regs_178_clock; // @[RegFile.scala 66:20:@36903.4]
  wire  regs_178_reset; // @[RegFile.scala 66:20:@36903.4]
  wire [63:0] regs_178_io_in; // @[RegFile.scala 66:20:@36903.4]
  wire  regs_178_io_reset; // @[RegFile.scala 66:20:@36903.4]
  wire [63:0] regs_178_io_out; // @[RegFile.scala 66:20:@36903.4]
  wire  regs_178_io_enable; // @[RegFile.scala 66:20:@36903.4]
  wire  regs_179_clock; // @[RegFile.scala 66:20:@36917.4]
  wire  regs_179_reset; // @[RegFile.scala 66:20:@36917.4]
  wire [63:0] regs_179_io_in; // @[RegFile.scala 66:20:@36917.4]
  wire  regs_179_io_reset; // @[RegFile.scala 66:20:@36917.4]
  wire [63:0] regs_179_io_out; // @[RegFile.scala 66:20:@36917.4]
  wire  regs_179_io_enable; // @[RegFile.scala 66:20:@36917.4]
  wire  regs_180_clock; // @[RegFile.scala 66:20:@36931.4]
  wire  regs_180_reset; // @[RegFile.scala 66:20:@36931.4]
  wire [63:0] regs_180_io_in; // @[RegFile.scala 66:20:@36931.4]
  wire  regs_180_io_reset; // @[RegFile.scala 66:20:@36931.4]
  wire [63:0] regs_180_io_out; // @[RegFile.scala 66:20:@36931.4]
  wire  regs_180_io_enable; // @[RegFile.scala 66:20:@36931.4]
  wire  regs_181_clock; // @[RegFile.scala 66:20:@36945.4]
  wire  regs_181_reset; // @[RegFile.scala 66:20:@36945.4]
  wire [63:0] regs_181_io_in; // @[RegFile.scala 66:20:@36945.4]
  wire  regs_181_io_reset; // @[RegFile.scala 66:20:@36945.4]
  wire [63:0] regs_181_io_out; // @[RegFile.scala 66:20:@36945.4]
  wire  regs_181_io_enable; // @[RegFile.scala 66:20:@36945.4]
  wire  regs_182_clock; // @[RegFile.scala 66:20:@36959.4]
  wire  regs_182_reset; // @[RegFile.scala 66:20:@36959.4]
  wire [63:0] regs_182_io_in; // @[RegFile.scala 66:20:@36959.4]
  wire  regs_182_io_reset; // @[RegFile.scala 66:20:@36959.4]
  wire [63:0] regs_182_io_out; // @[RegFile.scala 66:20:@36959.4]
  wire  regs_182_io_enable; // @[RegFile.scala 66:20:@36959.4]
  wire  regs_183_clock; // @[RegFile.scala 66:20:@36973.4]
  wire  regs_183_reset; // @[RegFile.scala 66:20:@36973.4]
  wire [63:0] regs_183_io_in; // @[RegFile.scala 66:20:@36973.4]
  wire  regs_183_io_reset; // @[RegFile.scala 66:20:@36973.4]
  wire [63:0] regs_183_io_out; // @[RegFile.scala 66:20:@36973.4]
  wire  regs_183_io_enable; // @[RegFile.scala 66:20:@36973.4]
  wire  regs_184_clock; // @[RegFile.scala 66:20:@36987.4]
  wire  regs_184_reset; // @[RegFile.scala 66:20:@36987.4]
  wire [63:0] regs_184_io_in; // @[RegFile.scala 66:20:@36987.4]
  wire  regs_184_io_reset; // @[RegFile.scala 66:20:@36987.4]
  wire [63:0] regs_184_io_out; // @[RegFile.scala 66:20:@36987.4]
  wire  regs_184_io_enable; // @[RegFile.scala 66:20:@36987.4]
  wire  regs_185_clock; // @[RegFile.scala 66:20:@37001.4]
  wire  regs_185_reset; // @[RegFile.scala 66:20:@37001.4]
  wire [63:0] regs_185_io_in; // @[RegFile.scala 66:20:@37001.4]
  wire  regs_185_io_reset; // @[RegFile.scala 66:20:@37001.4]
  wire [63:0] regs_185_io_out; // @[RegFile.scala 66:20:@37001.4]
  wire  regs_185_io_enable; // @[RegFile.scala 66:20:@37001.4]
  wire  regs_186_clock; // @[RegFile.scala 66:20:@37015.4]
  wire  regs_186_reset; // @[RegFile.scala 66:20:@37015.4]
  wire [63:0] regs_186_io_in; // @[RegFile.scala 66:20:@37015.4]
  wire  regs_186_io_reset; // @[RegFile.scala 66:20:@37015.4]
  wire [63:0] regs_186_io_out; // @[RegFile.scala 66:20:@37015.4]
  wire  regs_186_io_enable; // @[RegFile.scala 66:20:@37015.4]
  wire  regs_187_clock; // @[RegFile.scala 66:20:@37029.4]
  wire  regs_187_reset; // @[RegFile.scala 66:20:@37029.4]
  wire [63:0] regs_187_io_in; // @[RegFile.scala 66:20:@37029.4]
  wire  regs_187_io_reset; // @[RegFile.scala 66:20:@37029.4]
  wire [63:0] regs_187_io_out; // @[RegFile.scala 66:20:@37029.4]
  wire  regs_187_io_enable; // @[RegFile.scala 66:20:@37029.4]
  wire  regs_188_clock; // @[RegFile.scala 66:20:@37043.4]
  wire  regs_188_reset; // @[RegFile.scala 66:20:@37043.4]
  wire [63:0] regs_188_io_in; // @[RegFile.scala 66:20:@37043.4]
  wire  regs_188_io_reset; // @[RegFile.scala 66:20:@37043.4]
  wire [63:0] regs_188_io_out; // @[RegFile.scala 66:20:@37043.4]
  wire  regs_188_io_enable; // @[RegFile.scala 66:20:@37043.4]
  wire  regs_189_clock; // @[RegFile.scala 66:20:@37057.4]
  wire  regs_189_reset; // @[RegFile.scala 66:20:@37057.4]
  wire [63:0] regs_189_io_in; // @[RegFile.scala 66:20:@37057.4]
  wire  regs_189_io_reset; // @[RegFile.scala 66:20:@37057.4]
  wire [63:0] regs_189_io_out; // @[RegFile.scala 66:20:@37057.4]
  wire  regs_189_io_enable; // @[RegFile.scala 66:20:@37057.4]
  wire  regs_190_clock; // @[RegFile.scala 66:20:@37071.4]
  wire  regs_190_reset; // @[RegFile.scala 66:20:@37071.4]
  wire [63:0] regs_190_io_in; // @[RegFile.scala 66:20:@37071.4]
  wire  regs_190_io_reset; // @[RegFile.scala 66:20:@37071.4]
  wire [63:0] regs_190_io_out; // @[RegFile.scala 66:20:@37071.4]
  wire  regs_190_io_enable; // @[RegFile.scala 66:20:@37071.4]
  wire  regs_191_clock; // @[RegFile.scala 66:20:@37085.4]
  wire  regs_191_reset; // @[RegFile.scala 66:20:@37085.4]
  wire [63:0] regs_191_io_in; // @[RegFile.scala 66:20:@37085.4]
  wire  regs_191_io_reset; // @[RegFile.scala 66:20:@37085.4]
  wire [63:0] regs_191_io_out; // @[RegFile.scala 66:20:@37085.4]
  wire  regs_191_io_enable; // @[RegFile.scala 66:20:@37085.4]
  wire  regs_192_clock; // @[RegFile.scala 66:20:@37099.4]
  wire  regs_192_reset; // @[RegFile.scala 66:20:@37099.4]
  wire [63:0] regs_192_io_in; // @[RegFile.scala 66:20:@37099.4]
  wire  regs_192_io_reset; // @[RegFile.scala 66:20:@37099.4]
  wire [63:0] regs_192_io_out; // @[RegFile.scala 66:20:@37099.4]
  wire  regs_192_io_enable; // @[RegFile.scala 66:20:@37099.4]
  wire  regs_193_clock; // @[RegFile.scala 66:20:@37113.4]
  wire  regs_193_reset; // @[RegFile.scala 66:20:@37113.4]
  wire [63:0] regs_193_io_in; // @[RegFile.scala 66:20:@37113.4]
  wire  regs_193_io_reset; // @[RegFile.scala 66:20:@37113.4]
  wire [63:0] regs_193_io_out; // @[RegFile.scala 66:20:@37113.4]
  wire  regs_193_io_enable; // @[RegFile.scala 66:20:@37113.4]
  wire  regs_194_clock; // @[RegFile.scala 66:20:@37127.4]
  wire  regs_194_reset; // @[RegFile.scala 66:20:@37127.4]
  wire [63:0] regs_194_io_in; // @[RegFile.scala 66:20:@37127.4]
  wire  regs_194_io_reset; // @[RegFile.scala 66:20:@37127.4]
  wire [63:0] regs_194_io_out; // @[RegFile.scala 66:20:@37127.4]
  wire  regs_194_io_enable; // @[RegFile.scala 66:20:@37127.4]
  wire  regs_195_clock; // @[RegFile.scala 66:20:@37141.4]
  wire  regs_195_reset; // @[RegFile.scala 66:20:@37141.4]
  wire [63:0] regs_195_io_in; // @[RegFile.scala 66:20:@37141.4]
  wire  regs_195_io_reset; // @[RegFile.scala 66:20:@37141.4]
  wire [63:0] regs_195_io_out; // @[RegFile.scala 66:20:@37141.4]
  wire  regs_195_io_enable; // @[RegFile.scala 66:20:@37141.4]
  wire  regs_196_clock; // @[RegFile.scala 66:20:@37155.4]
  wire  regs_196_reset; // @[RegFile.scala 66:20:@37155.4]
  wire [63:0] regs_196_io_in; // @[RegFile.scala 66:20:@37155.4]
  wire  regs_196_io_reset; // @[RegFile.scala 66:20:@37155.4]
  wire [63:0] regs_196_io_out; // @[RegFile.scala 66:20:@37155.4]
  wire  regs_196_io_enable; // @[RegFile.scala 66:20:@37155.4]
  wire  regs_197_clock; // @[RegFile.scala 66:20:@37169.4]
  wire  regs_197_reset; // @[RegFile.scala 66:20:@37169.4]
  wire [63:0] regs_197_io_in; // @[RegFile.scala 66:20:@37169.4]
  wire  regs_197_io_reset; // @[RegFile.scala 66:20:@37169.4]
  wire [63:0] regs_197_io_out; // @[RegFile.scala 66:20:@37169.4]
  wire  regs_197_io_enable; // @[RegFile.scala 66:20:@37169.4]
  wire  regs_198_clock; // @[RegFile.scala 66:20:@37183.4]
  wire  regs_198_reset; // @[RegFile.scala 66:20:@37183.4]
  wire [63:0] regs_198_io_in; // @[RegFile.scala 66:20:@37183.4]
  wire  regs_198_io_reset; // @[RegFile.scala 66:20:@37183.4]
  wire [63:0] regs_198_io_out; // @[RegFile.scala 66:20:@37183.4]
  wire  regs_198_io_enable; // @[RegFile.scala 66:20:@37183.4]
  wire  regs_199_clock; // @[RegFile.scala 66:20:@37197.4]
  wire  regs_199_reset; // @[RegFile.scala 66:20:@37197.4]
  wire [63:0] regs_199_io_in; // @[RegFile.scala 66:20:@37197.4]
  wire  regs_199_io_reset; // @[RegFile.scala 66:20:@37197.4]
  wire [63:0] regs_199_io_out; // @[RegFile.scala 66:20:@37197.4]
  wire  regs_199_io_enable; // @[RegFile.scala 66:20:@37197.4]
  wire  regs_200_clock; // @[RegFile.scala 66:20:@37211.4]
  wire  regs_200_reset; // @[RegFile.scala 66:20:@37211.4]
  wire [63:0] regs_200_io_in; // @[RegFile.scala 66:20:@37211.4]
  wire  regs_200_io_reset; // @[RegFile.scala 66:20:@37211.4]
  wire [63:0] regs_200_io_out; // @[RegFile.scala 66:20:@37211.4]
  wire  regs_200_io_enable; // @[RegFile.scala 66:20:@37211.4]
  wire  regs_201_clock; // @[RegFile.scala 66:20:@37225.4]
  wire  regs_201_reset; // @[RegFile.scala 66:20:@37225.4]
  wire [63:0] regs_201_io_in; // @[RegFile.scala 66:20:@37225.4]
  wire  regs_201_io_reset; // @[RegFile.scala 66:20:@37225.4]
  wire [63:0] regs_201_io_out; // @[RegFile.scala 66:20:@37225.4]
  wire  regs_201_io_enable; // @[RegFile.scala 66:20:@37225.4]
  wire  regs_202_clock; // @[RegFile.scala 66:20:@37239.4]
  wire  regs_202_reset; // @[RegFile.scala 66:20:@37239.4]
  wire [63:0] regs_202_io_in; // @[RegFile.scala 66:20:@37239.4]
  wire  regs_202_io_reset; // @[RegFile.scala 66:20:@37239.4]
  wire [63:0] regs_202_io_out; // @[RegFile.scala 66:20:@37239.4]
  wire  regs_202_io_enable; // @[RegFile.scala 66:20:@37239.4]
  wire  regs_203_clock; // @[RegFile.scala 66:20:@37253.4]
  wire  regs_203_reset; // @[RegFile.scala 66:20:@37253.4]
  wire [63:0] regs_203_io_in; // @[RegFile.scala 66:20:@37253.4]
  wire  regs_203_io_reset; // @[RegFile.scala 66:20:@37253.4]
  wire [63:0] regs_203_io_out; // @[RegFile.scala 66:20:@37253.4]
  wire  regs_203_io_enable; // @[RegFile.scala 66:20:@37253.4]
  wire  regs_204_clock; // @[RegFile.scala 66:20:@37267.4]
  wire  regs_204_reset; // @[RegFile.scala 66:20:@37267.4]
  wire [63:0] regs_204_io_in; // @[RegFile.scala 66:20:@37267.4]
  wire  regs_204_io_reset; // @[RegFile.scala 66:20:@37267.4]
  wire [63:0] regs_204_io_out; // @[RegFile.scala 66:20:@37267.4]
  wire  regs_204_io_enable; // @[RegFile.scala 66:20:@37267.4]
  wire  regs_205_clock; // @[RegFile.scala 66:20:@37281.4]
  wire  regs_205_reset; // @[RegFile.scala 66:20:@37281.4]
  wire [63:0] regs_205_io_in; // @[RegFile.scala 66:20:@37281.4]
  wire  regs_205_io_reset; // @[RegFile.scala 66:20:@37281.4]
  wire [63:0] regs_205_io_out; // @[RegFile.scala 66:20:@37281.4]
  wire  regs_205_io_enable; // @[RegFile.scala 66:20:@37281.4]
  wire  regs_206_clock; // @[RegFile.scala 66:20:@37295.4]
  wire  regs_206_reset; // @[RegFile.scala 66:20:@37295.4]
  wire [63:0] regs_206_io_in; // @[RegFile.scala 66:20:@37295.4]
  wire  regs_206_io_reset; // @[RegFile.scala 66:20:@37295.4]
  wire [63:0] regs_206_io_out; // @[RegFile.scala 66:20:@37295.4]
  wire  regs_206_io_enable; // @[RegFile.scala 66:20:@37295.4]
  wire  regs_207_clock; // @[RegFile.scala 66:20:@37309.4]
  wire  regs_207_reset; // @[RegFile.scala 66:20:@37309.4]
  wire [63:0] regs_207_io_in; // @[RegFile.scala 66:20:@37309.4]
  wire  regs_207_io_reset; // @[RegFile.scala 66:20:@37309.4]
  wire [63:0] regs_207_io_out; // @[RegFile.scala 66:20:@37309.4]
  wire  regs_207_io_enable; // @[RegFile.scala 66:20:@37309.4]
  wire  regs_208_clock; // @[RegFile.scala 66:20:@37323.4]
  wire  regs_208_reset; // @[RegFile.scala 66:20:@37323.4]
  wire [63:0] regs_208_io_in; // @[RegFile.scala 66:20:@37323.4]
  wire  regs_208_io_reset; // @[RegFile.scala 66:20:@37323.4]
  wire [63:0] regs_208_io_out; // @[RegFile.scala 66:20:@37323.4]
  wire  regs_208_io_enable; // @[RegFile.scala 66:20:@37323.4]
  wire  regs_209_clock; // @[RegFile.scala 66:20:@37337.4]
  wire  regs_209_reset; // @[RegFile.scala 66:20:@37337.4]
  wire [63:0] regs_209_io_in; // @[RegFile.scala 66:20:@37337.4]
  wire  regs_209_io_reset; // @[RegFile.scala 66:20:@37337.4]
  wire [63:0] regs_209_io_out; // @[RegFile.scala 66:20:@37337.4]
  wire  regs_209_io_enable; // @[RegFile.scala 66:20:@37337.4]
  wire  regs_210_clock; // @[RegFile.scala 66:20:@37351.4]
  wire  regs_210_reset; // @[RegFile.scala 66:20:@37351.4]
  wire [63:0] regs_210_io_in; // @[RegFile.scala 66:20:@37351.4]
  wire  regs_210_io_reset; // @[RegFile.scala 66:20:@37351.4]
  wire [63:0] regs_210_io_out; // @[RegFile.scala 66:20:@37351.4]
  wire  regs_210_io_enable; // @[RegFile.scala 66:20:@37351.4]
  wire  regs_211_clock; // @[RegFile.scala 66:20:@37365.4]
  wire  regs_211_reset; // @[RegFile.scala 66:20:@37365.4]
  wire [63:0] regs_211_io_in; // @[RegFile.scala 66:20:@37365.4]
  wire  regs_211_io_reset; // @[RegFile.scala 66:20:@37365.4]
  wire [63:0] regs_211_io_out; // @[RegFile.scala 66:20:@37365.4]
  wire  regs_211_io_enable; // @[RegFile.scala 66:20:@37365.4]
  wire  regs_212_clock; // @[RegFile.scala 66:20:@37379.4]
  wire  regs_212_reset; // @[RegFile.scala 66:20:@37379.4]
  wire [63:0] regs_212_io_in; // @[RegFile.scala 66:20:@37379.4]
  wire  regs_212_io_reset; // @[RegFile.scala 66:20:@37379.4]
  wire [63:0] regs_212_io_out; // @[RegFile.scala 66:20:@37379.4]
  wire  regs_212_io_enable; // @[RegFile.scala 66:20:@37379.4]
  wire  regs_213_clock; // @[RegFile.scala 66:20:@37393.4]
  wire  regs_213_reset; // @[RegFile.scala 66:20:@37393.4]
  wire [63:0] regs_213_io_in; // @[RegFile.scala 66:20:@37393.4]
  wire  regs_213_io_reset; // @[RegFile.scala 66:20:@37393.4]
  wire [63:0] regs_213_io_out; // @[RegFile.scala 66:20:@37393.4]
  wire  regs_213_io_enable; // @[RegFile.scala 66:20:@37393.4]
  wire  regs_214_clock; // @[RegFile.scala 66:20:@37407.4]
  wire  regs_214_reset; // @[RegFile.scala 66:20:@37407.4]
  wire [63:0] regs_214_io_in; // @[RegFile.scala 66:20:@37407.4]
  wire  regs_214_io_reset; // @[RegFile.scala 66:20:@37407.4]
  wire [63:0] regs_214_io_out; // @[RegFile.scala 66:20:@37407.4]
  wire  regs_214_io_enable; // @[RegFile.scala 66:20:@37407.4]
  wire  regs_215_clock; // @[RegFile.scala 66:20:@37421.4]
  wire  regs_215_reset; // @[RegFile.scala 66:20:@37421.4]
  wire [63:0] regs_215_io_in; // @[RegFile.scala 66:20:@37421.4]
  wire  regs_215_io_reset; // @[RegFile.scala 66:20:@37421.4]
  wire [63:0] regs_215_io_out; // @[RegFile.scala 66:20:@37421.4]
  wire  regs_215_io_enable; // @[RegFile.scala 66:20:@37421.4]
  wire  regs_216_clock; // @[RegFile.scala 66:20:@37435.4]
  wire  regs_216_reset; // @[RegFile.scala 66:20:@37435.4]
  wire [63:0] regs_216_io_in; // @[RegFile.scala 66:20:@37435.4]
  wire  regs_216_io_reset; // @[RegFile.scala 66:20:@37435.4]
  wire [63:0] regs_216_io_out; // @[RegFile.scala 66:20:@37435.4]
  wire  regs_216_io_enable; // @[RegFile.scala 66:20:@37435.4]
  wire  regs_217_clock; // @[RegFile.scala 66:20:@37449.4]
  wire  regs_217_reset; // @[RegFile.scala 66:20:@37449.4]
  wire [63:0] regs_217_io_in; // @[RegFile.scala 66:20:@37449.4]
  wire  regs_217_io_reset; // @[RegFile.scala 66:20:@37449.4]
  wire [63:0] regs_217_io_out; // @[RegFile.scala 66:20:@37449.4]
  wire  regs_217_io_enable; // @[RegFile.scala 66:20:@37449.4]
  wire  regs_218_clock; // @[RegFile.scala 66:20:@37463.4]
  wire  regs_218_reset; // @[RegFile.scala 66:20:@37463.4]
  wire [63:0] regs_218_io_in; // @[RegFile.scala 66:20:@37463.4]
  wire  regs_218_io_reset; // @[RegFile.scala 66:20:@37463.4]
  wire [63:0] regs_218_io_out; // @[RegFile.scala 66:20:@37463.4]
  wire  regs_218_io_enable; // @[RegFile.scala 66:20:@37463.4]
  wire  regs_219_clock; // @[RegFile.scala 66:20:@37477.4]
  wire  regs_219_reset; // @[RegFile.scala 66:20:@37477.4]
  wire [63:0] regs_219_io_in; // @[RegFile.scala 66:20:@37477.4]
  wire  regs_219_io_reset; // @[RegFile.scala 66:20:@37477.4]
  wire [63:0] regs_219_io_out; // @[RegFile.scala 66:20:@37477.4]
  wire  regs_219_io_enable; // @[RegFile.scala 66:20:@37477.4]
  wire  regs_220_clock; // @[RegFile.scala 66:20:@37491.4]
  wire  regs_220_reset; // @[RegFile.scala 66:20:@37491.4]
  wire [63:0] regs_220_io_in; // @[RegFile.scala 66:20:@37491.4]
  wire  regs_220_io_reset; // @[RegFile.scala 66:20:@37491.4]
  wire [63:0] regs_220_io_out; // @[RegFile.scala 66:20:@37491.4]
  wire  regs_220_io_enable; // @[RegFile.scala 66:20:@37491.4]
  wire  regs_221_clock; // @[RegFile.scala 66:20:@37505.4]
  wire  regs_221_reset; // @[RegFile.scala 66:20:@37505.4]
  wire [63:0] regs_221_io_in; // @[RegFile.scala 66:20:@37505.4]
  wire  regs_221_io_reset; // @[RegFile.scala 66:20:@37505.4]
  wire [63:0] regs_221_io_out; // @[RegFile.scala 66:20:@37505.4]
  wire  regs_221_io_enable; // @[RegFile.scala 66:20:@37505.4]
  wire  regs_222_clock; // @[RegFile.scala 66:20:@37519.4]
  wire  regs_222_reset; // @[RegFile.scala 66:20:@37519.4]
  wire [63:0] regs_222_io_in; // @[RegFile.scala 66:20:@37519.4]
  wire  regs_222_io_reset; // @[RegFile.scala 66:20:@37519.4]
  wire [63:0] regs_222_io_out; // @[RegFile.scala 66:20:@37519.4]
  wire  regs_222_io_enable; // @[RegFile.scala 66:20:@37519.4]
  wire  regs_223_clock; // @[RegFile.scala 66:20:@37533.4]
  wire  regs_223_reset; // @[RegFile.scala 66:20:@37533.4]
  wire [63:0] regs_223_io_in; // @[RegFile.scala 66:20:@37533.4]
  wire  regs_223_io_reset; // @[RegFile.scala 66:20:@37533.4]
  wire [63:0] regs_223_io_out; // @[RegFile.scala 66:20:@37533.4]
  wire  regs_223_io_enable; // @[RegFile.scala 66:20:@37533.4]
  wire  regs_224_clock; // @[RegFile.scala 66:20:@37547.4]
  wire  regs_224_reset; // @[RegFile.scala 66:20:@37547.4]
  wire [63:0] regs_224_io_in; // @[RegFile.scala 66:20:@37547.4]
  wire  regs_224_io_reset; // @[RegFile.scala 66:20:@37547.4]
  wire [63:0] regs_224_io_out; // @[RegFile.scala 66:20:@37547.4]
  wire  regs_224_io_enable; // @[RegFile.scala 66:20:@37547.4]
  wire  regs_225_clock; // @[RegFile.scala 66:20:@37561.4]
  wire  regs_225_reset; // @[RegFile.scala 66:20:@37561.4]
  wire [63:0] regs_225_io_in; // @[RegFile.scala 66:20:@37561.4]
  wire  regs_225_io_reset; // @[RegFile.scala 66:20:@37561.4]
  wire [63:0] regs_225_io_out; // @[RegFile.scala 66:20:@37561.4]
  wire  regs_225_io_enable; // @[RegFile.scala 66:20:@37561.4]
  wire  regs_226_clock; // @[RegFile.scala 66:20:@37575.4]
  wire  regs_226_reset; // @[RegFile.scala 66:20:@37575.4]
  wire [63:0] regs_226_io_in; // @[RegFile.scala 66:20:@37575.4]
  wire  regs_226_io_reset; // @[RegFile.scala 66:20:@37575.4]
  wire [63:0] regs_226_io_out; // @[RegFile.scala 66:20:@37575.4]
  wire  regs_226_io_enable; // @[RegFile.scala 66:20:@37575.4]
  wire  regs_227_clock; // @[RegFile.scala 66:20:@37589.4]
  wire  regs_227_reset; // @[RegFile.scala 66:20:@37589.4]
  wire [63:0] regs_227_io_in; // @[RegFile.scala 66:20:@37589.4]
  wire  regs_227_io_reset; // @[RegFile.scala 66:20:@37589.4]
  wire [63:0] regs_227_io_out; // @[RegFile.scala 66:20:@37589.4]
  wire  regs_227_io_enable; // @[RegFile.scala 66:20:@37589.4]
  wire  regs_228_clock; // @[RegFile.scala 66:20:@37603.4]
  wire  regs_228_reset; // @[RegFile.scala 66:20:@37603.4]
  wire [63:0] regs_228_io_in; // @[RegFile.scala 66:20:@37603.4]
  wire  regs_228_io_reset; // @[RegFile.scala 66:20:@37603.4]
  wire [63:0] regs_228_io_out; // @[RegFile.scala 66:20:@37603.4]
  wire  regs_228_io_enable; // @[RegFile.scala 66:20:@37603.4]
  wire  regs_229_clock; // @[RegFile.scala 66:20:@37617.4]
  wire  regs_229_reset; // @[RegFile.scala 66:20:@37617.4]
  wire [63:0] regs_229_io_in; // @[RegFile.scala 66:20:@37617.4]
  wire  regs_229_io_reset; // @[RegFile.scala 66:20:@37617.4]
  wire [63:0] regs_229_io_out; // @[RegFile.scala 66:20:@37617.4]
  wire  regs_229_io_enable; // @[RegFile.scala 66:20:@37617.4]
  wire  regs_230_clock; // @[RegFile.scala 66:20:@37631.4]
  wire  regs_230_reset; // @[RegFile.scala 66:20:@37631.4]
  wire [63:0] regs_230_io_in; // @[RegFile.scala 66:20:@37631.4]
  wire  regs_230_io_reset; // @[RegFile.scala 66:20:@37631.4]
  wire [63:0] regs_230_io_out; // @[RegFile.scala 66:20:@37631.4]
  wire  regs_230_io_enable; // @[RegFile.scala 66:20:@37631.4]
  wire  regs_231_clock; // @[RegFile.scala 66:20:@37645.4]
  wire  regs_231_reset; // @[RegFile.scala 66:20:@37645.4]
  wire [63:0] regs_231_io_in; // @[RegFile.scala 66:20:@37645.4]
  wire  regs_231_io_reset; // @[RegFile.scala 66:20:@37645.4]
  wire [63:0] regs_231_io_out; // @[RegFile.scala 66:20:@37645.4]
  wire  regs_231_io_enable; // @[RegFile.scala 66:20:@37645.4]
  wire  regs_232_clock; // @[RegFile.scala 66:20:@37659.4]
  wire  regs_232_reset; // @[RegFile.scala 66:20:@37659.4]
  wire [63:0] regs_232_io_in; // @[RegFile.scala 66:20:@37659.4]
  wire  regs_232_io_reset; // @[RegFile.scala 66:20:@37659.4]
  wire [63:0] regs_232_io_out; // @[RegFile.scala 66:20:@37659.4]
  wire  regs_232_io_enable; // @[RegFile.scala 66:20:@37659.4]
  wire  regs_233_clock; // @[RegFile.scala 66:20:@37673.4]
  wire  regs_233_reset; // @[RegFile.scala 66:20:@37673.4]
  wire [63:0] regs_233_io_in; // @[RegFile.scala 66:20:@37673.4]
  wire  regs_233_io_reset; // @[RegFile.scala 66:20:@37673.4]
  wire [63:0] regs_233_io_out; // @[RegFile.scala 66:20:@37673.4]
  wire  regs_233_io_enable; // @[RegFile.scala 66:20:@37673.4]
  wire  regs_234_clock; // @[RegFile.scala 66:20:@37687.4]
  wire  regs_234_reset; // @[RegFile.scala 66:20:@37687.4]
  wire [63:0] regs_234_io_in; // @[RegFile.scala 66:20:@37687.4]
  wire  regs_234_io_reset; // @[RegFile.scala 66:20:@37687.4]
  wire [63:0] regs_234_io_out; // @[RegFile.scala 66:20:@37687.4]
  wire  regs_234_io_enable; // @[RegFile.scala 66:20:@37687.4]
  wire  regs_235_clock; // @[RegFile.scala 66:20:@37701.4]
  wire  regs_235_reset; // @[RegFile.scala 66:20:@37701.4]
  wire [63:0] regs_235_io_in; // @[RegFile.scala 66:20:@37701.4]
  wire  regs_235_io_reset; // @[RegFile.scala 66:20:@37701.4]
  wire [63:0] regs_235_io_out; // @[RegFile.scala 66:20:@37701.4]
  wire  regs_235_io_enable; // @[RegFile.scala 66:20:@37701.4]
  wire  regs_236_clock; // @[RegFile.scala 66:20:@37715.4]
  wire  regs_236_reset; // @[RegFile.scala 66:20:@37715.4]
  wire [63:0] regs_236_io_in; // @[RegFile.scala 66:20:@37715.4]
  wire  regs_236_io_reset; // @[RegFile.scala 66:20:@37715.4]
  wire [63:0] regs_236_io_out; // @[RegFile.scala 66:20:@37715.4]
  wire  regs_236_io_enable; // @[RegFile.scala 66:20:@37715.4]
  wire  regs_237_clock; // @[RegFile.scala 66:20:@37729.4]
  wire  regs_237_reset; // @[RegFile.scala 66:20:@37729.4]
  wire [63:0] regs_237_io_in; // @[RegFile.scala 66:20:@37729.4]
  wire  regs_237_io_reset; // @[RegFile.scala 66:20:@37729.4]
  wire [63:0] regs_237_io_out; // @[RegFile.scala 66:20:@37729.4]
  wire  regs_237_io_enable; // @[RegFile.scala 66:20:@37729.4]
  wire  regs_238_clock; // @[RegFile.scala 66:20:@37743.4]
  wire  regs_238_reset; // @[RegFile.scala 66:20:@37743.4]
  wire [63:0] regs_238_io_in; // @[RegFile.scala 66:20:@37743.4]
  wire  regs_238_io_reset; // @[RegFile.scala 66:20:@37743.4]
  wire [63:0] regs_238_io_out; // @[RegFile.scala 66:20:@37743.4]
  wire  regs_238_io_enable; // @[RegFile.scala 66:20:@37743.4]
  wire  regs_239_clock; // @[RegFile.scala 66:20:@37757.4]
  wire  regs_239_reset; // @[RegFile.scala 66:20:@37757.4]
  wire [63:0] regs_239_io_in; // @[RegFile.scala 66:20:@37757.4]
  wire  regs_239_io_reset; // @[RegFile.scala 66:20:@37757.4]
  wire [63:0] regs_239_io_out; // @[RegFile.scala 66:20:@37757.4]
  wire  regs_239_io_enable; // @[RegFile.scala 66:20:@37757.4]
  wire  regs_240_clock; // @[RegFile.scala 66:20:@37771.4]
  wire  regs_240_reset; // @[RegFile.scala 66:20:@37771.4]
  wire [63:0] regs_240_io_in; // @[RegFile.scala 66:20:@37771.4]
  wire  regs_240_io_reset; // @[RegFile.scala 66:20:@37771.4]
  wire [63:0] regs_240_io_out; // @[RegFile.scala 66:20:@37771.4]
  wire  regs_240_io_enable; // @[RegFile.scala 66:20:@37771.4]
  wire  regs_241_clock; // @[RegFile.scala 66:20:@37785.4]
  wire  regs_241_reset; // @[RegFile.scala 66:20:@37785.4]
  wire [63:0] regs_241_io_in; // @[RegFile.scala 66:20:@37785.4]
  wire  regs_241_io_reset; // @[RegFile.scala 66:20:@37785.4]
  wire [63:0] regs_241_io_out; // @[RegFile.scala 66:20:@37785.4]
  wire  regs_241_io_enable; // @[RegFile.scala 66:20:@37785.4]
  wire  regs_242_clock; // @[RegFile.scala 66:20:@37799.4]
  wire  regs_242_reset; // @[RegFile.scala 66:20:@37799.4]
  wire [63:0] regs_242_io_in; // @[RegFile.scala 66:20:@37799.4]
  wire  regs_242_io_reset; // @[RegFile.scala 66:20:@37799.4]
  wire [63:0] regs_242_io_out; // @[RegFile.scala 66:20:@37799.4]
  wire  regs_242_io_enable; // @[RegFile.scala 66:20:@37799.4]
  wire  regs_243_clock; // @[RegFile.scala 66:20:@37813.4]
  wire  regs_243_reset; // @[RegFile.scala 66:20:@37813.4]
  wire [63:0] regs_243_io_in; // @[RegFile.scala 66:20:@37813.4]
  wire  regs_243_io_reset; // @[RegFile.scala 66:20:@37813.4]
  wire [63:0] regs_243_io_out; // @[RegFile.scala 66:20:@37813.4]
  wire  regs_243_io_enable; // @[RegFile.scala 66:20:@37813.4]
  wire  regs_244_clock; // @[RegFile.scala 66:20:@37827.4]
  wire  regs_244_reset; // @[RegFile.scala 66:20:@37827.4]
  wire [63:0] regs_244_io_in; // @[RegFile.scala 66:20:@37827.4]
  wire  regs_244_io_reset; // @[RegFile.scala 66:20:@37827.4]
  wire [63:0] regs_244_io_out; // @[RegFile.scala 66:20:@37827.4]
  wire  regs_244_io_enable; // @[RegFile.scala 66:20:@37827.4]
  wire  regs_245_clock; // @[RegFile.scala 66:20:@37841.4]
  wire  regs_245_reset; // @[RegFile.scala 66:20:@37841.4]
  wire [63:0] regs_245_io_in; // @[RegFile.scala 66:20:@37841.4]
  wire  regs_245_io_reset; // @[RegFile.scala 66:20:@37841.4]
  wire [63:0] regs_245_io_out; // @[RegFile.scala 66:20:@37841.4]
  wire  regs_245_io_enable; // @[RegFile.scala 66:20:@37841.4]
  wire  regs_246_clock; // @[RegFile.scala 66:20:@37855.4]
  wire  regs_246_reset; // @[RegFile.scala 66:20:@37855.4]
  wire [63:0] regs_246_io_in; // @[RegFile.scala 66:20:@37855.4]
  wire  regs_246_io_reset; // @[RegFile.scala 66:20:@37855.4]
  wire [63:0] regs_246_io_out; // @[RegFile.scala 66:20:@37855.4]
  wire  regs_246_io_enable; // @[RegFile.scala 66:20:@37855.4]
  wire  regs_247_clock; // @[RegFile.scala 66:20:@37869.4]
  wire  regs_247_reset; // @[RegFile.scala 66:20:@37869.4]
  wire [63:0] regs_247_io_in; // @[RegFile.scala 66:20:@37869.4]
  wire  regs_247_io_reset; // @[RegFile.scala 66:20:@37869.4]
  wire [63:0] regs_247_io_out; // @[RegFile.scala 66:20:@37869.4]
  wire  regs_247_io_enable; // @[RegFile.scala 66:20:@37869.4]
  wire  regs_248_clock; // @[RegFile.scala 66:20:@37883.4]
  wire  regs_248_reset; // @[RegFile.scala 66:20:@37883.4]
  wire [63:0] regs_248_io_in; // @[RegFile.scala 66:20:@37883.4]
  wire  regs_248_io_reset; // @[RegFile.scala 66:20:@37883.4]
  wire [63:0] regs_248_io_out; // @[RegFile.scala 66:20:@37883.4]
  wire  regs_248_io_enable; // @[RegFile.scala 66:20:@37883.4]
  wire  regs_249_clock; // @[RegFile.scala 66:20:@37897.4]
  wire  regs_249_reset; // @[RegFile.scala 66:20:@37897.4]
  wire [63:0] regs_249_io_in; // @[RegFile.scala 66:20:@37897.4]
  wire  regs_249_io_reset; // @[RegFile.scala 66:20:@37897.4]
  wire [63:0] regs_249_io_out; // @[RegFile.scala 66:20:@37897.4]
  wire  regs_249_io_enable; // @[RegFile.scala 66:20:@37897.4]
  wire  regs_250_clock; // @[RegFile.scala 66:20:@37911.4]
  wire  regs_250_reset; // @[RegFile.scala 66:20:@37911.4]
  wire [63:0] regs_250_io_in; // @[RegFile.scala 66:20:@37911.4]
  wire  regs_250_io_reset; // @[RegFile.scala 66:20:@37911.4]
  wire [63:0] regs_250_io_out; // @[RegFile.scala 66:20:@37911.4]
  wire  regs_250_io_enable; // @[RegFile.scala 66:20:@37911.4]
  wire  regs_251_clock; // @[RegFile.scala 66:20:@37925.4]
  wire  regs_251_reset; // @[RegFile.scala 66:20:@37925.4]
  wire [63:0] regs_251_io_in; // @[RegFile.scala 66:20:@37925.4]
  wire  regs_251_io_reset; // @[RegFile.scala 66:20:@37925.4]
  wire [63:0] regs_251_io_out; // @[RegFile.scala 66:20:@37925.4]
  wire  regs_251_io_enable; // @[RegFile.scala 66:20:@37925.4]
  wire  regs_252_clock; // @[RegFile.scala 66:20:@37939.4]
  wire  regs_252_reset; // @[RegFile.scala 66:20:@37939.4]
  wire [63:0] regs_252_io_in; // @[RegFile.scala 66:20:@37939.4]
  wire  regs_252_io_reset; // @[RegFile.scala 66:20:@37939.4]
  wire [63:0] regs_252_io_out; // @[RegFile.scala 66:20:@37939.4]
  wire  regs_252_io_enable; // @[RegFile.scala 66:20:@37939.4]
  wire  regs_253_clock; // @[RegFile.scala 66:20:@37953.4]
  wire  regs_253_reset; // @[RegFile.scala 66:20:@37953.4]
  wire [63:0] regs_253_io_in; // @[RegFile.scala 66:20:@37953.4]
  wire  regs_253_io_reset; // @[RegFile.scala 66:20:@37953.4]
  wire [63:0] regs_253_io_out; // @[RegFile.scala 66:20:@37953.4]
  wire  regs_253_io_enable; // @[RegFile.scala 66:20:@37953.4]
  wire  regs_254_clock; // @[RegFile.scala 66:20:@37967.4]
  wire  regs_254_reset; // @[RegFile.scala 66:20:@37967.4]
  wire [63:0] regs_254_io_in; // @[RegFile.scala 66:20:@37967.4]
  wire  regs_254_io_reset; // @[RegFile.scala 66:20:@37967.4]
  wire [63:0] regs_254_io_out; // @[RegFile.scala 66:20:@37967.4]
  wire  regs_254_io_enable; // @[RegFile.scala 66:20:@37967.4]
  wire  regs_255_clock; // @[RegFile.scala 66:20:@37981.4]
  wire  regs_255_reset; // @[RegFile.scala 66:20:@37981.4]
  wire [63:0] regs_255_io_in; // @[RegFile.scala 66:20:@37981.4]
  wire  regs_255_io_reset; // @[RegFile.scala 66:20:@37981.4]
  wire [63:0] regs_255_io_out; // @[RegFile.scala 66:20:@37981.4]
  wire  regs_255_io_enable; // @[RegFile.scala 66:20:@37981.4]
  wire  regs_256_clock; // @[RegFile.scala 66:20:@37995.4]
  wire  regs_256_reset; // @[RegFile.scala 66:20:@37995.4]
  wire [63:0] regs_256_io_in; // @[RegFile.scala 66:20:@37995.4]
  wire  regs_256_io_reset; // @[RegFile.scala 66:20:@37995.4]
  wire [63:0] regs_256_io_out; // @[RegFile.scala 66:20:@37995.4]
  wire  regs_256_io_enable; // @[RegFile.scala 66:20:@37995.4]
  wire  regs_257_clock; // @[RegFile.scala 66:20:@38009.4]
  wire  regs_257_reset; // @[RegFile.scala 66:20:@38009.4]
  wire [63:0] regs_257_io_in; // @[RegFile.scala 66:20:@38009.4]
  wire  regs_257_io_reset; // @[RegFile.scala 66:20:@38009.4]
  wire [63:0] regs_257_io_out; // @[RegFile.scala 66:20:@38009.4]
  wire  regs_257_io_enable; // @[RegFile.scala 66:20:@38009.4]
  wire  regs_258_clock; // @[RegFile.scala 66:20:@38023.4]
  wire  regs_258_reset; // @[RegFile.scala 66:20:@38023.4]
  wire [63:0] regs_258_io_in; // @[RegFile.scala 66:20:@38023.4]
  wire  regs_258_io_reset; // @[RegFile.scala 66:20:@38023.4]
  wire [63:0] regs_258_io_out; // @[RegFile.scala 66:20:@38023.4]
  wire  regs_258_io_enable; // @[RegFile.scala 66:20:@38023.4]
  wire  regs_259_clock; // @[RegFile.scala 66:20:@38037.4]
  wire  regs_259_reset; // @[RegFile.scala 66:20:@38037.4]
  wire [63:0] regs_259_io_in; // @[RegFile.scala 66:20:@38037.4]
  wire  regs_259_io_reset; // @[RegFile.scala 66:20:@38037.4]
  wire [63:0] regs_259_io_out; // @[RegFile.scala 66:20:@38037.4]
  wire  regs_259_io_enable; // @[RegFile.scala 66:20:@38037.4]
  wire  regs_260_clock; // @[RegFile.scala 66:20:@38051.4]
  wire  regs_260_reset; // @[RegFile.scala 66:20:@38051.4]
  wire [63:0] regs_260_io_in; // @[RegFile.scala 66:20:@38051.4]
  wire  regs_260_io_reset; // @[RegFile.scala 66:20:@38051.4]
  wire [63:0] regs_260_io_out; // @[RegFile.scala 66:20:@38051.4]
  wire  regs_260_io_enable; // @[RegFile.scala 66:20:@38051.4]
  wire  regs_261_clock; // @[RegFile.scala 66:20:@38065.4]
  wire  regs_261_reset; // @[RegFile.scala 66:20:@38065.4]
  wire [63:0] regs_261_io_in; // @[RegFile.scala 66:20:@38065.4]
  wire  regs_261_io_reset; // @[RegFile.scala 66:20:@38065.4]
  wire [63:0] regs_261_io_out; // @[RegFile.scala 66:20:@38065.4]
  wire  regs_261_io_enable; // @[RegFile.scala 66:20:@38065.4]
  wire  regs_262_clock; // @[RegFile.scala 66:20:@38079.4]
  wire  regs_262_reset; // @[RegFile.scala 66:20:@38079.4]
  wire [63:0] regs_262_io_in; // @[RegFile.scala 66:20:@38079.4]
  wire  regs_262_io_reset; // @[RegFile.scala 66:20:@38079.4]
  wire [63:0] regs_262_io_out; // @[RegFile.scala 66:20:@38079.4]
  wire  regs_262_io_enable; // @[RegFile.scala 66:20:@38079.4]
  wire  regs_263_clock; // @[RegFile.scala 66:20:@38093.4]
  wire  regs_263_reset; // @[RegFile.scala 66:20:@38093.4]
  wire [63:0] regs_263_io_in; // @[RegFile.scala 66:20:@38093.4]
  wire  regs_263_io_reset; // @[RegFile.scala 66:20:@38093.4]
  wire [63:0] regs_263_io_out; // @[RegFile.scala 66:20:@38093.4]
  wire  regs_263_io_enable; // @[RegFile.scala 66:20:@38093.4]
  wire  regs_264_clock; // @[RegFile.scala 66:20:@38107.4]
  wire  regs_264_reset; // @[RegFile.scala 66:20:@38107.4]
  wire [63:0] regs_264_io_in; // @[RegFile.scala 66:20:@38107.4]
  wire  regs_264_io_reset; // @[RegFile.scala 66:20:@38107.4]
  wire [63:0] regs_264_io_out; // @[RegFile.scala 66:20:@38107.4]
  wire  regs_264_io_enable; // @[RegFile.scala 66:20:@38107.4]
  wire  regs_265_clock; // @[RegFile.scala 66:20:@38121.4]
  wire  regs_265_reset; // @[RegFile.scala 66:20:@38121.4]
  wire [63:0] regs_265_io_in; // @[RegFile.scala 66:20:@38121.4]
  wire  regs_265_io_reset; // @[RegFile.scala 66:20:@38121.4]
  wire [63:0] regs_265_io_out; // @[RegFile.scala 66:20:@38121.4]
  wire  regs_265_io_enable; // @[RegFile.scala 66:20:@38121.4]
  wire  regs_266_clock; // @[RegFile.scala 66:20:@38135.4]
  wire  regs_266_reset; // @[RegFile.scala 66:20:@38135.4]
  wire [63:0] regs_266_io_in; // @[RegFile.scala 66:20:@38135.4]
  wire  regs_266_io_reset; // @[RegFile.scala 66:20:@38135.4]
  wire [63:0] regs_266_io_out; // @[RegFile.scala 66:20:@38135.4]
  wire  regs_266_io_enable; // @[RegFile.scala 66:20:@38135.4]
  wire  regs_267_clock; // @[RegFile.scala 66:20:@38149.4]
  wire  regs_267_reset; // @[RegFile.scala 66:20:@38149.4]
  wire [63:0] regs_267_io_in; // @[RegFile.scala 66:20:@38149.4]
  wire  regs_267_io_reset; // @[RegFile.scala 66:20:@38149.4]
  wire [63:0] regs_267_io_out; // @[RegFile.scala 66:20:@38149.4]
  wire  regs_267_io_enable; // @[RegFile.scala 66:20:@38149.4]
  wire  regs_268_clock; // @[RegFile.scala 66:20:@38163.4]
  wire  regs_268_reset; // @[RegFile.scala 66:20:@38163.4]
  wire [63:0] regs_268_io_in; // @[RegFile.scala 66:20:@38163.4]
  wire  regs_268_io_reset; // @[RegFile.scala 66:20:@38163.4]
  wire [63:0] regs_268_io_out; // @[RegFile.scala 66:20:@38163.4]
  wire  regs_268_io_enable; // @[RegFile.scala 66:20:@38163.4]
  wire  regs_269_clock; // @[RegFile.scala 66:20:@38177.4]
  wire  regs_269_reset; // @[RegFile.scala 66:20:@38177.4]
  wire [63:0] regs_269_io_in; // @[RegFile.scala 66:20:@38177.4]
  wire  regs_269_io_reset; // @[RegFile.scala 66:20:@38177.4]
  wire [63:0] regs_269_io_out; // @[RegFile.scala 66:20:@38177.4]
  wire  regs_269_io_enable; // @[RegFile.scala 66:20:@38177.4]
  wire  regs_270_clock; // @[RegFile.scala 66:20:@38191.4]
  wire  regs_270_reset; // @[RegFile.scala 66:20:@38191.4]
  wire [63:0] regs_270_io_in; // @[RegFile.scala 66:20:@38191.4]
  wire  regs_270_io_reset; // @[RegFile.scala 66:20:@38191.4]
  wire [63:0] regs_270_io_out; // @[RegFile.scala 66:20:@38191.4]
  wire  regs_270_io_enable; // @[RegFile.scala 66:20:@38191.4]
  wire  regs_271_clock; // @[RegFile.scala 66:20:@38205.4]
  wire  regs_271_reset; // @[RegFile.scala 66:20:@38205.4]
  wire [63:0] regs_271_io_in; // @[RegFile.scala 66:20:@38205.4]
  wire  regs_271_io_reset; // @[RegFile.scala 66:20:@38205.4]
  wire [63:0] regs_271_io_out; // @[RegFile.scala 66:20:@38205.4]
  wire  regs_271_io_enable; // @[RegFile.scala 66:20:@38205.4]
  wire  regs_272_clock; // @[RegFile.scala 66:20:@38219.4]
  wire  regs_272_reset; // @[RegFile.scala 66:20:@38219.4]
  wire [63:0] regs_272_io_in; // @[RegFile.scala 66:20:@38219.4]
  wire  regs_272_io_reset; // @[RegFile.scala 66:20:@38219.4]
  wire [63:0] regs_272_io_out; // @[RegFile.scala 66:20:@38219.4]
  wire  regs_272_io_enable; // @[RegFile.scala 66:20:@38219.4]
  wire  regs_273_clock; // @[RegFile.scala 66:20:@38233.4]
  wire  regs_273_reset; // @[RegFile.scala 66:20:@38233.4]
  wire [63:0] regs_273_io_in; // @[RegFile.scala 66:20:@38233.4]
  wire  regs_273_io_reset; // @[RegFile.scala 66:20:@38233.4]
  wire [63:0] regs_273_io_out; // @[RegFile.scala 66:20:@38233.4]
  wire  regs_273_io_enable; // @[RegFile.scala 66:20:@38233.4]
  wire  regs_274_clock; // @[RegFile.scala 66:20:@38247.4]
  wire  regs_274_reset; // @[RegFile.scala 66:20:@38247.4]
  wire [63:0] regs_274_io_in; // @[RegFile.scala 66:20:@38247.4]
  wire  regs_274_io_reset; // @[RegFile.scala 66:20:@38247.4]
  wire [63:0] regs_274_io_out; // @[RegFile.scala 66:20:@38247.4]
  wire  regs_274_io_enable; // @[RegFile.scala 66:20:@38247.4]
  wire  regs_275_clock; // @[RegFile.scala 66:20:@38261.4]
  wire  regs_275_reset; // @[RegFile.scala 66:20:@38261.4]
  wire [63:0] regs_275_io_in; // @[RegFile.scala 66:20:@38261.4]
  wire  regs_275_io_reset; // @[RegFile.scala 66:20:@38261.4]
  wire [63:0] regs_275_io_out; // @[RegFile.scala 66:20:@38261.4]
  wire  regs_275_io_enable; // @[RegFile.scala 66:20:@38261.4]
  wire  regs_276_clock; // @[RegFile.scala 66:20:@38275.4]
  wire  regs_276_reset; // @[RegFile.scala 66:20:@38275.4]
  wire [63:0] regs_276_io_in; // @[RegFile.scala 66:20:@38275.4]
  wire  regs_276_io_reset; // @[RegFile.scala 66:20:@38275.4]
  wire [63:0] regs_276_io_out; // @[RegFile.scala 66:20:@38275.4]
  wire  regs_276_io_enable; // @[RegFile.scala 66:20:@38275.4]
  wire  regs_277_clock; // @[RegFile.scala 66:20:@38289.4]
  wire  regs_277_reset; // @[RegFile.scala 66:20:@38289.4]
  wire [63:0] regs_277_io_in; // @[RegFile.scala 66:20:@38289.4]
  wire  regs_277_io_reset; // @[RegFile.scala 66:20:@38289.4]
  wire [63:0] regs_277_io_out; // @[RegFile.scala 66:20:@38289.4]
  wire  regs_277_io_enable; // @[RegFile.scala 66:20:@38289.4]
  wire  regs_278_clock; // @[RegFile.scala 66:20:@38303.4]
  wire  regs_278_reset; // @[RegFile.scala 66:20:@38303.4]
  wire [63:0] regs_278_io_in; // @[RegFile.scala 66:20:@38303.4]
  wire  regs_278_io_reset; // @[RegFile.scala 66:20:@38303.4]
  wire [63:0] regs_278_io_out; // @[RegFile.scala 66:20:@38303.4]
  wire  regs_278_io_enable; // @[RegFile.scala 66:20:@38303.4]
  wire  regs_279_clock; // @[RegFile.scala 66:20:@38317.4]
  wire  regs_279_reset; // @[RegFile.scala 66:20:@38317.4]
  wire [63:0] regs_279_io_in; // @[RegFile.scala 66:20:@38317.4]
  wire  regs_279_io_reset; // @[RegFile.scala 66:20:@38317.4]
  wire [63:0] regs_279_io_out; // @[RegFile.scala 66:20:@38317.4]
  wire  regs_279_io_enable; // @[RegFile.scala 66:20:@38317.4]
  wire  regs_280_clock; // @[RegFile.scala 66:20:@38331.4]
  wire  regs_280_reset; // @[RegFile.scala 66:20:@38331.4]
  wire [63:0] regs_280_io_in; // @[RegFile.scala 66:20:@38331.4]
  wire  regs_280_io_reset; // @[RegFile.scala 66:20:@38331.4]
  wire [63:0] regs_280_io_out; // @[RegFile.scala 66:20:@38331.4]
  wire  regs_280_io_enable; // @[RegFile.scala 66:20:@38331.4]
  wire  regs_281_clock; // @[RegFile.scala 66:20:@38345.4]
  wire  regs_281_reset; // @[RegFile.scala 66:20:@38345.4]
  wire [63:0] regs_281_io_in; // @[RegFile.scala 66:20:@38345.4]
  wire  regs_281_io_reset; // @[RegFile.scala 66:20:@38345.4]
  wire [63:0] regs_281_io_out; // @[RegFile.scala 66:20:@38345.4]
  wire  regs_281_io_enable; // @[RegFile.scala 66:20:@38345.4]
  wire  regs_282_clock; // @[RegFile.scala 66:20:@38359.4]
  wire  regs_282_reset; // @[RegFile.scala 66:20:@38359.4]
  wire [63:0] regs_282_io_in; // @[RegFile.scala 66:20:@38359.4]
  wire  regs_282_io_reset; // @[RegFile.scala 66:20:@38359.4]
  wire [63:0] regs_282_io_out; // @[RegFile.scala 66:20:@38359.4]
  wire  regs_282_io_enable; // @[RegFile.scala 66:20:@38359.4]
  wire  regs_283_clock; // @[RegFile.scala 66:20:@38373.4]
  wire  regs_283_reset; // @[RegFile.scala 66:20:@38373.4]
  wire [63:0] regs_283_io_in; // @[RegFile.scala 66:20:@38373.4]
  wire  regs_283_io_reset; // @[RegFile.scala 66:20:@38373.4]
  wire [63:0] regs_283_io_out; // @[RegFile.scala 66:20:@38373.4]
  wire  regs_283_io_enable; // @[RegFile.scala 66:20:@38373.4]
  wire  regs_284_clock; // @[RegFile.scala 66:20:@38387.4]
  wire  regs_284_reset; // @[RegFile.scala 66:20:@38387.4]
  wire [63:0] regs_284_io_in; // @[RegFile.scala 66:20:@38387.4]
  wire  regs_284_io_reset; // @[RegFile.scala 66:20:@38387.4]
  wire [63:0] regs_284_io_out; // @[RegFile.scala 66:20:@38387.4]
  wire  regs_284_io_enable; // @[RegFile.scala 66:20:@38387.4]
  wire  regs_285_clock; // @[RegFile.scala 66:20:@38401.4]
  wire  regs_285_reset; // @[RegFile.scala 66:20:@38401.4]
  wire [63:0] regs_285_io_in; // @[RegFile.scala 66:20:@38401.4]
  wire  regs_285_io_reset; // @[RegFile.scala 66:20:@38401.4]
  wire [63:0] regs_285_io_out; // @[RegFile.scala 66:20:@38401.4]
  wire  regs_285_io_enable; // @[RegFile.scala 66:20:@38401.4]
  wire  regs_286_clock; // @[RegFile.scala 66:20:@38415.4]
  wire  regs_286_reset; // @[RegFile.scala 66:20:@38415.4]
  wire [63:0] regs_286_io_in; // @[RegFile.scala 66:20:@38415.4]
  wire  regs_286_io_reset; // @[RegFile.scala 66:20:@38415.4]
  wire [63:0] regs_286_io_out; // @[RegFile.scala 66:20:@38415.4]
  wire  regs_286_io_enable; // @[RegFile.scala 66:20:@38415.4]
  wire  regs_287_clock; // @[RegFile.scala 66:20:@38429.4]
  wire  regs_287_reset; // @[RegFile.scala 66:20:@38429.4]
  wire [63:0] regs_287_io_in; // @[RegFile.scala 66:20:@38429.4]
  wire  regs_287_io_reset; // @[RegFile.scala 66:20:@38429.4]
  wire [63:0] regs_287_io_out; // @[RegFile.scala 66:20:@38429.4]
  wire  regs_287_io_enable; // @[RegFile.scala 66:20:@38429.4]
  wire  regs_288_clock; // @[RegFile.scala 66:20:@38443.4]
  wire  regs_288_reset; // @[RegFile.scala 66:20:@38443.4]
  wire [63:0] regs_288_io_in; // @[RegFile.scala 66:20:@38443.4]
  wire  regs_288_io_reset; // @[RegFile.scala 66:20:@38443.4]
  wire [63:0] regs_288_io_out; // @[RegFile.scala 66:20:@38443.4]
  wire  regs_288_io_enable; // @[RegFile.scala 66:20:@38443.4]
  wire  regs_289_clock; // @[RegFile.scala 66:20:@38457.4]
  wire  regs_289_reset; // @[RegFile.scala 66:20:@38457.4]
  wire [63:0] regs_289_io_in; // @[RegFile.scala 66:20:@38457.4]
  wire  regs_289_io_reset; // @[RegFile.scala 66:20:@38457.4]
  wire [63:0] regs_289_io_out; // @[RegFile.scala 66:20:@38457.4]
  wire  regs_289_io_enable; // @[RegFile.scala 66:20:@38457.4]
  wire  regs_290_clock; // @[RegFile.scala 66:20:@38471.4]
  wire  regs_290_reset; // @[RegFile.scala 66:20:@38471.4]
  wire [63:0] regs_290_io_in; // @[RegFile.scala 66:20:@38471.4]
  wire  regs_290_io_reset; // @[RegFile.scala 66:20:@38471.4]
  wire [63:0] regs_290_io_out; // @[RegFile.scala 66:20:@38471.4]
  wire  regs_290_io_enable; // @[RegFile.scala 66:20:@38471.4]
  wire  regs_291_clock; // @[RegFile.scala 66:20:@38485.4]
  wire  regs_291_reset; // @[RegFile.scala 66:20:@38485.4]
  wire [63:0] regs_291_io_in; // @[RegFile.scala 66:20:@38485.4]
  wire  regs_291_io_reset; // @[RegFile.scala 66:20:@38485.4]
  wire [63:0] regs_291_io_out; // @[RegFile.scala 66:20:@38485.4]
  wire  regs_291_io_enable; // @[RegFile.scala 66:20:@38485.4]
  wire  regs_292_clock; // @[RegFile.scala 66:20:@38499.4]
  wire  regs_292_reset; // @[RegFile.scala 66:20:@38499.4]
  wire [63:0] regs_292_io_in; // @[RegFile.scala 66:20:@38499.4]
  wire  regs_292_io_reset; // @[RegFile.scala 66:20:@38499.4]
  wire [63:0] regs_292_io_out; // @[RegFile.scala 66:20:@38499.4]
  wire  regs_292_io_enable; // @[RegFile.scala 66:20:@38499.4]
  wire  regs_293_clock; // @[RegFile.scala 66:20:@38513.4]
  wire  regs_293_reset; // @[RegFile.scala 66:20:@38513.4]
  wire [63:0] regs_293_io_in; // @[RegFile.scala 66:20:@38513.4]
  wire  regs_293_io_reset; // @[RegFile.scala 66:20:@38513.4]
  wire [63:0] regs_293_io_out; // @[RegFile.scala 66:20:@38513.4]
  wire  regs_293_io_enable; // @[RegFile.scala 66:20:@38513.4]
  wire  regs_294_clock; // @[RegFile.scala 66:20:@38527.4]
  wire  regs_294_reset; // @[RegFile.scala 66:20:@38527.4]
  wire [63:0] regs_294_io_in; // @[RegFile.scala 66:20:@38527.4]
  wire  regs_294_io_reset; // @[RegFile.scala 66:20:@38527.4]
  wire [63:0] regs_294_io_out; // @[RegFile.scala 66:20:@38527.4]
  wire  regs_294_io_enable; // @[RegFile.scala 66:20:@38527.4]
  wire  regs_295_clock; // @[RegFile.scala 66:20:@38541.4]
  wire  regs_295_reset; // @[RegFile.scala 66:20:@38541.4]
  wire [63:0] regs_295_io_in; // @[RegFile.scala 66:20:@38541.4]
  wire  regs_295_io_reset; // @[RegFile.scala 66:20:@38541.4]
  wire [63:0] regs_295_io_out; // @[RegFile.scala 66:20:@38541.4]
  wire  regs_295_io_enable; // @[RegFile.scala 66:20:@38541.4]
  wire  regs_296_clock; // @[RegFile.scala 66:20:@38555.4]
  wire  regs_296_reset; // @[RegFile.scala 66:20:@38555.4]
  wire [63:0] regs_296_io_in; // @[RegFile.scala 66:20:@38555.4]
  wire  regs_296_io_reset; // @[RegFile.scala 66:20:@38555.4]
  wire [63:0] regs_296_io_out; // @[RegFile.scala 66:20:@38555.4]
  wire  regs_296_io_enable; // @[RegFile.scala 66:20:@38555.4]
  wire  regs_297_clock; // @[RegFile.scala 66:20:@38569.4]
  wire  regs_297_reset; // @[RegFile.scala 66:20:@38569.4]
  wire [63:0] regs_297_io_in; // @[RegFile.scala 66:20:@38569.4]
  wire  regs_297_io_reset; // @[RegFile.scala 66:20:@38569.4]
  wire [63:0] regs_297_io_out; // @[RegFile.scala 66:20:@38569.4]
  wire  regs_297_io_enable; // @[RegFile.scala 66:20:@38569.4]
  wire  regs_298_clock; // @[RegFile.scala 66:20:@38583.4]
  wire  regs_298_reset; // @[RegFile.scala 66:20:@38583.4]
  wire [63:0] regs_298_io_in; // @[RegFile.scala 66:20:@38583.4]
  wire  regs_298_io_reset; // @[RegFile.scala 66:20:@38583.4]
  wire [63:0] regs_298_io_out; // @[RegFile.scala 66:20:@38583.4]
  wire  regs_298_io_enable; // @[RegFile.scala 66:20:@38583.4]
  wire  regs_299_clock; // @[RegFile.scala 66:20:@38597.4]
  wire  regs_299_reset; // @[RegFile.scala 66:20:@38597.4]
  wire [63:0] regs_299_io_in; // @[RegFile.scala 66:20:@38597.4]
  wire  regs_299_io_reset; // @[RegFile.scala 66:20:@38597.4]
  wire [63:0] regs_299_io_out; // @[RegFile.scala 66:20:@38597.4]
  wire  regs_299_io_enable; // @[RegFile.scala 66:20:@38597.4]
  wire  regs_300_clock; // @[RegFile.scala 66:20:@38611.4]
  wire  regs_300_reset; // @[RegFile.scala 66:20:@38611.4]
  wire [63:0] regs_300_io_in; // @[RegFile.scala 66:20:@38611.4]
  wire  regs_300_io_reset; // @[RegFile.scala 66:20:@38611.4]
  wire [63:0] regs_300_io_out; // @[RegFile.scala 66:20:@38611.4]
  wire  regs_300_io_enable; // @[RegFile.scala 66:20:@38611.4]
  wire  regs_301_clock; // @[RegFile.scala 66:20:@38625.4]
  wire  regs_301_reset; // @[RegFile.scala 66:20:@38625.4]
  wire [63:0] regs_301_io_in; // @[RegFile.scala 66:20:@38625.4]
  wire  regs_301_io_reset; // @[RegFile.scala 66:20:@38625.4]
  wire [63:0] regs_301_io_out; // @[RegFile.scala 66:20:@38625.4]
  wire  regs_301_io_enable; // @[RegFile.scala 66:20:@38625.4]
  wire  regs_302_clock; // @[RegFile.scala 66:20:@38639.4]
  wire  regs_302_reset; // @[RegFile.scala 66:20:@38639.4]
  wire [63:0] regs_302_io_in; // @[RegFile.scala 66:20:@38639.4]
  wire  regs_302_io_reset; // @[RegFile.scala 66:20:@38639.4]
  wire [63:0] regs_302_io_out; // @[RegFile.scala 66:20:@38639.4]
  wire  regs_302_io_enable; // @[RegFile.scala 66:20:@38639.4]
  wire  regs_303_clock; // @[RegFile.scala 66:20:@38653.4]
  wire  regs_303_reset; // @[RegFile.scala 66:20:@38653.4]
  wire [63:0] regs_303_io_in; // @[RegFile.scala 66:20:@38653.4]
  wire  regs_303_io_reset; // @[RegFile.scala 66:20:@38653.4]
  wire [63:0] regs_303_io_out; // @[RegFile.scala 66:20:@38653.4]
  wire  regs_303_io_enable; // @[RegFile.scala 66:20:@38653.4]
  wire  regs_304_clock; // @[RegFile.scala 66:20:@38667.4]
  wire  regs_304_reset; // @[RegFile.scala 66:20:@38667.4]
  wire [63:0] regs_304_io_in; // @[RegFile.scala 66:20:@38667.4]
  wire  regs_304_io_reset; // @[RegFile.scala 66:20:@38667.4]
  wire [63:0] regs_304_io_out; // @[RegFile.scala 66:20:@38667.4]
  wire  regs_304_io_enable; // @[RegFile.scala 66:20:@38667.4]
  wire  regs_305_clock; // @[RegFile.scala 66:20:@38681.4]
  wire  regs_305_reset; // @[RegFile.scala 66:20:@38681.4]
  wire [63:0] regs_305_io_in; // @[RegFile.scala 66:20:@38681.4]
  wire  regs_305_io_reset; // @[RegFile.scala 66:20:@38681.4]
  wire [63:0] regs_305_io_out; // @[RegFile.scala 66:20:@38681.4]
  wire  regs_305_io_enable; // @[RegFile.scala 66:20:@38681.4]
  wire  regs_306_clock; // @[RegFile.scala 66:20:@38695.4]
  wire  regs_306_reset; // @[RegFile.scala 66:20:@38695.4]
  wire [63:0] regs_306_io_in; // @[RegFile.scala 66:20:@38695.4]
  wire  regs_306_io_reset; // @[RegFile.scala 66:20:@38695.4]
  wire [63:0] regs_306_io_out; // @[RegFile.scala 66:20:@38695.4]
  wire  regs_306_io_enable; // @[RegFile.scala 66:20:@38695.4]
  wire  regs_307_clock; // @[RegFile.scala 66:20:@38709.4]
  wire  regs_307_reset; // @[RegFile.scala 66:20:@38709.4]
  wire [63:0] regs_307_io_in; // @[RegFile.scala 66:20:@38709.4]
  wire  regs_307_io_reset; // @[RegFile.scala 66:20:@38709.4]
  wire [63:0] regs_307_io_out; // @[RegFile.scala 66:20:@38709.4]
  wire  regs_307_io_enable; // @[RegFile.scala 66:20:@38709.4]
  wire  regs_308_clock; // @[RegFile.scala 66:20:@38723.4]
  wire  regs_308_reset; // @[RegFile.scala 66:20:@38723.4]
  wire [63:0] regs_308_io_in; // @[RegFile.scala 66:20:@38723.4]
  wire  regs_308_io_reset; // @[RegFile.scala 66:20:@38723.4]
  wire [63:0] regs_308_io_out; // @[RegFile.scala 66:20:@38723.4]
  wire  regs_308_io_enable; // @[RegFile.scala 66:20:@38723.4]
  wire  regs_309_clock; // @[RegFile.scala 66:20:@38737.4]
  wire  regs_309_reset; // @[RegFile.scala 66:20:@38737.4]
  wire [63:0] regs_309_io_in; // @[RegFile.scala 66:20:@38737.4]
  wire  regs_309_io_reset; // @[RegFile.scala 66:20:@38737.4]
  wire [63:0] regs_309_io_out; // @[RegFile.scala 66:20:@38737.4]
  wire  regs_309_io_enable; // @[RegFile.scala 66:20:@38737.4]
  wire  regs_310_clock; // @[RegFile.scala 66:20:@38751.4]
  wire  regs_310_reset; // @[RegFile.scala 66:20:@38751.4]
  wire [63:0] regs_310_io_in; // @[RegFile.scala 66:20:@38751.4]
  wire  regs_310_io_reset; // @[RegFile.scala 66:20:@38751.4]
  wire [63:0] regs_310_io_out; // @[RegFile.scala 66:20:@38751.4]
  wire  regs_310_io_enable; // @[RegFile.scala 66:20:@38751.4]
  wire  regs_311_clock; // @[RegFile.scala 66:20:@38765.4]
  wire  regs_311_reset; // @[RegFile.scala 66:20:@38765.4]
  wire [63:0] regs_311_io_in; // @[RegFile.scala 66:20:@38765.4]
  wire  regs_311_io_reset; // @[RegFile.scala 66:20:@38765.4]
  wire [63:0] regs_311_io_out; // @[RegFile.scala 66:20:@38765.4]
  wire  regs_311_io_enable; // @[RegFile.scala 66:20:@38765.4]
  wire  regs_312_clock; // @[RegFile.scala 66:20:@38779.4]
  wire  regs_312_reset; // @[RegFile.scala 66:20:@38779.4]
  wire [63:0] regs_312_io_in; // @[RegFile.scala 66:20:@38779.4]
  wire  regs_312_io_reset; // @[RegFile.scala 66:20:@38779.4]
  wire [63:0] regs_312_io_out; // @[RegFile.scala 66:20:@38779.4]
  wire  regs_312_io_enable; // @[RegFile.scala 66:20:@38779.4]
  wire  regs_313_clock; // @[RegFile.scala 66:20:@38793.4]
  wire  regs_313_reset; // @[RegFile.scala 66:20:@38793.4]
  wire [63:0] regs_313_io_in; // @[RegFile.scala 66:20:@38793.4]
  wire  regs_313_io_reset; // @[RegFile.scala 66:20:@38793.4]
  wire [63:0] regs_313_io_out; // @[RegFile.scala 66:20:@38793.4]
  wire  regs_313_io_enable; // @[RegFile.scala 66:20:@38793.4]
  wire  regs_314_clock; // @[RegFile.scala 66:20:@38807.4]
  wire  regs_314_reset; // @[RegFile.scala 66:20:@38807.4]
  wire [63:0] regs_314_io_in; // @[RegFile.scala 66:20:@38807.4]
  wire  regs_314_io_reset; // @[RegFile.scala 66:20:@38807.4]
  wire [63:0] regs_314_io_out; // @[RegFile.scala 66:20:@38807.4]
  wire  regs_314_io_enable; // @[RegFile.scala 66:20:@38807.4]
  wire  regs_315_clock; // @[RegFile.scala 66:20:@38821.4]
  wire  regs_315_reset; // @[RegFile.scala 66:20:@38821.4]
  wire [63:0] regs_315_io_in; // @[RegFile.scala 66:20:@38821.4]
  wire  regs_315_io_reset; // @[RegFile.scala 66:20:@38821.4]
  wire [63:0] regs_315_io_out; // @[RegFile.scala 66:20:@38821.4]
  wire  regs_315_io_enable; // @[RegFile.scala 66:20:@38821.4]
  wire  regs_316_clock; // @[RegFile.scala 66:20:@38835.4]
  wire  regs_316_reset; // @[RegFile.scala 66:20:@38835.4]
  wire [63:0] regs_316_io_in; // @[RegFile.scala 66:20:@38835.4]
  wire  regs_316_io_reset; // @[RegFile.scala 66:20:@38835.4]
  wire [63:0] regs_316_io_out; // @[RegFile.scala 66:20:@38835.4]
  wire  regs_316_io_enable; // @[RegFile.scala 66:20:@38835.4]
  wire  regs_317_clock; // @[RegFile.scala 66:20:@38849.4]
  wire  regs_317_reset; // @[RegFile.scala 66:20:@38849.4]
  wire [63:0] regs_317_io_in; // @[RegFile.scala 66:20:@38849.4]
  wire  regs_317_io_reset; // @[RegFile.scala 66:20:@38849.4]
  wire [63:0] regs_317_io_out; // @[RegFile.scala 66:20:@38849.4]
  wire  regs_317_io_enable; // @[RegFile.scala 66:20:@38849.4]
  wire  regs_318_clock; // @[RegFile.scala 66:20:@38863.4]
  wire  regs_318_reset; // @[RegFile.scala 66:20:@38863.4]
  wire [63:0] regs_318_io_in; // @[RegFile.scala 66:20:@38863.4]
  wire  regs_318_io_reset; // @[RegFile.scala 66:20:@38863.4]
  wire [63:0] regs_318_io_out; // @[RegFile.scala 66:20:@38863.4]
  wire  regs_318_io_enable; // @[RegFile.scala 66:20:@38863.4]
  wire  regs_319_clock; // @[RegFile.scala 66:20:@38877.4]
  wire  regs_319_reset; // @[RegFile.scala 66:20:@38877.4]
  wire [63:0] regs_319_io_in; // @[RegFile.scala 66:20:@38877.4]
  wire  regs_319_io_reset; // @[RegFile.scala 66:20:@38877.4]
  wire [63:0] regs_319_io_out; // @[RegFile.scala 66:20:@38877.4]
  wire  regs_319_io_enable; // @[RegFile.scala 66:20:@38877.4]
  wire  regs_320_clock; // @[RegFile.scala 66:20:@38891.4]
  wire  regs_320_reset; // @[RegFile.scala 66:20:@38891.4]
  wire [63:0] regs_320_io_in; // @[RegFile.scala 66:20:@38891.4]
  wire  regs_320_io_reset; // @[RegFile.scala 66:20:@38891.4]
  wire [63:0] regs_320_io_out; // @[RegFile.scala 66:20:@38891.4]
  wire  regs_320_io_enable; // @[RegFile.scala 66:20:@38891.4]
  wire  regs_321_clock; // @[RegFile.scala 66:20:@38905.4]
  wire  regs_321_reset; // @[RegFile.scala 66:20:@38905.4]
  wire [63:0] regs_321_io_in; // @[RegFile.scala 66:20:@38905.4]
  wire  regs_321_io_reset; // @[RegFile.scala 66:20:@38905.4]
  wire [63:0] regs_321_io_out; // @[RegFile.scala 66:20:@38905.4]
  wire  regs_321_io_enable; // @[RegFile.scala 66:20:@38905.4]
  wire  regs_322_clock; // @[RegFile.scala 66:20:@38919.4]
  wire  regs_322_reset; // @[RegFile.scala 66:20:@38919.4]
  wire [63:0] regs_322_io_in; // @[RegFile.scala 66:20:@38919.4]
  wire  regs_322_io_reset; // @[RegFile.scala 66:20:@38919.4]
  wire [63:0] regs_322_io_out; // @[RegFile.scala 66:20:@38919.4]
  wire  regs_322_io_enable; // @[RegFile.scala 66:20:@38919.4]
  wire  regs_323_clock; // @[RegFile.scala 66:20:@38933.4]
  wire  regs_323_reset; // @[RegFile.scala 66:20:@38933.4]
  wire [63:0] regs_323_io_in; // @[RegFile.scala 66:20:@38933.4]
  wire  regs_323_io_reset; // @[RegFile.scala 66:20:@38933.4]
  wire [63:0] regs_323_io_out; // @[RegFile.scala 66:20:@38933.4]
  wire  regs_323_io_enable; // @[RegFile.scala 66:20:@38933.4]
  wire  regs_324_clock; // @[RegFile.scala 66:20:@38947.4]
  wire  regs_324_reset; // @[RegFile.scala 66:20:@38947.4]
  wire [63:0] regs_324_io_in; // @[RegFile.scala 66:20:@38947.4]
  wire  regs_324_io_reset; // @[RegFile.scala 66:20:@38947.4]
  wire [63:0] regs_324_io_out; // @[RegFile.scala 66:20:@38947.4]
  wire  regs_324_io_enable; // @[RegFile.scala 66:20:@38947.4]
  wire  regs_325_clock; // @[RegFile.scala 66:20:@38961.4]
  wire  regs_325_reset; // @[RegFile.scala 66:20:@38961.4]
  wire [63:0] regs_325_io_in; // @[RegFile.scala 66:20:@38961.4]
  wire  regs_325_io_reset; // @[RegFile.scala 66:20:@38961.4]
  wire [63:0] regs_325_io_out; // @[RegFile.scala 66:20:@38961.4]
  wire  regs_325_io_enable; // @[RegFile.scala 66:20:@38961.4]
  wire  regs_326_clock; // @[RegFile.scala 66:20:@38975.4]
  wire  regs_326_reset; // @[RegFile.scala 66:20:@38975.4]
  wire [63:0] regs_326_io_in; // @[RegFile.scala 66:20:@38975.4]
  wire  regs_326_io_reset; // @[RegFile.scala 66:20:@38975.4]
  wire [63:0] regs_326_io_out; // @[RegFile.scala 66:20:@38975.4]
  wire  regs_326_io_enable; // @[RegFile.scala 66:20:@38975.4]
  wire  regs_327_clock; // @[RegFile.scala 66:20:@38989.4]
  wire  regs_327_reset; // @[RegFile.scala 66:20:@38989.4]
  wire [63:0] regs_327_io_in; // @[RegFile.scala 66:20:@38989.4]
  wire  regs_327_io_reset; // @[RegFile.scala 66:20:@38989.4]
  wire [63:0] regs_327_io_out; // @[RegFile.scala 66:20:@38989.4]
  wire  regs_327_io_enable; // @[RegFile.scala 66:20:@38989.4]
  wire  regs_328_clock; // @[RegFile.scala 66:20:@39003.4]
  wire  regs_328_reset; // @[RegFile.scala 66:20:@39003.4]
  wire [63:0] regs_328_io_in; // @[RegFile.scala 66:20:@39003.4]
  wire  regs_328_io_reset; // @[RegFile.scala 66:20:@39003.4]
  wire [63:0] regs_328_io_out; // @[RegFile.scala 66:20:@39003.4]
  wire  regs_328_io_enable; // @[RegFile.scala 66:20:@39003.4]
  wire  regs_329_clock; // @[RegFile.scala 66:20:@39017.4]
  wire  regs_329_reset; // @[RegFile.scala 66:20:@39017.4]
  wire [63:0] regs_329_io_in; // @[RegFile.scala 66:20:@39017.4]
  wire  regs_329_io_reset; // @[RegFile.scala 66:20:@39017.4]
  wire [63:0] regs_329_io_out; // @[RegFile.scala 66:20:@39017.4]
  wire  regs_329_io_enable; // @[RegFile.scala 66:20:@39017.4]
  wire  regs_330_clock; // @[RegFile.scala 66:20:@39031.4]
  wire  regs_330_reset; // @[RegFile.scala 66:20:@39031.4]
  wire [63:0] regs_330_io_in; // @[RegFile.scala 66:20:@39031.4]
  wire  regs_330_io_reset; // @[RegFile.scala 66:20:@39031.4]
  wire [63:0] regs_330_io_out; // @[RegFile.scala 66:20:@39031.4]
  wire  regs_330_io_enable; // @[RegFile.scala 66:20:@39031.4]
  wire  regs_331_clock; // @[RegFile.scala 66:20:@39045.4]
  wire  regs_331_reset; // @[RegFile.scala 66:20:@39045.4]
  wire [63:0] regs_331_io_in; // @[RegFile.scala 66:20:@39045.4]
  wire  regs_331_io_reset; // @[RegFile.scala 66:20:@39045.4]
  wire [63:0] regs_331_io_out; // @[RegFile.scala 66:20:@39045.4]
  wire  regs_331_io_enable; // @[RegFile.scala 66:20:@39045.4]
  wire  regs_332_clock; // @[RegFile.scala 66:20:@39059.4]
  wire  regs_332_reset; // @[RegFile.scala 66:20:@39059.4]
  wire [63:0] regs_332_io_in; // @[RegFile.scala 66:20:@39059.4]
  wire  regs_332_io_reset; // @[RegFile.scala 66:20:@39059.4]
  wire [63:0] regs_332_io_out; // @[RegFile.scala 66:20:@39059.4]
  wire  regs_332_io_enable; // @[RegFile.scala 66:20:@39059.4]
  wire  regs_333_clock; // @[RegFile.scala 66:20:@39073.4]
  wire  regs_333_reset; // @[RegFile.scala 66:20:@39073.4]
  wire [63:0] regs_333_io_in; // @[RegFile.scala 66:20:@39073.4]
  wire  regs_333_io_reset; // @[RegFile.scala 66:20:@39073.4]
  wire [63:0] regs_333_io_out; // @[RegFile.scala 66:20:@39073.4]
  wire  regs_333_io_enable; // @[RegFile.scala 66:20:@39073.4]
  wire  regs_334_clock; // @[RegFile.scala 66:20:@39087.4]
  wire  regs_334_reset; // @[RegFile.scala 66:20:@39087.4]
  wire [63:0] regs_334_io_in; // @[RegFile.scala 66:20:@39087.4]
  wire  regs_334_io_reset; // @[RegFile.scala 66:20:@39087.4]
  wire [63:0] regs_334_io_out; // @[RegFile.scala 66:20:@39087.4]
  wire  regs_334_io_enable; // @[RegFile.scala 66:20:@39087.4]
  wire  regs_335_clock; // @[RegFile.scala 66:20:@39101.4]
  wire  regs_335_reset; // @[RegFile.scala 66:20:@39101.4]
  wire [63:0] regs_335_io_in; // @[RegFile.scala 66:20:@39101.4]
  wire  regs_335_io_reset; // @[RegFile.scala 66:20:@39101.4]
  wire [63:0] regs_335_io_out; // @[RegFile.scala 66:20:@39101.4]
  wire  regs_335_io_enable; // @[RegFile.scala 66:20:@39101.4]
  wire  regs_336_clock; // @[RegFile.scala 66:20:@39115.4]
  wire  regs_336_reset; // @[RegFile.scala 66:20:@39115.4]
  wire [63:0] regs_336_io_in; // @[RegFile.scala 66:20:@39115.4]
  wire  regs_336_io_reset; // @[RegFile.scala 66:20:@39115.4]
  wire [63:0] regs_336_io_out; // @[RegFile.scala 66:20:@39115.4]
  wire  regs_336_io_enable; // @[RegFile.scala 66:20:@39115.4]
  wire  regs_337_clock; // @[RegFile.scala 66:20:@39129.4]
  wire  regs_337_reset; // @[RegFile.scala 66:20:@39129.4]
  wire [63:0] regs_337_io_in; // @[RegFile.scala 66:20:@39129.4]
  wire  regs_337_io_reset; // @[RegFile.scala 66:20:@39129.4]
  wire [63:0] regs_337_io_out; // @[RegFile.scala 66:20:@39129.4]
  wire  regs_337_io_enable; // @[RegFile.scala 66:20:@39129.4]
  wire  regs_338_clock; // @[RegFile.scala 66:20:@39143.4]
  wire  regs_338_reset; // @[RegFile.scala 66:20:@39143.4]
  wire [63:0] regs_338_io_in; // @[RegFile.scala 66:20:@39143.4]
  wire  regs_338_io_reset; // @[RegFile.scala 66:20:@39143.4]
  wire [63:0] regs_338_io_out; // @[RegFile.scala 66:20:@39143.4]
  wire  regs_338_io_enable; // @[RegFile.scala 66:20:@39143.4]
  wire  regs_339_clock; // @[RegFile.scala 66:20:@39157.4]
  wire  regs_339_reset; // @[RegFile.scala 66:20:@39157.4]
  wire [63:0] regs_339_io_in; // @[RegFile.scala 66:20:@39157.4]
  wire  regs_339_io_reset; // @[RegFile.scala 66:20:@39157.4]
  wire [63:0] regs_339_io_out; // @[RegFile.scala 66:20:@39157.4]
  wire  regs_339_io_enable; // @[RegFile.scala 66:20:@39157.4]
  wire  regs_340_clock; // @[RegFile.scala 66:20:@39171.4]
  wire  regs_340_reset; // @[RegFile.scala 66:20:@39171.4]
  wire [63:0] regs_340_io_in; // @[RegFile.scala 66:20:@39171.4]
  wire  regs_340_io_reset; // @[RegFile.scala 66:20:@39171.4]
  wire [63:0] regs_340_io_out; // @[RegFile.scala 66:20:@39171.4]
  wire  regs_340_io_enable; // @[RegFile.scala 66:20:@39171.4]
  wire  regs_341_clock; // @[RegFile.scala 66:20:@39185.4]
  wire  regs_341_reset; // @[RegFile.scala 66:20:@39185.4]
  wire [63:0] regs_341_io_in; // @[RegFile.scala 66:20:@39185.4]
  wire  regs_341_io_reset; // @[RegFile.scala 66:20:@39185.4]
  wire [63:0] regs_341_io_out; // @[RegFile.scala 66:20:@39185.4]
  wire  regs_341_io_enable; // @[RegFile.scala 66:20:@39185.4]
  wire  regs_342_clock; // @[RegFile.scala 66:20:@39199.4]
  wire  regs_342_reset; // @[RegFile.scala 66:20:@39199.4]
  wire [63:0] regs_342_io_in; // @[RegFile.scala 66:20:@39199.4]
  wire  regs_342_io_reset; // @[RegFile.scala 66:20:@39199.4]
  wire [63:0] regs_342_io_out; // @[RegFile.scala 66:20:@39199.4]
  wire  regs_342_io_enable; // @[RegFile.scala 66:20:@39199.4]
  wire  regs_343_clock; // @[RegFile.scala 66:20:@39213.4]
  wire  regs_343_reset; // @[RegFile.scala 66:20:@39213.4]
  wire [63:0] regs_343_io_in; // @[RegFile.scala 66:20:@39213.4]
  wire  regs_343_io_reset; // @[RegFile.scala 66:20:@39213.4]
  wire [63:0] regs_343_io_out; // @[RegFile.scala 66:20:@39213.4]
  wire  regs_343_io_enable; // @[RegFile.scala 66:20:@39213.4]
  wire  regs_344_clock; // @[RegFile.scala 66:20:@39227.4]
  wire  regs_344_reset; // @[RegFile.scala 66:20:@39227.4]
  wire [63:0] regs_344_io_in; // @[RegFile.scala 66:20:@39227.4]
  wire  regs_344_io_reset; // @[RegFile.scala 66:20:@39227.4]
  wire [63:0] regs_344_io_out; // @[RegFile.scala 66:20:@39227.4]
  wire  regs_344_io_enable; // @[RegFile.scala 66:20:@39227.4]
  wire  regs_345_clock; // @[RegFile.scala 66:20:@39241.4]
  wire  regs_345_reset; // @[RegFile.scala 66:20:@39241.4]
  wire [63:0] regs_345_io_in; // @[RegFile.scala 66:20:@39241.4]
  wire  regs_345_io_reset; // @[RegFile.scala 66:20:@39241.4]
  wire [63:0] regs_345_io_out; // @[RegFile.scala 66:20:@39241.4]
  wire  regs_345_io_enable; // @[RegFile.scala 66:20:@39241.4]
  wire  regs_346_clock; // @[RegFile.scala 66:20:@39255.4]
  wire  regs_346_reset; // @[RegFile.scala 66:20:@39255.4]
  wire [63:0] regs_346_io_in; // @[RegFile.scala 66:20:@39255.4]
  wire  regs_346_io_reset; // @[RegFile.scala 66:20:@39255.4]
  wire [63:0] regs_346_io_out; // @[RegFile.scala 66:20:@39255.4]
  wire  regs_346_io_enable; // @[RegFile.scala 66:20:@39255.4]
  wire  regs_347_clock; // @[RegFile.scala 66:20:@39269.4]
  wire  regs_347_reset; // @[RegFile.scala 66:20:@39269.4]
  wire [63:0] regs_347_io_in; // @[RegFile.scala 66:20:@39269.4]
  wire  regs_347_io_reset; // @[RegFile.scala 66:20:@39269.4]
  wire [63:0] regs_347_io_out; // @[RegFile.scala 66:20:@39269.4]
  wire  regs_347_io_enable; // @[RegFile.scala 66:20:@39269.4]
  wire  regs_348_clock; // @[RegFile.scala 66:20:@39283.4]
  wire  regs_348_reset; // @[RegFile.scala 66:20:@39283.4]
  wire [63:0] regs_348_io_in; // @[RegFile.scala 66:20:@39283.4]
  wire  regs_348_io_reset; // @[RegFile.scala 66:20:@39283.4]
  wire [63:0] regs_348_io_out; // @[RegFile.scala 66:20:@39283.4]
  wire  regs_348_io_enable; // @[RegFile.scala 66:20:@39283.4]
  wire  regs_349_clock; // @[RegFile.scala 66:20:@39297.4]
  wire  regs_349_reset; // @[RegFile.scala 66:20:@39297.4]
  wire [63:0] regs_349_io_in; // @[RegFile.scala 66:20:@39297.4]
  wire  regs_349_io_reset; // @[RegFile.scala 66:20:@39297.4]
  wire [63:0] regs_349_io_out; // @[RegFile.scala 66:20:@39297.4]
  wire  regs_349_io_enable; // @[RegFile.scala 66:20:@39297.4]
  wire  regs_350_clock; // @[RegFile.scala 66:20:@39311.4]
  wire  regs_350_reset; // @[RegFile.scala 66:20:@39311.4]
  wire [63:0] regs_350_io_in; // @[RegFile.scala 66:20:@39311.4]
  wire  regs_350_io_reset; // @[RegFile.scala 66:20:@39311.4]
  wire [63:0] regs_350_io_out; // @[RegFile.scala 66:20:@39311.4]
  wire  regs_350_io_enable; // @[RegFile.scala 66:20:@39311.4]
  wire  regs_351_clock; // @[RegFile.scala 66:20:@39325.4]
  wire  regs_351_reset; // @[RegFile.scala 66:20:@39325.4]
  wire [63:0] regs_351_io_in; // @[RegFile.scala 66:20:@39325.4]
  wire  regs_351_io_reset; // @[RegFile.scala 66:20:@39325.4]
  wire [63:0] regs_351_io_out; // @[RegFile.scala 66:20:@39325.4]
  wire  regs_351_io_enable; // @[RegFile.scala 66:20:@39325.4]
  wire  regs_352_clock; // @[RegFile.scala 66:20:@39339.4]
  wire  regs_352_reset; // @[RegFile.scala 66:20:@39339.4]
  wire [63:0] regs_352_io_in; // @[RegFile.scala 66:20:@39339.4]
  wire  regs_352_io_reset; // @[RegFile.scala 66:20:@39339.4]
  wire [63:0] regs_352_io_out; // @[RegFile.scala 66:20:@39339.4]
  wire  regs_352_io_enable; // @[RegFile.scala 66:20:@39339.4]
  wire  regs_353_clock; // @[RegFile.scala 66:20:@39353.4]
  wire  regs_353_reset; // @[RegFile.scala 66:20:@39353.4]
  wire [63:0] regs_353_io_in; // @[RegFile.scala 66:20:@39353.4]
  wire  regs_353_io_reset; // @[RegFile.scala 66:20:@39353.4]
  wire [63:0] regs_353_io_out; // @[RegFile.scala 66:20:@39353.4]
  wire  regs_353_io_enable; // @[RegFile.scala 66:20:@39353.4]
  wire  regs_354_clock; // @[RegFile.scala 66:20:@39367.4]
  wire  regs_354_reset; // @[RegFile.scala 66:20:@39367.4]
  wire [63:0] regs_354_io_in; // @[RegFile.scala 66:20:@39367.4]
  wire  regs_354_io_reset; // @[RegFile.scala 66:20:@39367.4]
  wire [63:0] regs_354_io_out; // @[RegFile.scala 66:20:@39367.4]
  wire  regs_354_io_enable; // @[RegFile.scala 66:20:@39367.4]
  wire  regs_355_clock; // @[RegFile.scala 66:20:@39381.4]
  wire  regs_355_reset; // @[RegFile.scala 66:20:@39381.4]
  wire [63:0] regs_355_io_in; // @[RegFile.scala 66:20:@39381.4]
  wire  regs_355_io_reset; // @[RegFile.scala 66:20:@39381.4]
  wire [63:0] regs_355_io_out; // @[RegFile.scala 66:20:@39381.4]
  wire  regs_355_io_enable; // @[RegFile.scala 66:20:@39381.4]
  wire  regs_356_clock; // @[RegFile.scala 66:20:@39395.4]
  wire  regs_356_reset; // @[RegFile.scala 66:20:@39395.4]
  wire [63:0] regs_356_io_in; // @[RegFile.scala 66:20:@39395.4]
  wire  regs_356_io_reset; // @[RegFile.scala 66:20:@39395.4]
  wire [63:0] regs_356_io_out; // @[RegFile.scala 66:20:@39395.4]
  wire  regs_356_io_enable; // @[RegFile.scala 66:20:@39395.4]
  wire  regs_357_clock; // @[RegFile.scala 66:20:@39409.4]
  wire  regs_357_reset; // @[RegFile.scala 66:20:@39409.4]
  wire [63:0] regs_357_io_in; // @[RegFile.scala 66:20:@39409.4]
  wire  regs_357_io_reset; // @[RegFile.scala 66:20:@39409.4]
  wire [63:0] regs_357_io_out; // @[RegFile.scala 66:20:@39409.4]
  wire  regs_357_io_enable; // @[RegFile.scala 66:20:@39409.4]
  wire  regs_358_clock; // @[RegFile.scala 66:20:@39423.4]
  wire  regs_358_reset; // @[RegFile.scala 66:20:@39423.4]
  wire [63:0] regs_358_io_in; // @[RegFile.scala 66:20:@39423.4]
  wire  regs_358_io_reset; // @[RegFile.scala 66:20:@39423.4]
  wire [63:0] regs_358_io_out; // @[RegFile.scala 66:20:@39423.4]
  wire  regs_358_io_enable; // @[RegFile.scala 66:20:@39423.4]
  wire  regs_359_clock; // @[RegFile.scala 66:20:@39437.4]
  wire  regs_359_reset; // @[RegFile.scala 66:20:@39437.4]
  wire [63:0] regs_359_io_in; // @[RegFile.scala 66:20:@39437.4]
  wire  regs_359_io_reset; // @[RegFile.scala 66:20:@39437.4]
  wire [63:0] regs_359_io_out; // @[RegFile.scala 66:20:@39437.4]
  wire  regs_359_io_enable; // @[RegFile.scala 66:20:@39437.4]
  wire  regs_360_clock; // @[RegFile.scala 66:20:@39451.4]
  wire  regs_360_reset; // @[RegFile.scala 66:20:@39451.4]
  wire [63:0] regs_360_io_in; // @[RegFile.scala 66:20:@39451.4]
  wire  regs_360_io_reset; // @[RegFile.scala 66:20:@39451.4]
  wire [63:0] regs_360_io_out; // @[RegFile.scala 66:20:@39451.4]
  wire  regs_360_io_enable; // @[RegFile.scala 66:20:@39451.4]
  wire  regs_361_clock; // @[RegFile.scala 66:20:@39465.4]
  wire  regs_361_reset; // @[RegFile.scala 66:20:@39465.4]
  wire [63:0] regs_361_io_in; // @[RegFile.scala 66:20:@39465.4]
  wire  regs_361_io_reset; // @[RegFile.scala 66:20:@39465.4]
  wire [63:0] regs_361_io_out; // @[RegFile.scala 66:20:@39465.4]
  wire  regs_361_io_enable; // @[RegFile.scala 66:20:@39465.4]
  wire  regs_362_clock; // @[RegFile.scala 66:20:@39479.4]
  wire  regs_362_reset; // @[RegFile.scala 66:20:@39479.4]
  wire [63:0] regs_362_io_in; // @[RegFile.scala 66:20:@39479.4]
  wire  regs_362_io_reset; // @[RegFile.scala 66:20:@39479.4]
  wire [63:0] regs_362_io_out; // @[RegFile.scala 66:20:@39479.4]
  wire  regs_362_io_enable; // @[RegFile.scala 66:20:@39479.4]
  wire  regs_363_clock; // @[RegFile.scala 66:20:@39493.4]
  wire  regs_363_reset; // @[RegFile.scala 66:20:@39493.4]
  wire [63:0] regs_363_io_in; // @[RegFile.scala 66:20:@39493.4]
  wire  regs_363_io_reset; // @[RegFile.scala 66:20:@39493.4]
  wire [63:0] regs_363_io_out; // @[RegFile.scala 66:20:@39493.4]
  wire  regs_363_io_enable; // @[RegFile.scala 66:20:@39493.4]
  wire  regs_364_clock; // @[RegFile.scala 66:20:@39507.4]
  wire  regs_364_reset; // @[RegFile.scala 66:20:@39507.4]
  wire [63:0] regs_364_io_in; // @[RegFile.scala 66:20:@39507.4]
  wire  regs_364_io_reset; // @[RegFile.scala 66:20:@39507.4]
  wire [63:0] regs_364_io_out; // @[RegFile.scala 66:20:@39507.4]
  wire  regs_364_io_enable; // @[RegFile.scala 66:20:@39507.4]
  wire  regs_365_clock; // @[RegFile.scala 66:20:@39521.4]
  wire  regs_365_reset; // @[RegFile.scala 66:20:@39521.4]
  wire [63:0] regs_365_io_in; // @[RegFile.scala 66:20:@39521.4]
  wire  regs_365_io_reset; // @[RegFile.scala 66:20:@39521.4]
  wire [63:0] regs_365_io_out; // @[RegFile.scala 66:20:@39521.4]
  wire  regs_365_io_enable; // @[RegFile.scala 66:20:@39521.4]
  wire  regs_366_clock; // @[RegFile.scala 66:20:@39535.4]
  wire  regs_366_reset; // @[RegFile.scala 66:20:@39535.4]
  wire [63:0] regs_366_io_in; // @[RegFile.scala 66:20:@39535.4]
  wire  regs_366_io_reset; // @[RegFile.scala 66:20:@39535.4]
  wire [63:0] regs_366_io_out; // @[RegFile.scala 66:20:@39535.4]
  wire  regs_366_io_enable; // @[RegFile.scala 66:20:@39535.4]
  wire  regs_367_clock; // @[RegFile.scala 66:20:@39549.4]
  wire  regs_367_reset; // @[RegFile.scala 66:20:@39549.4]
  wire [63:0] regs_367_io_in; // @[RegFile.scala 66:20:@39549.4]
  wire  regs_367_io_reset; // @[RegFile.scala 66:20:@39549.4]
  wire [63:0] regs_367_io_out; // @[RegFile.scala 66:20:@39549.4]
  wire  regs_367_io_enable; // @[RegFile.scala 66:20:@39549.4]
  wire  regs_368_clock; // @[RegFile.scala 66:20:@39563.4]
  wire  regs_368_reset; // @[RegFile.scala 66:20:@39563.4]
  wire [63:0] regs_368_io_in; // @[RegFile.scala 66:20:@39563.4]
  wire  regs_368_io_reset; // @[RegFile.scala 66:20:@39563.4]
  wire [63:0] regs_368_io_out; // @[RegFile.scala 66:20:@39563.4]
  wire  regs_368_io_enable; // @[RegFile.scala 66:20:@39563.4]
  wire  regs_369_clock; // @[RegFile.scala 66:20:@39577.4]
  wire  regs_369_reset; // @[RegFile.scala 66:20:@39577.4]
  wire [63:0] regs_369_io_in; // @[RegFile.scala 66:20:@39577.4]
  wire  regs_369_io_reset; // @[RegFile.scala 66:20:@39577.4]
  wire [63:0] regs_369_io_out; // @[RegFile.scala 66:20:@39577.4]
  wire  regs_369_io_enable; // @[RegFile.scala 66:20:@39577.4]
  wire  regs_370_clock; // @[RegFile.scala 66:20:@39591.4]
  wire  regs_370_reset; // @[RegFile.scala 66:20:@39591.4]
  wire [63:0] regs_370_io_in; // @[RegFile.scala 66:20:@39591.4]
  wire  regs_370_io_reset; // @[RegFile.scala 66:20:@39591.4]
  wire [63:0] regs_370_io_out; // @[RegFile.scala 66:20:@39591.4]
  wire  regs_370_io_enable; // @[RegFile.scala 66:20:@39591.4]
  wire  regs_371_clock; // @[RegFile.scala 66:20:@39605.4]
  wire  regs_371_reset; // @[RegFile.scala 66:20:@39605.4]
  wire [63:0] regs_371_io_in; // @[RegFile.scala 66:20:@39605.4]
  wire  regs_371_io_reset; // @[RegFile.scala 66:20:@39605.4]
  wire [63:0] regs_371_io_out; // @[RegFile.scala 66:20:@39605.4]
  wire  regs_371_io_enable; // @[RegFile.scala 66:20:@39605.4]
  wire  regs_372_clock; // @[RegFile.scala 66:20:@39619.4]
  wire  regs_372_reset; // @[RegFile.scala 66:20:@39619.4]
  wire [63:0] regs_372_io_in; // @[RegFile.scala 66:20:@39619.4]
  wire  regs_372_io_reset; // @[RegFile.scala 66:20:@39619.4]
  wire [63:0] regs_372_io_out; // @[RegFile.scala 66:20:@39619.4]
  wire  regs_372_io_enable; // @[RegFile.scala 66:20:@39619.4]
  wire  regs_373_clock; // @[RegFile.scala 66:20:@39633.4]
  wire  regs_373_reset; // @[RegFile.scala 66:20:@39633.4]
  wire [63:0] regs_373_io_in; // @[RegFile.scala 66:20:@39633.4]
  wire  regs_373_io_reset; // @[RegFile.scala 66:20:@39633.4]
  wire [63:0] regs_373_io_out; // @[RegFile.scala 66:20:@39633.4]
  wire  regs_373_io_enable; // @[RegFile.scala 66:20:@39633.4]
  wire  regs_374_clock; // @[RegFile.scala 66:20:@39647.4]
  wire  regs_374_reset; // @[RegFile.scala 66:20:@39647.4]
  wire [63:0] regs_374_io_in; // @[RegFile.scala 66:20:@39647.4]
  wire  regs_374_io_reset; // @[RegFile.scala 66:20:@39647.4]
  wire [63:0] regs_374_io_out; // @[RegFile.scala 66:20:@39647.4]
  wire  regs_374_io_enable; // @[RegFile.scala 66:20:@39647.4]
  wire  regs_375_clock; // @[RegFile.scala 66:20:@39661.4]
  wire  regs_375_reset; // @[RegFile.scala 66:20:@39661.4]
  wire [63:0] regs_375_io_in; // @[RegFile.scala 66:20:@39661.4]
  wire  regs_375_io_reset; // @[RegFile.scala 66:20:@39661.4]
  wire [63:0] regs_375_io_out; // @[RegFile.scala 66:20:@39661.4]
  wire  regs_375_io_enable; // @[RegFile.scala 66:20:@39661.4]
  wire  regs_376_clock; // @[RegFile.scala 66:20:@39675.4]
  wire  regs_376_reset; // @[RegFile.scala 66:20:@39675.4]
  wire [63:0] regs_376_io_in; // @[RegFile.scala 66:20:@39675.4]
  wire  regs_376_io_reset; // @[RegFile.scala 66:20:@39675.4]
  wire [63:0] regs_376_io_out; // @[RegFile.scala 66:20:@39675.4]
  wire  regs_376_io_enable; // @[RegFile.scala 66:20:@39675.4]
  wire  regs_377_clock; // @[RegFile.scala 66:20:@39689.4]
  wire  regs_377_reset; // @[RegFile.scala 66:20:@39689.4]
  wire [63:0] regs_377_io_in; // @[RegFile.scala 66:20:@39689.4]
  wire  regs_377_io_reset; // @[RegFile.scala 66:20:@39689.4]
  wire [63:0] regs_377_io_out; // @[RegFile.scala 66:20:@39689.4]
  wire  regs_377_io_enable; // @[RegFile.scala 66:20:@39689.4]
  wire  regs_378_clock; // @[RegFile.scala 66:20:@39703.4]
  wire  regs_378_reset; // @[RegFile.scala 66:20:@39703.4]
  wire [63:0] regs_378_io_in; // @[RegFile.scala 66:20:@39703.4]
  wire  regs_378_io_reset; // @[RegFile.scala 66:20:@39703.4]
  wire [63:0] regs_378_io_out; // @[RegFile.scala 66:20:@39703.4]
  wire  regs_378_io_enable; // @[RegFile.scala 66:20:@39703.4]
  wire  regs_379_clock; // @[RegFile.scala 66:20:@39717.4]
  wire  regs_379_reset; // @[RegFile.scala 66:20:@39717.4]
  wire [63:0] regs_379_io_in; // @[RegFile.scala 66:20:@39717.4]
  wire  regs_379_io_reset; // @[RegFile.scala 66:20:@39717.4]
  wire [63:0] regs_379_io_out; // @[RegFile.scala 66:20:@39717.4]
  wire  regs_379_io_enable; // @[RegFile.scala 66:20:@39717.4]
  wire  regs_380_clock; // @[RegFile.scala 66:20:@39731.4]
  wire  regs_380_reset; // @[RegFile.scala 66:20:@39731.4]
  wire [63:0] regs_380_io_in; // @[RegFile.scala 66:20:@39731.4]
  wire  regs_380_io_reset; // @[RegFile.scala 66:20:@39731.4]
  wire [63:0] regs_380_io_out; // @[RegFile.scala 66:20:@39731.4]
  wire  regs_380_io_enable; // @[RegFile.scala 66:20:@39731.4]
  wire  regs_381_clock; // @[RegFile.scala 66:20:@39745.4]
  wire  regs_381_reset; // @[RegFile.scala 66:20:@39745.4]
  wire [63:0] regs_381_io_in; // @[RegFile.scala 66:20:@39745.4]
  wire  regs_381_io_reset; // @[RegFile.scala 66:20:@39745.4]
  wire [63:0] regs_381_io_out; // @[RegFile.scala 66:20:@39745.4]
  wire  regs_381_io_enable; // @[RegFile.scala 66:20:@39745.4]
  wire  regs_382_clock; // @[RegFile.scala 66:20:@39759.4]
  wire  regs_382_reset; // @[RegFile.scala 66:20:@39759.4]
  wire [63:0] regs_382_io_in; // @[RegFile.scala 66:20:@39759.4]
  wire  regs_382_io_reset; // @[RegFile.scala 66:20:@39759.4]
  wire [63:0] regs_382_io_out; // @[RegFile.scala 66:20:@39759.4]
  wire  regs_382_io_enable; // @[RegFile.scala 66:20:@39759.4]
  wire  regs_383_clock; // @[RegFile.scala 66:20:@39773.4]
  wire  regs_383_reset; // @[RegFile.scala 66:20:@39773.4]
  wire [63:0] regs_383_io_in; // @[RegFile.scala 66:20:@39773.4]
  wire  regs_383_io_reset; // @[RegFile.scala 66:20:@39773.4]
  wire [63:0] regs_383_io_out; // @[RegFile.scala 66:20:@39773.4]
  wire  regs_383_io_enable; // @[RegFile.scala 66:20:@39773.4]
  wire  regs_384_clock; // @[RegFile.scala 66:20:@39787.4]
  wire  regs_384_reset; // @[RegFile.scala 66:20:@39787.4]
  wire [63:0] regs_384_io_in; // @[RegFile.scala 66:20:@39787.4]
  wire  regs_384_io_reset; // @[RegFile.scala 66:20:@39787.4]
  wire [63:0] regs_384_io_out; // @[RegFile.scala 66:20:@39787.4]
  wire  regs_384_io_enable; // @[RegFile.scala 66:20:@39787.4]
  wire  regs_385_clock; // @[RegFile.scala 66:20:@39801.4]
  wire  regs_385_reset; // @[RegFile.scala 66:20:@39801.4]
  wire [63:0] regs_385_io_in; // @[RegFile.scala 66:20:@39801.4]
  wire  regs_385_io_reset; // @[RegFile.scala 66:20:@39801.4]
  wire [63:0] regs_385_io_out; // @[RegFile.scala 66:20:@39801.4]
  wire  regs_385_io_enable; // @[RegFile.scala 66:20:@39801.4]
  wire  regs_386_clock; // @[RegFile.scala 66:20:@39815.4]
  wire  regs_386_reset; // @[RegFile.scala 66:20:@39815.4]
  wire [63:0] regs_386_io_in; // @[RegFile.scala 66:20:@39815.4]
  wire  regs_386_io_reset; // @[RegFile.scala 66:20:@39815.4]
  wire [63:0] regs_386_io_out; // @[RegFile.scala 66:20:@39815.4]
  wire  regs_386_io_enable; // @[RegFile.scala 66:20:@39815.4]
  wire  regs_387_clock; // @[RegFile.scala 66:20:@39829.4]
  wire  regs_387_reset; // @[RegFile.scala 66:20:@39829.4]
  wire [63:0] regs_387_io_in; // @[RegFile.scala 66:20:@39829.4]
  wire  regs_387_io_reset; // @[RegFile.scala 66:20:@39829.4]
  wire [63:0] regs_387_io_out; // @[RegFile.scala 66:20:@39829.4]
  wire  regs_387_io_enable; // @[RegFile.scala 66:20:@39829.4]
  wire  regs_388_clock; // @[RegFile.scala 66:20:@39843.4]
  wire  regs_388_reset; // @[RegFile.scala 66:20:@39843.4]
  wire [63:0] regs_388_io_in; // @[RegFile.scala 66:20:@39843.4]
  wire  regs_388_io_reset; // @[RegFile.scala 66:20:@39843.4]
  wire [63:0] regs_388_io_out; // @[RegFile.scala 66:20:@39843.4]
  wire  regs_388_io_enable; // @[RegFile.scala 66:20:@39843.4]
  wire  regs_389_clock; // @[RegFile.scala 66:20:@39857.4]
  wire  regs_389_reset; // @[RegFile.scala 66:20:@39857.4]
  wire [63:0] regs_389_io_in; // @[RegFile.scala 66:20:@39857.4]
  wire  regs_389_io_reset; // @[RegFile.scala 66:20:@39857.4]
  wire [63:0] regs_389_io_out; // @[RegFile.scala 66:20:@39857.4]
  wire  regs_389_io_enable; // @[RegFile.scala 66:20:@39857.4]
  wire  regs_390_clock; // @[RegFile.scala 66:20:@39871.4]
  wire  regs_390_reset; // @[RegFile.scala 66:20:@39871.4]
  wire [63:0] regs_390_io_in; // @[RegFile.scala 66:20:@39871.4]
  wire  regs_390_io_reset; // @[RegFile.scala 66:20:@39871.4]
  wire [63:0] regs_390_io_out; // @[RegFile.scala 66:20:@39871.4]
  wire  regs_390_io_enable; // @[RegFile.scala 66:20:@39871.4]
  wire  regs_391_clock; // @[RegFile.scala 66:20:@39885.4]
  wire  regs_391_reset; // @[RegFile.scala 66:20:@39885.4]
  wire [63:0] regs_391_io_in; // @[RegFile.scala 66:20:@39885.4]
  wire  regs_391_io_reset; // @[RegFile.scala 66:20:@39885.4]
  wire [63:0] regs_391_io_out; // @[RegFile.scala 66:20:@39885.4]
  wire  regs_391_io_enable; // @[RegFile.scala 66:20:@39885.4]
  wire  regs_392_clock; // @[RegFile.scala 66:20:@39899.4]
  wire  regs_392_reset; // @[RegFile.scala 66:20:@39899.4]
  wire [63:0] regs_392_io_in; // @[RegFile.scala 66:20:@39899.4]
  wire  regs_392_io_reset; // @[RegFile.scala 66:20:@39899.4]
  wire [63:0] regs_392_io_out; // @[RegFile.scala 66:20:@39899.4]
  wire  regs_392_io_enable; // @[RegFile.scala 66:20:@39899.4]
  wire  regs_393_clock; // @[RegFile.scala 66:20:@39913.4]
  wire  regs_393_reset; // @[RegFile.scala 66:20:@39913.4]
  wire [63:0] regs_393_io_in; // @[RegFile.scala 66:20:@39913.4]
  wire  regs_393_io_reset; // @[RegFile.scala 66:20:@39913.4]
  wire [63:0] regs_393_io_out; // @[RegFile.scala 66:20:@39913.4]
  wire  regs_393_io_enable; // @[RegFile.scala 66:20:@39913.4]
  wire  regs_394_clock; // @[RegFile.scala 66:20:@39927.4]
  wire  regs_394_reset; // @[RegFile.scala 66:20:@39927.4]
  wire [63:0] regs_394_io_in; // @[RegFile.scala 66:20:@39927.4]
  wire  regs_394_io_reset; // @[RegFile.scala 66:20:@39927.4]
  wire [63:0] regs_394_io_out; // @[RegFile.scala 66:20:@39927.4]
  wire  regs_394_io_enable; // @[RegFile.scala 66:20:@39927.4]
  wire  regs_395_clock; // @[RegFile.scala 66:20:@39941.4]
  wire  regs_395_reset; // @[RegFile.scala 66:20:@39941.4]
  wire [63:0] regs_395_io_in; // @[RegFile.scala 66:20:@39941.4]
  wire  regs_395_io_reset; // @[RegFile.scala 66:20:@39941.4]
  wire [63:0] regs_395_io_out; // @[RegFile.scala 66:20:@39941.4]
  wire  regs_395_io_enable; // @[RegFile.scala 66:20:@39941.4]
  wire  regs_396_clock; // @[RegFile.scala 66:20:@39955.4]
  wire  regs_396_reset; // @[RegFile.scala 66:20:@39955.4]
  wire [63:0] regs_396_io_in; // @[RegFile.scala 66:20:@39955.4]
  wire  regs_396_io_reset; // @[RegFile.scala 66:20:@39955.4]
  wire [63:0] regs_396_io_out; // @[RegFile.scala 66:20:@39955.4]
  wire  regs_396_io_enable; // @[RegFile.scala 66:20:@39955.4]
  wire  regs_397_clock; // @[RegFile.scala 66:20:@39969.4]
  wire  regs_397_reset; // @[RegFile.scala 66:20:@39969.4]
  wire [63:0] regs_397_io_in; // @[RegFile.scala 66:20:@39969.4]
  wire  regs_397_io_reset; // @[RegFile.scala 66:20:@39969.4]
  wire [63:0] regs_397_io_out; // @[RegFile.scala 66:20:@39969.4]
  wire  regs_397_io_enable; // @[RegFile.scala 66:20:@39969.4]
  wire  regs_398_clock; // @[RegFile.scala 66:20:@39983.4]
  wire  regs_398_reset; // @[RegFile.scala 66:20:@39983.4]
  wire [63:0] regs_398_io_in; // @[RegFile.scala 66:20:@39983.4]
  wire  regs_398_io_reset; // @[RegFile.scala 66:20:@39983.4]
  wire [63:0] regs_398_io_out; // @[RegFile.scala 66:20:@39983.4]
  wire  regs_398_io_enable; // @[RegFile.scala 66:20:@39983.4]
  wire  regs_399_clock; // @[RegFile.scala 66:20:@39997.4]
  wire  regs_399_reset; // @[RegFile.scala 66:20:@39997.4]
  wire [63:0] regs_399_io_in; // @[RegFile.scala 66:20:@39997.4]
  wire  regs_399_io_reset; // @[RegFile.scala 66:20:@39997.4]
  wire [63:0] regs_399_io_out; // @[RegFile.scala 66:20:@39997.4]
  wire  regs_399_io_enable; // @[RegFile.scala 66:20:@39997.4]
  wire  regs_400_clock; // @[RegFile.scala 66:20:@40011.4]
  wire  regs_400_reset; // @[RegFile.scala 66:20:@40011.4]
  wire [63:0] regs_400_io_in; // @[RegFile.scala 66:20:@40011.4]
  wire  regs_400_io_reset; // @[RegFile.scala 66:20:@40011.4]
  wire [63:0] regs_400_io_out; // @[RegFile.scala 66:20:@40011.4]
  wire  regs_400_io_enable; // @[RegFile.scala 66:20:@40011.4]
  wire  regs_401_clock; // @[RegFile.scala 66:20:@40025.4]
  wire  regs_401_reset; // @[RegFile.scala 66:20:@40025.4]
  wire [63:0] regs_401_io_in; // @[RegFile.scala 66:20:@40025.4]
  wire  regs_401_io_reset; // @[RegFile.scala 66:20:@40025.4]
  wire [63:0] regs_401_io_out; // @[RegFile.scala 66:20:@40025.4]
  wire  regs_401_io_enable; // @[RegFile.scala 66:20:@40025.4]
  wire  regs_402_clock; // @[RegFile.scala 66:20:@40039.4]
  wire  regs_402_reset; // @[RegFile.scala 66:20:@40039.4]
  wire [63:0] regs_402_io_in; // @[RegFile.scala 66:20:@40039.4]
  wire  regs_402_io_reset; // @[RegFile.scala 66:20:@40039.4]
  wire [63:0] regs_402_io_out; // @[RegFile.scala 66:20:@40039.4]
  wire  regs_402_io_enable; // @[RegFile.scala 66:20:@40039.4]
  wire  regs_403_clock; // @[RegFile.scala 66:20:@40053.4]
  wire  regs_403_reset; // @[RegFile.scala 66:20:@40053.4]
  wire [63:0] regs_403_io_in; // @[RegFile.scala 66:20:@40053.4]
  wire  regs_403_io_reset; // @[RegFile.scala 66:20:@40053.4]
  wire [63:0] regs_403_io_out; // @[RegFile.scala 66:20:@40053.4]
  wire  regs_403_io_enable; // @[RegFile.scala 66:20:@40053.4]
  wire  regs_404_clock; // @[RegFile.scala 66:20:@40067.4]
  wire  regs_404_reset; // @[RegFile.scala 66:20:@40067.4]
  wire [63:0] regs_404_io_in; // @[RegFile.scala 66:20:@40067.4]
  wire  regs_404_io_reset; // @[RegFile.scala 66:20:@40067.4]
  wire [63:0] regs_404_io_out; // @[RegFile.scala 66:20:@40067.4]
  wire  regs_404_io_enable; // @[RegFile.scala 66:20:@40067.4]
  wire  regs_405_clock; // @[RegFile.scala 66:20:@40081.4]
  wire  regs_405_reset; // @[RegFile.scala 66:20:@40081.4]
  wire [63:0] regs_405_io_in; // @[RegFile.scala 66:20:@40081.4]
  wire  regs_405_io_reset; // @[RegFile.scala 66:20:@40081.4]
  wire [63:0] regs_405_io_out; // @[RegFile.scala 66:20:@40081.4]
  wire  regs_405_io_enable; // @[RegFile.scala 66:20:@40081.4]
  wire  regs_406_clock; // @[RegFile.scala 66:20:@40095.4]
  wire  regs_406_reset; // @[RegFile.scala 66:20:@40095.4]
  wire [63:0] regs_406_io_in; // @[RegFile.scala 66:20:@40095.4]
  wire  regs_406_io_reset; // @[RegFile.scala 66:20:@40095.4]
  wire [63:0] regs_406_io_out; // @[RegFile.scala 66:20:@40095.4]
  wire  regs_406_io_enable; // @[RegFile.scala 66:20:@40095.4]
  wire  regs_407_clock; // @[RegFile.scala 66:20:@40109.4]
  wire  regs_407_reset; // @[RegFile.scala 66:20:@40109.4]
  wire [63:0] regs_407_io_in; // @[RegFile.scala 66:20:@40109.4]
  wire  regs_407_io_reset; // @[RegFile.scala 66:20:@40109.4]
  wire [63:0] regs_407_io_out; // @[RegFile.scala 66:20:@40109.4]
  wire  regs_407_io_enable; // @[RegFile.scala 66:20:@40109.4]
  wire  regs_408_clock; // @[RegFile.scala 66:20:@40123.4]
  wire  regs_408_reset; // @[RegFile.scala 66:20:@40123.4]
  wire [63:0] regs_408_io_in; // @[RegFile.scala 66:20:@40123.4]
  wire  regs_408_io_reset; // @[RegFile.scala 66:20:@40123.4]
  wire [63:0] regs_408_io_out; // @[RegFile.scala 66:20:@40123.4]
  wire  regs_408_io_enable; // @[RegFile.scala 66:20:@40123.4]
  wire  regs_409_clock; // @[RegFile.scala 66:20:@40137.4]
  wire  regs_409_reset; // @[RegFile.scala 66:20:@40137.4]
  wire [63:0] regs_409_io_in; // @[RegFile.scala 66:20:@40137.4]
  wire  regs_409_io_reset; // @[RegFile.scala 66:20:@40137.4]
  wire [63:0] regs_409_io_out; // @[RegFile.scala 66:20:@40137.4]
  wire  regs_409_io_enable; // @[RegFile.scala 66:20:@40137.4]
  wire  regs_410_clock; // @[RegFile.scala 66:20:@40151.4]
  wire  regs_410_reset; // @[RegFile.scala 66:20:@40151.4]
  wire [63:0] regs_410_io_in; // @[RegFile.scala 66:20:@40151.4]
  wire  regs_410_io_reset; // @[RegFile.scala 66:20:@40151.4]
  wire [63:0] regs_410_io_out; // @[RegFile.scala 66:20:@40151.4]
  wire  regs_410_io_enable; // @[RegFile.scala 66:20:@40151.4]
  wire  regs_411_clock; // @[RegFile.scala 66:20:@40165.4]
  wire  regs_411_reset; // @[RegFile.scala 66:20:@40165.4]
  wire [63:0] regs_411_io_in; // @[RegFile.scala 66:20:@40165.4]
  wire  regs_411_io_reset; // @[RegFile.scala 66:20:@40165.4]
  wire [63:0] regs_411_io_out; // @[RegFile.scala 66:20:@40165.4]
  wire  regs_411_io_enable; // @[RegFile.scala 66:20:@40165.4]
  wire  regs_412_clock; // @[RegFile.scala 66:20:@40179.4]
  wire  regs_412_reset; // @[RegFile.scala 66:20:@40179.4]
  wire [63:0] regs_412_io_in; // @[RegFile.scala 66:20:@40179.4]
  wire  regs_412_io_reset; // @[RegFile.scala 66:20:@40179.4]
  wire [63:0] regs_412_io_out; // @[RegFile.scala 66:20:@40179.4]
  wire  regs_412_io_enable; // @[RegFile.scala 66:20:@40179.4]
  wire  regs_413_clock; // @[RegFile.scala 66:20:@40193.4]
  wire  regs_413_reset; // @[RegFile.scala 66:20:@40193.4]
  wire [63:0] regs_413_io_in; // @[RegFile.scala 66:20:@40193.4]
  wire  regs_413_io_reset; // @[RegFile.scala 66:20:@40193.4]
  wire [63:0] regs_413_io_out; // @[RegFile.scala 66:20:@40193.4]
  wire  regs_413_io_enable; // @[RegFile.scala 66:20:@40193.4]
  wire  regs_414_clock; // @[RegFile.scala 66:20:@40207.4]
  wire  regs_414_reset; // @[RegFile.scala 66:20:@40207.4]
  wire [63:0] regs_414_io_in; // @[RegFile.scala 66:20:@40207.4]
  wire  regs_414_io_reset; // @[RegFile.scala 66:20:@40207.4]
  wire [63:0] regs_414_io_out; // @[RegFile.scala 66:20:@40207.4]
  wire  regs_414_io_enable; // @[RegFile.scala 66:20:@40207.4]
  wire  regs_415_clock; // @[RegFile.scala 66:20:@40221.4]
  wire  regs_415_reset; // @[RegFile.scala 66:20:@40221.4]
  wire [63:0] regs_415_io_in; // @[RegFile.scala 66:20:@40221.4]
  wire  regs_415_io_reset; // @[RegFile.scala 66:20:@40221.4]
  wire [63:0] regs_415_io_out; // @[RegFile.scala 66:20:@40221.4]
  wire  regs_415_io_enable; // @[RegFile.scala 66:20:@40221.4]
  wire  regs_416_clock; // @[RegFile.scala 66:20:@40235.4]
  wire  regs_416_reset; // @[RegFile.scala 66:20:@40235.4]
  wire [63:0] regs_416_io_in; // @[RegFile.scala 66:20:@40235.4]
  wire  regs_416_io_reset; // @[RegFile.scala 66:20:@40235.4]
  wire [63:0] regs_416_io_out; // @[RegFile.scala 66:20:@40235.4]
  wire  regs_416_io_enable; // @[RegFile.scala 66:20:@40235.4]
  wire  regs_417_clock; // @[RegFile.scala 66:20:@40249.4]
  wire  regs_417_reset; // @[RegFile.scala 66:20:@40249.4]
  wire [63:0] regs_417_io_in; // @[RegFile.scala 66:20:@40249.4]
  wire  regs_417_io_reset; // @[RegFile.scala 66:20:@40249.4]
  wire [63:0] regs_417_io_out; // @[RegFile.scala 66:20:@40249.4]
  wire  regs_417_io_enable; // @[RegFile.scala 66:20:@40249.4]
  wire  regs_418_clock; // @[RegFile.scala 66:20:@40263.4]
  wire  regs_418_reset; // @[RegFile.scala 66:20:@40263.4]
  wire [63:0] regs_418_io_in; // @[RegFile.scala 66:20:@40263.4]
  wire  regs_418_io_reset; // @[RegFile.scala 66:20:@40263.4]
  wire [63:0] regs_418_io_out; // @[RegFile.scala 66:20:@40263.4]
  wire  regs_418_io_enable; // @[RegFile.scala 66:20:@40263.4]
  wire  regs_419_clock; // @[RegFile.scala 66:20:@40277.4]
  wire  regs_419_reset; // @[RegFile.scala 66:20:@40277.4]
  wire [63:0] regs_419_io_in; // @[RegFile.scala 66:20:@40277.4]
  wire  regs_419_io_reset; // @[RegFile.scala 66:20:@40277.4]
  wire [63:0] regs_419_io_out; // @[RegFile.scala 66:20:@40277.4]
  wire  regs_419_io_enable; // @[RegFile.scala 66:20:@40277.4]
  wire  regs_420_clock; // @[RegFile.scala 66:20:@40291.4]
  wire  regs_420_reset; // @[RegFile.scala 66:20:@40291.4]
  wire [63:0] regs_420_io_in; // @[RegFile.scala 66:20:@40291.4]
  wire  regs_420_io_reset; // @[RegFile.scala 66:20:@40291.4]
  wire [63:0] regs_420_io_out; // @[RegFile.scala 66:20:@40291.4]
  wire  regs_420_io_enable; // @[RegFile.scala 66:20:@40291.4]
  wire  regs_421_clock; // @[RegFile.scala 66:20:@40305.4]
  wire  regs_421_reset; // @[RegFile.scala 66:20:@40305.4]
  wire [63:0] regs_421_io_in; // @[RegFile.scala 66:20:@40305.4]
  wire  regs_421_io_reset; // @[RegFile.scala 66:20:@40305.4]
  wire [63:0] regs_421_io_out; // @[RegFile.scala 66:20:@40305.4]
  wire  regs_421_io_enable; // @[RegFile.scala 66:20:@40305.4]
  wire  regs_422_clock; // @[RegFile.scala 66:20:@40319.4]
  wire  regs_422_reset; // @[RegFile.scala 66:20:@40319.4]
  wire [63:0] regs_422_io_in; // @[RegFile.scala 66:20:@40319.4]
  wire  regs_422_io_reset; // @[RegFile.scala 66:20:@40319.4]
  wire [63:0] regs_422_io_out; // @[RegFile.scala 66:20:@40319.4]
  wire  regs_422_io_enable; // @[RegFile.scala 66:20:@40319.4]
  wire  regs_423_clock; // @[RegFile.scala 66:20:@40333.4]
  wire  regs_423_reset; // @[RegFile.scala 66:20:@40333.4]
  wire [63:0] regs_423_io_in; // @[RegFile.scala 66:20:@40333.4]
  wire  regs_423_io_reset; // @[RegFile.scala 66:20:@40333.4]
  wire [63:0] regs_423_io_out; // @[RegFile.scala 66:20:@40333.4]
  wire  regs_423_io_enable; // @[RegFile.scala 66:20:@40333.4]
  wire  regs_424_clock; // @[RegFile.scala 66:20:@40347.4]
  wire  regs_424_reset; // @[RegFile.scala 66:20:@40347.4]
  wire [63:0] regs_424_io_in; // @[RegFile.scala 66:20:@40347.4]
  wire  regs_424_io_reset; // @[RegFile.scala 66:20:@40347.4]
  wire [63:0] regs_424_io_out; // @[RegFile.scala 66:20:@40347.4]
  wire  regs_424_io_enable; // @[RegFile.scala 66:20:@40347.4]
  wire  regs_425_clock; // @[RegFile.scala 66:20:@40361.4]
  wire  regs_425_reset; // @[RegFile.scala 66:20:@40361.4]
  wire [63:0] regs_425_io_in; // @[RegFile.scala 66:20:@40361.4]
  wire  regs_425_io_reset; // @[RegFile.scala 66:20:@40361.4]
  wire [63:0] regs_425_io_out; // @[RegFile.scala 66:20:@40361.4]
  wire  regs_425_io_enable; // @[RegFile.scala 66:20:@40361.4]
  wire  regs_426_clock; // @[RegFile.scala 66:20:@40375.4]
  wire  regs_426_reset; // @[RegFile.scala 66:20:@40375.4]
  wire [63:0] regs_426_io_in; // @[RegFile.scala 66:20:@40375.4]
  wire  regs_426_io_reset; // @[RegFile.scala 66:20:@40375.4]
  wire [63:0] regs_426_io_out; // @[RegFile.scala 66:20:@40375.4]
  wire  regs_426_io_enable; // @[RegFile.scala 66:20:@40375.4]
  wire  regs_427_clock; // @[RegFile.scala 66:20:@40389.4]
  wire  regs_427_reset; // @[RegFile.scala 66:20:@40389.4]
  wire [63:0] regs_427_io_in; // @[RegFile.scala 66:20:@40389.4]
  wire  regs_427_io_reset; // @[RegFile.scala 66:20:@40389.4]
  wire [63:0] regs_427_io_out; // @[RegFile.scala 66:20:@40389.4]
  wire  regs_427_io_enable; // @[RegFile.scala 66:20:@40389.4]
  wire  regs_428_clock; // @[RegFile.scala 66:20:@40403.4]
  wire  regs_428_reset; // @[RegFile.scala 66:20:@40403.4]
  wire [63:0] regs_428_io_in; // @[RegFile.scala 66:20:@40403.4]
  wire  regs_428_io_reset; // @[RegFile.scala 66:20:@40403.4]
  wire [63:0] regs_428_io_out; // @[RegFile.scala 66:20:@40403.4]
  wire  regs_428_io_enable; // @[RegFile.scala 66:20:@40403.4]
  wire  regs_429_clock; // @[RegFile.scala 66:20:@40417.4]
  wire  regs_429_reset; // @[RegFile.scala 66:20:@40417.4]
  wire [63:0] regs_429_io_in; // @[RegFile.scala 66:20:@40417.4]
  wire  regs_429_io_reset; // @[RegFile.scala 66:20:@40417.4]
  wire [63:0] regs_429_io_out; // @[RegFile.scala 66:20:@40417.4]
  wire  regs_429_io_enable; // @[RegFile.scala 66:20:@40417.4]
  wire  regs_430_clock; // @[RegFile.scala 66:20:@40431.4]
  wire  regs_430_reset; // @[RegFile.scala 66:20:@40431.4]
  wire [63:0] regs_430_io_in; // @[RegFile.scala 66:20:@40431.4]
  wire  regs_430_io_reset; // @[RegFile.scala 66:20:@40431.4]
  wire [63:0] regs_430_io_out; // @[RegFile.scala 66:20:@40431.4]
  wire  regs_430_io_enable; // @[RegFile.scala 66:20:@40431.4]
  wire  regs_431_clock; // @[RegFile.scala 66:20:@40445.4]
  wire  regs_431_reset; // @[RegFile.scala 66:20:@40445.4]
  wire [63:0] regs_431_io_in; // @[RegFile.scala 66:20:@40445.4]
  wire  regs_431_io_reset; // @[RegFile.scala 66:20:@40445.4]
  wire [63:0] regs_431_io_out; // @[RegFile.scala 66:20:@40445.4]
  wire  regs_431_io_enable; // @[RegFile.scala 66:20:@40445.4]
  wire  regs_432_clock; // @[RegFile.scala 66:20:@40459.4]
  wire  regs_432_reset; // @[RegFile.scala 66:20:@40459.4]
  wire [63:0] regs_432_io_in; // @[RegFile.scala 66:20:@40459.4]
  wire  regs_432_io_reset; // @[RegFile.scala 66:20:@40459.4]
  wire [63:0] regs_432_io_out; // @[RegFile.scala 66:20:@40459.4]
  wire  regs_432_io_enable; // @[RegFile.scala 66:20:@40459.4]
  wire  regs_433_clock; // @[RegFile.scala 66:20:@40473.4]
  wire  regs_433_reset; // @[RegFile.scala 66:20:@40473.4]
  wire [63:0] regs_433_io_in; // @[RegFile.scala 66:20:@40473.4]
  wire  regs_433_io_reset; // @[RegFile.scala 66:20:@40473.4]
  wire [63:0] regs_433_io_out; // @[RegFile.scala 66:20:@40473.4]
  wire  regs_433_io_enable; // @[RegFile.scala 66:20:@40473.4]
  wire  regs_434_clock; // @[RegFile.scala 66:20:@40487.4]
  wire  regs_434_reset; // @[RegFile.scala 66:20:@40487.4]
  wire [63:0] regs_434_io_in; // @[RegFile.scala 66:20:@40487.4]
  wire  regs_434_io_reset; // @[RegFile.scala 66:20:@40487.4]
  wire [63:0] regs_434_io_out; // @[RegFile.scala 66:20:@40487.4]
  wire  regs_434_io_enable; // @[RegFile.scala 66:20:@40487.4]
  wire  regs_435_clock; // @[RegFile.scala 66:20:@40501.4]
  wire  regs_435_reset; // @[RegFile.scala 66:20:@40501.4]
  wire [63:0] regs_435_io_in; // @[RegFile.scala 66:20:@40501.4]
  wire  regs_435_io_reset; // @[RegFile.scala 66:20:@40501.4]
  wire [63:0] regs_435_io_out; // @[RegFile.scala 66:20:@40501.4]
  wire  regs_435_io_enable; // @[RegFile.scala 66:20:@40501.4]
  wire  regs_436_clock; // @[RegFile.scala 66:20:@40515.4]
  wire  regs_436_reset; // @[RegFile.scala 66:20:@40515.4]
  wire [63:0] regs_436_io_in; // @[RegFile.scala 66:20:@40515.4]
  wire  regs_436_io_reset; // @[RegFile.scala 66:20:@40515.4]
  wire [63:0] regs_436_io_out; // @[RegFile.scala 66:20:@40515.4]
  wire  regs_436_io_enable; // @[RegFile.scala 66:20:@40515.4]
  wire  regs_437_clock; // @[RegFile.scala 66:20:@40529.4]
  wire  regs_437_reset; // @[RegFile.scala 66:20:@40529.4]
  wire [63:0] regs_437_io_in; // @[RegFile.scala 66:20:@40529.4]
  wire  regs_437_io_reset; // @[RegFile.scala 66:20:@40529.4]
  wire [63:0] regs_437_io_out; // @[RegFile.scala 66:20:@40529.4]
  wire  regs_437_io_enable; // @[RegFile.scala 66:20:@40529.4]
  wire  regs_438_clock; // @[RegFile.scala 66:20:@40543.4]
  wire  regs_438_reset; // @[RegFile.scala 66:20:@40543.4]
  wire [63:0] regs_438_io_in; // @[RegFile.scala 66:20:@40543.4]
  wire  regs_438_io_reset; // @[RegFile.scala 66:20:@40543.4]
  wire [63:0] regs_438_io_out; // @[RegFile.scala 66:20:@40543.4]
  wire  regs_438_io_enable; // @[RegFile.scala 66:20:@40543.4]
  wire  regs_439_clock; // @[RegFile.scala 66:20:@40557.4]
  wire  regs_439_reset; // @[RegFile.scala 66:20:@40557.4]
  wire [63:0] regs_439_io_in; // @[RegFile.scala 66:20:@40557.4]
  wire  regs_439_io_reset; // @[RegFile.scala 66:20:@40557.4]
  wire [63:0] regs_439_io_out; // @[RegFile.scala 66:20:@40557.4]
  wire  regs_439_io_enable; // @[RegFile.scala 66:20:@40557.4]
  wire  regs_440_clock; // @[RegFile.scala 66:20:@40571.4]
  wire  regs_440_reset; // @[RegFile.scala 66:20:@40571.4]
  wire [63:0] regs_440_io_in; // @[RegFile.scala 66:20:@40571.4]
  wire  regs_440_io_reset; // @[RegFile.scala 66:20:@40571.4]
  wire [63:0] regs_440_io_out; // @[RegFile.scala 66:20:@40571.4]
  wire  regs_440_io_enable; // @[RegFile.scala 66:20:@40571.4]
  wire  regs_441_clock; // @[RegFile.scala 66:20:@40585.4]
  wire  regs_441_reset; // @[RegFile.scala 66:20:@40585.4]
  wire [63:0] regs_441_io_in; // @[RegFile.scala 66:20:@40585.4]
  wire  regs_441_io_reset; // @[RegFile.scala 66:20:@40585.4]
  wire [63:0] regs_441_io_out; // @[RegFile.scala 66:20:@40585.4]
  wire  regs_441_io_enable; // @[RegFile.scala 66:20:@40585.4]
  wire  regs_442_clock; // @[RegFile.scala 66:20:@40599.4]
  wire  regs_442_reset; // @[RegFile.scala 66:20:@40599.4]
  wire [63:0] regs_442_io_in; // @[RegFile.scala 66:20:@40599.4]
  wire  regs_442_io_reset; // @[RegFile.scala 66:20:@40599.4]
  wire [63:0] regs_442_io_out; // @[RegFile.scala 66:20:@40599.4]
  wire  regs_442_io_enable; // @[RegFile.scala 66:20:@40599.4]
  wire  regs_443_clock; // @[RegFile.scala 66:20:@40613.4]
  wire  regs_443_reset; // @[RegFile.scala 66:20:@40613.4]
  wire [63:0] regs_443_io_in; // @[RegFile.scala 66:20:@40613.4]
  wire  regs_443_io_reset; // @[RegFile.scala 66:20:@40613.4]
  wire [63:0] regs_443_io_out; // @[RegFile.scala 66:20:@40613.4]
  wire  regs_443_io_enable; // @[RegFile.scala 66:20:@40613.4]
  wire  regs_444_clock; // @[RegFile.scala 66:20:@40627.4]
  wire  regs_444_reset; // @[RegFile.scala 66:20:@40627.4]
  wire [63:0] regs_444_io_in; // @[RegFile.scala 66:20:@40627.4]
  wire  regs_444_io_reset; // @[RegFile.scala 66:20:@40627.4]
  wire [63:0] regs_444_io_out; // @[RegFile.scala 66:20:@40627.4]
  wire  regs_444_io_enable; // @[RegFile.scala 66:20:@40627.4]
  wire  regs_445_clock; // @[RegFile.scala 66:20:@40641.4]
  wire  regs_445_reset; // @[RegFile.scala 66:20:@40641.4]
  wire [63:0] regs_445_io_in; // @[RegFile.scala 66:20:@40641.4]
  wire  regs_445_io_reset; // @[RegFile.scala 66:20:@40641.4]
  wire [63:0] regs_445_io_out; // @[RegFile.scala 66:20:@40641.4]
  wire  regs_445_io_enable; // @[RegFile.scala 66:20:@40641.4]
  wire  regs_446_clock; // @[RegFile.scala 66:20:@40655.4]
  wire  regs_446_reset; // @[RegFile.scala 66:20:@40655.4]
  wire [63:0] regs_446_io_in; // @[RegFile.scala 66:20:@40655.4]
  wire  regs_446_io_reset; // @[RegFile.scala 66:20:@40655.4]
  wire [63:0] regs_446_io_out; // @[RegFile.scala 66:20:@40655.4]
  wire  regs_446_io_enable; // @[RegFile.scala 66:20:@40655.4]
  wire  regs_447_clock; // @[RegFile.scala 66:20:@40669.4]
  wire  regs_447_reset; // @[RegFile.scala 66:20:@40669.4]
  wire [63:0] regs_447_io_in; // @[RegFile.scala 66:20:@40669.4]
  wire  regs_447_io_reset; // @[RegFile.scala 66:20:@40669.4]
  wire [63:0] regs_447_io_out; // @[RegFile.scala 66:20:@40669.4]
  wire  regs_447_io_enable; // @[RegFile.scala 66:20:@40669.4]
  wire  regs_448_clock; // @[RegFile.scala 66:20:@40683.4]
  wire  regs_448_reset; // @[RegFile.scala 66:20:@40683.4]
  wire [63:0] regs_448_io_in; // @[RegFile.scala 66:20:@40683.4]
  wire  regs_448_io_reset; // @[RegFile.scala 66:20:@40683.4]
  wire [63:0] regs_448_io_out; // @[RegFile.scala 66:20:@40683.4]
  wire  regs_448_io_enable; // @[RegFile.scala 66:20:@40683.4]
  wire  regs_449_clock; // @[RegFile.scala 66:20:@40697.4]
  wire  regs_449_reset; // @[RegFile.scala 66:20:@40697.4]
  wire [63:0] regs_449_io_in; // @[RegFile.scala 66:20:@40697.4]
  wire  regs_449_io_reset; // @[RegFile.scala 66:20:@40697.4]
  wire [63:0] regs_449_io_out; // @[RegFile.scala 66:20:@40697.4]
  wire  regs_449_io_enable; // @[RegFile.scala 66:20:@40697.4]
  wire  regs_450_clock; // @[RegFile.scala 66:20:@40711.4]
  wire  regs_450_reset; // @[RegFile.scala 66:20:@40711.4]
  wire [63:0] regs_450_io_in; // @[RegFile.scala 66:20:@40711.4]
  wire  regs_450_io_reset; // @[RegFile.scala 66:20:@40711.4]
  wire [63:0] regs_450_io_out; // @[RegFile.scala 66:20:@40711.4]
  wire  regs_450_io_enable; // @[RegFile.scala 66:20:@40711.4]
  wire  regs_451_clock; // @[RegFile.scala 66:20:@40725.4]
  wire  regs_451_reset; // @[RegFile.scala 66:20:@40725.4]
  wire [63:0] regs_451_io_in; // @[RegFile.scala 66:20:@40725.4]
  wire  regs_451_io_reset; // @[RegFile.scala 66:20:@40725.4]
  wire [63:0] regs_451_io_out; // @[RegFile.scala 66:20:@40725.4]
  wire  regs_451_io_enable; // @[RegFile.scala 66:20:@40725.4]
  wire  regs_452_clock; // @[RegFile.scala 66:20:@40739.4]
  wire  regs_452_reset; // @[RegFile.scala 66:20:@40739.4]
  wire [63:0] regs_452_io_in; // @[RegFile.scala 66:20:@40739.4]
  wire  regs_452_io_reset; // @[RegFile.scala 66:20:@40739.4]
  wire [63:0] regs_452_io_out; // @[RegFile.scala 66:20:@40739.4]
  wire  regs_452_io_enable; // @[RegFile.scala 66:20:@40739.4]
  wire  regs_453_clock; // @[RegFile.scala 66:20:@40753.4]
  wire  regs_453_reset; // @[RegFile.scala 66:20:@40753.4]
  wire [63:0] regs_453_io_in; // @[RegFile.scala 66:20:@40753.4]
  wire  regs_453_io_reset; // @[RegFile.scala 66:20:@40753.4]
  wire [63:0] regs_453_io_out; // @[RegFile.scala 66:20:@40753.4]
  wire  regs_453_io_enable; // @[RegFile.scala 66:20:@40753.4]
  wire  regs_454_clock; // @[RegFile.scala 66:20:@40767.4]
  wire  regs_454_reset; // @[RegFile.scala 66:20:@40767.4]
  wire [63:0] regs_454_io_in; // @[RegFile.scala 66:20:@40767.4]
  wire  regs_454_io_reset; // @[RegFile.scala 66:20:@40767.4]
  wire [63:0] regs_454_io_out; // @[RegFile.scala 66:20:@40767.4]
  wire  regs_454_io_enable; // @[RegFile.scala 66:20:@40767.4]
  wire  regs_455_clock; // @[RegFile.scala 66:20:@40781.4]
  wire  regs_455_reset; // @[RegFile.scala 66:20:@40781.4]
  wire [63:0] regs_455_io_in; // @[RegFile.scala 66:20:@40781.4]
  wire  regs_455_io_reset; // @[RegFile.scala 66:20:@40781.4]
  wire [63:0] regs_455_io_out; // @[RegFile.scala 66:20:@40781.4]
  wire  regs_455_io_enable; // @[RegFile.scala 66:20:@40781.4]
  wire  regs_456_clock; // @[RegFile.scala 66:20:@40795.4]
  wire  regs_456_reset; // @[RegFile.scala 66:20:@40795.4]
  wire [63:0] regs_456_io_in; // @[RegFile.scala 66:20:@40795.4]
  wire  regs_456_io_reset; // @[RegFile.scala 66:20:@40795.4]
  wire [63:0] regs_456_io_out; // @[RegFile.scala 66:20:@40795.4]
  wire  regs_456_io_enable; // @[RegFile.scala 66:20:@40795.4]
  wire  regs_457_clock; // @[RegFile.scala 66:20:@40809.4]
  wire  regs_457_reset; // @[RegFile.scala 66:20:@40809.4]
  wire [63:0] regs_457_io_in; // @[RegFile.scala 66:20:@40809.4]
  wire  regs_457_io_reset; // @[RegFile.scala 66:20:@40809.4]
  wire [63:0] regs_457_io_out; // @[RegFile.scala 66:20:@40809.4]
  wire  regs_457_io_enable; // @[RegFile.scala 66:20:@40809.4]
  wire  regs_458_clock; // @[RegFile.scala 66:20:@40823.4]
  wire  regs_458_reset; // @[RegFile.scala 66:20:@40823.4]
  wire [63:0] regs_458_io_in; // @[RegFile.scala 66:20:@40823.4]
  wire  regs_458_io_reset; // @[RegFile.scala 66:20:@40823.4]
  wire [63:0] regs_458_io_out; // @[RegFile.scala 66:20:@40823.4]
  wire  regs_458_io_enable; // @[RegFile.scala 66:20:@40823.4]
  wire  regs_459_clock; // @[RegFile.scala 66:20:@40837.4]
  wire  regs_459_reset; // @[RegFile.scala 66:20:@40837.4]
  wire [63:0] regs_459_io_in; // @[RegFile.scala 66:20:@40837.4]
  wire  regs_459_io_reset; // @[RegFile.scala 66:20:@40837.4]
  wire [63:0] regs_459_io_out; // @[RegFile.scala 66:20:@40837.4]
  wire  regs_459_io_enable; // @[RegFile.scala 66:20:@40837.4]
  wire  regs_460_clock; // @[RegFile.scala 66:20:@40851.4]
  wire  regs_460_reset; // @[RegFile.scala 66:20:@40851.4]
  wire [63:0] regs_460_io_in; // @[RegFile.scala 66:20:@40851.4]
  wire  regs_460_io_reset; // @[RegFile.scala 66:20:@40851.4]
  wire [63:0] regs_460_io_out; // @[RegFile.scala 66:20:@40851.4]
  wire  regs_460_io_enable; // @[RegFile.scala 66:20:@40851.4]
  wire  regs_461_clock; // @[RegFile.scala 66:20:@40865.4]
  wire  regs_461_reset; // @[RegFile.scala 66:20:@40865.4]
  wire [63:0] regs_461_io_in; // @[RegFile.scala 66:20:@40865.4]
  wire  regs_461_io_reset; // @[RegFile.scala 66:20:@40865.4]
  wire [63:0] regs_461_io_out; // @[RegFile.scala 66:20:@40865.4]
  wire  regs_461_io_enable; // @[RegFile.scala 66:20:@40865.4]
  wire  regs_462_clock; // @[RegFile.scala 66:20:@40879.4]
  wire  regs_462_reset; // @[RegFile.scala 66:20:@40879.4]
  wire [63:0] regs_462_io_in; // @[RegFile.scala 66:20:@40879.4]
  wire  regs_462_io_reset; // @[RegFile.scala 66:20:@40879.4]
  wire [63:0] regs_462_io_out; // @[RegFile.scala 66:20:@40879.4]
  wire  regs_462_io_enable; // @[RegFile.scala 66:20:@40879.4]
  wire  regs_463_clock; // @[RegFile.scala 66:20:@40893.4]
  wire  regs_463_reset; // @[RegFile.scala 66:20:@40893.4]
  wire [63:0] regs_463_io_in; // @[RegFile.scala 66:20:@40893.4]
  wire  regs_463_io_reset; // @[RegFile.scala 66:20:@40893.4]
  wire [63:0] regs_463_io_out; // @[RegFile.scala 66:20:@40893.4]
  wire  regs_463_io_enable; // @[RegFile.scala 66:20:@40893.4]
  wire  regs_464_clock; // @[RegFile.scala 66:20:@40907.4]
  wire  regs_464_reset; // @[RegFile.scala 66:20:@40907.4]
  wire [63:0] regs_464_io_in; // @[RegFile.scala 66:20:@40907.4]
  wire  regs_464_io_reset; // @[RegFile.scala 66:20:@40907.4]
  wire [63:0] regs_464_io_out; // @[RegFile.scala 66:20:@40907.4]
  wire  regs_464_io_enable; // @[RegFile.scala 66:20:@40907.4]
  wire  regs_465_clock; // @[RegFile.scala 66:20:@40921.4]
  wire  regs_465_reset; // @[RegFile.scala 66:20:@40921.4]
  wire [63:0] regs_465_io_in; // @[RegFile.scala 66:20:@40921.4]
  wire  regs_465_io_reset; // @[RegFile.scala 66:20:@40921.4]
  wire [63:0] regs_465_io_out; // @[RegFile.scala 66:20:@40921.4]
  wire  regs_465_io_enable; // @[RegFile.scala 66:20:@40921.4]
  wire  regs_466_clock; // @[RegFile.scala 66:20:@40935.4]
  wire  regs_466_reset; // @[RegFile.scala 66:20:@40935.4]
  wire [63:0] regs_466_io_in; // @[RegFile.scala 66:20:@40935.4]
  wire  regs_466_io_reset; // @[RegFile.scala 66:20:@40935.4]
  wire [63:0] regs_466_io_out; // @[RegFile.scala 66:20:@40935.4]
  wire  regs_466_io_enable; // @[RegFile.scala 66:20:@40935.4]
  wire  regs_467_clock; // @[RegFile.scala 66:20:@40949.4]
  wire  regs_467_reset; // @[RegFile.scala 66:20:@40949.4]
  wire [63:0] regs_467_io_in; // @[RegFile.scala 66:20:@40949.4]
  wire  regs_467_io_reset; // @[RegFile.scala 66:20:@40949.4]
  wire [63:0] regs_467_io_out; // @[RegFile.scala 66:20:@40949.4]
  wire  regs_467_io_enable; // @[RegFile.scala 66:20:@40949.4]
  wire  regs_468_clock; // @[RegFile.scala 66:20:@40963.4]
  wire  regs_468_reset; // @[RegFile.scala 66:20:@40963.4]
  wire [63:0] regs_468_io_in; // @[RegFile.scala 66:20:@40963.4]
  wire  regs_468_io_reset; // @[RegFile.scala 66:20:@40963.4]
  wire [63:0] regs_468_io_out; // @[RegFile.scala 66:20:@40963.4]
  wire  regs_468_io_enable; // @[RegFile.scala 66:20:@40963.4]
  wire  regs_469_clock; // @[RegFile.scala 66:20:@40977.4]
  wire  regs_469_reset; // @[RegFile.scala 66:20:@40977.4]
  wire [63:0] regs_469_io_in; // @[RegFile.scala 66:20:@40977.4]
  wire  regs_469_io_reset; // @[RegFile.scala 66:20:@40977.4]
  wire [63:0] regs_469_io_out; // @[RegFile.scala 66:20:@40977.4]
  wire  regs_469_io_enable; // @[RegFile.scala 66:20:@40977.4]
  wire  regs_470_clock; // @[RegFile.scala 66:20:@40991.4]
  wire  regs_470_reset; // @[RegFile.scala 66:20:@40991.4]
  wire [63:0] regs_470_io_in; // @[RegFile.scala 66:20:@40991.4]
  wire  regs_470_io_reset; // @[RegFile.scala 66:20:@40991.4]
  wire [63:0] regs_470_io_out; // @[RegFile.scala 66:20:@40991.4]
  wire  regs_470_io_enable; // @[RegFile.scala 66:20:@40991.4]
  wire  regs_471_clock; // @[RegFile.scala 66:20:@41005.4]
  wire  regs_471_reset; // @[RegFile.scala 66:20:@41005.4]
  wire [63:0] regs_471_io_in; // @[RegFile.scala 66:20:@41005.4]
  wire  regs_471_io_reset; // @[RegFile.scala 66:20:@41005.4]
  wire [63:0] regs_471_io_out; // @[RegFile.scala 66:20:@41005.4]
  wire  regs_471_io_enable; // @[RegFile.scala 66:20:@41005.4]
  wire  regs_472_clock; // @[RegFile.scala 66:20:@41019.4]
  wire  regs_472_reset; // @[RegFile.scala 66:20:@41019.4]
  wire [63:0] regs_472_io_in; // @[RegFile.scala 66:20:@41019.4]
  wire  regs_472_io_reset; // @[RegFile.scala 66:20:@41019.4]
  wire [63:0] regs_472_io_out; // @[RegFile.scala 66:20:@41019.4]
  wire  regs_472_io_enable; // @[RegFile.scala 66:20:@41019.4]
  wire  regs_473_clock; // @[RegFile.scala 66:20:@41033.4]
  wire  regs_473_reset; // @[RegFile.scala 66:20:@41033.4]
  wire [63:0] regs_473_io_in; // @[RegFile.scala 66:20:@41033.4]
  wire  regs_473_io_reset; // @[RegFile.scala 66:20:@41033.4]
  wire [63:0] regs_473_io_out; // @[RegFile.scala 66:20:@41033.4]
  wire  regs_473_io_enable; // @[RegFile.scala 66:20:@41033.4]
  wire  regs_474_clock; // @[RegFile.scala 66:20:@41047.4]
  wire  regs_474_reset; // @[RegFile.scala 66:20:@41047.4]
  wire [63:0] regs_474_io_in; // @[RegFile.scala 66:20:@41047.4]
  wire  regs_474_io_reset; // @[RegFile.scala 66:20:@41047.4]
  wire [63:0] regs_474_io_out; // @[RegFile.scala 66:20:@41047.4]
  wire  regs_474_io_enable; // @[RegFile.scala 66:20:@41047.4]
  wire  regs_475_clock; // @[RegFile.scala 66:20:@41061.4]
  wire  regs_475_reset; // @[RegFile.scala 66:20:@41061.4]
  wire [63:0] regs_475_io_in; // @[RegFile.scala 66:20:@41061.4]
  wire  regs_475_io_reset; // @[RegFile.scala 66:20:@41061.4]
  wire [63:0] regs_475_io_out; // @[RegFile.scala 66:20:@41061.4]
  wire  regs_475_io_enable; // @[RegFile.scala 66:20:@41061.4]
  wire  regs_476_clock; // @[RegFile.scala 66:20:@41075.4]
  wire  regs_476_reset; // @[RegFile.scala 66:20:@41075.4]
  wire [63:0] regs_476_io_in; // @[RegFile.scala 66:20:@41075.4]
  wire  regs_476_io_reset; // @[RegFile.scala 66:20:@41075.4]
  wire [63:0] regs_476_io_out; // @[RegFile.scala 66:20:@41075.4]
  wire  regs_476_io_enable; // @[RegFile.scala 66:20:@41075.4]
  wire  regs_477_clock; // @[RegFile.scala 66:20:@41089.4]
  wire  regs_477_reset; // @[RegFile.scala 66:20:@41089.4]
  wire [63:0] regs_477_io_in; // @[RegFile.scala 66:20:@41089.4]
  wire  regs_477_io_reset; // @[RegFile.scala 66:20:@41089.4]
  wire [63:0] regs_477_io_out; // @[RegFile.scala 66:20:@41089.4]
  wire  regs_477_io_enable; // @[RegFile.scala 66:20:@41089.4]
  wire  regs_478_clock; // @[RegFile.scala 66:20:@41103.4]
  wire  regs_478_reset; // @[RegFile.scala 66:20:@41103.4]
  wire [63:0] regs_478_io_in; // @[RegFile.scala 66:20:@41103.4]
  wire  regs_478_io_reset; // @[RegFile.scala 66:20:@41103.4]
  wire [63:0] regs_478_io_out; // @[RegFile.scala 66:20:@41103.4]
  wire  regs_478_io_enable; // @[RegFile.scala 66:20:@41103.4]
  wire  regs_479_clock; // @[RegFile.scala 66:20:@41117.4]
  wire  regs_479_reset; // @[RegFile.scala 66:20:@41117.4]
  wire [63:0] regs_479_io_in; // @[RegFile.scala 66:20:@41117.4]
  wire  regs_479_io_reset; // @[RegFile.scala 66:20:@41117.4]
  wire [63:0] regs_479_io_out; // @[RegFile.scala 66:20:@41117.4]
  wire  regs_479_io_enable; // @[RegFile.scala 66:20:@41117.4]
  wire  regs_480_clock; // @[RegFile.scala 66:20:@41131.4]
  wire  regs_480_reset; // @[RegFile.scala 66:20:@41131.4]
  wire [63:0] regs_480_io_in; // @[RegFile.scala 66:20:@41131.4]
  wire  regs_480_io_reset; // @[RegFile.scala 66:20:@41131.4]
  wire [63:0] regs_480_io_out; // @[RegFile.scala 66:20:@41131.4]
  wire  regs_480_io_enable; // @[RegFile.scala 66:20:@41131.4]
  wire  regs_481_clock; // @[RegFile.scala 66:20:@41145.4]
  wire  regs_481_reset; // @[RegFile.scala 66:20:@41145.4]
  wire [63:0] regs_481_io_in; // @[RegFile.scala 66:20:@41145.4]
  wire  regs_481_io_reset; // @[RegFile.scala 66:20:@41145.4]
  wire [63:0] regs_481_io_out; // @[RegFile.scala 66:20:@41145.4]
  wire  regs_481_io_enable; // @[RegFile.scala 66:20:@41145.4]
  wire  regs_482_clock; // @[RegFile.scala 66:20:@41159.4]
  wire  regs_482_reset; // @[RegFile.scala 66:20:@41159.4]
  wire [63:0] regs_482_io_in; // @[RegFile.scala 66:20:@41159.4]
  wire  regs_482_io_reset; // @[RegFile.scala 66:20:@41159.4]
  wire [63:0] regs_482_io_out; // @[RegFile.scala 66:20:@41159.4]
  wire  regs_482_io_enable; // @[RegFile.scala 66:20:@41159.4]
  wire  regs_483_clock; // @[RegFile.scala 66:20:@41173.4]
  wire  regs_483_reset; // @[RegFile.scala 66:20:@41173.4]
  wire [63:0] regs_483_io_in; // @[RegFile.scala 66:20:@41173.4]
  wire  regs_483_io_reset; // @[RegFile.scala 66:20:@41173.4]
  wire [63:0] regs_483_io_out; // @[RegFile.scala 66:20:@41173.4]
  wire  regs_483_io_enable; // @[RegFile.scala 66:20:@41173.4]
  wire  regs_484_clock; // @[RegFile.scala 66:20:@41187.4]
  wire  regs_484_reset; // @[RegFile.scala 66:20:@41187.4]
  wire [63:0] regs_484_io_in; // @[RegFile.scala 66:20:@41187.4]
  wire  regs_484_io_reset; // @[RegFile.scala 66:20:@41187.4]
  wire [63:0] regs_484_io_out; // @[RegFile.scala 66:20:@41187.4]
  wire  regs_484_io_enable; // @[RegFile.scala 66:20:@41187.4]
  wire  regs_485_clock; // @[RegFile.scala 66:20:@41201.4]
  wire  regs_485_reset; // @[RegFile.scala 66:20:@41201.4]
  wire [63:0] regs_485_io_in; // @[RegFile.scala 66:20:@41201.4]
  wire  regs_485_io_reset; // @[RegFile.scala 66:20:@41201.4]
  wire [63:0] regs_485_io_out; // @[RegFile.scala 66:20:@41201.4]
  wire  regs_485_io_enable; // @[RegFile.scala 66:20:@41201.4]
  wire  regs_486_clock; // @[RegFile.scala 66:20:@41215.4]
  wire  regs_486_reset; // @[RegFile.scala 66:20:@41215.4]
  wire [63:0] regs_486_io_in; // @[RegFile.scala 66:20:@41215.4]
  wire  regs_486_io_reset; // @[RegFile.scala 66:20:@41215.4]
  wire [63:0] regs_486_io_out; // @[RegFile.scala 66:20:@41215.4]
  wire  regs_486_io_enable; // @[RegFile.scala 66:20:@41215.4]
  wire  regs_487_clock; // @[RegFile.scala 66:20:@41229.4]
  wire  regs_487_reset; // @[RegFile.scala 66:20:@41229.4]
  wire [63:0] regs_487_io_in; // @[RegFile.scala 66:20:@41229.4]
  wire  regs_487_io_reset; // @[RegFile.scala 66:20:@41229.4]
  wire [63:0] regs_487_io_out; // @[RegFile.scala 66:20:@41229.4]
  wire  regs_487_io_enable; // @[RegFile.scala 66:20:@41229.4]
  wire  regs_488_clock; // @[RegFile.scala 66:20:@41243.4]
  wire  regs_488_reset; // @[RegFile.scala 66:20:@41243.4]
  wire [63:0] regs_488_io_in; // @[RegFile.scala 66:20:@41243.4]
  wire  regs_488_io_reset; // @[RegFile.scala 66:20:@41243.4]
  wire [63:0] regs_488_io_out; // @[RegFile.scala 66:20:@41243.4]
  wire  regs_488_io_enable; // @[RegFile.scala 66:20:@41243.4]
  wire  regs_489_clock; // @[RegFile.scala 66:20:@41257.4]
  wire  regs_489_reset; // @[RegFile.scala 66:20:@41257.4]
  wire [63:0] regs_489_io_in; // @[RegFile.scala 66:20:@41257.4]
  wire  regs_489_io_reset; // @[RegFile.scala 66:20:@41257.4]
  wire [63:0] regs_489_io_out; // @[RegFile.scala 66:20:@41257.4]
  wire  regs_489_io_enable; // @[RegFile.scala 66:20:@41257.4]
  wire  regs_490_clock; // @[RegFile.scala 66:20:@41271.4]
  wire  regs_490_reset; // @[RegFile.scala 66:20:@41271.4]
  wire [63:0] regs_490_io_in; // @[RegFile.scala 66:20:@41271.4]
  wire  regs_490_io_reset; // @[RegFile.scala 66:20:@41271.4]
  wire [63:0] regs_490_io_out; // @[RegFile.scala 66:20:@41271.4]
  wire  regs_490_io_enable; // @[RegFile.scala 66:20:@41271.4]
  wire  regs_491_clock; // @[RegFile.scala 66:20:@41285.4]
  wire  regs_491_reset; // @[RegFile.scala 66:20:@41285.4]
  wire [63:0] regs_491_io_in; // @[RegFile.scala 66:20:@41285.4]
  wire  regs_491_io_reset; // @[RegFile.scala 66:20:@41285.4]
  wire [63:0] regs_491_io_out; // @[RegFile.scala 66:20:@41285.4]
  wire  regs_491_io_enable; // @[RegFile.scala 66:20:@41285.4]
  wire  regs_492_clock; // @[RegFile.scala 66:20:@41299.4]
  wire  regs_492_reset; // @[RegFile.scala 66:20:@41299.4]
  wire [63:0] regs_492_io_in; // @[RegFile.scala 66:20:@41299.4]
  wire  regs_492_io_reset; // @[RegFile.scala 66:20:@41299.4]
  wire [63:0] regs_492_io_out; // @[RegFile.scala 66:20:@41299.4]
  wire  regs_492_io_enable; // @[RegFile.scala 66:20:@41299.4]
  wire  regs_493_clock; // @[RegFile.scala 66:20:@41313.4]
  wire  regs_493_reset; // @[RegFile.scala 66:20:@41313.4]
  wire [63:0] regs_493_io_in; // @[RegFile.scala 66:20:@41313.4]
  wire  regs_493_io_reset; // @[RegFile.scala 66:20:@41313.4]
  wire [63:0] regs_493_io_out; // @[RegFile.scala 66:20:@41313.4]
  wire  regs_493_io_enable; // @[RegFile.scala 66:20:@41313.4]
  wire  regs_494_clock; // @[RegFile.scala 66:20:@41327.4]
  wire  regs_494_reset; // @[RegFile.scala 66:20:@41327.4]
  wire [63:0] regs_494_io_in; // @[RegFile.scala 66:20:@41327.4]
  wire  regs_494_io_reset; // @[RegFile.scala 66:20:@41327.4]
  wire [63:0] regs_494_io_out; // @[RegFile.scala 66:20:@41327.4]
  wire  regs_494_io_enable; // @[RegFile.scala 66:20:@41327.4]
  wire  regs_495_clock; // @[RegFile.scala 66:20:@41341.4]
  wire  regs_495_reset; // @[RegFile.scala 66:20:@41341.4]
  wire [63:0] regs_495_io_in; // @[RegFile.scala 66:20:@41341.4]
  wire  regs_495_io_reset; // @[RegFile.scala 66:20:@41341.4]
  wire [63:0] regs_495_io_out; // @[RegFile.scala 66:20:@41341.4]
  wire  regs_495_io_enable; // @[RegFile.scala 66:20:@41341.4]
  wire  regs_496_clock; // @[RegFile.scala 66:20:@41355.4]
  wire  regs_496_reset; // @[RegFile.scala 66:20:@41355.4]
  wire [63:0] regs_496_io_in; // @[RegFile.scala 66:20:@41355.4]
  wire  regs_496_io_reset; // @[RegFile.scala 66:20:@41355.4]
  wire [63:0] regs_496_io_out; // @[RegFile.scala 66:20:@41355.4]
  wire  regs_496_io_enable; // @[RegFile.scala 66:20:@41355.4]
  wire  regs_497_clock; // @[RegFile.scala 66:20:@41369.4]
  wire  regs_497_reset; // @[RegFile.scala 66:20:@41369.4]
  wire [63:0] regs_497_io_in; // @[RegFile.scala 66:20:@41369.4]
  wire  regs_497_io_reset; // @[RegFile.scala 66:20:@41369.4]
  wire [63:0] regs_497_io_out; // @[RegFile.scala 66:20:@41369.4]
  wire  regs_497_io_enable; // @[RegFile.scala 66:20:@41369.4]
  wire  regs_498_clock; // @[RegFile.scala 66:20:@41383.4]
  wire  regs_498_reset; // @[RegFile.scala 66:20:@41383.4]
  wire [63:0] regs_498_io_in; // @[RegFile.scala 66:20:@41383.4]
  wire  regs_498_io_reset; // @[RegFile.scala 66:20:@41383.4]
  wire [63:0] regs_498_io_out; // @[RegFile.scala 66:20:@41383.4]
  wire  regs_498_io_enable; // @[RegFile.scala 66:20:@41383.4]
  wire  regs_499_clock; // @[RegFile.scala 66:20:@41397.4]
  wire  regs_499_reset; // @[RegFile.scala 66:20:@41397.4]
  wire [63:0] regs_499_io_in; // @[RegFile.scala 66:20:@41397.4]
  wire  regs_499_io_reset; // @[RegFile.scala 66:20:@41397.4]
  wire [63:0] regs_499_io_out; // @[RegFile.scala 66:20:@41397.4]
  wire  regs_499_io_enable; // @[RegFile.scala 66:20:@41397.4]
  wire  regs_500_clock; // @[RegFile.scala 66:20:@41411.4]
  wire  regs_500_reset; // @[RegFile.scala 66:20:@41411.4]
  wire [63:0] regs_500_io_in; // @[RegFile.scala 66:20:@41411.4]
  wire  regs_500_io_reset; // @[RegFile.scala 66:20:@41411.4]
  wire [63:0] regs_500_io_out; // @[RegFile.scala 66:20:@41411.4]
  wire  regs_500_io_enable; // @[RegFile.scala 66:20:@41411.4]
  wire  regs_501_clock; // @[RegFile.scala 66:20:@41425.4]
  wire  regs_501_reset; // @[RegFile.scala 66:20:@41425.4]
  wire [63:0] regs_501_io_in; // @[RegFile.scala 66:20:@41425.4]
  wire  regs_501_io_reset; // @[RegFile.scala 66:20:@41425.4]
  wire [63:0] regs_501_io_out; // @[RegFile.scala 66:20:@41425.4]
  wire  regs_501_io_enable; // @[RegFile.scala 66:20:@41425.4]
  wire  regs_502_clock; // @[RegFile.scala 66:20:@41439.4]
  wire  regs_502_reset; // @[RegFile.scala 66:20:@41439.4]
  wire [63:0] regs_502_io_in; // @[RegFile.scala 66:20:@41439.4]
  wire  regs_502_io_reset; // @[RegFile.scala 66:20:@41439.4]
  wire [63:0] regs_502_io_out; // @[RegFile.scala 66:20:@41439.4]
  wire  regs_502_io_enable; // @[RegFile.scala 66:20:@41439.4]
  wire [63:0] rport_io_ins_0; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_1; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_2; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_3; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_4; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_5; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_6; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_7; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_8; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_9; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_10; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_11; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_12; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_13; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_14; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_15; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_16; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_17; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_18; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_19; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_20; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_21; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_22; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_23; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_24; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_25; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_26; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_27; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_28; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_29; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_30; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_31; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_32; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_33; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_34; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_35; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_36; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_37; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_38; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_39; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_40; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_41; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_42; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_43; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_44; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_45; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_46; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_47; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_48; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_49; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_50; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_51; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_52; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_53; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_54; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_55; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_56; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_57; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_58; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_59; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_60; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_61; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_62; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_63; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_64; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_65; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_66; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_67; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_68; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_69; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_70; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_71; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_72; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_73; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_74; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_75; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_76; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_77; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_78; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_79; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_80; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_81; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_82; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_83; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_84; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_85; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_86; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_87; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_88; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_89; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_90; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_91; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_92; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_93; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_94; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_95; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_96; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_97; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_98; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_99; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_100; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_101; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_102; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_103; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_104; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_105; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_106; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_107; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_108; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_109; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_110; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_111; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_112; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_113; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_114; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_115; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_116; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_117; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_118; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_119; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_120; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_121; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_122; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_123; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_124; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_125; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_126; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_127; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_128; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_129; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_130; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_131; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_132; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_133; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_134; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_135; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_136; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_137; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_138; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_139; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_140; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_141; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_142; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_143; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_144; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_145; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_146; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_147; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_148; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_149; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_150; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_151; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_152; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_153; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_154; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_155; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_156; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_157; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_158; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_159; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_160; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_161; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_162; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_163; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_164; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_165; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_166; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_167; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_168; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_169; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_170; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_171; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_172; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_173; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_174; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_175; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_176; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_177; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_178; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_179; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_180; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_181; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_182; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_183; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_184; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_185; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_186; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_187; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_188; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_189; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_190; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_191; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_192; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_193; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_194; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_195; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_196; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_197; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_198; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_199; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_200; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_201; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_202; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_203; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_204; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_205; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_206; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_207; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_208; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_209; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_210; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_211; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_212; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_213; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_214; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_215; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_216; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_217; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_218; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_219; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_220; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_221; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_222; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_223; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_224; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_225; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_226; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_227; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_228; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_229; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_230; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_231; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_232; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_233; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_234; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_235; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_236; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_237; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_238; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_239; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_240; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_241; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_242; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_243; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_244; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_245; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_246; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_247; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_248; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_249; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_250; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_251; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_252; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_253; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_254; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_255; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_256; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_257; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_258; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_259; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_260; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_261; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_262; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_263; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_264; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_265; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_266; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_267; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_268; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_269; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_270; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_271; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_272; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_273; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_274; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_275; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_276; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_277; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_278; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_279; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_280; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_281; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_282; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_283; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_284; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_285; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_286; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_287; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_288; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_289; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_290; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_291; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_292; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_293; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_294; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_295; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_296; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_297; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_298; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_299; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_300; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_301; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_302; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_303; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_304; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_305; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_306; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_307; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_308; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_309; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_310; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_311; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_312; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_313; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_314; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_315; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_316; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_317; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_318; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_319; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_320; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_321; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_322; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_323; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_324; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_325; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_326; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_327; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_328; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_329; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_330; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_331; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_332; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_333; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_334; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_335; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_336; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_337; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_338; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_339; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_340; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_341; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_342; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_343; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_344; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_345; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_346; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_347; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_348; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_349; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_350; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_351; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_352; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_353; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_354; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_355; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_356; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_357; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_358; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_359; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_360; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_361; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_362; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_363; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_364; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_365; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_366; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_367; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_368; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_369; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_370; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_371; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_372; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_373; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_374; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_375; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_376; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_377; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_378; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_379; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_380; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_381; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_382; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_383; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_384; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_385; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_386; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_387; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_388; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_389; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_390; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_391; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_392; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_393; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_394; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_395; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_396; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_397; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_398; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_399; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_400; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_401; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_402; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_403; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_404; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_405; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_406; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_407; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_408; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_409; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_410; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_411; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_412; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_413; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_414; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_415; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_416; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_417; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_418; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_419; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_420; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_421; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_422; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_423; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_424; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_425; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_426; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_427; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_428; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_429; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_430; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_431; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_432; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_433; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_434; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_435; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_436; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_437; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_438; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_439; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_440; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_441; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_442; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_443; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_444; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_445; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_446; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_447; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_448; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_449; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_450; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_451; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_452; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_453; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_454; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_455; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_456; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_457; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_458; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_459; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_460; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_461; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_462; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_463; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_464; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_465; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_466; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_467; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_468; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_469; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_470; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_471; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_472; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_473; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_474; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_475; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_476; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_477; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_478; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_479; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_480; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_481; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_482; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_483; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_484; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_485; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_486; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_487; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_488; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_489; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_490; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_491; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_492; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_493; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_494; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_495; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_496; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_497; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_498; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_499; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_500; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_501; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_ins_502; // @[RegFile.scala 95:21:@41453.4]
  wire [8:0] rport_io_sel; // @[RegFile.scala 95:21:@41453.4]
  wire [63:0] rport_io_out; // @[RegFile.scala 95:21:@41453.4]
  wire  _T_3076; // @[RegFile.scala 80:42:@34413.4]
  wire  _T_3082; // @[RegFile.scala 68:46:@34425.4]
  wire  _T_3083; // @[RegFile.scala 68:34:@34426.4]
  wire  _T_3096; // @[RegFile.scala 80:42:@34444.4]
  wire  _T_3102; // @[RegFile.scala 74:80:@34456.4]
  wire  _T_3103; // @[RegFile.scala 74:68:@34457.4]
  FringeFF regs_0 ( // @[RegFile.scala 66:20:@34410.4]
    .clock(regs_0_clock),
    .reset(regs_0_reset),
    .io_in(regs_0_io_in),
    .io_reset(regs_0_io_reset),
    .io_out(regs_0_io_out),
    .io_enable(regs_0_io_enable)
  );
  FringeFF regs_1 ( // @[RegFile.scala 66:20:@34422.4]
    .clock(regs_1_clock),
    .reset(regs_1_reset),
    .io_in(regs_1_io_in),
    .io_reset(regs_1_io_reset),
    .io_out(regs_1_io_out),
    .io_enable(regs_1_io_enable)
  );
  FringeFF regs_2 ( // @[RegFile.scala 66:20:@34441.4]
    .clock(regs_2_clock),
    .reset(regs_2_reset),
    .io_in(regs_2_io_in),
    .io_reset(regs_2_io_reset),
    .io_out(regs_2_io_out),
    .io_enable(regs_2_io_enable)
  );
  FringeFF regs_3 ( // @[RegFile.scala 66:20:@34453.4]
    .clock(regs_3_clock),
    .reset(regs_3_reset),
    .io_in(regs_3_io_in),
    .io_reset(regs_3_io_reset),
    .io_out(regs_3_io_out),
    .io_enable(regs_3_io_enable)
  );
  FringeFF regs_4 ( // @[RegFile.scala 66:20:@34467.4]
    .clock(regs_4_clock),
    .reset(regs_4_reset),
    .io_in(regs_4_io_in),
    .io_reset(regs_4_io_reset),
    .io_out(regs_4_io_out),
    .io_enable(regs_4_io_enable)
  );
  FringeFF regs_5 ( // @[RegFile.scala 66:20:@34481.4]
    .clock(regs_5_clock),
    .reset(regs_5_reset),
    .io_in(regs_5_io_in),
    .io_reset(regs_5_io_reset),
    .io_out(regs_5_io_out),
    .io_enable(regs_5_io_enable)
  );
  FringeFF regs_6 ( // @[RegFile.scala 66:20:@34495.4]
    .clock(regs_6_clock),
    .reset(regs_6_reset),
    .io_in(regs_6_io_in),
    .io_reset(regs_6_io_reset),
    .io_out(regs_6_io_out),
    .io_enable(regs_6_io_enable)
  );
  FringeFF regs_7 ( // @[RegFile.scala 66:20:@34509.4]
    .clock(regs_7_clock),
    .reset(regs_7_reset),
    .io_in(regs_7_io_in),
    .io_reset(regs_7_io_reset),
    .io_out(regs_7_io_out),
    .io_enable(regs_7_io_enable)
  );
  FringeFF regs_8 ( // @[RegFile.scala 66:20:@34523.4]
    .clock(regs_8_clock),
    .reset(regs_8_reset),
    .io_in(regs_8_io_in),
    .io_reset(regs_8_io_reset),
    .io_out(regs_8_io_out),
    .io_enable(regs_8_io_enable)
  );
  FringeFF regs_9 ( // @[RegFile.scala 66:20:@34537.4]
    .clock(regs_9_clock),
    .reset(regs_9_reset),
    .io_in(regs_9_io_in),
    .io_reset(regs_9_io_reset),
    .io_out(regs_9_io_out),
    .io_enable(regs_9_io_enable)
  );
  FringeFF regs_10 ( // @[RegFile.scala 66:20:@34551.4]
    .clock(regs_10_clock),
    .reset(regs_10_reset),
    .io_in(regs_10_io_in),
    .io_reset(regs_10_io_reset),
    .io_out(regs_10_io_out),
    .io_enable(regs_10_io_enable)
  );
  FringeFF regs_11 ( // @[RegFile.scala 66:20:@34565.4]
    .clock(regs_11_clock),
    .reset(regs_11_reset),
    .io_in(regs_11_io_in),
    .io_reset(regs_11_io_reset),
    .io_out(regs_11_io_out),
    .io_enable(regs_11_io_enable)
  );
  FringeFF regs_12 ( // @[RegFile.scala 66:20:@34579.4]
    .clock(regs_12_clock),
    .reset(regs_12_reset),
    .io_in(regs_12_io_in),
    .io_reset(regs_12_io_reset),
    .io_out(regs_12_io_out),
    .io_enable(regs_12_io_enable)
  );
  FringeFF regs_13 ( // @[RegFile.scala 66:20:@34593.4]
    .clock(regs_13_clock),
    .reset(regs_13_reset),
    .io_in(regs_13_io_in),
    .io_reset(regs_13_io_reset),
    .io_out(regs_13_io_out),
    .io_enable(regs_13_io_enable)
  );
  FringeFF regs_14 ( // @[RegFile.scala 66:20:@34607.4]
    .clock(regs_14_clock),
    .reset(regs_14_reset),
    .io_in(regs_14_io_in),
    .io_reset(regs_14_io_reset),
    .io_out(regs_14_io_out),
    .io_enable(regs_14_io_enable)
  );
  FringeFF regs_15 ( // @[RegFile.scala 66:20:@34621.4]
    .clock(regs_15_clock),
    .reset(regs_15_reset),
    .io_in(regs_15_io_in),
    .io_reset(regs_15_io_reset),
    .io_out(regs_15_io_out),
    .io_enable(regs_15_io_enable)
  );
  FringeFF regs_16 ( // @[RegFile.scala 66:20:@34635.4]
    .clock(regs_16_clock),
    .reset(regs_16_reset),
    .io_in(regs_16_io_in),
    .io_reset(regs_16_io_reset),
    .io_out(regs_16_io_out),
    .io_enable(regs_16_io_enable)
  );
  FringeFF regs_17 ( // @[RegFile.scala 66:20:@34649.4]
    .clock(regs_17_clock),
    .reset(regs_17_reset),
    .io_in(regs_17_io_in),
    .io_reset(regs_17_io_reset),
    .io_out(regs_17_io_out),
    .io_enable(regs_17_io_enable)
  );
  FringeFF regs_18 ( // @[RegFile.scala 66:20:@34663.4]
    .clock(regs_18_clock),
    .reset(regs_18_reset),
    .io_in(regs_18_io_in),
    .io_reset(regs_18_io_reset),
    .io_out(regs_18_io_out),
    .io_enable(regs_18_io_enable)
  );
  FringeFF regs_19 ( // @[RegFile.scala 66:20:@34677.4]
    .clock(regs_19_clock),
    .reset(regs_19_reset),
    .io_in(regs_19_io_in),
    .io_reset(regs_19_io_reset),
    .io_out(regs_19_io_out),
    .io_enable(regs_19_io_enable)
  );
  FringeFF regs_20 ( // @[RegFile.scala 66:20:@34691.4]
    .clock(regs_20_clock),
    .reset(regs_20_reset),
    .io_in(regs_20_io_in),
    .io_reset(regs_20_io_reset),
    .io_out(regs_20_io_out),
    .io_enable(regs_20_io_enable)
  );
  FringeFF regs_21 ( // @[RegFile.scala 66:20:@34705.4]
    .clock(regs_21_clock),
    .reset(regs_21_reset),
    .io_in(regs_21_io_in),
    .io_reset(regs_21_io_reset),
    .io_out(regs_21_io_out),
    .io_enable(regs_21_io_enable)
  );
  FringeFF regs_22 ( // @[RegFile.scala 66:20:@34719.4]
    .clock(regs_22_clock),
    .reset(regs_22_reset),
    .io_in(regs_22_io_in),
    .io_reset(regs_22_io_reset),
    .io_out(regs_22_io_out),
    .io_enable(regs_22_io_enable)
  );
  FringeFF regs_23 ( // @[RegFile.scala 66:20:@34733.4]
    .clock(regs_23_clock),
    .reset(regs_23_reset),
    .io_in(regs_23_io_in),
    .io_reset(regs_23_io_reset),
    .io_out(regs_23_io_out),
    .io_enable(regs_23_io_enable)
  );
  FringeFF regs_24 ( // @[RegFile.scala 66:20:@34747.4]
    .clock(regs_24_clock),
    .reset(regs_24_reset),
    .io_in(regs_24_io_in),
    .io_reset(regs_24_io_reset),
    .io_out(regs_24_io_out),
    .io_enable(regs_24_io_enable)
  );
  FringeFF regs_25 ( // @[RegFile.scala 66:20:@34761.4]
    .clock(regs_25_clock),
    .reset(regs_25_reset),
    .io_in(regs_25_io_in),
    .io_reset(regs_25_io_reset),
    .io_out(regs_25_io_out),
    .io_enable(regs_25_io_enable)
  );
  FringeFF regs_26 ( // @[RegFile.scala 66:20:@34775.4]
    .clock(regs_26_clock),
    .reset(regs_26_reset),
    .io_in(regs_26_io_in),
    .io_reset(regs_26_io_reset),
    .io_out(regs_26_io_out),
    .io_enable(regs_26_io_enable)
  );
  FringeFF regs_27 ( // @[RegFile.scala 66:20:@34789.4]
    .clock(regs_27_clock),
    .reset(regs_27_reset),
    .io_in(regs_27_io_in),
    .io_reset(regs_27_io_reset),
    .io_out(regs_27_io_out),
    .io_enable(regs_27_io_enable)
  );
  FringeFF regs_28 ( // @[RegFile.scala 66:20:@34803.4]
    .clock(regs_28_clock),
    .reset(regs_28_reset),
    .io_in(regs_28_io_in),
    .io_reset(regs_28_io_reset),
    .io_out(regs_28_io_out),
    .io_enable(regs_28_io_enable)
  );
  FringeFF regs_29 ( // @[RegFile.scala 66:20:@34817.4]
    .clock(regs_29_clock),
    .reset(regs_29_reset),
    .io_in(regs_29_io_in),
    .io_reset(regs_29_io_reset),
    .io_out(regs_29_io_out),
    .io_enable(regs_29_io_enable)
  );
  FringeFF regs_30 ( // @[RegFile.scala 66:20:@34831.4]
    .clock(regs_30_clock),
    .reset(regs_30_reset),
    .io_in(regs_30_io_in),
    .io_reset(regs_30_io_reset),
    .io_out(regs_30_io_out),
    .io_enable(regs_30_io_enable)
  );
  FringeFF regs_31 ( // @[RegFile.scala 66:20:@34845.4]
    .clock(regs_31_clock),
    .reset(regs_31_reset),
    .io_in(regs_31_io_in),
    .io_reset(regs_31_io_reset),
    .io_out(regs_31_io_out),
    .io_enable(regs_31_io_enable)
  );
  FringeFF regs_32 ( // @[RegFile.scala 66:20:@34859.4]
    .clock(regs_32_clock),
    .reset(regs_32_reset),
    .io_in(regs_32_io_in),
    .io_reset(regs_32_io_reset),
    .io_out(regs_32_io_out),
    .io_enable(regs_32_io_enable)
  );
  FringeFF regs_33 ( // @[RegFile.scala 66:20:@34873.4]
    .clock(regs_33_clock),
    .reset(regs_33_reset),
    .io_in(regs_33_io_in),
    .io_reset(regs_33_io_reset),
    .io_out(regs_33_io_out),
    .io_enable(regs_33_io_enable)
  );
  FringeFF regs_34 ( // @[RegFile.scala 66:20:@34887.4]
    .clock(regs_34_clock),
    .reset(regs_34_reset),
    .io_in(regs_34_io_in),
    .io_reset(regs_34_io_reset),
    .io_out(regs_34_io_out),
    .io_enable(regs_34_io_enable)
  );
  FringeFF regs_35 ( // @[RegFile.scala 66:20:@34901.4]
    .clock(regs_35_clock),
    .reset(regs_35_reset),
    .io_in(regs_35_io_in),
    .io_reset(regs_35_io_reset),
    .io_out(regs_35_io_out),
    .io_enable(regs_35_io_enable)
  );
  FringeFF regs_36 ( // @[RegFile.scala 66:20:@34915.4]
    .clock(regs_36_clock),
    .reset(regs_36_reset),
    .io_in(regs_36_io_in),
    .io_reset(regs_36_io_reset),
    .io_out(regs_36_io_out),
    .io_enable(regs_36_io_enable)
  );
  FringeFF regs_37 ( // @[RegFile.scala 66:20:@34929.4]
    .clock(regs_37_clock),
    .reset(regs_37_reset),
    .io_in(regs_37_io_in),
    .io_reset(regs_37_io_reset),
    .io_out(regs_37_io_out),
    .io_enable(regs_37_io_enable)
  );
  FringeFF regs_38 ( // @[RegFile.scala 66:20:@34943.4]
    .clock(regs_38_clock),
    .reset(regs_38_reset),
    .io_in(regs_38_io_in),
    .io_reset(regs_38_io_reset),
    .io_out(regs_38_io_out),
    .io_enable(regs_38_io_enable)
  );
  FringeFF regs_39 ( // @[RegFile.scala 66:20:@34957.4]
    .clock(regs_39_clock),
    .reset(regs_39_reset),
    .io_in(regs_39_io_in),
    .io_reset(regs_39_io_reset),
    .io_out(regs_39_io_out),
    .io_enable(regs_39_io_enable)
  );
  FringeFF regs_40 ( // @[RegFile.scala 66:20:@34971.4]
    .clock(regs_40_clock),
    .reset(regs_40_reset),
    .io_in(regs_40_io_in),
    .io_reset(regs_40_io_reset),
    .io_out(regs_40_io_out),
    .io_enable(regs_40_io_enable)
  );
  FringeFF regs_41 ( // @[RegFile.scala 66:20:@34985.4]
    .clock(regs_41_clock),
    .reset(regs_41_reset),
    .io_in(regs_41_io_in),
    .io_reset(regs_41_io_reset),
    .io_out(regs_41_io_out),
    .io_enable(regs_41_io_enable)
  );
  FringeFF regs_42 ( // @[RegFile.scala 66:20:@34999.4]
    .clock(regs_42_clock),
    .reset(regs_42_reset),
    .io_in(regs_42_io_in),
    .io_reset(regs_42_io_reset),
    .io_out(regs_42_io_out),
    .io_enable(regs_42_io_enable)
  );
  FringeFF regs_43 ( // @[RegFile.scala 66:20:@35013.4]
    .clock(regs_43_clock),
    .reset(regs_43_reset),
    .io_in(regs_43_io_in),
    .io_reset(regs_43_io_reset),
    .io_out(regs_43_io_out),
    .io_enable(regs_43_io_enable)
  );
  FringeFF regs_44 ( // @[RegFile.scala 66:20:@35027.4]
    .clock(regs_44_clock),
    .reset(regs_44_reset),
    .io_in(regs_44_io_in),
    .io_reset(regs_44_io_reset),
    .io_out(regs_44_io_out),
    .io_enable(regs_44_io_enable)
  );
  FringeFF regs_45 ( // @[RegFile.scala 66:20:@35041.4]
    .clock(regs_45_clock),
    .reset(regs_45_reset),
    .io_in(regs_45_io_in),
    .io_reset(regs_45_io_reset),
    .io_out(regs_45_io_out),
    .io_enable(regs_45_io_enable)
  );
  FringeFF regs_46 ( // @[RegFile.scala 66:20:@35055.4]
    .clock(regs_46_clock),
    .reset(regs_46_reset),
    .io_in(regs_46_io_in),
    .io_reset(regs_46_io_reset),
    .io_out(regs_46_io_out),
    .io_enable(regs_46_io_enable)
  );
  FringeFF regs_47 ( // @[RegFile.scala 66:20:@35069.4]
    .clock(regs_47_clock),
    .reset(regs_47_reset),
    .io_in(regs_47_io_in),
    .io_reset(regs_47_io_reset),
    .io_out(regs_47_io_out),
    .io_enable(regs_47_io_enable)
  );
  FringeFF regs_48 ( // @[RegFile.scala 66:20:@35083.4]
    .clock(regs_48_clock),
    .reset(regs_48_reset),
    .io_in(regs_48_io_in),
    .io_reset(regs_48_io_reset),
    .io_out(regs_48_io_out),
    .io_enable(regs_48_io_enable)
  );
  FringeFF regs_49 ( // @[RegFile.scala 66:20:@35097.4]
    .clock(regs_49_clock),
    .reset(regs_49_reset),
    .io_in(regs_49_io_in),
    .io_reset(regs_49_io_reset),
    .io_out(regs_49_io_out),
    .io_enable(regs_49_io_enable)
  );
  FringeFF regs_50 ( // @[RegFile.scala 66:20:@35111.4]
    .clock(regs_50_clock),
    .reset(regs_50_reset),
    .io_in(regs_50_io_in),
    .io_reset(regs_50_io_reset),
    .io_out(regs_50_io_out),
    .io_enable(regs_50_io_enable)
  );
  FringeFF regs_51 ( // @[RegFile.scala 66:20:@35125.4]
    .clock(regs_51_clock),
    .reset(regs_51_reset),
    .io_in(regs_51_io_in),
    .io_reset(regs_51_io_reset),
    .io_out(regs_51_io_out),
    .io_enable(regs_51_io_enable)
  );
  FringeFF regs_52 ( // @[RegFile.scala 66:20:@35139.4]
    .clock(regs_52_clock),
    .reset(regs_52_reset),
    .io_in(regs_52_io_in),
    .io_reset(regs_52_io_reset),
    .io_out(regs_52_io_out),
    .io_enable(regs_52_io_enable)
  );
  FringeFF regs_53 ( // @[RegFile.scala 66:20:@35153.4]
    .clock(regs_53_clock),
    .reset(regs_53_reset),
    .io_in(regs_53_io_in),
    .io_reset(regs_53_io_reset),
    .io_out(regs_53_io_out),
    .io_enable(regs_53_io_enable)
  );
  FringeFF regs_54 ( // @[RegFile.scala 66:20:@35167.4]
    .clock(regs_54_clock),
    .reset(regs_54_reset),
    .io_in(regs_54_io_in),
    .io_reset(regs_54_io_reset),
    .io_out(regs_54_io_out),
    .io_enable(regs_54_io_enable)
  );
  FringeFF regs_55 ( // @[RegFile.scala 66:20:@35181.4]
    .clock(regs_55_clock),
    .reset(regs_55_reset),
    .io_in(regs_55_io_in),
    .io_reset(regs_55_io_reset),
    .io_out(regs_55_io_out),
    .io_enable(regs_55_io_enable)
  );
  FringeFF regs_56 ( // @[RegFile.scala 66:20:@35195.4]
    .clock(regs_56_clock),
    .reset(regs_56_reset),
    .io_in(regs_56_io_in),
    .io_reset(regs_56_io_reset),
    .io_out(regs_56_io_out),
    .io_enable(regs_56_io_enable)
  );
  FringeFF regs_57 ( // @[RegFile.scala 66:20:@35209.4]
    .clock(regs_57_clock),
    .reset(regs_57_reset),
    .io_in(regs_57_io_in),
    .io_reset(regs_57_io_reset),
    .io_out(regs_57_io_out),
    .io_enable(regs_57_io_enable)
  );
  FringeFF regs_58 ( // @[RegFile.scala 66:20:@35223.4]
    .clock(regs_58_clock),
    .reset(regs_58_reset),
    .io_in(regs_58_io_in),
    .io_reset(regs_58_io_reset),
    .io_out(regs_58_io_out),
    .io_enable(regs_58_io_enable)
  );
  FringeFF regs_59 ( // @[RegFile.scala 66:20:@35237.4]
    .clock(regs_59_clock),
    .reset(regs_59_reset),
    .io_in(regs_59_io_in),
    .io_reset(regs_59_io_reset),
    .io_out(regs_59_io_out),
    .io_enable(regs_59_io_enable)
  );
  FringeFF regs_60 ( // @[RegFile.scala 66:20:@35251.4]
    .clock(regs_60_clock),
    .reset(regs_60_reset),
    .io_in(regs_60_io_in),
    .io_reset(regs_60_io_reset),
    .io_out(regs_60_io_out),
    .io_enable(regs_60_io_enable)
  );
  FringeFF regs_61 ( // @[RegFile.scala 66:20:@35265.4]
    .clock(regs_61_clock),
    .reset(regs_61_reset),
    .io_in(regs_61_io_in),
    .io_reset(regs_61_io_reset),
    .io_out(regs_61_io_out),
    .io_enable(regs_61_io_enable)
  );
  FringeFF regs_62 ( // @[RegFile.scala 66:20:@35279.4]
    .clock(regs_62_clock),
    .reset(regs_62_reset),
    .io_in(regs_62_io_in),
    .io_reset(regs_62_io_reset),
    .io_out(regs_62_io_out),
    .io_enable(regs_62_io_enable)
  );
  FringeFF regs_63 ( // @[RegFile.scala 66:20:@35293.4]
    .clock(regs_63_clock),
    .reset(regs_63_reset),
    .io_in(regs_63_io_in),
    .io_reset(regs_63_io_reset),
    .io_out(regs_63_io_out),
    .io_enable(regs_63_io_enable)
  );
  FringeFF regs_64 ( // @[RegFile.scala 66:20:@35307.4]
    .clock(regs_64_clock),
    .reset(regs_64_reset),
    .io_in(regs_64_io_in),
    .io_reset(regs_64_io_reset),
    .io_out(regs_64_io_out),
    .io_enable(regs_64_io_enable)
  );
  FringeFF regs_65 ( // @[RegFile.scala 66:20:@35321.4]
    .clock(regs_65_clock),
    .reset(regs_65_reset),
    .io_in(regs_65_io_in),
    .io_reset(regs_65_io_reset),
    .io_out(regs_65_io_out),
    .io_enable(regs_65_io_enable)
  );
  FringeFF regs_66 ( // @[RegFile.scala 66:20:@35335.4]
    .clock(regs_66_clock),
    .reset(regs_66_reset),
    .io_in(regs_66_io_in),
    .io_reset(regs_66_io_reset),
    .io_out(regs_66_io_out),
    .io_enable(regs_66_io_enable)
  );
  FringeFF regs_67 ( // @[RegFile.scala 66:20:@35349.4]
    .clock(regs_67_clock),
    .reset(regs_67_reset),
    .io_in(regs_67_io_in),
    .io_reset(regs_67_io_reset),
    .io_out(regs_67_io_out),
    .io_enable(regs_67_io_enable)
  );
  FringeFF regs_68 ( // @[RegFile.scala 66:20:@35363.4]
    .clock(regs_68_clock),
    .reset(regs_68_reset),
    .io_in(regs_68_io_in),
    .io_reset(regs_68_io_reset),
    .io_out(regs_68_io_out),
    .io_enable(regs_68_io_enable)
  );
  FringeFF regs_69 ( // @[RegFile.scala 66:20:@35377.4]
    .clock(regs_69_clock),
    .reset(regs_69_reset),
    .io_in(regs_69_io_in),
    .io_reset(regs_69_io_reset),
    .io_out(regs_69_io_out),
    .io_enable(regs_69_io_enable)
  );
  FringeFF regs_70 ( // @[RegFile.scala 66:20:@35391.4]
    .clock(regs_70_clock),
    .reset(regs_70_reset),
    .io_in(regs_70_io_in),
    .io_reset(regs_70_io_reset),
    .io_out(regs_70_io_out),
    .io_enable(regs_70_io_enable)
  );
  FringeFF regs_71 ( // @[RegFile.scala 66:20:@35405.4]
    .clock(regs_71_clock),
    .reset(regs_71_reset),
    .io_in(regs_71_io_in),
    .io_reset(regs_71_io_reset),
    .io_out(regs_71_io_out),
    .io_enable(regs_71_io_enable)
  );
  FringeFF regs_72 ( // @[RegFile.scala 66:20:@35419.4]
    .clock(regs_72_clock),
    .reset(regs_72_reset),
    .io_in(regs_72_io_in),
    .io_reset(regs_72_io_reset),
    .io_out(regs_72_io_out),
    .io_enable(regs_72_io_enable)
  );
  FringeFF regs_73 ( // @[RegFile.scala 66:20:@35433.4]
    .clock(regs_73_clock),
    .reset(regs_73_reset),
    .io_in(regs_73_io_in),
    .io_reset(regs_73_io_reset),
    .io_out(regs_73_io_out),
    .io_enable(regs_73_io_enable)
  );
  FringeFF regs_74 ( // @[RegFile.scala 66:20:@35447.4]
    .clock(regs_74_clock),
    .reset(regs_74_reset),
    .io_in(regs_74_io_in),
    .io_reset(regs_74_io_reset),
    .io_out(regs_74_io_out),
    .io_enable(regs_74_io_enable)
  );
  FringeFF regs_75 ( // @[RegFile.scala 66:20:@35461.4]
    .clock(regs_75_clock),
    .reset(regs_75_reset),
    .io_in(regs_75_io_in),
    .io_reset(regs_75_io_reset),
    .io_out(regs_75_io_out),
    .io_enable(regs_75_io_enable)
  );
  FringeFF regs_76 ( // @[RegFile.scala 66:20:@35475.4]
    .clock(regs_76_clock),
    .reset(regs_76_reset),
    .io_in(regs_76_io_in),
    .io_reset(regs_76_io_reset),
    .io_out(regs_76_io_out),
    .io_enable(regs_76_io_enable)
  );
  FringeFF regs_77 ( // @[RegFile.scala 66:20:@35489.4]
    .clock(regs_77_clock),
    .reset(regs_77_reset),
    .io_in(regs_77_io_in),
    .io_reset(regs_77_io_reset),
    .io_out(regs_77_io_out),
    .io_enable(regs_77_io_enable)
  );
  FringeFF regs_78 ( // @[RegFile.scala 66:20:@35503.4]
    .clock(regs_78_clock),
    .reset(regs_78_reset),
    .io_in(regs_78_io_in),
    .io_reset(regs_78_io_reset),
    .io_out(regs_78_io_out),
    .io_enable(regs_78_io_enable)
  );
  FringeFF regs_79 ( // @[RegFile.scala 66:20:@35517.4]
    .clock(regs_79_clock),
    .reset(regs_79_reset),
    .io_in(regs_79_io_in),
    .io_reset(regs_79_io_reset),
    .io_out(regs_79_io_out),
    .io_enable(regs_79_io_enable)
  );
  FringeFF regs_80 ( // @[RegFile.scala 66:20:@35531.4]
    .clock(regs_80_clock),
    .reset(regs_80_reset),
    .io_in(regs_80_io_in),
    .io_reset(regs_80_io_reset),
    .io_out(regs_80_io_out),
    .io_enable(regs_80_io_enable)
  );
  FringeFF regs_81 ( // @[RegFile.scala 66:20:@35545.4]
    .clock(regs_81_clock),
    .reset(regs_81_reset),
    .io_in(regs_81_io_in),
    .io_reset(regs_81_io_reset),
    .io_out(regs_81_io_out),
    .io_enable(regs_81_io_enable)
  );
  FringeFF regs_82 ( // @[RegFile.scala 66:20:@35559.4]
    .clock(regs_82_clock),
    .reset(regs_82_reset),
    .io_in(regs_82_io_in),
    .io_reset(regs_82_io_reset),
    .io_out(regs_82_io_out),
    .io_enable(regs_82_io_enable)
  );
  FringeFF regs_83 ( // @[RegFile.scala 66:20:@35573.4]
    .clock(regs_83_clock),
    .reset(regs_83_reset),
    .io_in(regs_83_io_in),
    .io_reset(regs_83_io_reset),
    .io_out(regs_83_io_out),
    .io_enable(regs_83_io_enable)
  );
  FringeFF regs_84 ( // @[RegFile.scala 66:20:@35587.4]
    .clock(regs_84_clock),
    .reset(regs_84_reset),
    .io_in(regs_84_io_in),
    .io_reset(regs_84_io_reset),
    .io_out(regs_84_io_out),
    .io_enable(regs_84_io_enable)
  );
  FringeFF regs_85 ( // @[RegFile.scala 66:20:@35601.4]
    .clock(regs_85_clock),
    .reset(regs_85_reset),
    .io_in(regs_85_io_in),
    .io_reset(regs_85_io_reset),
    .io_out(regs_85_io_out),
    .io_enable(regs_85_io_enable)
  );
  FringeFF regs_86 ( // @[RegFile.scala 66:20:@35615.4]
    .clock(regs_86_clock),
    .reset(regs_86_reset),
    .io_in(regs_86_io_in),
    .io_reset(regs_86_io_reset),
    .io_out(regs_86_io_out),
    .io_enable(regs_86_io_enable)
  );
  FringeFF regs_87 ( // @[RegFile.scala 66:20:@35629.4]
    .clock(regs_87_clock),
    .reset(regs_87_reset),
    .io_in(regs_87_io_in),
    .io_reset(regs_87_io_reset),
    .io_out(regs_87_io_out),
    .io_enable(regs_87_io_enable)
  );
  FringeFF regs_88 ( // @[RegFile.scala 66:20:@35643.4]
    .clock(regs_88_clock),
    .reset(regs_88_reset),
    .io_in(regs_88_io_in),
    .io_reset(regs_88_io_reset),
    .io_out(regs_88_io_out),
    .io_enable(regs_88_io_enable)
  );
  FringeFF regs_89 ( // @[RegFile.scala 66:20:@35657.4]
    .clock(regs_89_clock),
    .reset(regs_89_reset),
    .io_in(regs_89_io_in),
    .io_reset(regs_89_io_reset),
    .io_out(regs_89_io_out),
    .io_enable(regs_89_io_enable)
  );
  FringeFF regs_90 ( // @[RegFile.scala 66:20:@35671.4]
    .clock(regs_90_clock),
    .reset(regs_90_reset),
    .io_in(regs_90_io_in),
    .io_reset(regs_90_io_reset),
    .io_out(regs_90_io_out),
    .io_enable(regs_90_io_enable)
  );
  FringeFF regs_91 ( // @[RegFile.scala 66:20:@35685.4]
    .clock(regs_91_clock),
    .reset(regs_91_reset),
    .io_in(regs_91_io_in),
    .io_reset(regs_91_io_reset),
    .io_out(regs_91_io_out),
    .io_enable(regs_91_io_enable)
  );
  FringeFF regs_92 ( // @[RegFile.scala 66:20:@35699.4]
    .clock(regs_92_clock),
    .reset(regs_92_reset),
    .io_in(regs_92_io_in),
    .io_reset(regs_92_io_reset),
    .io_out(regs_92_io_out),
    .io_enable(regs_92_io_enable)
  );
  FringeFF regs_93 ( // @[RegFile.scala 66:20:@35713.4]
    .clock(regs_93_clock),
    .reset(regs_93_reset),
    .io_in(regs_93_io_in),
    .io_reset(regs_93_io_reset),
    .io_out(regs_93_io_out),
    .io_enable(regs_93_io_enable)
  );
  FringeFF regs_94 ( // @[RegFile.scala 66:20:@35727.4]
    .clock(regs_94_clock),
    .reset(regs_94_reset),
    .io_in(regs_94_io_in),
    .io_reset(regs_94_io_reset),
    .io_out(regs_94_io_out),
    .io_enable(regs_94_io_enable)
  );
  FringeFF regs_95 ( // @[RegFile.scala 66:20:@35741.4]
    .clock(regs_95_clock),
    .reset(regs_95_reset),
    .io_in(regs_95_io_in),
    .io_reset(regs_95_io_reset),
    .io_out(regs_95_io_out),
    .io_enable(regs_95_io_enable)
  );
  FringeFF regs_96 ( // @[RegFile.scala 66:20:@35755.4]
    .clock(regs_96_clock),
    .reset(regs_96_reset),
    .io_in(regs_96_io_in),
    .io_reset(regs_96_io_reset),
    .io_out(regs_96_io_out),
    .io_enable(regs_96_io_enable)
  );
  FringeFF regs_97 ( // @[RegFile.scala 66:20:@35769.4]
    .clock(regs_97_clock),
    .reset(regs_97_reset),
    .io_in(regs_97_io_in),
    .io_reset(regs_97_io_reset),
    .io_out(regs_97_io_out),
    .io_enable(regs_97_io_enable)
  );
  FringeFF regs_98 ( // @[RegFile.scala 66:20:@35783.4]
    .clock(regs_98_clock),
    .reset(regs_98_reset),
    .io_in(regs_98_io_in),
    .io_reset(regs_98_io_reset),
    .io_out(regs_98_io_out),
    .io_enable(regs_98_io_enable)
  );
  FringeFF regs_99 ( // @[RegFile.scala 66:20:@35797.4]
    .clock(regs_99_clock),
    .reset(regs_99_reset),
    .io_in(regs_99_io_in),
    .io_reset(regs_99_io_reset),
    .io_out(regs_99_io_out),
    .io_enable(regs_99_io_enable)
  );
  FringeFF regs_100 ( // @[RegFile.scala 66:20:@35811.4]
    .clock(regs_100_clock),
    .reset(regs_100_reset),
    .io_in(regs_100_io_in),
    .io_reset(regs_100_io_reset),
    .io_out(regs_100_io_out),
    .io_enable(regs_100_io_enable)
  );
  FringeFF regs_101 ( // @[RegFile.scala 66:20:@35825.4]
    .clock(regs_101_clock),
    .reset(regs_101_reset),
    .io_in(regs_101_io_in),
    .io_reset(regs_101_io_reset),
    .io_out(regs_101_io_out),
    .io_enable(regs_101_io_enable)
  );
  FringeFF regs_102 ( // @[RegFile.scala 66:20:@35839.4]
    .clock(regs_102_clock),
    .reset(regs_102_reset),
    .io_in(regs_102_io_in),
    .io_reset(regs_102_io_reset),
    .io_out(regs_102_io_out),
    .io_enable(regs_102_io_enable)
  );
  FringeFF regs_103 ( // @[RegFile.scala 66:20:@35853.4]
    .clock(regs_103_clock),
    .reset(regs_103_reset),
    .io_in(regs_103_io_in),
    .io_reset(regs_103_io_reset),
    .io_out(regs_103_io_out),
    .io_enable(regs_103_io_enable)
  );
  FringeFF regs_104 ( // @[RegFile.scala 66:20:@35867.4]
    .clock(regs_104_clock),
    .reset(regs_104_reset),
    .io_in(regs_104_io_in),
    .io_reset(regs_104_io_reset),
    .io_out(regs_104_io_out),
    .io_enable(regs_104_io_enable)
  );
  FringeFF regs_105 ( // @[RegFile.scala 66:20:@35881.4]
    .clock(regs_105_clock),
    .reset(regs_105_reset),
    .io_in(regs_105_io_in),
    .io_reset(regs_105_io_reset),
    .io_out(regs_105_io_out),
    .io_enable(regs_105_io_enable)
  );
  FringeFF regs_106 ( // @[RegFile.scala 66:20:@35895.4]
    .clock(regs_106_clock),
    .reset(regs_106_reset),
    .io_in(regs_106_io_in),
    .io_reset(regs_106_io_reset),
    .io_out(regs_106_io_out),
    .io_enable(regs_106_io_enable)
  );
  FringeFF regs_107 ( // @[RegFile.scala 66:20:@35909.4]
    .clock(regs_107_clock),
    .reset(regs_107_reset),
    .io_in(regs_107_io_in),
    .io_reset(regs_107_io_reset),
    .io_out(regs_107_io_out),
    .io_enable(regs_107_io_enable)
  );
  FringeFF regs_108 ( // @[RegFile.scala 66:20:@35923.4]
    .clock(regs_108_clock),
    .reset(regs_108_reset),
    .io_in(regs_108_io_in),
    .io_reset(regs_108_io_reset),
    .io_out(regs_108_io_out),
    .io_enable(regs_108_io_enable)
  );
  FringeFF regs_109 ( // @[RegFile.scala 66:20:@35937.4]
    .clock(regs_109_clock),
    .reset(regs_109_reset),
    .io_in(regs_109_io_in),
    .io_reset(regs_109_io_reset),
    .io_out(regs_109_io_out),
    .io_enable(regs_109_io_enable)
  );
  FringeFF regs_110 ( // @[RegFile.scala 66:20:@35951.4]
    .clock(regs_110_clock),
    .reset(regs_110_reset),
    .io_in(regs_110_io_in),
    .io_reset(regs_110_io_reset),
    .io_out(regs_110_io_out),
    .io_enable(regs_110_io_enable)
  );
  FringeFF regs_111 ( // @[RegFile.scala 66:20:@35965.4]
    .clock(regs_111_clock),
    .reset(regs_111_reset),
    .io_in(regs_111_io_in),
    .io_reset(regs_111_io_reset),
    .io_out(regs_111_io_out),
    .io_enable(regs_111_io_enable)
  );
  FringeFF regs_112 ( // @[RegFile.scala 66:20:@35979.4]
    .clock(regs_112_clock),
    .reset(regs_112_reset),
    .io_in(regs_112_io_in),
    .io_reset(regs_112_io_reset),
    .io_out(regs_112_io_out),
    .io_enable(regs_112_io_enable)
  );
  FringeFF regs_113 ( // @[RegFile.scala 66:20:@35993.4]
    .clock(regs_113_clock),
    .reset(regs_113_reset),
    .io_in(regs_113_io_in),
    .io_reset(regs_113_io_reset),
    .io_out(regs_113_io_out),
    .io_enable(regs_113_io_enable)
  );
  FringeFF regs_114 ( // @[RegFile.scala 66:20:@36007.4]
    .clock(regs_114_clock),
    .reset(regs_114_reset),
    .io_in(regs_114_io_in),
    .io_reset(regs_114_io_reset),
    .io_out(regs_114_io_out),
    .io_enable(regs_114_io_enable)
  );
  FringeFF regs_115 ( // @[RegFile.scala 66:20:@36021.4]
    .clock(regs_115_clock),
    .reset(regs_115_reset),
    .io_in(regs_115_io_in),
    .io_reset(regs_115_io_reset),
    .io_out(regs_115_io_out),
    .io_enable(regs_115_io_enable)
  );
  FringeFF regs_116 ( // @[RegFile.scala 66:20:@36035.4]
    .clock(regs_116_clock),
    .reset(regs_116_reset),
    .io_in(regs_116_io_in),
    .io_reset(regs_116_io_reset),
    .io_out(regs_116_io_out),
    .io_enable(regs_116_io_enable)
  );
  FringeFF regs_117 ( // @[RegFile.scala 66:20:@36049.4]
    .clock(regs_117_clock),
    .reset(regs_117_reset),
    .io_in(regs_117_io_in),
    .io_reset(regs_117_io_reset),
    .io_out(regs_117_io_out),
    .io_enable(regs_117_io_enable)
  );
  FringeFF regs_118 ( // @[RegFile.scala 66:20:@36063.4]
    .clock(regs_118_clock),
    .reset(regs_118_reset),
    .io_in(regs_118_io_in),
    .io_reset(regs_118_io_reset),
    .io_out(regs_118_io_out),
    .io_enable(regs_118_io_enable)
  );
  FringeFF regs_119 ( // @[RegFile.scala 66:20:@36077.4]
    .clock(regs_119_clock),
    .reset(regs_119_reset),
    .io_in(regs_119_io_in),
    .io_reset(regs_119_io_reset),
    .io_out(regs_119_io_out),
    .io_enable(regs_119_io_enable)
  );
  FringeFF regs_120 ( // @[RegFile.scala 66:20:@36091.4]
    .clock(regs_120_clock),
    .reset(regs_120_reset),
    .io_in(regs_120_io_in),
    .io_reset(regs_120_io_reset),
    .io_out(regs_120_io_out),
    .io_enable(regs_120_io_enable)
  );
  FringeFF regs_121 ( // @[RegFile.scala 66:20:@36105.4]
    .clock(regs_121_clock),
    .reset(regs_121_reset),
    .io_in(regs_121_io_in),
    .io_reset(regs_121_io_reset),
    .io_out(regs_121_io_out),
    .io_enable(regs_121_io_enable)
  );
  FringeFF regs_122 ( // @[RegFile.scala 66:20:@36119.4]
    .clock(regs_122_clock),
    .reset(regs_122_reset),
    .io_in(regs_122_io_in),
    .io_reset(regs_122_io_reset),
    .io_out(regs_122_io_out),
    .io_enable(regs_122_io_enable)
  );
  FringeFF regs_123 ( // @[RegFile.scala 66:20:@36133.4]
    .clock(regs_123_clock),
    .reset(regs_123_reset),
    .io_in(regs_123_io_in),
    .io_reset(regs_123_io_reset),
    .io_out(regs_123_io_out),
    .io_enable(regs_123_io_enable)
  );
  FringeFF regs_124 ( // @[RegFile.scala 66:20:@36147.4]
    .clock(regs_124_clock),
    .reset(regs_124_reset),
    .io_in(regs_124_io_in),
    .io_reset(regs_124_io_reset),
    .io_out(regs_124_io_out),
    .io_enable(regs_124_io_enable)
  );
  FringeFF regs_125 ( // @[RegFile.scala 66:20:@36161.4]
    .clock(regs_125_clock),
    .reset(regs_125_reset),
    .io_in(regs_125_io_in),
    .io_reset(regs_125_io_reset),
    .io_out(regs_125_io_out),
    .io_enable(regs_125_io_enable)
  );
  FringeFF regs_126 ( // @[RegFile.scala 66:20:@36175.4]
    .clock(regs_126_clock),
    .reset(regs_126_reset),
    .io_in(regs_126_io_in),
    .io_reset(regs_126_io_reset),
    .io_out(regs_126_io_out),
    .io_enable(regs_126_io_enable)
  );
  FringeFF regs_127 ( // @[RegFile.scala 66:20:@36189.4]
    .clock(regs_127_clock),
    .reset(regs_127_reset),
    .io_in(regs_127_io_in),
    .io_reset(regs_127_io_reset),
    .io_out(regs_127_io_out),
    .io_enable(regs_127_io_enable)
  );
  FringeFF regs_128 ( // @[RegFile.scala 66:20:@36203.4]
    .clock(regs_128_clock),
    .reset(regs_128_reset),
    .io_in(regs_128_io_in),
    .io_reset(regs_128_io_reset),
    .io_out(regs_128_io_out),
    .io_enable(regs_128_io_enable)
  );
  FringeFF regs_129 ( // @[RegFile.scala 66:20:@36217.4]
    .clock(regs_129_clock),
    .reset(regs_129_reset),
    .io_in(regs_129_io_in),
    .io_reset(regs_129_io_reset),
    .io_out(regs_129_io_out),
    .io_enable(regs_129_io_enable)
  );
  FringeFF regs_130 ( // @[RegFile.scala 66:20:@36231.4]
    .clock(regs_130_clock),
    .reset(regs_130_reset),
    .io_in(regs_130_io_in),
    .io_reset(regs_130_io_reset),
    .io_out(regs_130_io_out),
    .io_enable(regs_130_io_enable)
  );
  FringeFF regs_131 ( // @[RegFile.scala 66:20:@36245.4]
    .clock(regs_131_clock),
    .reset(regs_131_reset),
    .io_in(regs_131_io_in),
    .io_reset(regs_131_io_reset),
    .io_out(regs_131_io_out),
    .io_enable(regs_131_io_enable)
  );
  FringeFF regs_132 ( // @[RegFile.scala 66:20:@36259.4]
    .clock(regs_132_clock),
    .reset(regs_132_reset),
    .io_in(regs_132_io_in),
    .io_reset(regs_132_io_reset),
    .io_out(regs_132_io_out),
    .io_enable(regs_132_io_enable)
  );
  FringeFF regs_133 ( // @[RegFile.scala 66:20:@36273.4]
    .clock(regs_133_clock),
    .reset(regs_133_reset),
    .io_in(regs_133_io_in),
    .io_reset(regs_133_io_reset),
    .io_out(regs_133_io_out),
    .io_enable(regs_133_io_enable)
  );
  FringeFF regs_134 ( // @[RegFile.scala 66:20:@36287.4]
    .clock(regs_134_clock),
    .reset(regs_134_reset),
    .io_in(regs_134_io_in),
    .io_reset(regs_134_io_reset),
    .io_out(regs_134_io_out),
    .io_enable(regs_134_io_enable)
  );
  FringeFF regs_135 ( // @[RegFile.scala 66:20:@36301.4]
    .clock(regs_135_clock),
    .reset(regs_135_reset),
    .io_in(regs_135_io_in),
    .io_reset(regs_135_io_reset),
    .io_out(regs_135_io_out),
    .io_enable(regs_135_io_enable)
  );
  FringeFF regs_136 ( // @[RegFile.scala 66:20:@36315.4]
    .clock(regs_136_clock),
    .reset(regs_136_reset),
    .io_in(regs_136_io_in),
    .io_reset(regs_136_io_reset),
    .io_out(regs_136_io_out),
    .io_enable(regs_136_io_enable)
  );
  FringeFF regs_137 ( // @[RegFile.scala 66:20:@36329.4]
    .clock(regs_137_clock),
    .reset(regs_137_reset),
    .io_in(regs_137_io_in),
    .io_reset(regs_137_io_reset),
    .io_out(regs_137_io_out),
    .io_enable(regs_137_io_enable)
  );
  FringeFF regs_138 ( // @[RegFile.scala 66:20:@36343.4]
    .clock(regs_138_clock),
    .reset(regs_138_reset),
    .io_in(regs_138_io_in),
    .io_reset(regs_138_io_reset),
    .io_out(regs_138_io_out),
    .io_enable(regs_138_io_enable)
  );
  FringeFF regs_139 ( // @[RegFile.scala 66:20:@36357.4]
    .clock(regs_139_clock),
    .reset(regs_139_reset),
    .io_in(regs_139_io_in),
    .io_reset(regs_139_io_reset),
    .io_out(regs_139_io_out),
    .io_enable(regs_139_io_enable)
  );
  FringeFF regs_140 ( // @[RegFile.scala 66:20:@36371.4]
    .clock(regs_140_clock),
    .reset(regs_140_reset),
    .io_in(regs_140_io_in),
    .io_reset(regs_140_io_reset),
    .io_out(regs_140_io_out),
    .io_enable(regs_140_io_enable)
  );
  FringeFF regs_141 ( // @[RegFile.scala 66:20:@36385.4]
    .clock(regs_141_clock),
    .reset(regs_141_reset),
    .io_in(regs_141_io_in),
    .io_reset(regs_141_io_reset),
    .io_out(regs_141_io_out),
    .io_enable(regs_141_io_enable)
  );
  FringeFF regs_142 ( // @[RegFile.scala 66:20:@36399.4]
    .clock(regs_142_clock),
    .reset(regs_142_reset),
    .io_in(regs_142_io_in),
    .io_reset(regs_142_io_reset),
    .io_out(regs_142_io_out),
    .io_enable(regs_142_io_enable)
  );
  FringeFF regs_143 ( // @[RegFile.scala 66:20:@36413.4]
    .clock(regs_143_clock),
    .reset(regs_143_reset),
    .io_in(regs_143_io_in),
    .io_reset(regs_143_io_reset),
    .io_out(regs_143_io_out),
    .io_enable(regs_143_io_enable)
  );
  FringeFF regs_144 ( // @[RegFile.scala 66:20:@36427.4]
    .clock(regs_144_clock),
    .reset(regs_144_reset),
    .io_in(regs_144_io_in),
    .io_reset(regs_144_io_reset),
    .io_out(regs_144_io_out),
    .io_enable(regs_144_io_enable)
  );
  FringeFF regs_145 ( // @[RegFile.scala 66:20:@36441.4]
    .clock(regs_145_clock),
    .reset(regs_145_reset),
    .io_in(regs_145_io_in),
    .io_reset(regs_145_io_reset),
    .io_out(regs_145_io_out),
    .io_enable(regs_145_io_enable)
  );
  FringeFF regs_146 ( // @[RegFile.scala 66:20:@36455.4]
    .clock(regs_146_clock),
    .reset(regs_146_reset),
    .io_in(regs_146_io_in),
    .io_reset(regs_146_io_reset),
    .io_out(regs_146_io_out),
    .io_enable(regs_146_io_enable)
  );
  FringeFF regs_147 ( // @[RegFile.scala 66:20:@36469.4]
    .clock(regs_147_clock),
    .reset(regs_147_reset),
    .io_in(regs_147_io_in),
    .io_reset(regs_147_io_reset),
    .io_out(regs_147_io_out),
    .io_enable(regs_147_io_enable)
  );
  FringeFF regs_148 ( // @[RegFile.scala 66:20:@36483.4]
    .clock(regs_148_clock),
    .reset(regs_148_reset),
    .io_in(regs_148_io_in),
    .io_reset(regs_148_io_reset),
    .io_out(regs_148_io_out),
    .io_enable(regs_148_io_enable)
  );
  FringeFF regs_149 ( // @[RegFile.scala 66:20:@36497.4]
    .clock(regs_149_clock),
    .reset(regs_149_reset),
    .io_in(regs_149_io_in),
    .io_reset(regs_149_io_reset),
    .io_out(regs_149_io_out),
    .io_enable(regs_149_io_enable)
  );
  FringeFF regs_150 ( // @[RegFile.scala 66:20:@36511.4]
    .clock(regs_150_clock),
    .reset(regs_150_reset),
    .io_in(regs_150_io_in),
    .io_reset(regs_150_io_reset),
    .io_out(regs_150_io_out),
    .io_enable(regs_150_io_enable)
  );
  FringeFF regs_151 ( // @[RegFile.scala 66:20:@36525.4]
    .clock(regs_151_clock),
    .reset(regs_151_reset),
    .io_in(regs_151_io_in),
    .io_reset(regs_151_io_reset),
    .io_out(regs_151_io_out),
    .io_enable(regs_151_io_enable)
  );
  FringeFF regs_152 ( // @[RegFile.scala 66:20:@36539.4]
    .clock(regs_152_clock),
    .reset(regs_152_reset),
    .io_in(regs_152_io_in),
    .io_reset(regs_152_io_reset),
    .io_out(regs_152_io_out),
    .io_enable(regs_152_io_enable)
  );
  FringeFF regs_153 ( // @[RegFile.scala 66:20:@36553.4]
    .clock(regs_153_clock),
    .reset(regs_153_reset),
    .io_in(regs_153_io_in),
    .io_reset(regs_153_io_reset),
    .io_out(regs_153_io_out),
    .io_enable(regs_153_io_enable)
  );
  FringeFF regs_154 ( // @[RegFile.scala 66:20:@36567.4]
    .clock(regs_154_clock),
    .reset(regs_154_reset),
    .io_in(regs_154_io_in),
    .io_reset(regs_154_io_reset),
    .io_out(regs_154_io_out),
    .io_enable(regs_154_io_enable)
  );
  FringeFF regs_155 ( // @[RegFile.scala 66:20:@36581.4]
    .clock(regs_155_clock),
    .reset(regs_155_reset),
    .io_in(regs_155_io_in),
    .io_reset(regs_155_io_reset),
    .io_out(regs_155_io_out),
    .io_enable(regs_155_io_enable)
  );
  FringeFF regs_156 ( // @[RegFile.scala 66:20:@36595.4]
    .clock(regs_156_clock),
    .reset(regs_156_reset),
    .io_in(regs_156_io_in),
    .io_reset(regs_156_io_reset),
    .io_out(regs_156_io_out),
    .io_enable(regs_156_io_enable)
  );
  FringeFF regs_157 ( // @[RegFile.scala 66:20:@36609.4]
    .clock(regs_157_clock),
    .reset(regs_157_reset),
    .io_in(regs_157_io_in),
    .io_reset(regs_157_io_reset),
    .io_out(regs_157_io_out),
    .io_enable(regs_157_io_enable)
  );
  FringeFF regs_158 ( // @[RegFile.scala 66:20:@36623.4]
    .clock(regs_158_clock),
    .reset(regs_158_reset),
    .io_in(regs_158_io_in),
    .io_reset(regs_158_io_reset),
    .io_out(regs_158_io_out),
    .io_enable(regs_158_io_enable)
  );
  FringeFF regs_159 ( // @[RegFile.scala 66:20:@36637.4]
    .clock(regs_159_clock),
    .reset(regs_159_reset),
    .io_in(regs_159_io_in),
    .io_reset(regs_159_io_reset),
    .io_out(regs_159_io_out),
    .io_enable(regs_159_io_enable)
  );
  FringeFF regs_160 ( // @[RegFile.scala 66:20:@36651.4]
    .clock(regs_160_clock),
    .reset(regs_160_reset),
    .io_in(regs_160_io_in),
    .io_reset(regs_160_io_reset),
    .io_out(regs_160_io_out),
    .io_enable(regs_160_io_enable)
  );
  FringeFF regs_161 ( // @[RegFile.scala 66:20:@36665.4]
    .clock(regs_161_clock),
    .reset(regs_161_reset),
    .io_in(regs_161_io_in),
    .io_reset(regs_161_io_reset),
    .io_out(regs_161_io_out),
    .io_enable(regs_161_io_enable)
  );
  FringeFF regs_162 ( // @[RegFile.scala 66:20:@36679.4]
    .clock(regs_162_clock),
    .reset(regs_162_reset),
    .io_in(regs_162_io_in),
    .io_reset(regs_162_io_reset),
    .io_out(regs_162_io_out),
    .io_enable(regs_162_io_enable)
  );
  FringeFF regs_163 ( // @[RegFile.scala 66:20:@36693.4]
    .clock(regs_163_clock),
    .reset(regs_163_reset),
    .io_in(regs_163_io_in),
    .io_reset(regs_163_io_reset),
    .io_out(regs_163_io_out),
    .io_enable(regs_163_io_enable)
  );
  FringeFF regs_164 ( // @[RegFile.scala 66:20:@36707.4]
    .clock(regs_164_clock),
    .reset(regs_164_reset),
    .io_in(regs_164_io_in),
    .io_reset(regs_164_io_reset),
    .io_out(regs_164_io_out),
    .io_enable(regs_164_io_enable)
  );
  FringeFF regs_165 ( // @[RegFile.scala 66:20:@36721.4]
    .clock(regs_165_clock),
    .reset(regs_165_reset),
    .io_in(regs_165_io_in),
    .io_reset(regs_165_io_reset),
    .io_out(regs_165_io_out),
    .io_enable(regs_165_io_enable)
  );
  FringeFF regs_166 ( // @[RegFile.scala 66:20:@36735.4]
    .clock(regs_166_clock),
    .reset(regs_166_reset),
    .io_in(regs_166_io_in),
    .io_reset(regs_166_io_reset),
    .io_out(regs_166_io_out),
    .io_enable(regs_166_io_enable)
  );
  FringeFF regs_167 ( // @[RegFile.scala 66:20:@36749.4]
    .clock(regs_167_clock),
    .reset(regs_167_reset),
    .io_in(regs_167_io_in),
    .io_reset(regs_167_io_reset),
    .io_out(regs_167_io_out),
    .io_enable(regs_167_io_enable)
  );
  FringeFF regs_168 ( // @[RegFile.scala 66:20:@36763.4]
    .clock(regs_168_clock),
    .reset(regs_168_reset),
    .io_in(regs_168_io_in),
    .io_reset(regs_168_io_reset),
    .io_out(regs_168_io_out),
    .io_enable(regs_168_io_enable)
  );
  FringeFF regs_169 ( // @[RegFile.scala 66:20:@36777.4]
    .clock(regs_169_clock),
    .reset(regs_169_reset),
    .io_in(regs_169_io_in),
    .io_reset(regs_169_io_reset),
    .io_out(regs_169_io_out),
    .io_enable(regs_169_io_enable)
  );
  FringeFF regs_170 ( // @[RegFile.scala 66:20:@36791.4]
    .clock(regs_170_clock),
    .reset(regs_170_reset),
    .io_in(regs_170_io_in),
    .io_reset(regs_170_io_reset),
    .io_out(regs_170_io_out),
    .io_enable(regs_170_io_enable)
  );
  FringeFF regs_171 ( // @[RegFile.scala 66:20:@36805.4]
    .clock(regs_171_clock),
    .reset(regs_171_reset),
    .io_in(regs_171_io_in),
    .io_reset(regs_171_io_reset),
    .io_out(regs_171_io_out),
    .io_enable(regs_171_io_enable)
  );
  FringeFF regs_172 ( // @[RegFile.scala 66:20:@36819.4]
    .clock(regs_172_clock),
    .reset(regs_172_reset),
    .io_in(regs_172_io_in),
    .io_reset(regs_172_io_reset),
    .io_out(regs_172_io_out),
    .io_enable(regs_172_io_enable)
  );
  FringeFF regs_173 ( // @[RegFile.scala 66:20:@36833.4]
    .clock(regs_173_clock),
    .reset(regs_173_reset),
    .io_in(regs_173_io_in),
    .io_reset(regs_173_io_reset),
    .io_out(regs_173_io_out),
    .io_enable(regs_173_io_enable)
  );
  FringeFF regs_174 ( // @[RegFile.scala 66:20:@36847.4]
    .clock(regs_174_clock),
    .reset(regs_174_reset),
    .io_in(regs_174_io_in),
    .io_reset(regs_174_io_reset),
    .io_out(regs_174_io_out),
    .io_enable(regs_174_io_enable)
  );
  FringeFF regs_175 ( // @[RegFile.scala 66:20:@36861.4]
    .clock(regs_175_clock),
    .reset(regs_175_reset),
    .io_in(regs_175_io_in),
    .io_reset(regs_175_io_reset),
    .io_out(regs_175_io_out),
    .io_enable(regs_175_io_enable)
  );
  FringeFF regs_176 ( // @[RegFile.scala 66:20:@36875.4]
    .clock(regs_176_clock),
    .reset(regs_176_reset),
    .io_in(regs_176_io_in),
    .io_reset(regs_176_io_reset),
    .io_out(regs_176_io_out),
    .io_enable(regs_176_io_enable)
  );
  FringeFF regs_177 ( // @[RegFile.scala 66:20:@36889.4]
    .clock(regs_177_clock),
    .reset(regs_177_reset),
    .io_in(regs_177_io_in),
    .io_reset(regs_177_io_reset),
    .io_out(regs_177_io_out),
    .io_enable(regs_177_io_enable)
  );
  FringeFF regs_178 ( // @[RegFile.scala 66:20:@36903.4]
    .clock(regs_178_clock),
    .reset(regs_178_reset),
    .io_in(regs_178_io_in),
    .io_reset(regs_178_io_reset),
    .io_out(regs_178_io_out),
    .io_enable(regs_178_io_enable)
  );
  FringeFF regs_179 ( // @[RegFile.scala 66:20:@36917.4]
    .clock(regs_179_clock),
    .reset(regs_179_reset),
    .io_in(regs_179_io_in),
    .io_reset(regs_179_io_reset),
    .io_out(regs_179_io_out),
    .io_enable(regs_179_io_enable)
  );
  FringeFF regs_180 ( // @[RegFile.scala 66:20:@36931.4]
    .clock(regs_180_clock),
    .reset(regs_180_reset),
    .io_in(regs_180_io_in),
    .io_reset(regs_180_io_reset),
    .io_out(regs_180_io_out),
    .io_enable(regs_180_io_enable)
  );
  FringeFF regs_181 ( // @[RegFile.scala 66:20:@36945.4]
    .clock(regs_181_clock),
    .reset(regs_181_reset),
    .io_in(regs_181_io_in),
    .io_reset(regs_181_io_reset),
    .io_out(regs_181_io_out),
    .io_enable(regs_181_io_enable)
  );
  FringeFF regs_182 ( // @[RegFile.scala 66:20:@36959.4]
    .clock(regs_182_clock),
    .reset(regs_182_reset),
    .io_in(regs_182_io_in),
    .io_reset(regs_182_io_reset),
    .io_out(regs_182_io_out),
    .io_enable(regs_182_io_enable)
  );
  FringeFF regs_183 ( // @[RegFile.scala 66:20:@36973.4]
    .clock(regs_183_clock),
    .reset(regs_183_reset),
    .io_in(regs_183_io_in),
    .io_reset(regs_183_io_reset),
    .io_out(regs_183_io_out),
    .io_enable(regs_183_io_enable)
  );
  FringeFF regs_184 ( // @[RegFile.scala 66:20:@36987.4]
    .clock(regs_184_clock),
    .reset(regs_184_reset),
    .io_in(regs_184_io_in),
    .io_reset(regs_184_io_reset),
    .io_out(regs_184_io_out),
    .io_enable(regs_184_io_enable)
  );
  FringeFF regs_185 ( // @[RegFile.scala 66:20:@37001.4]
    .clock(regs_185_clock),
    .reset(regs_185_reset),
    .io_in(regs_185_io_in),
    .io_reset(regs_185_io_reset),
    .io_out(regs_185_io_out),
    .io_enable(regs_185_io_enable)
  );
  FringeFF regs_186 ( // @[RegFile.scala 66:20:@37015.4]
    .clock(regs_186_clock),
    .reset(regs_186_reset),
    .io_in(regs_186_io_in),
    .io_reset(regs_186_io_reset),
    .io_out(regs_186_io_out),
    .io_enable(regs_186_io_enable)
  );
  FringeFF regs_187 ( // @[RegFile.scala 66:20:@37029.4]
    .clock(regs_187_clock),
    .reset(regs_187_reset),
    .io_in(regs_187_io_in),
    .io_reset(regs_187_io_reset),
    .io_out(regs_187_io_out),
    .io_enable(regs_187_io_enable)
  );
  FringeFF regs_188 ( // @[RegFile.scala 66:20:@37043.4]
    .clock(regs_188_clock),
    .reset(regs_188_reset),
    .io_in(regs_188_io_in),
    .io_reset(regs_188_io_reset),
    .io_out(regs_188_io_out),
    .io_enable(regs_188_io_enable)
  );
  FringeFF regs_189 ( // @[RegFile.scala 66:20:@37057.4]
    .clock(regs_189_clock),
    .reset(regs_189_reset),
    .io_in(regs_189_io_in),
    .io_reset(regs_189_io_reset),
    .io_out(regs_189_io_out),
    .io_enable(regs_189_io_enable)
  );
  FringeFF regs_190 ( // @[RegFile.scala 66:20:@37071.4]
    .clock(regs_190_clock),
    .reset(regs_190_reset),
    .io_in(regs_190_io_in),
    .io_reset(regs_190_io_reset),
    .io_out(regs_190_io_out),
    .io_enable(regs_190_io_enable)
  );
  FringeFF regs_191 ( // @[RegFile.scala 66:20:@37085.4]
    .clock(regs_191_clock),
    .reset(regs_191_reset),
    .io_in(regs_191_io_in),
    .io_reset(regs_191_io_reset),
    .io_out(regs_191_io_out),
    .io_enable(regs_191_io_enable)
  );
  FringeFF regs_192 ( // @[RegFile.scala 66:20:@37099.4]
    .clock(regs_192_clock),
    .reset(regs_192_reset),
    .io_in(regs_192_io_in),
    .io_reset(regs_192_io_reset),
    .io_out(regs_192_io_out),
    .io_enable(regs_192_io_enable)
  );
  FringeFF regs_193 ( // @[RegFile.scala 66:20:@37113.4]
    .clock(regs_193_clock),
    .reset(regs_193_reset),
    .io_in(regs_193_io_in),
    .io_reset(regs_193_io_reset),
    .io_out(regs_193_io_out),
    .io_enable(regs_193_io_enable)
  );
  FringeFF regs_194 ( // @[RegFile.scala 66:20:@37127.4]
    .clock(regs_194_clock),
    .reset(regs_194_reset),
    .io_in(regs_194_io_in),
    .io_reset(regs_194_io_reset),
    .io_out(regs_194_io_out),
    .io_enable(regs_194_io_enable)
  );
  FringeFF regs_195 ( // @[RegFile.scala 66:20:@37141.4]
    .clock(regs_195_clock),
    .reset(regs_195_reset),
    .io_in(regs_195_io_in),
    .io_reset(regs_195_io_reset),
    .io_out(regs_195_io_out),
    .io_enable(regs_195_io_enable)
  );
  FringeFF regs_196 ( // @[RegFile.scala 66:20:@37155.4]
    .clock(regs_196_clock),
    .reset(regs_196_reset),
    .io_in(regs_196_io_in),
    .io_reset(regs_196_io_reset),
    .io_out(regs_196_io_out),
    .io_enable(regs_196_io_enable)
  );
  FringeFF regs_197 ( // @[RegFile.scala 66:20:@37169.4]
    .clock(regs_197_clock),
    .reset(regs_197_reset),
    .io_in(regs_197_io_in),
    .io_reset(regs_197_io_reset),
    .io_out(regs_197_io_out),
    .io_enable(regs_197_io_enable)
  );
  FringeFF regs_198 ( // @[RegFile.scala 66:20:@37183.4]
    .clock(regs_198_clock),
    .reset(regs_198_reset),
    .io_in(regs_198_io_in),
    .io_reset(regs_198_io_reset),
    .io_out(regs_198_io_out),
    .io_enable(regs_198_io_enable)
  );
  FringeFF regs_199 ( // @[RegFile.scala 66:20:@37197.4]
    .clock(regs_199_clock),
    .reset(regs_199_reset),
    .io_in(regs_199_io_in),
    .io_reset(regs_199_io_reset),
    .io_out(regs_199_io_out),
    .io_enable(regs_199_io_enable)
  );
  FringeFF regs_200 ( // @[RegFile.scala 66:20:@37211.4]
    .clock(regs_200_clock),
    .reset(regs_200_reset),
    .io_in(regs_200_io_in),
    .io_reset(regs_200_io_reset),
    .io_out(regs_200_io_out),
    .io_enable(regs_200_io_enable)
  );
  FringeFF regs_201 ( // @[RegFile.scala 66:20:@37225.4]
    .clock(regs_201_clock),
    .reset(regs_201_reset),
    .io_in(regs_201_io_in),
    .io_reset(regs_201_io_reset),
    .io_out(regs_201_io_out),
    .io_enable(regs_201_io_enable)
  );
  FringeFF regs_202 ( // @[RegFile.scala 66:20:@37239.4]
    .clock(regs_202_clock),
    .reset(regs_202_reset),
    .io_in(regs_202_io_in),
    .io_reset(regs_202_io_reset),
    .io_out(regs_202_io_out),
    .io_enable(regs_202_io_enable)
  );
  FringeFF regs_203 ( // @[RegFile.scala 66:20:@37253.4]
    .clock(regs_203_clock),
    .reset(regs_203_reset),
    .io_in(regs_203_io_in),
    .io_reset(regs_203_io_reset),
    .io_out(regs_203_io_out),
    .io_enable(regs_203_io_enable)
  );
  FringeFF regs_204 ( // @[RegFile.scala 66:20:@37267.4]
    .clock(regs_204_clock),
    .reset(regs_204_reset),
    .io_in(regs_204_io_in),
    .io_reset(regs_204_io_reset),
    .io_out(regs_204_io_out),
    .io_enable(regs_204_io_enable)
  );
  FringeFF regs_205 ( // @[RegFile.scala 66:20:@37281.4]
    .clock(regs_205_clock),
    .reset(regs_205_reset),
    .io_in(regs_205_io_in),
    .io_reset(regs_205_io_reset),
    .io_out(regs_205_io_out),
    .io_enable(regs_205_io_enable)
  );
  FringeFF regs_206 ( // @[RegFile.scala 66:20:@37295.4]
    .clock(regs_206_clock),
    .reset(regs_206_reset),
    .io_in(regs_206_io_in),
    .io_reset(regs_206_io_reset),
    .io_out(regs_206_io_out),
    .io_enable(regs_206_io_enable)
  );
  FringeFF regs_207 ( // @[RegFile.scala 66:20:@37309.4]
    .clock(regs_207_clock),
    .reset(regs_207_reset),
    .io_in(regs_207_io_in),
    .io_reset(regs_207_io_reset),
    .io_out(regs_207_io_out),
    .io_enable(regs_207_io_enable)
  );
  FringeFF regs_208 ( // @[RegFile.scala 66:20:@37323.4]
    .clock(regs_208_clock),
    .reset(regs_208_reset),
    .io_in(regs_208_io_in),
    .io_reset(regs_208_io_reset),
    .io_out(regs_208_io_out),
    .io_enable(regs_208_io_enable)
  );
  FringeFF regs_209 ( // @[RegFile.scala 66:20:@37337.4]
    .clock(regs_209_clock),
    .reset(regs_209_reset),
    .io_in(regs_209_io_in),
    .io_reset(regs_209_io_reset),
    .io_out(regs_209_io_out),
    .io_enable(regs_209_io_enable)
  );
  FringeFF regs_210 ( // @[RegFile.scala 66:20:@37351.4]
    .clock(regs_210_clock),
    .reset(regs_210_reset),
    .io_in(regs_210_io_in),
    .io_reset(regs_210_io_reset),
    .io_out(regs_210_io_out),
    .io_enable(regs_210_io_enable)
  );
  FringeFF regs_211 ( // @[RegFile.scala 66:20:@37365.4]
    .clock(regs_211_clock),
    .reset(regs_211_reset),
    .io_in(regs_211_io_in),
    .io_reset(regs_211_io_reset),
    .io_out(regs_211_io_out),
    .io_enable(regs_211_io_enable)
  );
  FringeFF regs_212 ( // @[RegFile.scala 66:20:@37379.4]
    .clock(regs_212_clock),
    .reset(regs_212_reset),
    .io_in(regs_212_io_in),
    .io_reset(regs_212_io_reset),
    .io_out(regs_212_io_out),
    .io_enable(regs_212_io_enable)
  );
  FringeFF regs_213 ( // @[RegFile.scala 66:20:@37393.4]
    .clock(regs_213_clock),
    .reset(regs_213_reset),
    .io_in(regs_213_io_in),
    .io_reset(regs_213_io_reset),
    .io_out(regs_213_io_out),
    .io_enable(regs_213_io_enable)
  );
  FringeFF regs_214 ( // @[RegFile.scala 66:20:@37407.4]
    .clock(regs_214_clock),
    .reset(regs_214_reset),
    .io_in(regs_214_io_in),
    .io_reset(regs_214_io_reset),
    .io_out(regs_214_io_out),
    .io_enable(regs_214_io_enable)
  );
  FringeFF regs_215 ( // @[RegFile.scala 66:20:@37421.4]
    .clock(regs_215_clock),
    .reset(regs_215_reset),
    .io_in(regs_215_io_in),
    .io_reset(regs_215_io_reset),
    .io_out(regs_215_io_out),
    .io_enable(regs_215_io_enable)
  );
  FringeFF regs_216 ( // @[RegFile.scala 66:20:@37435.4]
    .clock(regs_216_clock),
    .reset(regs_216_reset),
    .io_in(regs_216_io_in),
    .io_reset(regs_216_io_reset),
    .io_out(regs_216_io_out),
    .io_enable(regs_216_io_enable)
  );
  FringeFF regs_217 ( // @[RegFile.scala 66:20:@37449.4]
    .clock(regs_217_clock),
    .reset(regs_217_reset),
    .io_in(regs_217_io_in),
    .io_reset(regs_217_io_reset),
    .io_out(regs_217_io_out),
    .io_enable(regs_217_io_enable)
  );
  FringeFF regs_218 ( // @[RegFile.scala 66:20:@37463.4]
    .clock(regs_218_clock),
    .reset(regs_218_reset),
    .io_in(regs_218_io_in),
    .io_reset(regs_218_io_reset),
    .io_out(regs_218_io_out),
    .io_enable(regs_218_io_enable)
  );
  FringeFF regs_219 ( // @[RegFile.scala 66:20:@37477.4]
    .clock(regs_219_clock),
    .reset(regs_219_reset),
    .io_in(regs_219_io_in),
    .io_reset(regs_219_io_reset),
    .io_out(regs_219_io_out),
    .io_enable(regs_219_io_enable)
  );
  FringeFF regs_220 ( // @[RegFile.scala 66:20:@37491.4]
    .clock(regs_220_clock),
    .reset(regs_220_reset),
    .io_in(regs_220_io_in),
    .io_reset(regs_220_io_reset),
    .io_out(regs_220_io_out),
    .io_enable(regs_220_io_enable)
  );
  FringeFF regs_221 ( // @[RegFile.scala 66:20:@37505.4]
    .clock(regs_221_clock),
    .reset(regs_221_reset),
    .io_in(regs_221_io_in),
    .io_reset(regs_221_io_reset),
    .io_out(regs_221_io_out),
    .io_enable(regs_221_io_enable)
  );
  FringeFF regs_222 ( // @[RegFile.scala 66:20:@37519.4]
    .clock(regs_222_clock),
    .reset(regs_222_reset),
    .io_in(regs_222_io_in),
    .io_reset(regs_222_io_reset),
    .io_out(regs_222_io_out),
    .io_enable(regs_222_io_enable)
  );
  FringeFF regs_223 ( // @[RegFile.scala 66:20:@37533.4]
    .clock(regs_223_clock),
    .reset(regs_223_reset),
    .io_in(regs_223_io_in),
    .io_reset(regs_223_io_reset),
    .io_out(regs_223_io_out),
    .io_enable(regs_223_io_enable)
  );
  FringeFF regs_224 ( // @[RegFile.scala 66:20:@37547.4]
    .clock(regs_224_clock),
    .reset(regs_224_reset),
    .io_in(regs_224_io_in),
    .io_reset(regs_224_io_reset),
    .io_out(regs_224_io_out),
    .io_enable(regs_224_io_enable)
  );
  FringeFF regs_225 ( // @[RegFile.scala 66:20:@37561.4]
    .clock(regs_225_clock),
    .reset(regs_225_reset),
    .io_in(regs_225_io_in),
    .io_reset(regs_225_io_reset),
    .io_out(regs_225_io_out),
    .io_enable(regs_225_io_enable)
  );
  FringeFF regs_226 ( // @[RegFile.scala 66:20:@37575.4]
    .clock(regs_226_clock),
    .reset(regs_226_reset),
    .io_in(regs_226_io_in),
    .io_reset(regs_226_io_reset),
    .io_out(regs_226_io_out),
    .io_enable(regs_226_io_enable)
  );
  FringeFF regs_227 ( // @[RegFile.scala 66:20:@37589.4]
    .clock(regs_227_clock),
    .reset(regs_227_reset),
    .io_in(regs_227_io_in),
    .io_reset(regs_227_io_reset),
    .io_out(regs_227_io_out),
    .io_enable(regs_227_io_enable)
  );
  FringeFF regs_228 ( // @[RegFile.scala 66:20:@37603.4]
    .clock(regs_228_clock),
    .reset(regs_228_reset),
    .io_in(regs_228_io_in),
    .io_reset(regs_228_io_reset),
    .io_out(regs_228_io_out),
    .io_enable(regs_228_io_enable)
  );
  FringeFF regs_229 ( // @[RegFile.scala 66:20:@37617.4]
    .clock(regs_229_clock),
    .reset(regs_229_reset),
    .io_in(regs_229_io_in),
    .io_reset(regs_229_io_reset),
    .io_out(regs_229_io_out),
    .io_enable(regs_229_io_enable)
  );
  FringeFF regs_230 ( // @[RegFile.scala 66:20:@37631.4]
    .clock(regs_230_clock),
    .reset(regs_230_reset),
    .io_in(regs_230_io_in),
    .io_reset(regs_230_io_reset),
    .io_out(regs_230_io_out),
    .io_enable(regs_230_io_enable)
  );
  FringeFF regs_231 ( // @[RegFile.scala 66:20:@37645.4]
    .clock(regs_231_clock),
    .reset(regs_231_reset),
    .io_in(regs_231_io_in),
    .io_reset(regs_231_io_reset),
    .io_out(regs_231_io_out),
    .io_enable(regs_231_io_enable)
  );
  FringeFF regs_232 ( // @[RegFile.scala 66:20:@37659.4]
    .clock(regs_232_clock),
    .reset(regs_232_reset),
    .io_in(regs_232_io_in),
    .io_reset(regs_232_io_reset),
    .io_out(regs_232_io_out),
    .io_enable(regs_232_io_enable)
  );
  FringeFF regs_233 ( // @[RegFile.scala 66:20:@37673.4]
    .clock(regs_233_clock),
    .reset(regs_233_reset),
    .io_in(regs_233_io_in),
    .io_reset(regs_233_io_reset),
    .io_out(regs_233_io_out),
    .io_enable(regs_233_io_enable)
  );
  FringeFF regs_234 ( // @[RegFile.scala 66:20:@37687.4]
    .clock(regs_234_clock),
    .reset(regs_234_reset),
    .io_in(regs_234_io_in),
    .io_reset(regs_234_io_reset),
    .io_out(regs_234_io_out),
    .io_enable(regs_234_io_enable)
  );
  FringeFF regs_235 ( // @[RegFile.scala 66:20:@37701.4]
    .clock(regs_235_clock),
    .reset(regs_235_reset),
    .io_in(regs_235_io_in),
    .io_reset(regs_235_io_reset),
    .io_out(regs_235_io_out),
    .io_enable(regs_235_io_enable)
  );
  FringeFF regs_236 ( // @[RegFile.scala 66:20:@37715.4]
    .clock(regs_236_clock),
    .reset(regs_236_reset),
    .io_in(regs_236_io_in),
    .io_reset(regs_236_io_reset),
    .io_out(regs_236_io_out),
    .io_enable(regs_236_io_enable)
  );
  FringeFF regs_237 ( // @[RegFile.scala 66:20:@37729.4]
    .clock(regs_237_clock),
    .reset(regs_237_reset),
    .io_in(regs_237_io_in),
    .io_reset(regs_237_io_reset),
    .io_out(regs_237_io_out),
    .io_enable(regs_237_io_enable)
  );
  FringeFF regs_238 ( // @[RegFile.scala 66:20:@37743.4]
    .clock(regs_238_clock),
    .reset(regs_238_reset),
    .io_in(regs_238_io_in),
    .io_reset(regs_238_io_reset),
    .io_out(regs_238_io_out),
    .io_enable(regs_238_io_enable)
  );
  FringeFF regs_239 ( // @[RegFile.scala 66:20:@37757.4]
    .clock(regs_239_clock),
    .reset(regs_239_reset),
    .io_in(regs_239_io_in),
    .io_reset(regs_239_io_reset),
    .io_out(regs_239_io_out),
    .io_enable(regs_239_io_enable)
  );
  FringeFF regs_240 ( // @[RegFile.scala 66:20:@37771.4]
    .clock(regs_240_clock),
    .reset(regs_240_reset),
    .io_in(regs_240_io_in),
    .io_reset(regs_240_io_reset),
    .io_out(regs_240_io_out),
    .io_enable(regs_240_io_enable)
  );
  FringeFF regs_241 ( // @[RegFile.scala 66:20:@37785.4]
    .clock(regs_241_clock),
    .reset(regs_241_reset),
    .io_in(regs_241_io_in),
    .io_reset(regs_241_io_reset),
    .io_out(regs_241_io_out),
    .io_enable(regs_241_io_enable)
  );
  FringeFF regs_242 ( // @[RegFile.scala 66:20:@37799.4]
    .clock(regs_242_clock),
    .reset(regs_242_reset),
    .io_in(regs_242_io_in),
    .io_reset(regs_242_io_reset),
    .io_out(regs_242_io_out),
    .io_enable(regs_242_io_enable)
  );
  FringeFF regs_243 ( // @[RegFile.scala 66:20:@37813.4]
    .clock(regs_243_clock),
    .reset(regs_243_reset),
    .io_in(regs_243_io_in),
    .io_reset(regs_243_io_reset),
    .io_out(regs_243_io_out),
    .io_enable(regs_243_io_enable)
  );
  FringeFF regs_244 ( // @[RegFile.scala 66:20:@37827.4]
    .clock(regs_244_clock),
    .reset(regs_244_reset),
    .io_in(regs_244_io_in),
    .io_reset(regs_244_io_reset),
    .io_out(regs_244_io_out),
    .io_enable(regs_244_io_enable)
  );
  FringeFF regs_245 ( // @[RegFile.scala 66:20:@37841.4]
    .clock(regs_245_clock),
    .reset(regs_245_reset),
    .io_in(regs_245_io_in),
    .io_reset(regs_245_io_reset),
    .io_out(regs_245_io_out),
    .io_enable(regs_245_io_enable)
  );
  FringeFF regs_246 ( // @[RegFile.scala 66:20:@37855.4]
    .clock(regs_246_clock),
    .reset(regs_246_reset),
    .io_in(regs_246_io_in),
    .io_reset(regs_246_io_reset),
    .io_out(regs_246_io_out),
    .io_enable(regs_246_io_enable)
  );
  FringeFF regs_247 ( // @[RegFile.scala 66:20:@37869.4]
    .clock(regs_247_clock),
    .reset(regs_247_reset),
    .io_in(regs_247_io_in),
    .io_reset(regs_247_io_reset),
    .io_out(regs_247_io_out),
    .io_enable(regs_247_io_enable)
  );
  FringeFF regs_248 ( // @[RegFile.scala 66:20:@37883.4]
    .clock(regs_248_clock),
    .reset(regs_248_reset),
    .io_in(regs_248_io_in),
    .io_reset(regs_248_io_reset),
    .io_out(regs_248_io_out),
    .io_enable(regs_248_io_enable)
  );
  FringeFF regs_249 ( // @[RegFile.scala 66:20:@37897.4]
    .clock(regs_249_clock),
    .reset(regs_249_reset),
    .io_in(regs_249_io_in),
    .io_reset(regs_249_io_reset),
    .io_out(regs_249_io_out),
    .io_enable(regs_249_io_enable)
  );
  FringeFF regs_250 ( // @[RegFile.scala 66:20:@37911.4]
    .clock(regs_250_clock),
    .reset(regs_250_reset),
    .io_in(regs_250_io_in),
    .io_reset(regs_250_io_reset),
    .io_out(regs_250_io_out),
    .io_enable(regs_250_io_enable)
  );
  FringeFF regs_251 ( // @[RegFile.scala 66:20:@37925.4]
    .clock(regs_251_clock),
    .reset(regs_251_reset),
    .io_in(regs_251_io_in),
    .io_reset(regs_251_io_reset),
    .io_out(regs_251_io_out),
    .io_enable(regs_251_io_enable)
  );
  FringeFF regs_252 ( // @[RegFile.scala 66:20:@37939.4]
    .clock(regs_252_clock),
    .reset(regs_252_reset),
    .io_in(regs_252_io_in),
    .io_reset(regs_252_io_reset),
    .io_out(regs_252_io_out),
    .io_enable(regs_252_io_enable)
  );
  FringeFF regs_253 ( // @[RegFile.scala 66:20:@37953.4]
    .clock(regs_253_clock),
    .reset(regs_253_reset),
    .io_in(regs_253_io_in),
    .io_reset(regs_253_io_reset),
    .io_out(regs_253_io_out),
    .io_enable(regs_253_io_enable)
  );
  FringeFF regs_254 ( // @[RegFile.scala 66:20:@37967.4]
    .clock(regs_254_clock),
    .reset(regs_254_reset),
    .io_in(regs_254_io_in),
    .io_reset(regs_254_io_reset),
    .io_out(regs_254_io_out),
    .io_enable(regs_254_io_enable)
  );
  FringeFF regs_255 ( // @[RegFile.scala 66:20:@37981.4]
    .clock(regs_255_clock),
    .reset(regs_255_reset),
    .io_in(regs_255_io_in),
    .io_reset(regs_255_io_reset),
    .io_out(regs_255_io_out),
    .io_enable(regs_255_io_enable)
  );
  FringeFF regs_256 ( // @[RegFile.scala 66:20:@37995.4]
    .clock(regs_256_clock),
    .reset(regs_256_reset),
    .io_in(regs_256_io_in),
    .io_reset(regs_256_io_reset),
    .io_out(regs_256_io_out),
    .io_enable(regs_256_io_enable)
  );
  FringeFF regs_257 ( // @[RegFile.scala 66:20:@38009.4]
    .clock(regs_257_clock),
    .reset(regs_257_reset),
    .io_in(regs_257_io_in),
    .io_reset(regs_257_io_reset),
    .io_out(regs_257_io_out),
    .io_enable(regs_257_io_enable)
  );
  FringeFF regs_258 ( // @[RegFile.scala 66:20:@38023.4]
    .clock(regs_258_clock),
    .reset(regs_258_reset),
    .io_in(regs_258_io_in),
    .io_reset(regs_258_io_reset),
    .io_out(regs_258_io_out),
    .io_enable(regs_258_io_enable)
  );
  FringeFF regs_259 ( // @[RegFile.scala 66:20:@38037.4]
    .clock(regs_259_clock),
    .reset(regs_259_reset),
    .io_in(regs_259_io_in),
    .io_reset(regs_259_io_reset),
    .io_out(regs_259_io_out),
    .io_enable(regs_259_io_enable)
  );
  FringeFF regs_260 ( // @[RegFile.scala 66:20:@38051.4]
    .clock(regs_260_clock),
    .reset(regs_260_reset),
    .io_in(regs_260_io_in),
    .io_reset(regs_260_io_reset),
    .io_out(regs_260_io_out),
    .io_enable(regs_260_io_enable)
  );
  FringeFF regs_261 ( // @[RegFile.scala 66:20:@38065.4]
    .clock(regs_261_clock),
    .reset(regs_261_reset),
    .io_in(regs_261_io_in),
    .io_reset(regs_261_io_reset),
    .io_out(regs_261_io_out),
    .io_enable(regs_261_io_enable)
  );
  FringeFF regs_262 ( // @[RegFile.scala 66:20:@38079.4]
    .clock(regs_262_clock),
    .reset(regs_262_reset),
    .io_in(regs_262_io_in),
    .io_reset(regs_262_io_reset),
    .io_out(regs_262_io_out),
    .io_enable(regs_262_io_enable)
  );
  FringeFF regs_263 ( // @[RegFile.scala 66:20:@38093.4]
    .clock(regs_263_clock),
    .reset(regs_263_reset),
    .io_in(regs_263_io_in),
    .io_reset(regs_263_io_reset),
    .io_out(regs_263_io_out),
    .io_enable(regs_263_io_enable)
  );
  FringeFF regs_264 ( // @[RegFile.scala 66:20:@38107.4]
    .clock(regs_264_clock),
    .reset(regs_264_reset),
    .io_in(regs_264_io_in),
    .io_reset(regs_264_io_reset),
    .io_out(regs_264_io_out),
    .io_enable(regs_264_io_enable)
  );
  FringeFF regs_265 ( // @[RegFile.scala 66:20:@38121.4]
    .clock(regs_265_clock),
    .reset(regs_265_reset),
    .io_in(regs_265_io_in),
    .io_reset(regs_265_io_reset),
    .io_out(regs_265_io_out),
    .io_enable(regs_265_io_enable)
  );
  FringeFF regs_266 ( // @[RegFile.scala 66:20:@38135.4]
    .clock(regs_266_clock),
    .reset(regs_266_reset),
    .io_in(regs_266_io_in),
    .io_reset(regs_266_io_reset),
    .io_out(regs_266_io_out),
    .io_enable(regs_266_io_enable)
  );
  FringeFF regs_267 ( // @[RegFile.scala 66:20:@38149.4]
    .clock(regs_267_clock),
    .reset(regs_267_reset),
    .io_in(regs_267_io_in),
    .io_reset(regs_267_io_reset),
    .io_out(regs_267_io_out),
    .io_enable(regs_267_io_enable)
  );
  FringeFF regs_268 ( // @[RegFile.scala 66:20:@38163.4]
    .clock(regs_268_clock),
    .reset(regs_268_reset),
    .io_in(regs_268_io_in),
    .io_reset(regs_268_io_reset),
    .io_out(regs_268_io_out),
    .io_enable(regs_268_io_enable)
  );
  FringeFF regs_269 ( // @[RegFile.scala 66:20:@38177.4]
    .clock(regs_269_clock),
    .reset(regs_269_reset),
    .io_in(regs_269_io_in),
    .io_reset(regs_269_io_reset),
    .io_out(regs_269_io_out),
    .io_enable(regs_269_io_enable)
  );
  FringeFF regs_270 ( // @[RegFile.scala 66:20:@38191.4]
    .clock(regs_270_clock),
    .reset(regs_270_reset),
    .io_in(regs_270_io_in),
    .io_reset(regs_270_io_reset),
    .io_out(regs_270_io_out),
    .io_enable(regs_270_io_enable)
  );
  FringeFF regs_271 ( // @[RegFile.scala 66:20:@38205.4]
    .clock(regs_271_clock),
    .reset(regs_271_reset),
    .io_in(regs_271_io_in),
    .io_reset(regs_271_io_reset),
    .io_out(regs_271_io_out),
    .io_enable(regs_271_io_enable)
  );
  FringeFF regs_272 ( // @[RegFile.scala 66:20:@38219.4]
    .clock(regs_272_clock),
    .reset(regs_272_reset),
    .io_in(regs_272_io_in),
    .io_reset(regs_272_io_reset),
    .io_out(regs_272_io_out),
    .io_enable(regs_272_io_enable)
  );
  FringeFF regs_273 ( // @[RegFile.scala 66:20:@38233.4]
    .clock(regs_273_clock),
    .reset(regs_273_reset),
    .io_in(regs_273_io_in),
    .io_reset(regs_273_io_reset),
    .io_out(regs_273_io_out),
    .io_enable(regs_273_io_enable)
  );
  FringeFF regs_274 ( // @[RegFile.scala 66:20:@38247.4]
    .clock(regs_274_clock),
    .reset(regs_274_reset),
    .io_in(regs_274_io_in),
    .io_reset(regs_274_io_reset),
    .io_out(regs_274_io_out),
    .io_enable(regs_274_io_enable)
  );
  FringeFF regs_275 ( // @[RegFile.scala 66:20:@38261.4]
    .clock(regs_275_clock),
    .reset(regs_275_reset),
    .io_in(regs_275_io_in),
    .io_reset(regs_275_io_reset),
    .io_out(regs_275_io_out),
    .io_enable(regs_275_io_enable)
  );
  FringeFF regs_276 ( // @[RegFile.scala 66:20:@38275.4]
    .clock(regs_276_clock),
    .reset(regs_276_reset),
    .io_in(regs_276_io_in),
    .io_reset(regs_276_io_reset),
    .io_out(regs_276_io_out),
    .io_enable(regs_276_io_enable)
  );
  FringeFF regs_277 ( // @[RegFile.scala 66:20:@38289.4]
    .clock(regs_277_clock),
    .reset(regs_277_reset),
    .io_in(regs_277_io_in),
    .io_reset(regs_277_io_reset),
    .io_out(regs_277_io_out),
    .io_enable(regs_277_io_enable)
  );
  FringeFF regs_278 ( // @[RegFile.scala 66:20:@38303.4]
    .clock(regs_278_clock),
    .reset(regs_278_reset),
    .io_in(regs_278_io_in),
    .io_reset(regs_278_io_reset),
    .io_out(regs_278_io_out),
    .io_enable(regs_278_io_enable)
  );
  FringeFF regs_279 ( // @[RegFile.scala 66:20:@38317.4]
    .clock(regs_279_clock),
    .reset(regs_279_reset),
    .io_in(regs_279_io_in),
    .io_reset(regs_279_io_reset),
    .io_out(regs_279_io_out),
    .io_enable(regs_279_io_enable)
  );
  FringeFF regs_280 ( // @[RegFile.scala 66:20:@38331.4]
    .clock(regs_280_clock),
    .reset(regs_280_reset),
    .io_in(regs_280_io_in),
    .io_reset(regs_280_io_reset),
    .io_out(regs_280_io_out),
    .io_enable(regs_280_io_enable)
  );
  FringeFF regs_281 ( // @[RegFile.scala 66:20:@38345.4]
    .clock(regs_281_clock),
    .reset(regs_281_reset),
    .io_in(regs_281_io_in),
    .io_reset(regs_281_io_reset),
    .io_out(regs_281_io_out),
    .io_enable(regs_281_io_enable)
  );
  FringeFF regs_282 ( // @[RegFile.scala 66:20:@38359.4]
    .clock(regs_282_clock),
    .reset(regs_282_reset),
    .io_in(regs_282_io_in),
    .io_reset(regs_282_io_reset),
    .io_out(regs_282_io_out),
    .io_enable(regs_282_io_enable)
  );
  FringeFF regs_283 ( // @[RegFile.scala 66:20:@38373.4]
    .clock(regs_283_clock),
    .reset(regs_283_reset),
    .io_in(regs_283_io_in),
    .io_reset(regs_283_io_reset),
    .io_out(regs_283_io_out),
    .io_enable(regs_283_io_enable)
  );
  FringeFF regs_284 ( // @[RegFile.scala 66:20:@38387.4]
    .clock(regs_284_clock),
    .reset(regs_284_reset),
    .io_in(regs_284_io_in),
    .io_reset(regs_284_io_reset),
    .io_out(regs_284_io_out),
    .io_enable(regs_284_io_enable)
  );
  FringeFF regs_285 ( // @[RegFile.scala 66:20:@38401.4]
    .clock(regs_285_clock),
    .reset(regs_285_reset),
    .io_in(regs_285_io_in),
    .io_reset(regs_285_io_reset),
    .io_out(regs_285_io_out),
    .io_enable(regs_285_io_enable)
  );
  FringeFF regs_286 ( // @[RegFile.scala 66:20:@38415.4]
    .clock(regs_286_clock),
    .reset(regs_286_reset),
    .io_in(regs_286_io_in),
    .io_reset(regs_286_io_reset),
    .io_out(regs_286_io_out),
    .io_enable(regs_286_io_enable)
  );
  FringeFF regs_287 ( // @[RegFile.scala 66:20:@38429.4]
    .clock(regs_287_clock),
    .reset(regs_287_reset),
    .io_in(regs_287_io_in),
    .io_reset(regs_287_io_reset),
    .io_out(regs_287_io_out),
    .io_enable(regs_287_io_enable)
  );
  FringeFF regs_288 ( // @[RegFile.scala 66:20:@38443.4]
    .clock(regs_288_clock),
    .reset(regs_288_reset),
    .io_in(regs_288_io_in),
    .io_reset(regs_288_io_reset),
    .io_out(regs_288_io_out),
    .io_enable(regs_288_io_enable)
  );
  FringeFF regs_289 ( // @[RegFile.scala 66:20:@38457.4]
    .clock(regs_289_clock),
    .reset(regs_289_reset),
    .io_in(regs_289_io_in),
    .io_reset(regs_289_io_reset),
    .io_out(regs_289_io_out),
    .io_enable(regs_289_io_enable)
  );
  FringeFF regs_290 ( // @[RegFile.scala 66:20:@38471.4]
    .clock(regs_290_clock),
    .reset(regs_290_reset),
    .io_in(regs_290_io_in),
    .io_reset(regs_290_io_reset),
    .io_out(regs_290_io_out),
    .io_enable(regs_290_io_enable)
  );
  FringeFF regs_291 ( // @[RegFile.scala 66:20:@38485.4]
    .clock(regs_291_clock),
    .reset(regs_291_reset),
    .io_in(regs_291_io_in),
    .io_reset(regs_291_io_reset),
    .io_out(regs_291_io_out),
    .io_enable(regs_291_io_enable)
  );
  FringeFF regs_292 ( // @[RegFile.scala 66:20:@38499.4]
    .clock(regs_292_clock),
    .reset(regs_292_reset),
    .io_in(regs_292_io_in),
    .io_reset(regs_292_io_reset),
    .io_out(regs_292_io_out),
    .io_enable(regs_292_io_enable)
  );
  FringeFF regs_293 ( // @[RegFile.scala 66:20:@38513.4]
    .clock(regs_293_clock),
    .reset(regs_293_reset),
    .io_in(regs_293_io_in),
    .io_reset(regs_293_io_reset),
    .io_out(regs_293_io_out),
    .io_enable(regs_293_io_enable)
  );
  FringeFF regs_294 ( // @[RegFile.scala 66:20:@38527.4]
    .clock(regs_294_clock),
    .reset(regs_294_reset),
    .io_in(regs_294_io_in),
    .io_reset(regs_294_io_reset),
    .io_out(regs_294_io_out),
    .io_enable(regs_294_io_enable)
  );
  FringeFF regs_295 ( // @[RegFile.scala 66:20:@38541.4]
    .clock(regs_295_clock),
    .reset(regs_295_reset),
    .io_in(regs_295_io_in),
    .io_reset(regs_295_io_reset),
    .io_out(regs_295_io_out),
    .io_enable(regs_295_io_enable)
  );
  FringeFF regs_296 ( // @[RegFile.scala 66:20:@38555.4]
    .clock(regs_296_clock),
    .reset(regs_296_reset),
    .io_in(regs_296_io_in),
    .io_reset(regs_296_io_reset),
    .io_out(regs_296_io_out),
    .io_enable(regs_296_io_enable)
  );
  FringeFF regs_297 ( // @[RegFile.scala 66:20:@38569.4]
    .clock(regs_297_clock),
    .reset(regs_297_reset),
    .io_in(regs_297_io_in),
    .io_reset(regs_297_io_reset),
    .io_out(regs_297_io_out),
    .io_enable(regs_297_io_enable)
  );
  FringeFF regs_298 ( // @[RegFile.scala 66:20:@38583.4]
    .clock(regs_298_clock),
    .reset(regs_298_reset),
    .io_in(regs_298_io_in),
    .io_reset(regs_298_io_reset),
    .io_out(regs_298_io_out),
    .io_enable(regs_298_io_enable)
  );
  FringeFF regs_299 ( // @[RegFile.scala 66:20:@38597.4]
    .clock(regs_299_clock),
    .reset(regs_299_reset),
    .io_in(regs_299_io_in),
    .io_reset(regs_299_io_reset),
    .io_out(regs_299_io_out),
    .io_enable(regs_299_io_enable)
  );
  FringeFF regs_300 ( // @[RegFile.scala 66:20:@38611.4]
    .clock(regs_300_clock),
    .reset(regs_300_reset),
    .io_in(regs_300_io_in),
    .io_reset(regs_300_io_reset),
    .io_out(regs_300_io_out),
    .io_enable(regs_300_io_enable)
  );
  FringeFF regs_301 ( // @[RegFile.scala 66:20:@38625.4]
    .clock(regs_301_clock),
    .reset(regs_301_reset),
    .io_in(regs_301_io_in),
    .io_reset(regs_301_io_reset),
    .io_out(regs_301_io_out),
    .io_enable(regs_301_io_enable)
  );
  FringeFF regs_302 ( // @[RegFile.scala 66:20:@38639.4]
    .clock(regs_302_clock),
    .reset(regs_302_reset),
    .io_in(regs_302_io_in),
    .io_reset(regs_302_io_reset),
    .io_out(regs_302_io_out),
    .io_enable(regs_302_io_enable)
  );
  FringeFF regs_303 ( // @[RegFile.scala 66:20:@38653.4]
    .clock(regs_303_clock),
    .reset(regs_303_reset),
    .io_in(regs_303_io_in),
    .io_reset(regs_303_io_reset),
    .io_out(regs_303_io_out),
    .io_enable(regs_303_io_enable)
  );
  FringeFF regs_304 ( // @[RegFile.scala 66:20:@38667.4]
    .clock(regs_304_clock),
    .reset(regs_304_reset),
    .io_in(regs_304_io_in),
    .io_reset(regs_304_io_reset),
    .io_out(regs_304_io_out),
    .io_enable(regs_304_io_enable)
  );
  FringeFF regs_305 ( // @[RegFile.scala 66:20:@38681.4]
    .clock(regs_305_clock),
    .reset(regs_305_reset),
    .io_in(regs_305_io_in),
    .io_reset(regs_305_io_reset),
    .io_out(regs_305_io_out),
    .io_enable(regs_305_io_enable)
  );
  FringeFF regs_306 ( // @[RegFile.scala 66:20:@38695.4]
    .clock(regs_306_clock),
    .reset(regs_306_reset),
    .io_in(regs_306_io_in),
    .io_reset(regs_306_io_reset),
    .io_out(regs_306_io_out),
    .io_enable(regs_306_io_enable)
  );
  FringeFF regs_307 ( // @[RegFile.scala 66:20:@38709.4]
    .clock(regs_307_clock),
    .reset(regs_307_reset),
    .io_in(regs_307_io_in),
    .io_reset(regs_307_io_reset),
    .io_out(regs_307_io_out),
    .io_enable(regs_307_io_enable)
  );
  FringeFF regs_308 ( // @[RegFile.scala 66:20:@38723.4]
    .clock(regs_308_clock),
    .reset(regs_308_reset),
    .io_in(regs_308_io_in),
    .io_reset(regs_308_io_reset),
    .io_out(regs_308_io_out),
    .io_enable(regs_308_io_enable)
  );
  FringeFF regs_309 ( // @[RegFile.scala 66:20:@38737.4]
    .clock(regs_309_clock),
    .reset(regs_309_reset),
    .io_in(regs_309_io_in),
    .io_reset(regs_309_io_reset),
    .io_out(regs_309_io_out),
    .io_enable(regs_309_io_enable)
  );
  FringeFF regs_310 ( // @[RegFile.scala 66:20:@38751.4]
    .clock(regs_310_clock),
    .reset(regs_310_reset),
    .io_in(regs_310_io_in),
    .io_reset(regs_310_io_reset),
    .io_out(regs_310_io_out),
    .io_enable(regs_310_io_enable)
  );
  FringeFF regs_311 ( // @[RegFile.scala 66:20:@38765.4]
    .clock(regs_311_clock),
    .reset(regs_311_reset),
    .io_in(regs_311_io_in),
    .io_reset(regs_311_io_reset),
    .io_out(regs_311_io_out),
    .io_enable(regs_311_io_enable)
  );
  FringeFF regs_312 ( // @[RegFile.scala 66:20:@38779.4]
    .clock(regs_312_clock),
    .reset(regs_312_reset),
    .io_in(regs_312_io_in),
    .io_reset(regs_312_io_reset),
    .io_out(regs_312_io_out),
    .io_enable(regs_312_io_enable)
  );
  FringeFF regs_313 ( // @[RegFile.scala 66:20:@38793.4]
    .clock(regs_313_clock),
    .reset(regs_313_reset),
    .io_in(regs_313_io_in),
    .io_reset(regs_313_io_reset),
    .io_out(regs_313_io_out),
    .io_enable(regs_313_io_enable)
  );
  FringeFF regs_314 ( // @[RegFile.scala 66:20:@38807.4]
    .clock(regs_314_clock),
    .reset(regs_314_reset),
    .io_in(regs_314_io_in),
    .io_reset(regs_314_io_reset),
    .io_out(regs_314_io_out),
    .io_enable(regs_314_io_enable)
  );
  FringeFF regs_315 ( // @[RegFile.scala 66:20:@38821.4]
    .clock(regs_315_clock),
    .reset(regs_315_reset),
    .io_in(regs_315_io_in),
    .io_reset(regs_315_io_reset),
    .io_out(regs_315_io_out),
    .io_enable(regs_315_io_enable)
  );
  FringeFF regs_316 ( // @[RegFile.scala 66:20:@38835.4]
    .clock(regs_316_clock),
    .reset(regs_316_reset),
    .io_in(regs_316_io_in),
    .io_reset(regs_316_io_reset),
    .io_out(regs_316_io_out),
    .io_enable(regs_316_io_enable)
  );
  FringeFF regs_317 ( // @[RegFile.scala 66:20:@38849.4]
    .clock(regs_317_clock),
    .reset(regs_317_reset),
    .io_in(regs_317_io_in),
    .io_reset(regs_317_io_reset),
    .io_out(regs_317_io_out),
    .io_enable(regs_317_io_enable)
  );
  FringeFF regs_318 ( // @[RegFile.scala 66:20:@38863.4]
    .clock(regs_318_clock),
    .reset(regs_318_reset),
    .io_in(regs_318_io_in),
    .io_reset(regs_318_io_reset),
    .io_out(regs_318_io_out),
    .io_enable(regs_318_io_enable)
  );
  FringeFF regs_319 ( // @[RegFile.scala 66:20:@38877.4]
    .clock(regs_319_clock),
    .reset(regs_319_reset),
    .io_in(regs_319_io_in),
    .io_reset(regs_319_io_reset),
    .io_out(regs_319_io_out),
    .io_enable(regs_319_io_enable)
  );
  FringeFF regs_320 ( // @[RegFile.scala 66:20:@38891.4]
    .clock(regs_320_clock),
    .reset(regs_320_reset),
    .io_in(regs_320_io_in),
    .io_reset(regs_320_io_reset),
    .io_out(regs_320_io_out),
    .io_enable(regs_320_io_enable)
  );
  FringeFF regs_321 ( // @[RegFile.scala 66:20:@38905.4]
    .clock(regs_321_clock),
    .reset(regs_321_reset),
    .io_in(regs_321_io_in),
    .io_reset(regs_321_io_reset),
    .io_out(regs_321_io_out),
    .io_enable(regs_321_io_enable)
  );
  FringeFF regs_322 ( // @[RegFile.scala 66:20:@38919.4]
    .clock(regs_322_clock),
    .reset(regs_322_reset),
    .io_in(regs_322_io_in),
    .io_reset(regs_322_io_reset),
    .io_out(regs_322_io_out),
    .io_enable(regs_322_io_enable)
  );
  FringeFF regs_323 ( // @[RegFile.scala 66:20:@38933.4]
    .clock(regs_323_clock),
    .reset(regs_323_reset),
    .io_in(regs_323_io_in),
    .io_reset(regs_323_io_reset),
    .io_out(regs_323_io_out),
    .io_enable(regs_323_io_enable)
  );
  FringeFF regs_324 ( // @[RegFile.scala 66:20:@38947.4]
    .clock(regs_324_clock),
    .reset(regs_324_reset),
    .io_in(regs_324_io_in),
    .io_reset(regs_324_io_reset),
    .io_out(regs_324_io_out),
    .io_enable(regs_324_io_enable)
  );
  FringeFF regs_325 ( // @[RegFile.scala 66:20:@38961.4]
    .clock(regs_325_clock),
    .reset(regs_325_reset),
    .io_in(regs_325_io_in),
    .io_reset(regs_325_io_reset),
    .io_out(regs_325_io_out),
    .io_enable(regs_325_io_enable)
  );
  FringeFF regs_326 ( // @[RegFile.scala 66:20:@38975.4]
    .clock(regs_326_clock),
    .reset(regs_326_reset),
    .io_in(regs_326_io_in),
    .io_reset(regs_326_io_reset),
    .io_out(regs_326_io_out),
    .io_enable(regs_326_io_enable)
  );
  FringeFF regs_327 ( // @[RegFile.scala 66:20:@38989.4]
    .clock(regs_327_clock),
    .reset(regs_327_reset),
    .io_in(regs_327_io_in),
    .io_reset(regs_327_io_reset),
    .io_out(regs_327_io_out),
    .io_enable(regs_327_io_enable)
  );
  FringeFF regs_328 ( // @[RegFile.scala 66:20:@39003.4]
    .clock(regs_328_clock),
    .reset(regs_328_reset),
    .io_in(regs_328_io_in),
    .io_reset(regs_328_io_reset),
    .io_out(regs_328_io_out),
    .io_enable(regs_328_io_enable)
  );
  FringeFF regs_329 ( // @[RegFile.scala 66:20:@39017.4]
    .clock(regs_329_clock),
    .reset(regs_329_reset),
    .io_in(regs_329_io_in),
    .io_reset(regs_329_io_reset),
    .io_out(regs_329_io_out),
    .io_enable(regs_329_io_enable)
  );
  FringeFF regs_330 ( // @[RegFile.scala 66:20:@39031.4]
    .clock(regs_330_clock),
    .reset(regs_330_reset),
    .io_in(regs_330_io_in),
    .io_reset(regs_330_io_reset),
    .io_out(regs_330_io_out),
    .io_enable(regs_330_io_enable)
  );
  FringeFF regs_331 ( // @[RegFile.scala 66:20:@39045.4]
    .clock(regs_331_clock),
    .reset(regs_331_reset),
    .io_in(regs_331_io_in),
    .io_reset(regs_331_io_reset),
    .io_out(regs_331_io_out),
    .io_enable(regs_331_io_enable)
  );
  FringeFF regs_332 ( // @[RegFile.scala 66:20:@39059.4]
    .clock(regs_332_clock),
    .reset(regs_332_reset),
    .io_in(regs_332_io_in),
    .io_reset(regs_332_io_reset),
    .io_out(regs_332_io_out),
    .io_enable(regs_332_io_enable)
  );
  FringeFF regs_333 ( // @[RegFile.scala 66:20:@39073.4]
    .clock(regs_333_clock),
    .reset(regs_333_reset),
    .io_in(regs_333_io_in),
    .io_reset(regs_333_io_reset),
    .io_out(regs_333_io_out),
    .io_enable(regs_333_io_enable)
  );
  FringeFF regs_334 ( // @[RegFile.scala 66:20:@39087.4]
    .clock(regs_334_clock),
    .reset(regs_334_reset),
    .io_in(regs_334_io_in),
    .io_reset(regs_334_io_reset),
    .io_out(regs_334_io_out),
    .io_enable(regs_334_io_enable)
  );
  FringeFF regs_335 ( // @[RegFile.scala 66:20:@39101.4]
    .clock(regs_335_clock),
    .reset(regs_335_reset),
    .io_in(regs_335_io_in),
    .io_reset(regs_335_io_reset),
    .io_out(regs_335_io_out),
    .io_enable(regs_335_io_enable)
  );
  FringeFF regs_336 ( // @[RegFile.scala 66:20:@39115.4]
    .clock(regs_336_clock),
    .reset(regs_336_reset),
    .io_in(regs_336_io_in),
    .io_reset(regs_336_io_reset),
    .io_out(regs_336_io_out),
    .io_enable(regs_336_io_enable)
  );
  FringeFF regs_337 ( // @[RegFile.scala 66:20:@39129.4]
    .clock(regs_337_clock),
    .reset(regs_337_reset),
    .io_in(regs_337_io_in),
    .io_reset(regs_337_io_reset),
    .io_out(regs_337_io_out),
    .io_enable(regs_337_io_enable)
  );
  FringeFF regs_338 ( // @[RegFile.scala 66:20:@39143.4]
    .clock(regs_338_clock),
    .reset(regs_338_reset),
    .io_in(regs_338_io_in),
    .io_reset(regs_338_io_reset),
    .io_out(regs_338_io_out),
    .io_enable(regs_338_io_enable)
  );
  FringeFF regs_339 ( // @[RegFile.scala 66:20:@39157.4]
    .clock(regs_339_clock),
    .reset(regs_339_reset),
    .io_in(regs_339_io_in),
    .io_reset(regs_339_io_reset),
    .io_out(regs_339_io_out),
    .io_enable(regs_339_io_enable)
  );
  FringeFF regs_340 ( // @[RegFile.scala 66:20:@39171.4]
    .clock(regs_340_clock),
    .reset(regs_340_reset),
    .io_in(regs_340_io_in),
    .io_reset(regs_340_io_reset),
    .io_out(regs_340_io_out),
    .io_enable(regs_340_io_enable)
  );
  FringeFF regs_341 ( // @[RegFile.scala 66:20:@39185.4]
    .clock(regs_341_clock),
    .reset(regs_341_reset),
    .io_in(regs_341_io_in),
    .io_reset(regs_341_io_reset),
    .io_out(regs_341_io_out),
    .io_enable(regs_341_io_enable)
  );
  FringeFF regs_342 ( // @[RegFile.scala 66:20:@39199.4]
    .clock(regs_342_clock),
    .reset(regs_342_reset),
    .io_in(regs_342_io_in),
    .io_reset(regs_342_io_reset),
    .io_out(regs_342_io_out),
    .io_enable(regs_342_io_enable)
  );
  FringeFF regs_343 ( // @[RegFile.scala 66:20:@39213.4]
    .clock(regs_343_clock),
    .reset(regs_343_reset),
    .io_in(regs_343_io_in),
    .io_reset(regs_343_io_reset),
    .io_out(regs_343_io_out),
    .io_enable(regs_343_io_enable)
  );
  FringeFF regs_344 ( // @[RegFile.scala 66:20:@39227.4]
    .clock(regs_344_clock),
    .reset(regs_344_reset),
    .io_in(regs_344_io_in),
    .io_reset(regs_344_io_reset),
    .io_out(regs_344_io_out),
    .io_enable(regs_344_io_enable)
  );
  FringeFF regs_345 ( // @[RegFile.scala 66:20:@39241.4]
    .clock(regs_345_clock),
    .reset(regs_345_reset),
    .io_in(regs_345_io_in),
    .io_reset(regs_345_io_reset),
    .io_out(regs_345_io_out),
    .io_enable(regs_345_io_enable)
  );
  FringeFF regs_346 ( // @[RegFile.scala 66:20:@39255.4]
    .clock(regs_346_clock),
    .reset(regs_346_reset),
    .io_in(regs_346_io_in),
    .io_reset(regs_346_io_reset),
    .io_out(regs_346_io_out),
    .io_enable(regs_346_io_enable)
  );
  FringeFF regs_347 ( // @[RegFile.scala 66:20:@39269.4]
    .clock(regs_347_clock),
    .reset(regs_347_reset),
    .io_in(regs_347_io_in),
    .io_reset(regs_347_io_reset),
    .io_out(regs_347_io_out),
    .io_enable(regs_347_io_enable)
  );
  FringeFF regs_348 ( // @[RegFile.scala 66:20:@39283.4]
    .clock(regs_348_clock),
    .reset(regs_348_reset),
    .io_in(regs_348_io_in),
    .io_reset(regs_348_io_reset),
    .io_out(regs_348_io_out),
    .io_enable(regs_348_io_enable)
  );
  FringeFF regs_349 ( // @[RegFile.scala 66:20:@39297.4]
    .clock(regs_349_clock),
    .reset(regs_349_reset),
    .io_in(regs_349_io_in),
    .io_reset(regs_349_io_reset),
    .io_out(regs_349_io_out),
    .io_enable(regs_349_io_enable)
  );
  FringeFF regs_350 ( // @[RegFile.scala 66:20:@39311.4]
    .clock(regs_350_clock),
    .reset(regs_350_reset),
    .io_in(regs_350_io_in),
    .io_reset(regs_350_io_reset),
    .io_out(regs_350_io_out),
    .io_enable(regs_350_io_enable)
  );
  FringeFF regs_351 ( // @[RegFile.scala 66:20:@39325.4]
    .clock(regs_351_clock),
    .reset(regs_351_reset),
    .io_in(regs_351_io_in),
    .io_reset(regs_351_io_reset),
    .io_out(regs_351_io_out),
    .io_enable(regs_351_io_enable)
  );
  FringeFF regs_352 ( // @[RegFile.scala 66:20:@39339.4]
    .clock(regs_352_clock),
    .reset(regs_352_reset),
    .io_in(regs_352_io_in),
    .io_reset(regs_352_io_reset),
    .io_out(regs_352_io_out),
    .io_enable(regs_352_io_enable)
  );
  FringeFF regs_353 ( // @[RegFile.scala 66:20:@39353.4]
    .clock(regs_353_clock),
    .reset(regs_353_reset),
    .io_in(regs_353_io_in),
    .io_reset(regs_353_io_reset),
    .io_out(regs_353_io_out),
    .io_enable(regs_353_io_enable)
  );
  FringeFF regs_354 ( // @[RegFile.scala 66:20:@39367.4]
    .clock(regs_354_clock),
    .reset(regs_354_reset),
    .io_in(regs_354_io_in),
    .io_reset(regs_354_io_reset),
    .io_out(regs_354_io_out),
    .io_enable(regs_354_io_enable)
  );
  FringeFF regs_355 ( // @[RegFile.scala 66:20:@39381.4]
    .clock(regs_355_clock),
    .reset(regs_355_reset),
    .io_in(regs_355_io_in),
    .io_reset(regs_355_io_reset),
    .io_out(regs_355_io_out),
    .io_enable(regs_355_io_enable)
  );
  FringeFF regs_356 ( // @[RegFile.scala 66:20:@39395.4]
    .clock(regs_356_clock),
    .reset(regs_356_reset),
    .io_in(regs_356_io_in),
    .io_reset(regs_356_io_reset),
    .io_out(regs_356_io_out),
    .io_enable(regs_356_io_enable)
  );
  FringeFF regs_357 ( // @[RegFile.scala 66:20:@39409.4]
    .clock(regs_357_clock),
    .reset(regs_357_reset),
    .io_in(regs_357_io_in),
    .io_reset(regs_357_io_reset),
    .io_out(regs_357_io_out),
    .io_enable(regs_357_io_enable)
  );
  FringeFF regs_358 ( // @[RegFile.scala 66:20:@39423.4]
    .clock(regs_358_clock),
    .reset(regs_358_reset),
    .io_in(regs_358_io_in),
    .io_reset(regs_358_io_reset),
    .io_out(regs_358_io_out),
    .io_enable(regs_358_io_enable)
  );
  FringeFF regs_359 ( // @[RegFile.scala 66:20:@39437.4]
    .clock(regs_359_clock),
    .reset(regs_359_reset),
    .io_in(regs_359_io_in),
    .io_reset(regs_359_io_reset),
    .io_out(regs_359_io_out),
    .io_enable(regs_359_io_enable)
  );
  FringeFF regs_360 ( // @[RegFile.scala 66:20:@39451.4]
    .clock(regs_360_clock),
    .reset(regs_360_reset),
    .io_in(regs_360_io_in),
    .io_reset(regs_360_io_reset),
    .io_out(regs_360_io_out),
    .io_enable(regs_360_io_enable)
  );
  FringeFF regs_361 ( // @[RegFile.scala 66:20:@39465.4]
    .clock(regs_361_clock),
    .reset(regs_361_reset),
    .io_in(regs_361_io_in),
    .io_reset(regs_361_io_reset),
    .io_out(regs_361_io_out),
    .io_enable(regs_361_io_enable)
  );
  FringeFF regs_362 ( // @[RegFile.scala 66:20:@39479.4]
    .clock(regs_362_clock),
    .reset(regs_362_reset),
    .io_in(regs_362_io_in),
    .io_reset(regs_362_io_reset),
    .io_out(regs_362_io_out),
    .io_enable(regs_362_io_enable)
  );
  FringeFF regs_363 ( // @[RegFile.scala 66:20:@39493.4]
    .clock(regs_363_clock),
    .reset(regs_363_reset),
    .io_in(regs_363_io_in),
    .io_reset(regs_363_io_reset),
    .io_out(regs_363_io_out),
    .io_enable(regs_363_io_enable)
  );
  FringeFF regs_364 ( // @[RegFile.scala 66:20:@39507.4]
    .clock(regs_364_clock),
    .reset(regs_364_reset),
    .io_in(regs_364_io_in),
    .io_reset(regs_364_io_reset),
    .io_out(regs_364_io_out),
    .io_enable(regs_364_io_enable)
  );
  FringeFF regs_365 ( // @[RegFile.scala 66:20:@39521.4]
    .clock(regs_365_clock),
    .reset(regs_365_reset),
    .io_in(regs_365_io_in),
    .io_reset(regs_365_io_reset),
    .io_out(regs_365_io_out),
    .io_enable(regs_365_io_enable)
  );
  FringeFF regs_366 ( // @[RegFile.scala 66:20:@39535.4]
    .clock(regs_366_clock),
    .reset(regs_366_reset),
    .io_in(regs_366_io_in),
    .io_reset(regs_366_io_reset),
    .io_out(regs_366_io_out),
    .io_enable(regs_366_io_enable)
  );
  FringeFF regs_367 ( // @[RegFile.scala 66:20:@39549.4]
    .clock(regs_367_clock),
    .reset(regs_367_reset),
    .io_in(regs_367_io_in),
    .io_reset(regs_367_io_reset),
    .io_out(regs_367_io_out),
    .io_enable(regs_367_io_enable)
  );
  FringeFF regs_368 ( // @[RegFile.scala 66:20:@39563.4]
    .clock(regs_368_clock),
    .reset(regs_368_reset),
    .io_in(regs_368_io_in),
    .io_reset(regs_368_io_reset),
    .io_out(regs_368_io_out),
    .io_enable(regs_368_io_enable)
  );
  FringeFF regs_369 ( // @[RegFile.scala 66:20:@39577.4]
    .clock(regs_369_clock),
    .reset(regs_369_reset),
    .io_in(regs_369_io_in),
    .io_reset(regs_369_io_reset),
    .io_out(regs_369_io_out),
    .io_enable(regs_369_io_enable)
  );
  FringeFF regs_370 ( // @[RegFile.scala 66:20:@39591.4]
    .clock(regs_370_clock),
    .reset(regs_370_reset),
    .io_in(regs_370_io_in),
    .io_reset(regs_370_io_reset),
    .io_out(regs_370_io_out),
    .io_enable(regs_370_io_enable)
  );
  FringeFF regs_371 ( // @[RegFile.scala 66:20:@39605.4]
    .clock(regs_371_clock),
    .reset(regs_371_reset),
    .io_in(regs_371_io_in),
    .io_reset(regs_371_io_reset),
    .io_out(regs_371_io_out),
    .io_enable(regs_371_io_enable)
  );
  FringeFF regs_372 ( // @[RegFile.scala 66:20:@39619.4]
    .clock(regs_372_clock),
    .reset(regs_372_reset),
    .io_in(regs_372_io_in),
    .io_reset(regs_372_io_reset),
    .io_out(regs_372_io_out),
    .io_enable(regs_372_io_enable)
  );
  FringeFF regs_373 ( // @[RegFile.scala 66:20:@39633.4]
    .clock(regs_373_clock),
    .reset(regs_373_reset),
    .io_in(regs_373_io_in),
    .io_reset(regs_373_io_reset),
    .io_out(regs_373_io_out),
    .io_enable(regs_373_io_enable)
  );
  FringeFF regs_374 ( // @[RegFile.scala 66:20:@39647.4]
    .clock(regs_374_clock),
    .reset(regs_374_reset),
    .io_in(regs_374_io_in),
    .io_reset(regs_374_io_reset),
    .io_out(regs_374_io_out),
    .io_enable(regs_374_io_enable)
  );
  FringeFF regs_375 ( // @[RegFile.scala 66:20:@39661.4]
    .clock(regs_375_clock),
    .reset(regs_375_reset),
    .io_in(regs_375_io_in),
    .io_reset(regs_375_io_reset),
    .io_out(regs_375_io_out),
    .io_enable(regs_375_io_enable)
  );
  FringeFF regs_376 ( // @[RegFile.scala 66:20:@39675.4]
    .clock(regs_376_clock),
    .reset(regs_376_reset),
    .io_in(regs_376_io_in),
    .io_reset(regs_376_io_reset),
    .io_out(regs_376_io_out),
    .io_enable(regs_376_io_enable)
  );
  FringeFF regs_377 ( // @[RegFile.scala 66:20:@39689.4]
    .clock(regs_377_clock),
    .reset(regs_377_reset),
    .io_in(regs_377_io_in),
    .io_reset(regs_377_io_reset),
    .io_out(regs_377_io_out),
    .io_enable(regs_377_io_enable)
  );
  FringeFF regs_378 ( // @[RegFile.scala 66:20:@39703.4]
    .clock(regs_378_clock),
    .reset(regs_378_reset),
    .io_in(regs_378_io_in),
    .io_reset(regs_378_io_reset),
    .io_out(regs_378_io_out),
    .io_enable(regs_378_io_enable)
  );
  FringeFF regs_379 ( // @[RegFile.scala 66:20:@39717.4]
    .clock(regs_379_clock),
    .reset(regs_379_reset),
    .io_in(regs_379_io_in),
    .io_reset(regs_379_io_reset),
    .io_out(regs_379_io_out),
    .io_enable(regs_379_io_enable)
  );
  FringeFF regs_380 ( // @[RegFile.scala 66:20:@39731.4]
    .clock(regs_380_clock),
    .reset(regs_380_reset),
    .io_in(regs_380_io_in),
    .io_reset(regs_380_io_reset),
    .io_out(regs_380_io_out),
    .io_enable(regs_380_io_enable)
  );
  FringeFF regs_381 ( // @[RegFile.scala 66:20:@39745.4]
    .clock(regs_381_clock),
    .reset(regs_381_reset),
    .io_in(regs_381_io_in),
    .io_reset(regs_381_io_reset),
    .io_out(regs_381_io_out),
    .io_enable(regs_381_io_enable)
  );
  FringeFF regs_382 ( // @[RegFile.scala 66:20:@39759.4]
    .clock(regs_382_clock),
    .reset(regs_382_reset),
    .io_in(regs_382_io_in),
    .io_reset(regs_382_io_reset),
    .io_out(regs_382_io_out),
    .io_enable(regs_382_io_enable)
  );
  FringeFF regs_383 ( // @[RegFile.scala 66:20:@39773.4]
    .clock(regs_383_clock),
    .reset(regs_383_reset),
    .io_in(regs_383_io_in),
    .io_reset(regs_383_io_reset),
    .io_out(regs_383_io_out),
    .io_enable(regs_383_io_enable)
  );
  FringeFF regs_384 ( // @[RegFile.scala 66:20:@39787.4]
    .clock(regs_384_clock),
    .reset(regs_384_reset),
    .io_in(regs_384_io_in),
    .io_reset(regs_384_io_reset),
    .io_out(regs_384_io_out),
    .io_enable(regs_384_io_enable)
  );
  FringeFF regs_385 ( // @[RegFile.scala 66:20:@39801.4]
    .clock(regs_385_clock),
    .reset(regs_385_reset),
    .io_in(regs_385_io_in),
    .io_reset(regs_385_io_reset),
    .io_out(regs_385_io_out),
    .io_enable(regs_385_io_enable)
  );
  FringeFF regs_386 ( // @[RegFile.scala 66:20:@39815.4]
    .clock(regs_386_clock),
    .reset(regs_386_reset),
    .io_in(regs_386_io_in),
    .io_reset(regs_386_io_reset),
    .io_out(regs_386_io_out),
    .io_enable(regs_386_io_enable)
  );
  FringeFF regs_387 ( // @[RegFile.scala 66:20:@39829.4]
    .clock(regs_387_clock),
    .reset(regs_387_reset),
    .io_in(regs_387_io_in),
    .io_reset(regs_387_io_reset),
    .io_out(regs_387_io_out),
    .io_enable(regs_387_io_enable)
  );
  FringeFF regs_388 ( // @[RegFile.scala 66:20:@39843.4]
    .clock(regs_388_clock),
    .reset(regs_388_reset),
    .io_in(regs_388_io_in),
    .io_reset(regs_388_io_reset),
    .io_out(regs_388_io_out),
    .io_enable(regs_388_io_enable)
  );
  FringeFF regs_389 ( // @[RegFile.scala 66:20:@39857.4]
    .clock(regs_389_clock),
    .reset(regs_389_reset),
    .io_in(regs_389_io_in),
    .io_reset(regs_389_io_reset),
    .io_out(regs_389_io_out),
    .io_enable(regs_389_io_enable)
  );
  FringeFF regs_390 ( // @[RegFile.scala 66:20:@39871.4]
    .clock(regs_390_clock),
    .reset(regs_390_reset),
    .io_in(regs_390_io_in),
    .io_reset(regs_390_io_reset),
    .io_out(regs_390_io_out),
    .io_enable(regs_390_io_enable)
  );
  FringeFF regs_391 ( // @[RegFile.scala 66:20:@39885.4]
    .clock(regs_391_clock),
    .reset(regs_391_reset),
    .io_in(regs_391_io_in),
    .io_reset(regs_391_io_reset),
    .io_out(regs_391_io_out),
    .io_enable(regs_391_io_enable)
  );
  FringeFF regs_392 ( // @[RegFile.scala 66:20:@39899.4]
    .clock(regs_392_clock),
    .reset(regs_392_reset),
    .io_in(regs_392_io_in),
    .io_reset(regs_392_io_reset),
    .io_out(regs_392_io_out),
    .io_enable(regs_392_io_enable)
  );
  FringeFF regs_393 ( // @[RegFile.scala 66:20:@39913.4]
    .clock(regs_393_clock),
    .reset(regs_393_reset),
    .io_in(regs_393_io_in),
    .io_reset(regs_393_io_reset),
    .io_out(regs_393_io_out),
    .io_enable(regs_393_io_enable)
  );
  FringeFF regs_394 ( // @[RegFile.scala 66:20:@39927.4]
    .clock(regs_394_clock),
    .reset(regs_394_reset),
    .io_in(regs_394_io_in),
    .io_reset(regs_394_io_reset),
    .io_out(regs_394_io_out),
    .io_enable(regs_394_io_enable)
  );
  FringeFF regs_395 ( // @[RegFile.scala 66:20:@39941.4]
    .clock(regs_395_clock),
    .reset(regs_395_reset),
    .io_in(regs_395_io_in),
    .io_reset(regs_395_io_reset),
    .io_out(regs_395_io_out),
    .io_enable(regs_395_io_enable)
  );
  FringeFF regs_396 ( // @[RegFile.scala 66:20:@39955.4]
    .clock(regs_396_clock),
    .reset(regs_396_reset),
    .io_in(regs_396_io_in),
    .io_reset(regs_396_io_reset),
    .io_out(regs_396_io_out),
    .io_enable(regs_396_io_enable)
  );
  FringeFF regs_397 ( // @[RegFile.scala 66:20:@39969.4]
    .clock(regs_397_clock),
    .reset(regs_397_reset),
    .io_in(regs_397_io_in),
    .io_reset(regs_397_io_reset),
    .io_out(regs_397_io_out),
    .io_enable(regs_397_io_enable)
  );
  FringeFF regs_398 ( // @[RegFile.scala 66:20:@39983.4]
    .clock(regs_398_clock),
    .reset(regs_398_reset),
    .io_in(regs_398_io_in),
    .io_reset(regs_398_io_reset),
    .io_out(regs_398_io_out),
    .io_enable(regs_398_io_enable)
  );
  FringeFF regs_399 ( // @[RegFile.scala 66:20:@39997.4]
    .clock(regs_399_clock),
    .reset(regs_399_reset),
    .io_in(regs_399_io_in),
    .io_reset(regs_399_io_reset),
    .io_out(regs_399_io_out),
    .io_enable(regs_399_io_enable)
  );
  FringeFF regs_400 ( // @[RegFile.scala 66:20:@40011.4]
    .clock(regs_400_clock),
    .reset(regs_400_reset),
    .io_in(regs_400_io_in),
    .io_reset(regs_400_io_reset),
    .io_out(regs_400_io_out),
    .io_enable(regs_400_io_enable)
  );
  FringeFF regs_401 ( // @[RegFile.scala 66:20:@40025.4]
    .clock(regs_401_clock),
    .reset(regs_401_reset),
    .io_in(regs_401_io_in),
    .io_reset(regs_401_io_reset),
    .io_out(regs_401_io_out),
    .io_enable(regs_401_io_enable)
  );
  FringeFF regs_402 ( // @[RegFile.scala 66:20:@40039.4]
    .clock(regs_402_clock),
    .reset(regs_402_reset),
    .io_in(regs_402_io_in),
    .io_reset(regs_402_io_reset),
    .io_out(regs_402_io_out),
    .io_enable(regs_402_io_enable)
  );
  FringeFF regs_403 ( // @[RegFile.scala 66:20:@40053.4]
    .clock(regs_403_clock),
    .reset(regs_403_reset),
    .io_in(regs_403_io_in),
    .io_reset(regs_403_io_reset),
    .io_out(regs_403_io_out),
    .io_enable(regs_403_io_enable)
  );
  FringeFF regs_404 ( // @[RegFile.scala 66:20:@40067.4]
    .clock(regs_404_clock),
    .reset(regs_404_reset),
    .io_in(regs_404_io_in),
    .io_reset(regs_404_io_reset),
    .io_out(regs_404_io_out),
    .io_enable(regs_404_io_enable)
  );
  FringeFF regs_405 ( // @[RegFile.scala 66:20:@40081.4]
    .clock(regs_405_clock),
    .reset(regs_405_reset),
    .io_in(regs_405_io_in),
    .io_reset(regs_405_io_reset),
    .io_out(regs_405_io_out),
    .io_enable(regs_405_io_enable)
  );
  FringeFF regs_406 ( // @[RegFile.scala 66:20:@40095.4]
    .clock(regs_406_clock),
    .reset(regs_406_reset),
    .io_in(regs_406_io_in),
    .io_reset(regs_406_io_reset),
    .io_out(regs_406_io_out),
    .io_enable(regs_406_io_enable)
  );
  FringeFF regs_407 ( // @[RegFile.scala 66:20:@40109.4]
    .clock(regs_407_clock),
    .reset(regs_407_reset),
    .io_in(regs_407_io_in),
    .io_reset(regs_407_io_reset),
    .io_out(regs_407_io_out),
    .io_enable(regs_407_io_enable)
  );
  FringeFF regs_408 ( // @[RegFile.scala 66:20:@40123.4]
    .clock(regs_408_clock),
    .reset(regs_408_reset),
    .io_in(regs_408_io_in),
    .io_reset(regs_408_io_reset),
    .io_out(regs_408_io_out),
    .io_enable(regs_408_io_enable)
  );
  FringeFF regs_409 ( // @[RegFile.scala 66:20:@40137.4]
    .clock(regs_409_clock),
    .reset(regs_409_reset),
    .io_in(regs_409_io_in),
    .io_reset(regs_409_io_reset),
    .io_out(regs_409_io_out),
    .io_enable(regs_409_io_enable)
  );
  FringeFF regs_410 ( // @[RegFile.scala 66:20:@40151.4]
    .clock(regs_410_clock),
    .reset(regs_410_reset),
    .io_in(regs_410_io_in),
    .io_reset(regs_410_io_reset),
    .io_out(regs_410_io_out),
    .io_enable(regs_410_io_enable)
  );
  FringeFF regs_411 ( // @[RegFile.scala 66:20:@40165.4]
    .clock(regs_411_clock),
    .reset(regs_411_reset),
    .io_in(regs_411_io_in),
    .io_reset(regs_411_io_reset),
    .io_out(regs_411_io_out),
    .io_enable(regs_411_io_enable)
  );
  FringeFF regs_412 ( // @[RegFile.scala 66:20:@40179.4]
    .clock(regs_412_clock),
    .reset(regs_412_reset),
    .io_in(regs_412_io_in),
    .io_reset(regs_412_io_reset),
    .io_out(regs_412_io_out),
    .io_enable(regs_412_io_enable)
  );
  FringeFF regs_413 ( // @[RegFile.scala 66:20:@40193.4]
    .clock(regs_413_clock),
    .reset(regs_413_reset),
    .io_in(regs_413_io_in),
    .io_reset(regs_413_io_reset),
    .io_out(regs_413_io_out),
    .io_enable(regs_413_io_enable)
  );
  FringeFF regs_414 ( // @[RegFile.scala 66:20:@40207.4]
    .clock(regs_414_clock),
    .reset(regs_414_reset),
    .io_in(regs_414_io_in),
    .io_reset(regs_414_io_reset),
    .io_out(regs_414_io_out),
    .io_enable(regs_414_io_enable)
  );
  FringeFF regs_415 ( // @[RegFile.scala 66:20:@40221.4]
    .clock(regs_415_clock),
    .reset(regs_415_reset),
    .io_in(regs_415_io_in),
    .io_reset(regs_415_io_reset),
    .io_out(regs_415_io_out),
    .io_enable(regs_415_io_enable)
  );
  FringeFF regs_416 ( // @[RegFile.scala 66:20:@40235.4]
    .clock(regs_416_clock),
    .reset(regs_416_reset),
    .io_in(regs_416_io_in),
    .io_reset(regs_416_io_reset),
    .io_out(regs_416_io_out),
    .io_enable(regs_416_io_enable)
  );
  FringeFF regs_417 ( // @[RegFile.scala 66:20:@40249.4]
    .clock(regs_417_clock),
    .reset(regs_417_reset),
    .io_in(regs_417_io_in),
    .io_reset(regs_417_io_reset),
    .io_out(regs_417_io_out),
    .io_enable(regs_417_io_enable)
  );
  FringeFF regs_418 ( // @[RegFile.scala 66:20:@40263.4]
    .clock(regs_418_clock),
    .reset(regs_418_reset),
    .io_in(regs_418_io_in),
    .io_reset(regs_418_io_reset),
    .io_out(regs_418_io_out),
    .io_enable(regs_418_io_enable)
  );
  FringeFF regs_419 ( // @[RegFile.scala 66:20:@40277.4]
    .clock(regs_419_clock),
    .reset(regs_419_reset),
    .io_in(regs_419_io_in),
    .io_reset(regs_419_io_reset),
    .io_out(regs_419_io_out),
    .io_enable(regs_419_io_enable)
  );
  FringeFF regs_420 ( // @[RegFile.scala 66:20:@40291.4]
    .clock(regs_420_clock),
    .reset(regs_420_reset),
    .io_in(regs_420_io_in),
    .io_reset(regs_420_io_reset),
    .io_out(regs_420_io_out),
    .io_enable(regs_420_io_enable)
  );
  FringeFF regs_421 ( // @[RegFile.scala 66:20:@40305.4]
    .clock(regs_421_clock),
    .reset(regs_421_reset),
    .io_in(regs_421_io_in),
    .io_reset(regs_421_io_reset),
    .io_out(regs_421_io_out),
    .io_enable(regs_421_io_enable)
  );
  FringeFF regs_422 ( // @[RegFile.scala 66:20:@40319.4]
    .clock(regs_422_clock),
    .reset(regs_422_reset),
    .io_in(regs_422_io_in),
    .io_reset(regs_422_io_reset),
    .io_out(regs_422_io_out),
    .io_enable(regs_422_io_enable)
  );
  FringeFF regs_423 ( // @[RegFile.scala 66:20:@40333.4]
    .clock(regs_423_clock),
    .reset(regs_423_reset),
    .io_in(regs_423_io_in),
    .io_reset(regs_423_io_reset),
    .io_out(regs_423_io_out),
    .io_enable(regs_423_io_enable)
  );
  FringeFF regs_424 ( // @[RegFile.scala 66:20:@40347.4]
    .clock(regs_424_clock),
    .reset(regs_424_reset),
    .io_in(regs_424_io_in),
    .io_reset(regs_424_io_reset),
    .io_out(regs_424_io_out),
    .io_enable(regs_424_io_enable)
  );
  FringeFF regs_425 ( // @[RegFile.scala 66:20:@40361.4]
    .clock(regs_425_clock),
    .reset(regs_425_reset),
    .io_in(regs_425_io_in),
    .io_reset(regs_425_io_reset),
    .io_out(regs_425_io_out),
    .io_enable(regs_425_io_enable)
  );
  FringeFF regs_426 ( // @[RegFile.scala 66:20:@40375.4]
    .clock(regs_426_clock),
    .reset(regs_426_reset),
    .io_in(regs_426_io_in),
    .io_reset(regs_426_io_reset),
    .io_out(regs_426_io_out),
    .io_enable(regs_426_io_enable)
  );
  FringeFF regs_427 ( // @[RegFile.scala 66:20:@40389.4]
    .clock(regs_427_clock),
    .reset(regs_427_reset),
    .io_in(regs_427_io_in),
    .io_reset(regs_427_io_reset),
    .io_out(regs_427_io_out),
    .io_enable(regs_427_io_enable)
  );
  FringeFF regs_428 ( // @[RegFile.scala 66:20:@40403.4]
    .clock(regs_428_clock),
    .reset(regs_428_reset),
    .io_in(regs_428_io_in),
    .io_reset(regs_428_io_reset),
    .io_out(regs_428_io_out),
    .io_enable(regs_428_io_enable)
  );
  FringeFF regs_429 ( // @[RegFile.scala 66:20:@40417.4]
    .clock(regs_429_clock),
    .reset(regs_429_reset),
    .io_in(regs_429_io_in),
    .io_reset(regs_429_io_reset),
    .io_out(regs_429_io_out),
    .io_enable(regs_429_io_enable)
  );
  FringeFF regs_430 ( // @[RegFile.scala 66:20:@40431.4]
    .clock(regs_430_clock),
    .reset(regs_430_reset),
    .io_in(regs_430_io_in),
    .io_reset(regs_430_io_reset),
    .io_out(regs_430_io_out),
    .io_enable(regs_430_io_enable)
  );
  FringeFF regs_431 ( // @[RegFile.scala 66:20:@40445.4]
    .clock(regs_431_clock),
    .reset(regs_431_reset),
    .io_in(regs_431_io_in),
    .io_reset(regs_431_io_reset),
    .io_out(regs_431_io_out),
    .io_enable(regs_431_io_enable)
  );
  FringeFF regs_432 ( // @[RegFile.scala 66:20:@40459.4]
    .clock(regs_432_clock),
    .reset(regs_432_reset),
    .io_in(regs_432_io_in),
    .io_reset(regs_432_io_reset),
    .io_out(regs_432_io_out),
    .io_enable(regs_432_io_enable)
  );
  FringeFF regs_433 ( // @[RegFile.scala 66:20:@40473.4]
    .clock(regs_433_clock),
    .reset(regs_433_reset),
    .io_in(regs_433_io_in),
    .io_reset(regs_433_io_reset),
    .io_out(regs_433_io_out),
    .io_enable(regs_433_io_enable)
  );
  FringeFF regs_434 ( // @[RegFile.scala 66:20:@40487.4]
    .clock(regs_434_clock),
    .reset(regs_434_reset),
    .io_in(regs_434_io_in),
    .io_reset(regs_434_io_reset),
    .io_out(regs_434_io_out),
    .io_enable(regs_434_io_enable)
  );
  FringeFF regs_435 ( // @[RegFile.scala 66:20:@40501.4]
    .clock(regs_435_clock),
    .reset(regs_435_reset),
    .io_in(regs_435_io_in),
    .io_reset(regs_435_io_reset),
    .io_out(regs_435_io_out),
    .io_enable(regs_435_io_enable)
  );
  FringeFF regs_436 ( // @[RegFile.scala 66:20:@40515.4]
    .clock(regs_436_clock),
    .reset(regs_436_reset),
    .io_in(regs_436_io_in),
    .io_reset(regs_436_io_reset),
    .io_out(regs_436_io_out),
    .io_enable(regs_436_io_enable)
  );
  FringeFF regs_437 ( // @[RegFile.scala 66:20:@40529.4]
    .clock(regs_437_clock),
    .reset(regs_437_reset),
    .io_in(regs_437_io_in),
    .io_reset(regs_437_io_reset),
    .io_out(regs_437_io_out),
    .io_enable(regs_437_io_enable)
  );
  FringeFF regs_438 ( // @[RegFile.scala 66:20:@40543.4]
    .clock(regs_438_clock),
    .reset(regs_438_reset),
    .io_in(regs_438_io_in),
    .io_reset(regs_438_io_reset),
    .io_out(regs_438_io_out),
    .io_enable(regs_438_io_enable)
  );
  FringeFF regs_439 ( // @[RegFile.scala 66:20:@40557.4]
    .clock(regs_439_clock),
    .reset(regs_439_reset),
    .io_in(regs_439_io_in),
    .io_reset(regs_439_io_reset),
    .io_out(regs_439_io_out),
    .io_enable(regs_439_io_enable)
  );
  FringeFF regs_440 ( // @[RegFile.scala 66:20:@40571.4]
    .clock(regs_440_clock),
    .reset(regs_440_reset),
    .io_in(regs_440_io_in),
    .io_reset(regs_440_io_reset),
    .io_out(regs_440_io_out),
    .io_enable(regs_440_io_enable)
  );
  FringeFF regs_441 ( // @[RegFile.scala 66:20:@40585.4]
    .clock(regs_441_clock),
    .reset(regs_441_reset),
    .io_in(regs_441_io_in),
    .io_reset(regs_441_io_reset),
    .io_out(regs_441_io_out),
    .io_enable(regs_441_io_enable)
  );
  FringeFF regs_442 ( // @[RegFile.scala 66:20:@40599.4]
    .clock(regs_442_clock),
    .reset(regs_442_reset),
    .io_in(regs_442_io_in),
    .io_reset(regs_442_io_reset),
    .io_out(regs_442_io_out),
    .io_enable(regs_442_io_enable)
  );
  FringeFF regs_443 ( // @[RegFile.scala 66:20:@40613.4]
    .clock(regs_443_clock),
    .reset(regs_443_reset),
    .io_in(regs_443_io_in),
    .io_reset(regs_443_io_reset),
    .io_out(regs_443_io_out),
    .io_enable(regs_443_io_enable)
  );
  FringeFF regs_444 ( // @[RegFile.scala 66:20:@40627.4]
    .clock(regs_444_clock),
    .reset(regs_444_reset),
    .io_in(regs_444_io_in),
    .io_reset(regs_444_io_reset),
    .io_out(regs_444_io_out),
    .io_enable(regs_444_io_enable)
  );
  FringeFF regs_445 ( // @[RegFile.scala 66:20:@40641.4]
    .clock(regs_445_clock),
    .reset(regs_445_reset),
    .io_in(regs_445_io_in),
    .io_reset(regs_445_io_reset),
    .io_out(regs_445_io_out),
    .io_enable(regs_445_io_enable)
  );
  FringeFF regs_446 ( // @[RegFile.scala 66:20:@40655.4]
    .clock(regs_446_clock),
    .reset(regs_446_reset),
    .io_in(regs_446_io_in),
    .io_reset(regs_446_io_reset),
    .io_out(regs_446_io_out),
    .io_enable(regs_446_io_enable)
  );
  FringeFF regs_447 ( // @[RegFile.scala 66:20:@40669.4]
    .clock(regs_447_clock),
    .reset(regs_447_reset),
    .io_in(regs_447_io_in),
    .io_reset(regs_447_io_reset),
    .io_out(regs_447_io_out),
    .io_enable(regs_447_io_enable)
  );
  FringeFF regs_448 ( // @[RegFile.scala 66:20:@40683.4]
    .clock(regs_448_clock),
    .reset(regs_448_reset),
    .io_in(regs_448_io_in),
    .io_reset(regs_448_io_reset),
    .io_out(regs_448_io_out),
    .io_enable(regs_448_io_enable)
  );
  FringeFF regs_449 ( // @[RegFile.scala 66:20:@40697.4]
    .clock(regs_449_clock),
    .reset(regs_449_reset),
    .io_in(regs_449_io_in),
    .io_reset(regs_449_io_reset),
    .io_out(regs_449_io_out),
    .io_enable(regs_449_io_enable)
  );
  FringeFF regs_450 ( // @[RegFile.scala 66:20:@40711.4]
    .clock(regs_450_clock),
    .reset(regs_450_reset),
    .io_in(regs_450_io_in),
    .io_reset(regs_450_io_reset),
    .io_out(regs_450_io_out),
    .io_enable(regs_450_io_enable)
  );
  FringeFF regs_451 ( // @[RegFile.scala 66:20:@40725.4]
    .clock(regs_451_clock),
    .reset(regs_451_reset),
    .io_in(regs_451_io_in),
    .io_reset(regs_451_io_reset),
    .io_out(regs_451_io_out),
    .io_enable(regs_451_io_enable)
  );
  FringeFF regs_452 ( // @[RegFile.scala 66:20:@40739.4]
    .clock(regs_452_clock),
    .reset(regs_452_reset),
    .io_in(regs_452_io_in),
    .io_reset(regs_452_io_reset),
    .io_out(regs_452_io_out),
    .io_enable(regs_452_io_enable)
  );
  FringeFF regs_453 ( // @[RegFile.scala 66:20:@40753.4]
    .clock(regs_453_clock),
    .reset(regs_453_reset),
    .io_in(regs_453_io_in),
    .io_reset(regs_453_io_reset),
    .io_out(regs_453_io_out),
    .io_enable(regs_453_io_enable)
  );
  FringeFF regs_454 ( // @[RegFile.scala 66:20:@40767.4]
    .clock(regs_454_clock),
    .reset(regs_454_reset),
    .io_in(regs_454_io_in),
    .io_reset(regs_454_io_reset),
    .io_out(regs_454_io_out),
    .io_enable(regs_454_io_enable)
  );
  FringeFF regs_455 ( // @[RegFile.scala 66:20:@40781.4]
    .clock(regs_455_clock),
    .reset(regs_455_reset),
    .io_in(regs_455_io_in),
    .io_reset(regs_455_io_reset),
    .io_out(regs_455_io_out),
    .io_enable(regs_455_io_enable)
  );
  FringeFF regs_456 ( // @[RegFile.scala 66:20:@40795.4]
    .clock(regs_456_clock),
    .reset(regs_456_reset),
    .io_in(regs_456_io_in),
    .io_reset(regs_456_io_reset),
    .io_out(regs_456_io_out),
    .io_enable(regs_456_io_enable)
  );
  FringeFF regs_457 ( // @[RegFile.scala 66:20:@40809.4]
    .clock(regs_457_clock),
    .reset(regs_457_reset),
    .io_in(regs_457_io_in),
    .io_reset(regs_457_io_reset),
    .io_out(regs_457_io_out),
    .io_enable(regs_457_io_enable)
  );
  FringeFF regs_458 ( // @[RegFile.scala 66:20:@40823.4]
    .clock(regs_458_clock),
    .reset(regs_458_reset),
    .io_in(regs_458_io_in),
    .io_reset(regs_458_io_reset),
    .io_out(regs_458_io_out),
    .io_enable(regs_458_io_enable)
  );
  FringeFF regs_459 ( // @[RegFile.scala 66:20:@40837.4]
    .clock(regs_459_clock),
    .reset(regs_459_reset),
    .io_in(regs_459_io_in),
    .io_reset(regs_459_io_reset),
    .io_out(regs_459_io_out),
    .io_enable(regs_459_io_enable)
  );
  FringeFF regs_460 ( // @[RegFile.scala 66:20:@40851.4]
    .clock(regs_460_clock),
    .reset(regs_460_reset),
    .io_in(regs_460_io_in),
    .io_reset(regs_460_io_reset),
    .io_out(regs_460_io_out),
    .io_enable(regs_460_io_enable)
  );
  FringeFF regs_461 ( // @[RegFile.scala 66:20:@40865.4]
    .clock(regs_461_clock),
    .reset(regs_461_reset),
    .io_in(regs_461_io_in),
    .io_reset(regs_461_io_reset),
    .io_out(regs_461_io_out),
    .io_enable(regs_461_io_enable)
  );
  FringeFF regs_462 ( // @[RegFile.scala 66:20:@40879.4]
    .clock(regs_462_clock),
    .reset(regs_462_reset),
    .io_in(regs_462_io_in),
    .io_reset(regs_462_io_reset),
    .io_out(regs_462_io_out),
    .io_enable(regs_462_io_enable)
  );
  FringeFF regs_463 ( // @[RegFile.scala 66:20:@40893.4]
    .clock(regs_463_clock),
    .reset(regs_463_reset),
    .io_in(regs_463_io_in),
    .io_reset(regs_463_io_reset),
    .io_out(regs_463_io_out),
    .io_enable(regs_463_io_enable)
  );
  FringeFF regs_464 ( // @[RegFile.scala 66:20:@40907.4]
    .clock(regs_464_clock),
    .reset(regs_464_reset),
    .io_in(regs_464_io_in),
    .io_reset(regs_464_io_reset),
    .io_out(regs_464_io_out),
    .io_enable(regs_464_io_enable)
  );
  FringeFF regs_465 ( // @[RegFile.scala 66:20:@40921.4]
    .clock(regs_465_clock),
    .reset(regs_465_reset),
    .io_in(regs_465_io_in),
    .io_reset(regs_465_io_reset),
    .io_out(regs_465_io_out),
    .io_enable(regs_465_io_enable)
  );
  FringeFF regs_466 ( // @[RegFile.scala 66:20:@40935.4]
    .clock(regs_466_clock),
    .reset(regs_466_reset),
    .io_in(regs_466_io_in),
    .io_reset(regs_466_io_reset),
    .io_out(regs_466_io_out),
    .io_enable(regs_466_io_enable)
  );
  FringeFF regs_467 ( // @[RegFile.scala 66:20:@40949.4]
    .clock(regs_467_clock),
    .reset(regs_467_reset),
    .io_in(regs_467_io_in),
    .io_reset(regs_467_io_reset),
    .io_out(regs_467_io_out),
    .io_enable(regs_467_io_enable)
  );
  FringeFF regs_468 ( // @[RegFile.scala 66:20:@40963.4]
    .clock(regs_468_clock),
    .reset(regs_468_reset),
    .io_in(regs_468_io_in),
    .io_reset(regs_468_io_reset),
    .io_out(regs_468_io_out),
    .io_enable(regs_468_io_enable)
  );
  FringeFF regs_469 ( // @[RegFile.scala 66:20:@40977.4]
    .clock(regs_469_clock),
    .reset(regs_469_reset),
    .io_in(regs_469_io_in),
    .io_reset(regs_469_io_reset),
    .io_out(regs_469_io_out),
    .io_enable(regs_469_io_enable)
  );
  FringeFF regs_470 ( // @[RegFile.scala 66:20:@40991.4]
    .clock(regs_470_clock),
    .reset(regs_470_reset),
    .io_in(regs_470_io_in),
    .io_reset(regs_470_io_reset),
    .io_out(regs_470_io_out),
    .io_enable(regs_470_io_enable)
  );
  FringeFF regs_471 ( // @[RegFile.scala 66:20:@41005.4]
    .clock(regs_471_clock),
    .reset(regs_471_reset),
    .io_in(regs_471_io_in),
    .io_reset(regs_471_io_reset),
    .io_out(regs_471_io_out),
    .io_enable(regs_471_io_enable)
  );
  FringeFF regs_472 ( // @[RegFile.scala 66:20:@41019.4]
    .clock(regs_472_clock),
    .reset(regs_472_reset),
    .io_in(regs_472_io_in),
    .io_reset(regs_472_io_reset),
    .io_out(regs_472_io_out),
    .io_enable(regs_472_io_enable)
  );
  FringeFF regs_473 ( // @[RegFile.scala 66:20:@41033.4]
    .clock(regs_473_clock),
    .reset(regs_473_reset),
    .io_in(regs_473_io_in),
    .io_reset(regs_473_io_reset),
    .io_out(regs_473_io_out),
    .io_enable(regs_473_io_enable)
  );
  FringeFF regs_474 ( // @[RegFile.scala 66:20:@41047.4]
    .clock(regs_474_clock),
    .reset(regs_474_reset),
    .io_in(regs_474_io_in),
    .io_reset(regs_474_io_reset),
    .io_out(regs_474_io_out),
    .io_enable(regs_474_io_enable)
  );
  FringeFF regs_475 ( // @[RegFile.scala 66:20:@41061.4]
    .clock(regs_475_clock),
    .reset(regs_475_reset),
    .io_in(regs_475_io_in),
    .io_reset(regs_475_io_reset),
    .io_out(regs_475_io_out),
    .io_enable(regs_475_io_enable)
  );
  FringeFF regs_476 ( // @[RegFile.scala 66:20:@41075.4]
    .clock(regs_476_clock),
    .reset(regs_476_reset),
    .io_in(regs_476_io_in),
    .io_reset(regs_476_io_reset),
    .io_out(regs_476_io_out),
    .io_enable(regs_476_io_enable)
  );
  FringeFF regs_477 ( // @[RegFile.scala 66:20:@41089.4]
    .clock(regs_477_clock),
    .reset(regs_477_reset),
    .io_in(regs_477_io_in),
    .io_reset(regs_477_io_reset),
    .io_out(regs_477_io_out),
    .io_enable(regs_477_io_enable)
  );
  FringeFF regs_478 ( // @[RegFile.scala 66:20:@41103.4]
    .clock(regs_478_clock),
    .reset(regs_478_reset),
    .io_in(regs_478_io_in),
    .io_reset(regs_478_io_reset),
    .io_out(regs_478_io_out),
    .io_enable(regs_478_io_enable)
  );
  FringeFF regs_479 ( // @[RegFile.scala 66:20:@41117.4]
    .clock(regs_479_clock),
    .reset(regs_479_reset),
    .io_in(regs_479_io_in),
    .io_reset(regs_479_io_reset),
    .io_out(regs_479_io_out),
    .io_enable(regs_479_io_enable)
  );
  FringeFF regs_480 ( // @[RegFile.scala 66:20:@41131.4]
    .clock(regs_480_clock),
    .reset(regs_480_reset),
    .io_in(regs_480_io_in),
    .io_reset(regs_480_io_reset),
    .io_out(regs_480_io_out),
    .io_enable(regs_480_io_enable)
  );
  FringeFF regs_481 ( // @[RegFile.scala 66:20:@41145.4]
    .clock(regs_481_clock),
    .reset(regs_481_reset),
    .io_in(regs_481_io_in),
    .io_reset(regs_481_io_reset),
    .io_out(regs_481_io_out),
    .io_enable(regs_481_io_enable)
  );
  FringeFF regs_482 ( // @[RegFile.scala 66:20:@41159.4]
    .clock(regs_482_clock),
    .reset(regs_482_reset),
    .io_in(regs_482_io_in),
    .io_reset(regs_482_io_reset),
    .io_out(regs_482_io_out),
    .io_enable(regs_482_io_enable)
  );
  FringeFF regs_483 ( // @[RegFile.scala 66:20:@41173.4]
    .clock(regs_483_clock),
    .reset(regs_483_reset),
    .io_in(regs_483_io_in),
    .io_reset(regs_483_io_reset),
    .io_out(regs_483_io_out),
    .io_enable(regs_483_io_enable)
  );
  FringeFF regs_484 ( // @[RegFile.scala 66:20:@41187.4]
    .clock(regs_484_clock),
    .reset(regs_484_reset),
    .io_in(regs_484_io_in),
    .io_reset(regs_484_io_reset),
    .io_out(regs_484_io_out),
    .io_enable(regs_484_io_enable)
  );
  FringeFF regs_485 ( // @[RegFile.scala 66:20:@41201.4]
    .clock(regs_485_clock),
    .reset(regs_485_reset),
    .io_in(regs_485_io_in),
    .io_reset(regs_485_io_reset),
    .io_out(regs_485_io_out),
    .io_enable(regs_485_io_enable)
  );
  FringeFF regs_486 ( // @[RegFile.scala 66:20:@41215.4]
    .clock(regs_486_clock),
    .reset(regs_486_reset),
    .io_in(regs_486_io_in),
    .io_reset(regs_486_io_reset),
    .io_out(regs_486_io_out),
    .io_enable(regs_486_io_enable)
  );
  FringeFF regs_487 ( // @[RegFile.scala 66:20:@41229.4]
    .clock(regs_487_clock),
    .reset(regs_487_reset),
    .io_in(regs_487_io_in),
    .io_reset(regs_487_io_reset),
    .io_out(regs_487_io_out),
    .io_enable(regs_487_io_enable)
  );
  FringeFF regs_488 ( // @[RegFile.scala 66:20:@41243.4]
    .clock(regs_488_clock),
    .reset(regs_488_reset),
    .io_in(regs_488_io_in),
    .io_reset(regs_488_io_reset),
    .io_out(regs_488_io_out),
    .io_enable(regs_488_io_enable)
  );
  FringeFF regs_489 ( // @[RegFile.scala 66:20:@41257.4]
    .clock(regs_489_clock),
    .reset(regs_489_reset),
    .io_in(regs_489_io_in),
    .io_reset(regs_489_io_reset),
    .io_out(regs_489_io_out),
    .io_enable(regs_489_io_enable)
  );
  FringeFF regs_490 ( // @[RegFile.scala 66:20:@41271.4]
    .clock(regs_490_clock),
    .reset(regs_490_reset),
    .io_in(regs_490_io_in),
    .io_reset(regs_490_io_reset),
    .io_out(regs_490_io_out),
    .io_enable(regs_490_io_enable)
  );
  FringeFF regs_491 ( // @[RegFile.scala 66:20:@41285.4]
    .clock(regs_491_clock),
    .reset(regs_491_reset),
    .io_in(regs_491_io_in),
    .io_reset(regs_491_io_reset),
    .io_out(regs_491_io_out),
    .io_enable(regs_491_io_enable)
  );
  FringeFF regs_492 ( // @[RegFile.scala 66:20:@41299.4]
    .clock(regs_492_clock),
    .reset(regs_492_reset),
    .io_in(regs_492_io_in),
    .io_reset(regs_492_io_reset),
    .io_out(regs_492_io_out),
    .io_enable(regs_492_io_enable)
  );
  FringeFF regs_493 ( // @[RegFile.scala 66:20:@41313.4]
    .clock(regs_493_clock),
    .reset(regs_493_reset),
    .io_in(regs_493_io_in),
    .io_reset(regs_493_io_reset),
    .io_out(regs_493_io_out),
    .io_enable(regs_493_io_enable)
  );
  FringeFF regs_494 ( // @[RegFile.scala 66:20:@41327.4]
    .clock(regs_494_clock),
    .reset(regs_494_reset),
    .io_in(regs_494_io_in),
    .io_reset(regs_494_io_reset),
    .io_out(regs_494_io_out),
    .io_enable(regs_494_io_enable)
  );
  FringeFF regs_495 ( // @[RegFile.scala 66:20:@41341.4]
    .clock(regs_495_clock),
    .reset(regs_495_reset),
    .io_in(regs_495_io_in),
    .io_reset(regs_495_io_reset),
    .io_out(regs_495_io_out),
    .io_enable(regs_495_io_enable)
  );
  FringeFF regs_496 ( // @[RegFile.scala 66:20:@41355.4]
    .clock(regs_496_clock),
    .reset(regs_496_reset),
    .io_in(regs_496_io_in),
    .io_reset(regs_496_io_reset),
    .io_out(regs_496_io_out),
    .io_enable(regs_496_io_enable)
  );
  FringeFF regs_497 ( // @[RegFile.scala 66:20:@41369.4]
    .clock(regs_497_clock),
    .reset(regs_497_reset),
    .io_in(regs_497_io_in),
    .io_reset(regs_497_io_reset),
    .io_out(regs_497_io_out),
    .io_enable(regs_497_io_enable)
  );
  FringeFF regs_498 ( // @[RegFile.scala 66:20:@41383.4]
    .clock(regs_498_clock),
    .reset(regs_498_reset),
    .io_in(regs_498_io_in),
    .io_reset(regs_498_io_reset),
    .io_out(regs_498_io_out),
    .io_enable(regs_498_io_enable)
  );
  FringeFF regs_499 ( // @[RegFile.scala 66:20:@41397.4]
    .clock(regs_499_clock),
    .reset(regs_499_reset),
    .io_in(regs_499_io_in),
    .io_reset(regs_499_io_reset),
    .io_out(regs_499_io_out),
    .io_enable(regs_499_io_enable)
  );
  FringeFF regs_500 ( // @[RegFile.scala 66:20:@41411.4]
    .clock(regs_500_clock),
    .reset(regs_500_reset),
    .io_in(regs_500_io_in),
    .io_reset(regs_500_io_reset),
    .io_out(regs_500_io_out),
    .io_enable(regs_500_io_enable)
  );
  FringeFF regs_501 ( // @[RegFile.scala 66:20:@41425.4]
    .clock(regs_501_clock),
    .reset(regs_501_reset),
    .io_in(regs_501_io_in),
    .io_reset(regs_501_io_reset),
    .io_out(regs_501_io_out),
    .io_enable(regs_501_io_enable)
  );
  FringeFF regs_502 ( // @[RegFile.scala 66:20:@41439.4]
    .clock(regs_502_clock),
    .reset(regs_502_reset),
    .io_in(regs_502_io_in),
    .io_reset(regs_502_io_reset),
    .io_out(regs_502_io_out),
    .io_enable(regs_502_io_enable)
  );
  MuxN rport ( // @[RegFile.scala 95:21:@41453.4]
    .io_ins_0(rport_io_ins_0),
    .io_ins_1(rport_io_ins_1),
    .io_ins_2(rport_io_ins_2),
    .io_ins_3(rport_io_ins_3),
    .io_ins_4(rport_io_ins_4),
    .io_ins_5(rport_io_ins_5),
    .io_ins_6(rport_io_ins_6),
    .io_ins_7(rport_io_ins_7),
    .io_ins_8(rport_io_ins_8),
    .io_ins_9(rport_io_ins_9),
    .io_ins_10(rport_io_ins_10),
    .io_ins_11(rport_io_ins_11),
    .io_ins_12(rport_io_ins_12),
    .io_ins_13(rport_io_ins_13),
    .io_ins_14(rport_io_ins_14),
    .io_ins_15(rport_io_ins_15),
    .io_ins_16(rport_io_ins_16),
    .io_ins_17(rport_io_ins_17),
    .io_ins_18(rport_io_ins_18),
    .io_ins_19(rport_io_ins_19),
    .io_ins_20(rport_io_ins_20),
    .io_ins_21(rport_io_ins_21),
    .io_ins_22(rport_io_ins_22),
    .io_ins_23(rport_io_ins_23),
    .io_ins_24(rport_io_ins_24),
    .io_ins_25(rport_io_ins_25),
    .io_ins_26(rport_io_ins_26),
    .io_ins_27(rport_io_ins_27),
    .io_ins_28(rport_io_ins_28),
    .io_ins_29(rport_io_ins_29),
    .io_ins_30(rport_io_ins_30),
    .io_ins_31(rport_io_ins_31),
    .io_ins_32(rport_io_ins_32),
    .io_ins_33(rport_io_ins_33),
    .io_ins_34(rport_io_ins_34),
    .io_ins_35(rport_io_ins_35),
    .io_ins_36(rport_io_ins_36),
    .io_ins_37(rport_io_ins_37),
    .io_ins_38(rport_io_ins_38),
    .io_ins_39(rport_io_ins_39),
    .io_ins_40(rport_io_ins_40),
    .io_ins_41(rport_io_ins_41),
    .io_ins_42(rport_io_ins_42),
    .io_ins_43(rport_io_ins_43),
    .io_ins_44(rport_io_ins_44),
    .io_ins_45(rport_io_ins_45),
    .io_ins_46(rport_io_ins_46),
    .io_ins_47(rport_io_ins_47),
    .io_ins_48(rport_io_ins_48),
    .io_ins_49(rport_io_ins_49),
    .io_ins_50(rport_io_ins_50),
    .io_ins_51(rport_io_ins_51),
    .io_ins_52(rport_io_ins_52),
    .io_ins_53(rport_io_ins_53),
    .io_ins_54(rport_io_ins_54),
    .io_ins_55(rport_io_ins_55),
    .io_ins_56(rport_io_ins_56),
    .io_ins_57(rport_io_ins_57),
    .io_ins_58(rport_io_ins_58),
    .io_ins_59(rport_io_ins_59),
    .io_ins_60(rport_io_ins_60),
    .io_ins_61(rport_io_ins_61),
    .io_ins_62(rport_io_ins_62),
    .io_ins_63(rport_io_ins_63),
    .io_ins_64(rport_io_ins_64),
    .io_ins_65(rport_io_ins_65),
    .io_ins_66(rport_io_ins_66),
    .io_ins_67(rport_io_ins_67),
    .io_ins_68(rport_io_ins_68),
    .io_ins_69(rport_io_ins_69),
    .io_ins_70(rport_io_ins_70),
    .io_ins_71(rport_io_ins_71),
    .io_ins_72(rport_io_ins_72),
    .io_ins_73(rport_io_ins_73),
    .io_ins_74(rport_io_ins_74),
    .io_ins_75(rport_io_ins_75),
    .io_ins_76(rport_io_ins_76),
    .io_ins_77(rport_io_ins_77),
    .io_ins_78(rport_io_ins_78),
    .io_ins_79(rport_io_ins_79),
    .io_ins_80(rport_io_ins_80),
    .io_ins_81(rport_io_ins_81),
    .io_ins_82(rport_io_ins_82),
    .io_ins_83(rport_io_ins_83),
    .io_ins_84(rport_io_ins_84),
    .io_ins_85(rport_io_ins_85),
    .io_ins_86(rport_io_ins_86),
    .io_ins_87(rport_io_ins_87),
    .io_ins_88(rport_io_ins_88),
    .io_ins_89(rport_io_ins_89),
    .io_ins_90(rport_io_ins_90),
    .io_ins_91(rport_io_ins_91),
    .io_ins_92(rport_io_ins_92),
    .io_ins_93(rport_io_ins_93),
    .io_ins_94(rport_io_ins_94),
    .io_ins_95(rport_io_ins_95),
    .io_ins_96(rport_io_ins_96),
    .io_ins_97(rport_io_ins_97),
    .io_ins_98(rport_io_ins_98),
    .io_ins_99(rport_io_ins_99),
    .io_ins_100(rport_io_ins_100),
    .io_ins_101(rport_io_ins_101),
    .io_ins_102(rport_io_ins_102),
    .io_ins_103(rport_io_ins_103),
    .io_ins_104(rport_io_ins_104),
    .io_ins_105(rport_io_ins_105),
    .io_ins_106(rport_io_ins_106),
    .io_ins_107(rport_io_ins_107),
    .io_ins_108(rport_io_ins_108),
    .io_ins_109(rport_io_ins_109),
    .io_ins_110(rport_io_ins_110),
    .io_ins_111(rport_io_ins_111),
    .io_ins_112(rport_io_ins_112),
    .io_ins_113(rport_io_ins_113),
    .io_ins_114(rport_io_ins_114),
    .io_ins_115(rport_io_ins_115),
    .io_ins_116(rport_io_ins_116),
    .io_ins_117(rport_io_ins_117),
    .io_ins_118(rport_io_ins_118),
    .io_ins_119(rport_io_ins_119),
    .io_ins_120(rport_io_ins_120),
    .io_ins_121(rport_io_ins_121),
    .io_ins_122(rport_io_ins_122),
    .io_ins_123(rport_io_ins_123),
    .io_ins_124(rport_io_ins_124),
    .io_ins_125(rport_io_ins_125),
    .io_ins_126(rport_io_ins_126),
    .io_ins_127(rport_io_ins_127),
    .io_ins_128(rport_io_ins_128),
    .io_ins_129(rport_io_ins_129),
    .io_ins_130(rport_io_ins_130),
    .io_ins_131(rport_io_ins_131),
    .io_ins_132(rport_io_ins_132),
    .io_ins_133(rport_io_ins_133),
    .io_ins_134(rport_io_ins_134),
    .io_ins_135(rport_io_ins_135),
    .io_ins_136(rport_io_ins_136),
    .io_ins_137(rport_io_ins_137),
    .io_ins_138(rport_io_ins_138),
    .io_ins_139(rport_io_ins_139),
    .io_ins_140(rport_io_ins_140),
    .io_ins_141(rport_io_ins_141),
    .io_ins_142(rport_io_ins_142),
    .io_ins_143(rport_io_ins_143),
    .io_ins_144(rport_io_ins_144),
    .io_ins_145(rport_io_ins_145),
    .io_ins_146(rport_io_ins_146),
    .io_ins_147(rport_io_ins_147),
    .io_ins_148(rport_io_ins_148),
    .io_ins_149(rport_io_ins_149),
    .io_ins_150(rport_io_ins_150),
    .io_ins_151(rport_io_ins_151),
    .io_ins_152(rport_io_ins_152),
    .io_ins_153(rport_io_ins_153),
    .io_ins_154(rport_io_ins_154),
    .io_ins_155(rport_io_ins_155),
    .io_ins_156(rport_io_ins_156),
    .io_ins_157(rport_io_ins_157),
    .io_ins_158(rport_io_ins_158),
    .io_ins_159(rport_io_ins_159),
    .io_ins_160(rport_io_ins_160),
    .io_ins_161(rport_io_ins_161),
    .io_ins_162(rport_io_ins_162),
    .io_ins_163(rport_io_ins_163),
    .io_ins_164(rport_io_ins_164),
    .io_ins_165(rport_io_ins_165),
    .io_ins_166(rport_io_ins_166),
    .io_ins_167(rport_io_ins_167),
    .io_ins_168(rport_io_ins_168),
    .io_ins_169(rport_io_ins_169),
    .io_ins_170(rport_io_ins_170),
    .io_ins_171(rport_io_ins_171),
    .io_ins_172(rport_io_ins_172),
    .io_ins_173(rport_io_ins_173),
    .io_ins_174(rport_io_ins_174),
    .io_ins_175(rport_io_ins_175),
    .io_ins_176(rport_io_ins_176),
    .io_ins_177(rport_io_ins_177),
    .io_ins_178(rport_io_ins_178),
    .io_ins_179(rport_io_ins_179),
    .io_ins_180(rport_io_ins_180),
    .io_ins_181(rport_io_ins_181),
    .io_ins_182(rport_io_ins_182),
    .io_ins_183(rport_io_ins_183),
    .io_ins_184(rport_io_ins_184),
    .io_ins_185(rport_io_ins_185),
    .io_ins_186(rport_io_ins_186),
    .io_ins_187(rport_io_ins_187),
    .io_ins_188(rport_io_ins_188),
    .io_ins_189(rport_io_ins_189),
    .io_ins_190(rport_io_ins_190),
    .io_ins_191(rport_io_ins_191),
    .io_ins_192(rport_io_ins_192),
    .io_ins_193(rport_io_ins_193),
    .io_ins_194(rport_io_ins_194),
    .io_ins_195(rport_io_ins_195),
    .io_ins_196(rport_io_ins_196),
    .io_ins_197(rport_io_ins_197),
    .io_ins_198(rport_io_ins_198),
    .io_ins_199(rport_io_ins_199),
    .io_ins_200(rport_io_ins_200),
    .io_ins_201(rport_io_ins_201),
    .io_ins_202(rport_io_ins_202),
    .io_ins_203(rport_io_ins_203),
    .io_ins_204(rport_io_ins_204),
    .io_ins_205(rport_io_ins_205),
    .io_ins_206(rport_io_ins_206),
    .io_ins_207(rport_io_ins_207),
    .io_ins_208(rport_io_ins_208),
    .io_ins_209(rport_io_ins_209),
    .io_ins_210(rport_io_ins_210),
    .io_ins_211(rport_io_ins_211),
    .io_ins_212(rport_io_ins_212),
    .io_ins_213(rport_io_ins_213),
    .io_ins_214(rport_io_ins_214),
    .io_ins_215(rport_io_ins_215),
    .io_ins_216(rport_io_ins_216),
    .io_ins_217(rport_io_ins_217),
    .io_ins_218(rport_io_ins_218),
    .io_ins_219(rport_io_ins_219),
    .io_ins_220(rport_io_ins_220),
    .io_ins_221(rport_io_ins_221),
    .io_ins_222(rport_io_ins_222),
    .io_ins_223(rport_io_ins_223),
    .io_ins_224(rport_io_ins_224),
    .io_ins_225(rport_io_ins_225),
    .io_ins_226(rport_io_ins_226),
    .io_ins_227(rport_io_ins_227),
    .io_ins_228(rport_io_ins_228),
    .io_ins_229(rport_io_ins_229),
    .io_ins_230(rport_io_ins_230),
    .io_ins_231(rport_io_ins_231),
    .io_ins_232(rport_io_ins_232),
    .io_ins_233(rport_io_ins_233),
    .io_ins_234(rport_io_ins_234),
    .io_ins_235(rport_io_ins_235),
    .io_ins_236(rport_io_ins_236),
    .io_ins_237(rport_io_ins_237),
    .io_ins_238(rport_io_ins_238),
    .io_ins_239(rport_io_ins_239),
    .io_ins_240(rport_io_ins_240),
    .io_ins_241(rport_io_ins_241),
    .io_ins_242(rport_io_ins_242),
    .io_ins_243(rport_io_ins_243),
    .io_ins_244(rport_io_ins_244),
    .io_ins_245(rport_io_ins_245),
    .io_ins_246(rport_io_ins_246),
    .io_ins_247(rport_io_ins_247),
    .io_ins_248(rport_io_ins_248),
    .io_ins_249(rport_io_ins_249),
    .io_ins_250(rport_io_ins_250),
    .io_ins_251(rport_io_ins_251),
    .io_ins_252(rport_io_ins_252),
    .io_ins_253(rport_io_ins_253),
    .io_ins_254(rport_io_ins_254),
    .io_ins_255(rport_io_ins_255),
    .io_ins_256(rport_io_ins_256),
    .io_ins_257(rport_io_ins_257),
    .io_ins_258(rport_io_ins_258),
    .io_ins_259(rport_io_ins_259),
    .io_ins_260(rport_io_ins_260),
    .io_ins_261(rport_io_ins_261),
    .io_ins_262(rport_io_ins_262),
    .io_ins_263(rport_io_ins_263),
    .io_ins_264(rport_io_ins_264),
    .io_ins_265(rport_io_ins_265),
    .io_ins_266(rport_io_ins_266),
    .io_ins_267(rport_io_ins_267),
    .io_ins_268(rport_io_ins_268),
    .io_ins_269(rport_io_ins_269),
    .io_ins_270(rport_io_ins_270),
    .io_ins_271(rport_io_ins_271),
    .io_ins_272(rport_io_ins_272),
    .io_ins_273(rport_io_ins_273),
    .io_ins_274(rport_io_ins_274),
    .io_ins_275(rport_io_ins_275),
    .io_ins_276(rport_io_ins_276),
    .io_ins_277(rport_io_ins_277),
    .io_ins_278(rport_io_ins_278),
    .io_ins_279(rport_io_ins_279),
    .io_ins_280(rport_io_ins_280),
    .io_ins_281(rport_io_ins_281),
    .io_ins_282(rport_io_ins_282),
    .io_ins_283(rport_io_ins_283),
    .io_ins_284(rport_io_ins_284),
    .io_ins_285(rport_io_ins_285),
    .io_ins_286(rport_io_ins_286),
    .io_ins_287(rport_io_ins_287),
    .io_ins_288(rport_io_ins_288),
    .io_ins_289(rport_io_ins_289),
    .io_ins_290(rport_io_ins_290),
    .io_ins_291(rport_io_ins_291),
    .io_ins_292(rport_io_ins_292),
    .io_ins_293(rport_io_ins_293),
    .io_ins_294(rport_io_ins_294),
    .io_ins_295(rport_io_ins_295),
    .io_ins_296(rport_io_ins_296),
    .io_ins_297(rport_io_ins_297),
    .io_ins_298(rport_io_ins_298),
    .io_ins_299(rport_io_ins_299),
    .io_ins_300(rport_io_ins_300),
    .io_ins_301(rport_io_ins_301),
    .io_ins_302(rport_io_ins_302),
    .io_ins_303(rport_io_ins_303),
    .io_ins_304(rport_io_ins_304),
    .io_ins_305(rport_io_ins_305),
    .io_ins_306(rport_io_ins_306),
    .io_ins_307(rport_io_ins_307),
    .io_ins_308(rport_io_ins_308),
    .io_ins_309(rport_io_ins_309),
    .io_ins_310(rport_io_ins_310),
    .io_ins_311(rport_io_ins_311),
    .io_ins_312(rport_io_ins_312),
    .io_ins_313(rport_io_ins_313),
    .io_ins_314(rport_io_ins_314),
    .io_ins_315(rport_io_ins_315),
    .io_ins_316(rport_io_ins_316),
    .io_ins_317(rport_io_ins_317),
    .io_ins_318(rport_io_ins_318),
    .io_ins_319(rport_io_ins_319),
    .io_ins_320(rport_io_ins_320),
    .io_ins_321(rport_io_ins_321),
    .io_ins_322(rport_io_ins_322),
    .io_ins_323(rport_io_ins_323),
    .io_ins_324(rport_io_ins_324),
    .io_ins_325(rport_io_ins_325),
    .io_ins_326(rport_io_ins_326),
    .io_ins_327(rport_io_ins_327),
    .io_ins_328(rport_io_ins_328),
    .io_ins_329(rport_io_ins_329),
    .io_ins_330(rport_io_ins_330),
    .io_ins_331(rport_io_ins_331),
    .io_ins_332(rport_io_ins_332),
    .io_ins_333(rport_io_ins_333),
    .io_ins_334(rport_io_ins_334),
    .io_ins_335(rport_io_ins_335),
    .io_ins_336(rport_io_ins_336),
    .io_ins_337(rport_io_ins_337),
    .io_ins_338(rport_io_ins_338),
    .io_ins_339(rport_io_ins_339),
    .io_ins_340(rport_io_ins_340),
    .io_ins_341(rport_io_ins_341),
    .io_ins_342(rport_io_ins_342),
    .io_ins_343(rport_io_ins_343),
    .io_ins_344(rport_io_ins_344),
    .io_ins_345(rport_io_ins_345),
    .io_ins_346(rport_io_ins_346),
    .io_ins_347(rport_io_ins_347),
    .io_ins_348(rport_io_ins_348),
    .io_ins_349(rport_io_ins_349),
    .io_ins_350(rport_io_ins_350),
    .io_ins_351(rport_io_ins_351),
    .io_ins_352(rport_io_ins_352),
    .io_ins_353(rport_io_ins_353),
    .io_ins_354(rport_io_ins_354),
    .io_ins_355(rport_io_ins_355),
    .io_ins_356(rport_io_ins_356),
    .io_ins_357(rport_io_ins_357),
    .io_ins_358(rport_io_ins_358),
    .io_ins_359(rport_io_ins_359),
    .io_ins_360(rport_io_ins_360),
    .io_ins_361(rport_io_ins_361),
    .io_ins_362(rport_io_ins_362),
    .io_ins_363(rport_io_ins_363),
    .io_ins_364(rport_io_ins_364),
    .io_ins_365(rport_io_ins_365),
    .io_ins_366(rport_io_ins_366),
    .io_ins_367(rport_io_ins_367),
    .io_ins_368(rport_io_ins_368),
    .io_ins_369(rport_io_ins_369),
    .io_ins_370(rport_io_ins_370),
    .io_ins_371(rport_io_ins_371),
    .io_ins_372(rport_io_ins_372),
    .io_ins_373(rport_io_ins_373),
    .io_ins_374(rport_io_ins_374),
    .io_ins_375(rport_io_ins_375),
    .io_ins_376(rport_io_ins_376),
    .io_ins_377(rport_io_ins_377),
    .io_ins_378(rport_io_ins_378),
    .io_ins_379(rport_io_ins_379),
    .io_ins_380(rport_io_ins_380),
    .io_ins_381(rport_io_ins_381),
    .io_ins_382(rport_io_ins_382),
    .io_ins_383(rport_io_ins_383),
    .io_ins_384(rport_io_ins_384),
    .io_ins_385(rport_io_ins_385),
    .io_ins_386(rport_io_ins_386),
    .io_ins_387(rport_io_ins_387),
    .io_ins_388(rport_io_ins_388),
    .io_ins_389(rport_io_ins_389),
    .io_ins_390(rport_io_ins_390),
    .io_ins_391(rport_io_ins_391),
    .io_ins_392(rport_io_ins_392),
    .io_ins_393(rport_io_ins_393),
    .io_ins_394(rport_io_ins_394),
    .io_ins_395(rport_io_ins_395),
    .io_ins_396(rport_io_ins_396),
    .io_ins_397(rport_io_ins_397),
    .io_ins_398(rport_io_ins_398),
    .io_ins_399(rport_io_ins_399),
    .io_ins_400(rport_io_ins_400),
    .io_ins_401(rport_io_ins_401),
    .io_ins_402(rport_io_ins_402),
    .io_ins_403(rport_io_ins_403),
    .io_ins_404(rport_io_ins_404),
    .io_ins_405(rport_io_ins_405),
    .io_ins_406(rport_io_ins_406),
    .io_ins_407(rport_io_ins_407),
    .io_ins_408(rport_io_ins_408),
    .io_ins_409(rport_io_ins_409),
    .io_ins_410(rport_io_ins_410),
    .io_ins_411(rport_io_ins_411),
    .io_ins_412(rport_io_ins_412),
    .io_ins_413(rport_io_ins_413),
    .io_ins_414(rport_io_ins_414),
    .io_ins_415(rport_io_ins_415),
    .io_ins_416(rport_io_ins_416),
    .io_ins_417(rport_io_ins_417),
    .io_ins_418(rport_io_ins_418),
    .io_ins_419(rport_io_ins_419),
    .io_ins_420(rport_io_ins_420),
    .io_ins_421(rport_io_ins_421),
    .io_ins_422(rport_io_ins_422),
    .io_ins_423(rport_io_ins_423),
    .io_ins_424(rport_io_ins_424),
    .io_ins_425(rport_io_ins_425),
    .io_ins_426(rport_io_ins_426),
    .io_ins_427(rport_io_ins_427),
    .io_ins_428(rport_io_ins_428),
    .io_ins_429(rport_io_ins_429),
    .io_ins_430(rport_io_ins_430),
    .io_ins_431(rport_io_ins_431),
    .io_ins_432(rport_io_ins_432),
    .io_ins_433(rport_io_ins_433),
    .io_ins_434(rport_io_ins_434),
    .io_ins_435(rport_io_ins_435),
    .io_ins_436(rport_io_ins_436),
    .io_ins_437(rport_io_ins_437),
    .io_ins_438(rport_io_ins_438),
    .io_ins_439(rport_io_ins_439),
    .io_ins_440(rport_io_ins_440),
    .io_ins_441(rport_io_ins_441),
    .io_ins_442(rport_io_ins_442),
    .io_ins_443(rport_io_ins_443),
    .io_ins_444(rport_io_ins_444),
    .io_ins_445(rport_io_ins_445),
    .io_ins_446(rport_io_ins_446),
    .io_ins_447(rport_io_ins_447),
    .io_ins_448(rport_io_ins_448),
    .io_ins_449(rport_io_ins_449),
    .io_ins_450(rport_io_ins_450),
    .io_ins_451(rport_io_ins_451),
    .io_ins_452(rport_io_ins_452),
    .io_ins_453(rport_io_ins_453),
    .io_ins_454(rport_io_ins_454),
    .io_ins_455(rport_io_ins_455),
    .io_ins_456(rport_io_ins_456),
    .io_ins_457(rport_io_ins_457),
    .io_ins_458(rport_io_ins_458),
    .io_ins_459(rport_io_ins_459),
    .io_ins_460(rport_io_ins_460),
    .io_ins_461(rport_io_ins_461),
    .io_ins_462(rport_io_ins_462),
    .io_ins_463(rport_io_ins_463),
    .io_ins_464(rport_io_ins_464),
    .io_ins_465(rport_io_ins_465),
    .io_ins_466(rport_io_ins_466),
    .io_ins_467(rport_io_ins_467),
    .io_ins_468(rport_io_ins_468),
    .io_ins_469(rport_io_ins_469),
    .io_ins_470(rport_io_ins_470),
    .io_ins_471(rport_io_ins_471),
    .io_ins_472(rport_io_ins_472),
    .io_ins_473(rport_io_ins_473),
    .io_ins_474(rport_io_ins_474),
    .io_ins_475(rport_io_ins_475),
    .io_ins_476(rport_io_ins_476),
    .io_ins_477(rport_io_ins_477),
    .io_ins_478(rport_io_ins_478),
    .io_ins_479(rport_io_ins_479),
    .io_ins_480(rport_io_ins_480),
    .io_ins_481(rport_io_ins_481),
    .io_ins_482(rport_io_ins_482),
    .io_ins_483(rport_io_ins_483),
    .io_ins_484(rport_io_ins_484),
    .io_ins_485(rport_io_ins_485),
    .io_ins_486(rport_io_ins_486),
    .io_ins_487(rport_io_ins_487),
    .io_ins_488(rport_io_ins_488),
    .io_ins_489(rport_io_ins_489),
    .io_ins_490(rport_io_ins_490),
    .io_ins_491(rport_io_ins_491),
    .io_ins_492(rport_io_ins_492),
    .io_ins_493(rport_io_ins_493),
    .io_ins_494(rport_io_ins_494),
    .io_ins_495(rport_io_ins_495),
    .io_ins_496(rport_io_ins_496),
    .io_ins_497(rport_io_ins_497),
    .io_ins_498(rport_io_ins_498),
    .io_ins_499(rport_io_ins_499),
    .io_ins_500(rport_io_ins_500),
    .io_ins_501(rport_io_ins_501),
    .io_ins_502(rport_io_ins_502),
    .io_sel(rport_io_sel),
    .io_out(rport_io_out)
  );
  assign _T_3076 = io_waddr == 10'h0; // @[RegFile.scala 80:42:@34413.4]
  assign _T_3082 = io_waddr == 10'h1; // @[RegFile.scala 68:46:@34425.4]
  assign _T_3083 = io_wen & _T_3082; // @[RegFile.scala 68:34:@34426.4]
  assign _T_3096 = io_waddr == 10'h2; // @[RegFile.scala 80:42:@34444.4]
  assign _T_3102 = io_waddr == 10'h3; // @[RegFile.scala 74:80:@34456.4]
  assign _T_3103 = io_wen & _T_3102; // @[RegFile.scala 74:68:@34457.4]
  assign io_rdata = rport_io_out; // @[RegFile.scala 107:14:@42464.4]
  assign io_argIns_0 = regs_0_io_out; // @[RegFile.scala 111:13:@42469.4]
  assign io_argIns_1 = regs_1_io_out; // @[RegFile.scala 111:13:@42470.4]
  assign io_argIns_2 = regs_2_io_out; // @[RegFile.scala 111:13:@42471.4]
  assign io_argEchos_1 = regs_3_io_out; // @[RegFile.scala 77:37:@34463.4]
  assign regs_0_clock = clock; // @[:@34411.4]
  assign regs_0_reset = reset; // @[:@34412.4 RegFile.scala 82:16:@34418.4]
  assign regs_0_io_in = io_wdata; // @[RegFile.scala 81:16:@34416.4]
  assign regs_0_io_reset = reset; // @[RegFile.scala 83:19:@34420.4]
  assign regs_0_io_enable = io_wen & _T_3076; // @[RegFile.scala 80:20:@34415.4]
  assign regs_1_clock = clock; // @[:@34423.4]
  assign regs_1_reset = reset; // @[:@34424.4 RegFile.scala 70:16:@34436.4]
  assign regs_1_io_in = _T_3083 ? io_wdata : io_argOuts_0_bits; // @[RegFile.scala 69:16:@34434.4]
  assign regs_1_io_reset = reset; // @[RegFile.scala 72:19:@34439.4]
  assign regs_1_io_enable = _T_3083 ? _T_3083 : io_argOuts_0_valid; // @[RegFile.scala 68:20:@34430.4]
  assign regs_2_clock = clock; // @[:@34442.4]
  assign regs_2_reset = reset; // @[:@34443.4 RegFile.scala 82:16:@34449.4]
  assign regs_2_io_in = io_wdata; // @[RegFile.scala 81:16:@34447.4]
  assign regs_2_io_reset = reset; // @[RegFile.scala 83:19:@34451.4]
  assign regs_2_io_enable = io_wen & _T_3096; // @[RegFile.scala 80:20:@34446.4]
  assign regs_3_clock = clock; // @[:@34454.4]
  assign regs_3_reset = io_reset; // @[:@34455.4 RegFile.scala 76:16:@34462.4]
  assign regs_3_io_in = io_argOuts_1_valid ? io_argOuts_1_bits : io_wdata; // @[RegFile.scala 75:16:@34461.4]
  assign regs_3_io_reset = reset; // @[RegFile.scala 78:19:@34465.4]
  assign regs_3_io_enable = io_argOuts_1_valid | _T_3103; // @[RegFile.scala 74:20:@34459.4]
  assign regs_4_clock = clock; // @[:@34468.4]
  assign regs_4_reset = io_reset; // @[:@34469.4 RegFile.scala 76:16:@34476.4]
  assign regs_4_io_in = 64'h0; // @[RegFile.scala 75:16:@34475.4]
  assign regs_4_io_reset = reset; // @[RegFile.scala 78:19:@34479.4]
  assign regs_4_io_enable = 1'h1; // @[RegFile.scala 74:20:@34473.4]
  assign regs_5_clock = clock; // @[:@34482.4]
  assign regs_5_reset = io_reset; // @[:@34483.4 RegFile.scala 76:16:@34490.4]
  assign regs_5_io_in = 64'h0; // @[RegFile.scala 75:16:@34489.4]
  assign regs_5_io_reset = reset; // @[RegFile.scala 78:19:@34493.4]
  assign regs_5_io_enable = 1'h1; // @[RegFile.scala 74:20:@34487.4]
  assign regs_6_clock = clock; // @[:@34496.4]
  assign regs_6_reset = io_reset; // @[:@34497.4 RegFile.scala 76:16:@34504.4]
  assign regs_6_io_in = 64'h0; // @[RegFile.scala 75:16:@34503.4]
  assign regs_6_io_reset = reset; // @[RegFile.scala 78:19:@34507.4]
  assign regs_6_io_enable = 1'h1; // @[RegFile.scala 74:20:@34501.4]
  assign regs_7_clock = clock; // @[:@34510.4]
  assign regs_7_reset = io_reset; // @[:@34511.4 RegFile.scala 76:16:@34518.4]
  assign regs_7_io_in = 64'h0; // @[RegFile.scala 75:16:@34517.4]
  assign regs_7_io_reset = reset; // @[RegFile.scala 78:19:@34521.4]
  assign regs_7_io_enable = 1'h1; // @[RegFile.scala 74:20:@34515.4]
  assign regs_8_clock = clock; // @[:@34524.4]
  assign regs_8_reset = io_reset; // @[:@34525.4 RegFile.scala 76:16:@34532.4]
  assign regs_8_io_in = 64'h0; // @[RegFile.scala 75:16:@34531.4]
  assign regs_8_io_reset = reset; // @[RegFile.scala 78:19:@34535.4]
  assign regs_8_io_enable = 1'h1; // @[RegFile.scala 74:20:@34529.4]
  assign regs_9_clock = clock; // @[:@34538.4]
  assign regs_9_reset = io_reset; // @[:@34539.4 RegFile.scala 76:16:@34546.4]
  assign regs_9_io_in = 64'h0; // @[RegFile.scala 75:16:@34545.4]
  assign regs_9_io_reset = reset; // @[RegFile.scala 78:19:@34549.4]
  assign regs_9_io_enable = 1'h1; // @[RegFile.scala 74:20:@34543.4]
  assign regs_10_clock = clock; // @[:@34552.4]
  assign regs_10_reset = io_reset; // @[:@34553.4 RegFile.scala 76:16:@34560.4]
  assign regs_10_io_in = 64'h0; // @[RegFile.scala 75:16:@34559.4]
  assign regs_10_io_reset = reset; // @[RegFile.scala 78:19:@34563.4]
  assign regs_10_io_enable = 1'h1; // @[RegFile.scala 74:20:@34557.4]
  assign regs_11_clock = clock; // @[:@34566.4]
  assign regs_11_reset = io_reset; // @[:@34567.4 RegFile.scala 76:16:@34574.4]
  assign regs_11_io_in = 64'h0; // @[RegFile.scala 75:16:@34573.4]
  assign regs_11_io_reset = reset; // @[RegFile.scala 78:19:@34577.4]
  assign regs_11_io_enable = 1'h1; // @[RegFile.scala 74:20:@34571.4]
  assign regs_12_clock = clock; // @[:@34580.4]
  assign regs_12_reset = io_reset; // @[:@34581.4 RegFile.scala 76:16:@34588.4]
  assign regs_12_io_in = 64'h0; // @[RegFile.scala 75:16:@34587.4]
  assign regs_12_io_reset = reset; // @[RegFile.scala 78:19:@34591.4]
  assign regs_12_io_enable = 1'h1; // @[RegFile.scala 74:20:@34585.4]
  assign regs_13_clock = clock; // @[:@34594.4]
  assign regs_13_reset = io_reset; // @[:@34595.4 RegFile.scala 76:16:@34602.4]
  assign regs_13_io_in = 64'h0; // @[RegFile.scala 75:16:@34601.4]
  assign regs_13_io_reset = reset; // @[RegFile.scala 78:19:@34605.4]
  assign regs_13_io_enable = 1'h1; // @[RegFile.scala 74:20:@34599.4]
  assign regs_14_clock = clock; // @[:@34608.4]
  assign regs_14_reset = io_reset; // @[:@34609.4 RegFile.scala 76:16:@34616.4]
  assign regs_14_io_in = 64'h0; // @[RegFile.scala 75:16:@34615.4]
  assign regs_14_io_reset = reset; // @[RegFile.scala 78:19:@34619.4]
  assign regs_14_io_enable = 1'h1; // @[RegFile.scala 74:20:@34613.4]
  assign regs_15_clock = clock; // @[:@34622.4]
  assign regs_15_reset = io_reset; // @[:@34623.4 RegFile.scala 76:16:@34630.4]
  assign regs_15_io_in = 64'h0; // @[RegFile.scala 75:16:@34629.4]
  assign regs_15_io_reset = reset; // @[RegFile.scala 78:19:@34633.4]
  assign regs_15_io_enable = 1'h1; // @[RegFile.scala 74:20:@34627.4]
  assign regs_16_clock = clock; // @[:@34636.4]
  assign regs_16_reset = io_reset; // @[:@34637.4 RegFile.scala 76:16:@34644.4]
  assign regs_16_io_in = 64'h0; // @[RegFile.scala 75:16:@34643.4]
  assign regs_16_io_reset = reset; // @[RegFile.scala 78:19:@34647.4]
  assign regs_16_io_enable = 1'h1; // @[RegFile.scala 74:20:@34641.4]
  assign regs_17_clock = clock; // @[:@34650.4]
  assign regs_17_reset = io_reset; // @[:@34651.4 RegFile.scala 76:16:@34658.4]
  assign regs_17_io_in = 64'h0; // @[RegFile.scala 75:16:@34657.4]
  assign regs_17_io_reset = reset; // @[RegFile.scala 78:19:@34661.4]
  assign regs_17_io_enable = 1'h1; // @[RegFile.scala 74:20:@34655.4]
  assign regs_18_clock = clock; // @[:@34664.4]
  assign regs_18_reset = io_reset; // @[:@34665.4 RegFile.scala 76:16:@34672.4]
  assign regs_18_io_in = 64'h0; // @[RegFile.scala 75:16:@34671.4]
  assign regs_18_io_reset = reset; // @[RegFile.scala 78:19:@34675.4]
  assign regs_18_io_enable = 1'h1; // @[RegFile.scala 74:20:@34669.4]
  assign regs_19_clock = clock; // @[:@34678.4]
  assign regs_19_reset = io_reset; // @[:@34679.4 RegFile.scala 76:16:@34686.4]
  assign regs_19_io_in = 64'h0; // @[RegFile.scala 75:16:@34685.4]
  assign regs_19_io_reset = reset; // @[RegFile.scala 78:19:@34689.4]
  assign regs_19_io_enable = 1'h1; // @[RegFile.scala 74:20:@34683.4]
  assign regs_20_clock = clock; // @[:@34692.4]
  assign regs_20_reset = io_reset; // @[:@34693.4 RegFile.scala 76:16:@34700.4]
  assign regs_20_io_in = 64'h0; // @[RegFile.scala 75:16:@34699.4]
  assign regs_20_io_reset = reset; // @[RegFile.scala 78:19:@34703.4]
  assign regs_20_io_enable = 1'h1; // @[RegFile.scala 74:20:@34697.4]
  assign regs_21_clock = clock; // @[:@34706.4]
  assign regs_21_reset = io_reset; // @[:@34707.4 RegFile.scala 76:16:@34714.4]
  assign regs_21_io_in = 64'h0; // @[RegFile.scala 75:16:@34713.4]
  assign regs_21_io_reset = reset; // @[RegFile.scala 78:19:@34717.4]
  assign regs_21_io_enable = 1'h1; // @[RegFile.scala 74:20:@34711.4]
  assign regs_22_clock = clock; // @[:@34720.4]
  assign regs_22_reset = io_reset; // @[:@34721.4 RegFile.scala 76:16:@34728.4]
  assign regs_22_io_in = 64'h0; // @[RegFile.scala 75:16:@34727.4]
  assign regs_22_io_reset = reset; // @[RegFile.scala 78:19:@34731.4]
  assign regs_22_io_enable = 1'h1; // @[RegFile.scala 74:20:@34725.4]
  assign regs_23_clock = clock; // @[:@34734.4]
  assign regs_23_reset = io_reset; // @[:@34735.4 RegFile.scala 76:16:@34742.4]
  assign regs_23_io_in = 64'h0; // @[RegFile.scala 75:16:@34741.4]
  assign regs_23_io_reset = reset; // @[RegFile.scala 78:19:@34745.4]
  assign regs_23_io_enable = 1'h1; // @[RegFile.scala 74:20:@34739.4]
  assign regs_24_clock = clock; // @[:@34748.4]
  assign regs_24_reset = io_reset; // @[:@34749.4 RegFile.scala 76:16:@34756.4]
  assign regs_24_io_in = 64'h0; // @[RegFile.scala 75:16:@34755.4]
  assign regs_24_io_reset = reset; // @[RegFile.scala 78:19:@34759.4]
  assign regs_24_io_enable = 1'h1; // @[RegFile.scala 74:20:@34753.4]
  assign regs_25_clock = clock; // @[:@34762.4]
  assign regs_25_reset = io_reset; // @[:@34763.4 RegFile.scala 76:16:@34770.4]
  assign regs_25_io_in = 64'h0; // @[RegFile.scala 75:16:@34769.4]
  assign regs_25_io_reset = reset; // @[RegFile.scala 78:19:@34773.4]
  assign regs_25_io_enable = 1'h1; // @[RegFile.scala 74:20:@34767.4]
  assign regs_26_clock = clock; // @[:@34776.4]
  assign regs_26_reset = io_reset; // @[:@34777.4 RegFile.scala 76:16:@34784.4]
  assign regs_26_io_in = 64'h0; // @[RegFile.scala 75:16:@34783.4]
  assign regs_26_io_reset = reset; // @[RegFile.scala 78:19:@34787.4]
  assign regs_26_io_enable = 1'h1; // @[RegFile.scala 74:20:@34781.4]
  assign regs_27_clock = clock; // @[:@34790.4]
  assign regs_27_reset = io_reset; // @[:@34791.4 RegFile.scala 76:16:@34798.4]
  assign regs_27_io_in = 64'h0; // @[RegFile.scala 75:16:@34797.4]
  assign regs_27_io_reset = reset; // @[RegFile.scala 78:19:@34801.4]
  assign regs_27_io_enable = 1'h1; // @[RegFile.scala 74:20:@34795.4]
  assign regs_28_clock = clock; // @[:@34804.4]
  assign regs_28_reset = io_reset; // @[:@34805.4 RegFile.scala 76:16:@34812.4]
  assign regs_28_io_in = 64'h0; // @[RegFile.scala 75:16:@34811.4]
  assign regs_28_io_reset = reset; // @[RegFile.scala 78:19:@34815.4]
  assign regs_28_io_enable = 1'h1; // @[RegFile.scala 74:20:@34809.4]
  assign regs_29_clock = clock; // @[:@34818.4]
  assign regs_29_reset = io_reset; // @[:@34819.4 RegFile.scala 76:16:@34826.4]
  assign regs_29_io_in = 64'h0; // @[RegFile.scala 75:16:@34825.4]
  assign regs_29_io_reset = reset; // @[RegFile.scala 78:19:@34829.4]
  assign regs_29_io_enable = 1'h1; // @[RegFile.scala 74:20:@34823.4]
  assign regs_30_clock = clock; // @[:@34832.4]
  assign regs_30_reset = io_reset; // @[:@34833.4 RegFile.scala 76:16:@34840.4]
  assign regs_30_io_in = 64'h0; // @[RegFile.scala 75:16:@34839.4]
  assign regs_30_io_reset = reset; // @[RegFile.scala 78:19:@34843.4]
  assign regs_30_io_enable = 1'h1; // @[RegFile.scala 74:20:@34837.4]
  assign regs_31_clock = clock; // @[:@34846.4]
  assign regs_31_reset = io_reset; // @[:@34847.4 RegFile.scala 76:16:@34854.4]
  assign regs_31_io_in = 64'h0; // @[RegFile.scala 75:16:@34853.4]
  assign regs_31_io_reset = reset; // @[RegFile.scala 78:19:@34857.4]
  assign regs_31_io_enable = 1'h1; // @[RegFile.scala 74:20:@34851.4]
  assign regs_32_clock = clock; // @[:@34860.4]
  assign regs_32_reset = io_reset; // @[:@34861.4 RegFile.scala 76:16:@34868.4]
  assign regs_32_io_in = 64'h0; // @[RegFile.scala 75:16:@34867.4]
  assign regs_32_io_reset = reset; // @[RegFile.scala 78:19:@34871.4]
  assign regs_32_io_enable = 1'h1; // @[RegFile.scala 74:20:@34865.4]
  assign regs_33_clock = clock; // @[:@34874.4]
  assign regs_33_reset = io_reset; // @[:@34875.4 RegFile.scala 76:16:@34882.4]
  assign regs_33_io_in = 64'h0; // @[RegFile.scala 75:16:@34881.4]
  assign regs_33_io_reset = reset; // @[RegFile.scala 78:19:@34885.4]
  assign regs_33_io_enable = 1'h1; // @[RegFile.scala 74:20:@34879.4]
  assign regs_34_clock = clock; // @[:@34888.4]
  assign regs_34_reset = io_reset; // @[:@34889.4 RegFile.scala 76:16:@34896.4]
  assign regs_34_io_in = 64'h0; // @[RegFile.scala 75:16:@34895.4]
  assign regs_34_io_reset = reset; // @[RegFile.scala 78:19:@34899.4]
  assign regs_34_io_enable = 1'h1; // @[RegFile.scala 74:20:@34893.4]
  assign regs_35_clock = clock; // @[:@34902.4]
  assign regs_35_reset = io_reset; // @[:@34903.4 RegFile.scala 76:16:@34910.4]
  assign regs_35_io_in = 64'h0; // @[RegFile.scala 75:16:@34909.4]
  assign regs_35_io_reset = reset; // @[RegFile.scala 78:19:@34913.4]
  assign regs_35_io_enable = 1'h1; // @[RegFile.scala 74:20:@34907.4]
  assign regs_36_clock = clock; // @[:@34916.4]
  assign regs_36_reset = io_reset; // @[:@34917.4 RegFile.scala 76:16:@34924.4]
  assign regs_36_io_in = 64'h0; // @[RegFile.scala 75:16:@34923.4]
  assign regs_36_io_reset = reset; // @[RegFile.scala 78:19:@34927.4]
  assign regs_36_io_enable = 1'h1; // @[RegFile.scala 74:20:@34921.4]
  assign regs_37_clock = clock; // @[:@34930.4]
  assign regs_37_reset = io_reset; // @[:@34931.4 RegFile.scala 76:16:@34938.4]
  assign regs_37_io_in = 64'h0; // @[RegFile.scala 75:16:@34937.4]
  assign regs_37_io_reset = reset; // @[RegFile.scala 78:19:@34941.4]
  assign regs_37_io_enable = 1'h1; // @[RegFile.scala 74:20:@34935.4]
  assign regs_38_clock = clock; // @[:@34944.4]
  assign regs_38_reset = io_reset; // @[:@34945.4 RegFile.scala 76:16:@34952.4]
  assign regs_38_io_in = 64'h0; // @[RegFile.scala 75:16:@34951.4]
  assign regs_38_io_reset = reset; // @[RegFile.scala 78:19:@34955.4]
  assign regs_38_io_enable = 1'h1; // @[RegFile.scala 74:20:@34949.4]
  assign regs_39_clock = clock; // @[:@34958.4]
  assign regs_39_reset = io_reset; // @[:@34959.4 RegFile.scala 76:16:@34966.4]
  assign regs_39_io_in = 64'h0; // @[RegFile.scala 75:16:@34965.4]
  assign regs_39_io_reset = reset; // @[RegFile.scala 78:19:@34969.4]
  assign regs_39_io_enable = 1'h1; // @[RegFile.scala 74:20:@34963.4]
  assign regs_40_clock = clock; // @[:@34972.4]
  assign regs_40_reset = io_reset; // @[:@34973.4 RegFile.scala 76:16:@34980.4]
  assign regs_40_io_in = 64'h0; // @[RegFile.scala 75:16:@34979.4]
  assign regs_40_io_reset = reset; // @[RegFile.scala 78:19:@34983.4]
  assign regs_40_io_enable = 1'h1; // @[RegFile.scala 74:20:@34977.4]
  assign regs_41_clock = clock; // @[:@34986.4]
  assign regs_41_reset = io_reset; // @[:@34987.4 RegFile.scala 76:16:@34994.4]
  assign regs_41_io_in = 64'h0; // @[RegFile.scala 75:16:@34993.4]
  assign regs_41_io_reset = reset; // @[RegFile.scala 78:19:@34997.4]
  assign regs_41_io_enable = 1'h1; // @[RegFile.scala 74:20:@34991.4]
  assign regs_42_clock = clock; // @[:@35000.4]
  assign regs_42_reset = io_reset; // @[:@35001.4 RegFile.scala 76:16:@35008.4]
  assign regs_42_io_in = 64'h0; // @[RegFile.scala 75:16:@35007.4]
  assign regs_42_io_reset = reset; // @[RegFile.scala 78:19:@35011.4]
  assign regs_42_io_enable = 1'h1; // @[RegFile.scala 74:20:@35005.4]
  assign regs_43_clock = clock; // @[:@35014.4]
  assign regs_43_reset = io_reset; // @[:@35015.4 RegFile.scala 76:16:@35022.4]
  assign regs_43_io_in = 64'h0; // @[RegFile.scala 75:16:@35021.4]
  assign regs_43_io_reset = reset; // @[RegFile.scala 78:19:@35025.4]
  assign regs_43_io_enable = 1'h1; // @[RegFile.scala 74:20:@35019.4]
  assign regs_44_clock = clock; // @[:@35028.4]
  assign regs_44_reset = io_reset; // @[:@35029.4 RegFile.scala 76:16:@35036.4]
  assign regs_44_io_in = 64'h0; // @[RegFile.scala 75:16:@35035.4]
  assign regs_44_io_reset = reset; // @[RegFile.scala 78:19:@35039.4]
  assign regs_44_io_enable = 1'h1; // @[RegFile.scala 74:20:@35033.4]
  assign regs_45_clock = clock; // @[:@35042.4]
  assign regs_45_reset = io_reset; // @[:@35043.4 RegFile.scala 76:16:@35050.4]
  assign regs_45_io_in = 64'h0; // @[RegFile.scala 75:16:@35049.4]
  assign regs_45_io_reset = reset; // @[RegFile.scala 78:19:@35053.4]
  assign regs_45_io_enable = 1'h1; // @[RegFile.scala 74:20:@35047.4]
  assign regs_46_clock = clock; // @[:@35056.4]
  assign regs_46_reset = io_reset; // @[:@35057.4 RegFile.scala 76:16:@35064.4]
  assign regs_46_io_in = 64'h0; // @[RegFile.scala 75:16:@35063.4]
  assign regs_46_io_reset = reset; // @[RegFile.scala 78:19:@35067.4]
  assign regs_46_io_enable = 1'h1; // @[RegFile.scala 74:20:@35061.4]
  assign regs_47_clock = clock; // @[:@35070.4]
  assign regs_47_reset = io_reset; // @[:@35071.4 RegFile.scala 76:16:@35078.4]
  assign regs_47_io_in = 64'h0; // @[RegFile.scala 75:16:@35077.4]
  assign regs_47_io_reset = reset; // @[RegFile.scala 78:19:@35081.4]
  assign regs_47_io_enable = 1'h1; // @[RegFile.scala 74:20:@35075.4]
  assign regs_48_clock = clock; // @[:@35084.4]
  assign regs_48_reset = io_reset; // @[:@35085.4 RegFile.scala 76:16:@35092.4]
  assign regs_48_io_in = 64'h0; // @[RegFile.scala 75:16:@35091.4]
  assign regs_48_io_reset = reset; // @[RegFile.scala 78:19:@35095.4]
  assign regs_48_io_enable = 1'h1; // @[RegFile.scala 74:20:@35089.4]
  assign regs_49_clock = clock; // @[:@35098.4]
  assign regs_49_reset = io_reset; // @[:@35099.4 RegFile.scala 76:16:@35106.4]
  assign regs_49_io_in = 64'h0; // @[RegFile.scala 75:16:@35105.4]
  assign regs_49_io_reset = reset; // @[RegFile.scala 78:19:@35109.4]
  assign regs_49_io_enable = 1'h1; // @[RegFile.scala 74:20:@35103.4]
  assign regs_50_clock = clock; // @[:@35112.4]
  assign regs_50_reset = io_reset; // @[:@35113.4 RegFile.scala 76:16:@35120.4]
  assign regs_50_io_in = 64'h0; // @[RegFile.scala 75:16:@35119.4]
  assign regs_50_io_reset = reset; // @[RegFile.scala 78:19:@35123.4]
  assign regs_50_io_enable = 1'h1; // @[RegFile.scala 74:20:@35117.4]
  assign regs_51_clock = clock; // @[:@35126.4]
  assign regs_51_reset = io_reset; // @[:@35127.4 RegFile.scala 76:16:@35134.4]
  assign regs_51_io_in = 64'h0; // @[RegFile.scala 75:16:@35133.4]
  assign regs_51_io_reset = reset; // @[RegFile.scala 78:19:@35137.4]
  assign regs_51_io_enable = 1'h1; // @[RegFile.scala 74:20:@35131.4]
  assign regs_52_clock = clock; // @[:@35140.4]
  assign regs_52_reset = io_reset; // @[:@35141.4 RegFile.scala 76:16:@35148.4]
  assign regs_52_io_in = 64'h0; // @[RegFile.scala 75:16:@35147.4]
  assign regs_52_io_reset = reset; // @[RegFile.scala 78:19:@35151.4]
  assign regs_52_io_enable = 1'h1; // @[RegFile.scala 74:20:@35145.4]
  assign regs_53_clock = clock; // @[:@35154.4]
  assign regs_53_reset = io_reset; // @[:@35155.4 RegFile.scala 76:16:@35162.4]
  assign regs_53_io_in = 64'h0; // @[RegFile.scala 75:16:@35161.4]
  assign regs_53_io_reset = reset; // @[RegFile.scala 78:19:@35165.4]
  assign regs_53_io_enable = 1'h1; // @[RegFile.scala 74:20:@35159.4]
  assign regs_54_clock = clock; // @[:@35168.4]
  assign regs_54_reset = io_reset; // @[:@35169.4 RegFile.scala 76:16:@35176.4]
  assign regs_54_io_in = 64'h0; // @[RegFile.scala 75:16:@35175.4]
  assign regs_54_io_reset = reset; // @[RegFile.scala 78:19:@35179.4]
  assign regs_54_io_enable = 1'h1; // @[RegFile.scala 74:20:@35173.4]
  assign regs_55_clock = clock; // @[:@35182.4]
  assign regs_55_reset = io_reset; // @[:@35183.4 RegFile.scala 76:16:@35190.4]
  assign regs_55_io_in = 64'h0; // @[RegFile.scala 75:16:@35189.4]
  assign regs_55_io_reset = reset; // @[RegFile.scala 78:19:@35193.4]
  assign regs_55_io_enable = 1'h1; // @[RegFile.scala 74:20:@35187.4]
  assign regs_56_clock = clock; // @[:@35196.4]
  assign regs_56_reset = io_reset; // @[:@35197.4 RegFile.scala 76:16:@35204.4]
  assign regs_56_io_in = 64'h0; // @[RegFile.scala 75:16:@35203.4]
  assign regs_56_io_reset = reset; // @[RegFile.scala 78:19:@35207.4]
  assign regs_56_io_enable = 1'h1; // @[RegFile.scala 74:20:@35201.4]
  assign regs_57_clock = clock; // @[:@35210.4]
  assign regs_57_reset = io_reset; // @[:@35211.4 RegFile.scala 76:16:@35218.4]
  assign regs_57_io_in = 64'h0; // @[RegFile.scala 75:16:@35217.4]
  assign regs_57_io_reset = reset; // @[RegFile.scala 78:19:@35221.4]
  assign regs_57_io_enable = 1'h1; // @[RegFile.scala 74:20:@35215.4]
  assign regs_58_clock = clock; // @[:@35224.4]
  assign regs_58_reset = io_reset; // @[:@35225.4 RegFile.scala 76:16:@35232.4]
  assign regs_58_io_in = 64'h0; // @[RegFile.scala 75:16:@35231.4]
  assign regs_58_io_reset = reset; // @[RegFile.scala 78:19:@35235.4]
  assign regs_58_io_enable = 1'h1; // @[RegFile.scala 74:20:@35229.4]
  assign regs_59_clock = clock; // @[:@35238.4]
  assign regs_59_reset = io_reset; // @[:@35239.4 RegFile.scala 76:16:@35246.4]
  assign regs_59_io_in = 64'h0; // @[RegFile.scala 75:16:@35245.4]
  assign regs_59_io_reset = reset; // @[RegFile.scala 78:19:@35249.4]
  assign regs_59_io_enable = 1'h1; // @[RegFile.scala 74:20:@35243.4]
  assign regs_60_clock = clock; // @[:@35252.4]
  assign regs_60_reset = io_reset; // @[:@35253.4 RegFile.scala 76:16:@35260.4]
  assign regs_60_io_in = 64'h0; // @[RegFile.scala 75:16:@35259.4]
  assign regs_60_io_reset = reset; // @[RegFile.scala 78:19:@35263.4]
  assign regs_60_io_enable = 1'h1; // @[RegFile.scala 74:20:@35257.4]
  assign regs_61_clock = clock; // @[:@35266.4]
  assign regs_61_reset = io_reset; // @[:@35267.4 RegFile.scala 76:16:@35274.4]
  assign regs_61_io_in = 64'h0; // @[RegFile.scala 75:16:@35273.4]
  assign regs_61_io_reset = reset; // @[RegFile.scala 78:19:@35277.4]
  assign regs_61_io_enable = 1'h1; // @[RegFile.scala 74:20:@35271.4]
  assign regs_62_clock = clock; // @[:@35280.4]
  assign regs_62_reset = io_reset; // @[:@35281.4 RegFile.scala 76:16:@35288.4]
  assign regs_62_io_in = 64'h0; // @[RegFile.scala 75:16:@35287.4]
  assign regs_62_io_reset = reset; // @[RegFile.scala 78:19:@35291.4]
  assign regs_62_io_enable = 1'h1; // @[RegFile.scala 74:20:@35285.4]
  assign regs_63_clock = clock; // @[:@35294.4]
  assign regs_63_reset = io_reset; // @[:@35295.4 RegFile.scala 76:16:@35302.4]
  assign regs_63_io_in = 64'h0; // @[RegFile.scala 75:16:@35301.4]
  assign regs_63_io_reset = reset; // @[RegFile.scala 78:19:@35305.4]
  assign regs_63_io_enable = 1'h1; // @[RegFile.scala 74:20:@35299.4]
  assign regs_64_clock = clock; // @[:@35308.4]
  assign regs_64_reset = io_reset; // @[:@35309.4 RegFile.scala 76:16:@35316.4]
  assign regs_64_io_in = 64'h0; // @[RegFile.scala 75:16:@35315.4]
  assign regs_64_io_reset = reset; // @[RegFile.scala 78:19:@35319.4]
  assign regs_64_io_enable = 1'h1; // @[RegFile.scala 74:20:@35313.4]
  assign regs_65_clock = clock; // @[:@35322.4]
  assign regs_65_reset = io_reset; // @[:@35323.4 RegFile.scala 76:16:@35330.4]
  assign regs_65_io_in = 64'h0; // @[RegFile.scala 75:16:@35329.4]
  assign regs_65_io_reset = reset; // @[RegFile.scala 78:19:@35333.4]
  assign regs_65_io_enable = 1'h1; // @[RegFile.scala 74:20:@35327.4]
  assign regs_66_clock = clock; // @[:@35336.4]
  assign regs_66_reset = io_reset; // @[:@35337.4 RegFile.scala 76:16:@35344.4]
  assign regs_66_io_in = 64'h0; // @[RegFile.scala 75:16:@35343.4]
  assign regs_66_io_reset = reset; // @[RegFile.scala 78:19:@35347.4]
  assign regs_66_io_enable = 1'h1; // @[RegFile.scala 74:20:@35341.4]
  assign regs_67_clock = clock; // @[:@35350.4]
  assign regs_67_reset = io_reset; // @[:@35351.4 RegFile.scala 76:16:@35358.4]
  assign regs_67_io_in = 64'h0; // @[RegFile.scala 75:16:@35357.4]
  assign regs_67_io_reset = reset; // @[RegFile.scala 78:19:@35361.4]
  assign regs_67_io_enable = 1'h1; // @[RegFile.scala 74:20:@35355.4]
  assign regs_68_clock = clock; // @[:@35364.4]
  assign regs_68_reset = io_reset; // @[:@35365.4 RegFile.scala 76:16:@35372.4]
  assign regs_68_io_in = 64'h0; // @[RegFile.scala 75:16:@35371.4]
  assign regs_68_io_reset = reset; // @[RegFile.scala 78:19:@35375.4]
  assign regs_68_io_enable = 1'h1; // @[RegFile.scala 74:20:@35369.4]
  assign regs_69_clock = clock; // @[:@35378.4]
  assign regs_69_reset = io_reset; // @[:@35379.4 RegFile.scala 76:16:@35386.4]
  assign regs_69_io_in = 64'h0; // @[RegFile.scala 75:16:@35385.4]
  assign regs_69_io_reset = reset; // @[RegFile.scala 78:19:@35389.4]
  assign regs_69_io_enable = 1'h1; // @[RegFile.scala 74:20:@35383.4]
  assign regs_70_clock = clock; // @[:@35392.4]
  assign regs_70_reset = io_reset; // @[:@35393.4 RegFile.scala 76:16:@35400.4]
  assign regs_70_io_in = 64'h0; // @[RegFile.scala 75:16:@35399.4]
  assign regs_70_io_reset = reset; // @[RegFile.scala 78:19:@35403.4]
  assign regs_70_io_enable = 1'h1; // @[RegFile.scala 74:20:@35397.4]
  assign regs_71_clock = clock; // @[:@35406.4]
  assign regs_71_reset = io_reset; // @[:@35407.4 RegFile.scala 76:16:@35414.4]
  assign regs_71_io_in = 64'h0; // @[RegFile.scala 75:16:@35413.4]
  assign regs_71_io_reset = reset; // @[RegFile.scala 78:19:@35417.4]
  assign regs_71_io_enable = 1'h1; // @[RegFile.scala 74:20:@35411.4]
  assign regs_72_clock = clock; // @[:@35420.4]
  assign regs_72_reset = io_reset; // @[:@35421.4 RegFile.scala 76:16:@35428.4]
  assign regs_72_io_in = 64'h0; // @[RegFile.scala 75:16:@35427.4]
  assign regs_72_io_reset = reset; // @[RegFile.scala 78:19:@35431.4]
  assign regs_72_io_enable = 1'h1; // @[RegFile.scala 74:20:@35425.4]
  assign regs_73_clock = clock; // @[:@35434.4]
  assign regs_73_reset = io_reset; // @[:@35435.4 RegFile.scala 76:16:@35442.4]
  assign regs_73_io_in = 64'h0; // @[RegFile.scala 75:16:@35441.4]
  assign regs_73_io_reset = reset; // @[RegFile.scala 78:19:@35445.4]
  assign regs_73_io_enable = 1'h1; // @[RegFile.scala 74:20:@35439.4]
  assign regs_74_clock = clock; // @[:@35448.4]
  assign regs_74_reset = io_reset; // @[:@35449.4 RegFile.scala 76:16:@35456.4]
  assign regs_74_io_in = 64'h0; // @[RegFile.scala 75:16:@35455.4]
  assign regs_74_io_reset = reset; // @[RegFile.scala 78:19:@35459.4]
  assign regs_74_io_enable = 1'h1; // @[RegFile.scala 74:20:@35453.4]
  assign regs_75_clock = clock; // @[:@35462.4]
  assign regs_75_reset = io_reset; // @[:@35463.4 RegFile.scala 76:16:@35470.4]
  assign regs_75_io_in = 64'h0; // @[RegFile.scala 75:16:@35469.4]
  assign regs_75_io_reset = reset; // @[RegFile.scala 78:19:@35473.4]
  assign regs_75_io_enable = 1'h1; // @[RegFile.scala 74:20:@35467.4]
  assign regs_76_clock = clock; // @[:@35476.4]
  assign regs_76_reset = io_reset; // @[:@35477.4 RegFile.scala 76:16:@35484.4]
  assign regs_76_io_in = 64'h0; // @[RegFile.scala 75:16:@35483.4]
  assign regs_76_io_reset = reset; // @[RegFile.scala 78:19:@35487.4]
  assign regs_76_io_enable = 1'h1; // @[RegFile.scala 74:20:@35481.4]
  assign regs_77_clock = clock; // @[:@35490.4]
  assign regs_77_reset = io_reset; // @[:@35491.4 RegFile.scala 76:16:@35498.4]
  assign regs_77_io_in = 64'h0; // @[RegFile.scala 75:16:@35497.4]
  assign regs_77_io_reset = reset; // @[RegFile.scala 78:19:@35501.4]
  assign regs_77_io_enable = 1'h1; // @[RegFile.scala 74:20:@35495.4]
  assign regs_78_clock = clock; // @[:@35504.4]
  assign regs_78_reset = io_reset; // @[:@35505.4 RegFile.scala 76:16:@35512.4]
  assign regs_78_io_in = 64'h0; // @[RegFile.scala 75:16:@35511.4]
  assign regs_78_io_reset = reset; // @[RegFile.scala 78:19:@35515.4]
  assign regs_78_io_enable = 1'h1; // @[RegFile.scala 74:20:@35509.4]
  assign regs_79_clock = clock; // @[:@35518.4]
  assign regs_79_reset = io_reset; // @[:@35519.4 RegFile.scala 76:16:@35526.4]
  assign regs_79_io_in = 64'h0; // @[RegFile.scala 75:16:@35525.4]
  assign regs_79_io_reset = reset; // @[RegFile.scala 78:19:@35529.4]
  assign regs_79_io_enable = 1'h1; // @[RegFile.scala 74:20:@35523.4]
  assign regs_80_clock = clock; // @[:@35532.4]
  assign regs_80_reset = io_reset; // @[:@35533.4 RegFile.scala 76:16:@35540.4]
  assign regs_80_io_in = 64'h0; // @[RegFile.scala 75:16:@35539.4]
  assign regs_80_io_reset = reset; // @[RegFile.scala 78:19:@35543.4]
  assign regs_80_io_enable = 1'h1; // @[RegFile.scala 74:20:@35537.4]
  assign regs_81_clock = clock; // @[:@35546.4]
  assign regs_81_reset = io_reset; // @[:@35547.4 RegFile.scala 76:16:@35554.4]
  assign regs_81_io_in = 64'h0; // @[RegFile.scala 75:16:@35553.4]
  assign regs_81_io_reset = reset; // @[RegFile.scala 78:19:@35557.4]
  assign regs_81_io_enable = 1'h1; // @[RegFile.scala 74:20:@35551.4]
  assign regs_82_clock = clock; // @[:@35560.4]
  assign regs_82_reset = io_reset; // @[:@35561.4 RegFile.scala 76:16:@35568.4]
  assign regs_82_io_in = 64'h0; // @[RegFile.scala 75:16:@35567.4]
  assign regs_82_io_reset = reset; // @[RegFile.scala 78:19:@35571.4]
  assign regs_82_io_enable = 1'h1; // @[RegFile.scala 74:20:@35565.4]
  assign regs_83_clock = clock; // @[:@35574.4]
  assign regs_83_reset = io_reset; // @[:@35575.4 RegFile.scala 76:16:@35582.4]
  assign regs_83_io_in = 64'h0; // @[RegFile.scala 75:16:@35581.4]
  assign regs_83_io_reset = reset; // @[RegFile.scala 78:19:@35585.4]
  assign regs_83_io_enable = 1'h1; // @[RegFile.scala 74:20:@35579.4]
  assign regs_84_clock = clock; // @[:@35588.4]
  assign regs_84_reset = io_reset; // @[:@35589.4 RegFile.scala 76:16:@35596.4]
  assign regs_84_io_in = 64'h0; // @[RegFile.scala 75:16:@35595.4]
  assign regs_84_io_reset = reset; // @[RegFile.scala 78:19:@35599.4]
  assign regs_84_io_enable = 1'h1; // @[RegFile.scala 74:20:@35593.4]
  assign regs_85_clock = clock; // @[:@35602.4]
  assign regs_85_reset = io_reset; // @[:@35603.4 RegFile.scala 76:16:@35610.4]
  assign regs_85_io_in = 64'h0; // @[RegFile.scala 75:16:@35609.4]
  assign regs_85_io_reset = reset; // @[RegFile.scala 78:19:@35613.4]
  assign regs_85_io_enable = 1'h1; // @[RegFile.scala 74:20:@35607.4]
  assign regs_86_clock = clock; // @[:@35616.4]
  assign regs_86_reset = io_reset; // @[:@35617.4 RegFile.scala 76:16:@35624.4]
  assign regs_86_io_in = 64'h0; // @[RegFile.scala 75:16:@35623.4]
  assign regs_86_io_reset = reset; // @[RegFile.scala 78:19:@35627.4]
  assign regs_86_io_enable = 1'h1; // @[RegFile.scala 74:20:@35621.4]
  assign regs_87_clock = clock; // @[:@35630.4]
  assign regs_87_reset = io_reset; // @[:@35631.4 RegFile.scala 76:16:@35638.4]
  assign regs_87_io_in = 64'h0; // @[RegFile.scala 75:16:@35637.4]
  assign regs_87_io_reset = reset; // @[RegFile.scala 78:19:@35641.4]
  assign regs_87_io_enable = 1'h1; // @[RegFile.scala 74:20:@35635.4]
  assign regs_88_clock = clock; // @[:@35644.4]
  assign regs_88_reset = io_reset; // @[:@35645.4 RegFile.scala 76:16:@35652.4]
  assign regs_88_io_in = 64'h0; // @[RegFile.scala 75:16:@35651.4]
  assign regs_88_io_reset = reset; // @[RegFile.scala 78:19:@35655.4]
  assign regs_88_io_enable = 1'h1; // @[RegFile.scala 74:20:@35649.4]
  assign regs_89_clock = clock; // @[:@35658.4]
  assign regs_89_reset = io_reset; // @[:@35659.4 RegFile.scala 76:16:@35666.4]
  assign regs_89_io_in = 64'h0; // @[RegFile.scala 75:16:@35665.4]
  assign regs_89_io_reset = reset; // @[RegFile.scala 78:19:@35669.4]
  assign regs_89_io_enable = 1'h1; // @[RegFile.scala 74:20:@35663.4]
  assign regs_90_clock = clock; // @[:@35672.4]
  assign regs_90_reset = io_reset; // @[:@35673.4 RegFile.scala 76:16:@35680.4]
  assign regs_90_io_in = 64'h0; // @[RegFile.scala 75:16:@35679.4]
  assign regs_90_io_reset = reset; // @[RegFile.scala 78:19:@35683.4]
  assign regs_90_io_enable = 1'h1; // @[RegFile.scala 74:20:@35677.4]
  assign regs_91_clock = clock; // @[:@35686.4]
  assign regs_91_reset = io_reset; // @[:@35687.4 RegFile.scala 76:16:@35694.4]
  assign regs_91_io_in = 64'h0; // @[RegFile.scala 75:16:@35693.4]
  assign regs_91_io_reset = reset; // @[RegFile.scala 78:19:@35697.4]
  assign regs_91_io_enable = 1'h1; // @[RegFile.scala 74:20:@35691.4]
  assign regs_92_clock = clock; // @[:@35700.4]
  assign regs_92_reset = io_reset; // @[:@35701.4 RegFile.scala 76:16:@35708.4]
  assign regs_92_io_in = 64'h0; // @[RegFile.scala 75:16:@35707.4]
  assign regs_92_io_reset = reset; // @[RegFile.scala 78:19:@35711.4]
  assign regs_92_io_enable = 1'h1; // @[RegFile.scala 74:20:@35705.4]
  assign regs_93_clock = clock; // @[:@35714.4]
  assign regs_93_reset = io_reset; // @[:@35715.4 RegFile.scala 76:16:@35722.4]
  assign regs_93_io_in = 64'h0; // @[RegFile.scala 75:16:@35721.4]
  assign regs_93_io_reset = reset; // @[RegFile.scala 78:19:@35725.4]
  assign regs_93_io_enable = 1'h1; // @[RegFile.scala 74:20:@35719.4]
  assign regs_94_clock = clock; // @[:@35728.4]
  assign regs_94_reset = io_reset; // @[:@35729.4 RegFile.scala 76:16:@35736.4]
  assign regs_94_io_in = 64'h0; // @[RegFile.scala 75:16:@35735.4]
  assign regs_94_io_reset = reset; // @[RegFile.scala 78:19:@35739.4]
  assign regs_94_io_enable = 1'h1; // @[RegFile.scala 74:20:@35733.4]
  assign regs_95_clock = clock; // @[:@35742.4]
  assign regs_95_reset = io_reset; // @[:@35743.4 RegFile.scala 76:16:@35750.4]
  assign regs_95_io_in = 64'h0; // @[RegFile.scala 75:16:@35749.4]
  assign regs_95_io_reset = reset; // @[RegFile.scala 78:19:@35753.4]
  assign regs_95_io_enable = 1'h1; // @[RegFile.scala 74:20:@35747.4]
  assign regs_96_clock = clock; // @[:@35756.4]
  assign regs_96_reset = io_reset; // @[:@35757.4 RegFile.scala 76:16:@35764.4]
  assign regs_96_io_in = 64'h0; // @[RegFile.scala 75:16:@35763.4]
  assign regs_96_io_reset = reset; // @[RegFile.scala 78:19:@35767.4]
  assign regs_96_io_enable = 1'h1; // @[RegFile.scala 74:20:@35761.4]
  assign regs_97_clock = clock; // @[:@35770.4]
  assign regs_97_reset = io_reset; // @[:@35771.4 RegFile.scala 76:16:@35778.4]
  assign regs_97_io_in = 64'h0; // @[RegFile.scala 75:16:@35777.4]
  assign regs_97_io_reset = reset; // @[RegFile.scala 78:19:@35781.4]
  assign regs_97_io_enable = 1'h1; // @[RegFile.scala 74:20:@35775.4]
  assign regs_98_clock = clock; // @[:@35784.4]
  assign regs_98_reset = io_reset; // @[:@35785.4 RegFile.scala 76:16:@35792.4]
  assign regs_98_io_in = 64'h0; // @[RegFile.scala 75:16:@35791.4]
  assign regs_98_io_reset = reset; // @[RegFile.scala 78:19:@35795.4]
  assign regs_98_io_enable = 1'h1; // @[RegFile.scala 74:20:@35789.4]
  assign regs_99_clock = clock; // @[:@35798.4]
  assign regs_99_reset = io_reset; // @[:@35799.4 RegFile.scala 76:16:@35806.4]
  assign regs_99_io_in = 64'h0; // @[RegFile.scala 75:16:@35805.4]
  assign regs_99_io_reset = reset; // @[RegFile.scala 78:19:@35809.4]
  assign regs_99_io_enable = 1'h1; // @[RegFile.scala 74:20:@35803.4]
  assign regs_100_clock = clock; // @[:@35812.4]
  assign regs_100_reset = io_reset; // @[:@35813.4 RegFile.scala 76:16:@35820.4]
  assign regs_100_io_in = 64'h0; // @[RegFile.scala 75:16:@35819.4]
  assign regs_100_io_reset = reset; // @[RegFile.scala 78:19:@35823.4]
  assign regs_100_io_enable = 1'h1; // @[RegFile.scala 74:20:@35817.4]
  assign regs_101_clock = clock; // @[:@35826.4]
  assign regs_101_reset = io_reset; // @[:@35827.4 RegFile.scala 76:16:@35834.4]
  assign regs_101_io_in = 64'h0; // @[RegFile.scala 75:16:@35833.4]
  assign regs_101_io_reset = reset; // @[RegFile.scala 78:19:@35837.4]
  assign regs_101_io_enable = 1'h1; // @[RegFile.scala 74:20:@35831.4]
  assign regs_102_clock = clock; // @[:@35840.4]
  assign regs_102_reset = io_reset; // @[:@35841.4 RegFile.scala 76:16:@35848.4]
  assign regs_102_io_in = 64'h0; // @[RegFile.scala 75:16:@35847.4]
  assign regs_102_io_reset = reset; // @[RegFile.scala 78:19:@35851.4]
  assign regs_102_io_enable = 1'h1; // @[RegFile.scala 74:20:@35845.4]
  assign regs_103_clock = clock; // @[:@35854.4]
  assign regs_103_reset = io_reset; // @[:@35855.4 RegFile.scala 76:16:@35862.4]
  assign regs_103_io_in = 64'h0; // @[RegFile.scala 75:16:@35861.4]
  assign regs_103_io_reset = reset; // @[RegFile.scala 78:19:@35865.4]
  assign regs_103_io_enable = 1'h1; // @[RegFile.scala 74:20:@35859.4]
  assign regs_104_clock = clock; // @[:@35868.4]
  assign regs_104_reset = io_reset; // @[:@35869.4 RegFile.scala 76:16:@35876.4]
  assign regs_104_io_in = 64'h0; // @[RegFile.scala 75:16:@35875.4]
  assign regs_104_io_reset = reset; // @[RegFile.scala 78:19:@35879.4]
  assign regs_104_io_enable = 1'h1; // @[RegFile.scala 74:20:@35873.4]
  assign regs_105_clock = clock; // @[:@35882.4]
  assign regs_105_reset = io_reset; // @[:@35883.4 RegFile.scala 76:16:@35890.4]
  assign regs_105_io_in = 64'h0; // @[RegFile.scala 75:16:@35889.4]
  assign regs_105_io_reset = reset; // @[RegFile.scala 78:19:@35893.4]
  assign regs_105_io_enable = 1'h1; // @[RegFile.scala 74:20:@35887.4]
  assign regs_106_clock = clock; // @[:@35896.4]
  assign regs_106_reset = io_reset; // @[:@35897.4 RegFile.scala 76:16:@35904.4]
  assign regs_106_io_in = 64'h0; // @[RegFile.scala 75:16:@35903.4]
  assign regs_106_io_reset = reset; // @[RegFile.scala 78:19:@35907.4]
  assign regs_106_io_enable = 1'h1; // @[RegFile.scala 74:20:@35901.4]
  assign regs_107_clock = clock; // @[:@35910.4]
  assign regs_107_reset = io_reset; // @[:@35911.4 RegFile.scala 76:16:@35918.4]
  assign regs_107_io_in = 64'h0; // @[RegFile.scala 75:16:@35917.4]
  assign regs_107_io_reset = reset; // @[RegFile.scala 78:19:@35921.4]
  assign regs_107_io_enable = 1'h1; // @[RegFile.scala 74:20:@35915.4]
  assign regs_108_clock = clock; // @[:@35924.4]
  assign regs_108_reset = io_reset; // @[:@35925.4 RegFile.scala 76:16:@35932.4]
  assign regs_108_io_in = 64'h0; // @[RegFile.scala 75:16:@35931.4]
  assign regs_108_io_reset = reset; // @[RegFile.scala 78:19:@35935.4]
  assign regs_108_io_enable = 1'h1; // @[RegFile.scala 74:20:@35929.4]
  assign regs_109_clock = clock; // @[:@35938.4]
  assign regs_109_reset = io_reset; // @[:@35939.4 RegFile.scala 76:16:@35946.4]
  assign regs_109_io_in = 64'h0; // @[RegFile.scala 75:16:@35945.4]
  assign regs_109_io_reset = reset; // @[RegFile.scala 78:19:@35949.4]
  assign regs_109_io_enable = 1'h1; // @[RegFile.scala 74:20:@35943.4]
  assign regs_110_clock = clock; // @[:@35952.4]
  assign regs_110_reset = io_reset; // @[:@35953.4 RegFile.scala 76:16:@35960.4]
  assign regs_110_io_in = 64'h0; // @[RegFile.scala 75:16:@35959.4]
  assign regs_110_io_reset = reset; // @[RegFile.scala 78:19:@35963.4]
  assign regs_110_io_enable = 1'h1; // @[RegFile.scala 74:20:@35957.4]
  assign regs_111_clock = clock; // @[:@35966.4]
  assign regs_111_reset = io_reset; // @[:@35967.4 RegFile.scala 76:16:@35974.4]
  assign regs_111_io_in = 64'h0; // @[RegFile.scala 75:16:@35973.4]
  assign regs_111_io_reset = reset; // @[RegFile.scala 78:19:@35977.4]
  assign regs_111_io_enable = 1'h1; // @[RegFile.scala 74:20:@35971.4]
  assign regs_112_clock = clock; // @[:@35980.4]
  assign regs_112_reset = io_reset; // @[:@35981.4 RegFile.scala 76:16:@35988.4]
  assign regs_112_io_in = 64'h0; // @[RegFile.scala 75:16:@35987.4]
  assign regs_112_io_reset = reset; // @[RegFile.scala 78:19:@35991.4]
  assign regs_112_io_enable = 1'h1; // @[RegFile.scala 74:20:@35985.4]
  assign regs_113_clock = clock; // @[:@35994.4]
  assign regs_113_reset = io_reset; // @[:@35995.4 RegFile.scala 76:16:@36002.4]
  assign regs_113_io_in = 64'h0; // @[RegFile.scala 75:16:@36001.4]
  assign regs_113_io_reset = reset; // @[RegFile.scala 78:19:@36005.4]
  assign regs_113_io_enable = 1'h1; // @[RegFile.scala 74:20:@35999.4]
  assign regs_114_clock = clock; // @[:@36008.4]
  assign regs_114_reset = io_reset; // @[:@36009.4 RegFile.scala 76:16:@36016.4]
  assign regs_114_io_in = 64'h0; // @[RegFile.scala 75:16:@36015.4]
  assign regs_114_io_reset = reset; // @[RegFile.scala 78:19:@36019.4]
  assign regs_114_io_enable = 1'h1; // @[RegFile.scala 74:20:@36013.4]
  assign regs_115_clock = clock; // @[:@36022.4]
  assign regs_115_reset = io_reset; // @[:@36023.4 RegFile.scala 76:16:@36030.4]
  assign regs_115_io_in = 64'h0; // @[RegFile.scala 75:16:@36029.4]
  assign regs_115_io_reset = reset; // @[RegFile.scala 78:19:@36033.4]
  assign regs_115_io_enable = 1'h1; // @[RegFile.scala 74:20:@36027.4]
  assign regs_116_clock = clock; // @[:@36036.4]
  assign regs_116_reset = io_reset; // @[:@36037.4 RegFile.scala 76:16:@36044.4]
  assign regs_116_io_in = 64'h0; // @[RegFile.scala 75:16:@36043.4]
  assign regs_116_io_reset = reset; // @[RegFile.scala 78:19:@36047.4]
  assign regs_116_io_enable = 1'h1; // @[RegFile.scala 74:20:@36041.4]
  assign regs_117_clock = clock; // @[:@36050.4]
  assign regs_117_reset = io_reset; // @[:@36051.4 RegFile.scala 76:16:@36058.4]
  assign regs_117_io_in = 64'h0; // @[RegFile.scala 75:16:@36057.4]
  assign regs_117_io_reset = reset; // @[RegFile.scala 78:19:@36061.4]
  assign regs_117_io_enable = 1'h1; // @[RegFile.scala 74:20:@36055.4]
  assign regs_118_clock = clock; // @[:@36064.4]
  assign regs_118_reset = io_reset; // @[:@36065.4 RegFile.scala 76:16:@36072.4]
  assign regs_118_io_in = 64'h0; // @[RegFile.scala 75:16:@36071.4]
  assign regs_118_io_reset = reset; // @[RegFile.scala 78:19:@36075.4]
  assign regs_118_io_enable = 1'h1; // @[RegFile.scala 74:20:@36069.4]
  assign regs_119_clock = clock; // @[:@36078.4]
  assign regs_119_reset = io_reset; // @[:@36079.4 RegFile.scala 76:16:@36086.4]
  assign regs_119_io_in = 64'h0; // @[RegFile.scala 75:16:@36085.4]
  assign regs_119_io_reset = reset; // @[RegFile.scala 78:19:@36089.4]
  assign regs_119_io_enable = 1'h1; // @[RegFile.scala 74:20:@36083.4]
  assign regs_120_clock = clock; // @[:@36092.4]
  assign regs_120_reset = io_reset; // @[:@36093.4 RegFile.scala 76:16:@36100.4]
  assign regs_120_io_in = 64'h0; // @[RegFile.scala 75:16:@36099.4]
  assign regs_120_io_reset = reset; // @[RegFile.scala 78:19:@36103.4]
  assign regs_120_io_enable = 1'h1; // @[RegFile.scala 74:20:@36097.4]
  assign regs_121_clock = clock; // @[:@36106.4]
  assign regs_121_reset = io_reset; // @[:@36107.4 RegFile.scala 76:16:@36114.4]
  assign regs_121_io_in = 64'h0; // @[RegFile.scala 75:16:@36113.4]
  assign regs_121_io_reset = reset; // @[RegFile.scala 78:19:@36117.4]
  assign regs_121_io_enable = 1'h1; // @[RegFile.scala 74:20:@36111.4]
  assign regs_122_clock = clock; // @[:@36120.4]
  assign regs_122_reset = io_reset; // @[:@36121.4 RegFile.scala 76:16:@36128.4]
  assign regs_122_io_in = 64'h0; // @[RegFile.scala 75:16:@36127.4]
  assign regs_122_io_reset = reset; // @[RegFile.scala 78:19:@36131.4]
  assign regs_122_io_enable = 1'h1; // @[RegFile.scala 74:20:@36125.4]
  assign regs_123_clock = clock; // @[:@36134.4]
  assign regs_123_reset = io_reset; // @[:@36135.4 RegFile.scala 76:16:@36142.4]
  assign regs_123_io_in = 64'h0; // @[RegFile.scala 75:16:@36141.4]
  assign regs_123_io_reset = reset; // @[RegFile.scala 78:19:@36145.4]
  assign regs_123_io_enable = 1'h1; // @[RegFile.scala 74:20:@36139.4]
  assign regs_124_clock = clock; // @[:@36148.4]
  assign regs_124_reset = io_reset; // @[:@36149.4 RegFile.scala 76:16:@36156.4]
  assign regs_124_io_in = 64'h0; // @[RegFile.scala 75:16:@36155.4]
  assign regs_124_io_reset = reset; // @[RegFile.scala 78:19:@36159.4]
  assign regs_124_io_enable = 1'h1; // @[RegFile.scala 74:20:@36153.4]
  assign regs_125_clock = clock; // @[:@36162.4]
  assign regs_125_reset = io_reset; // @[:@36163.4 RegFile.scala 76:16:@36170.4]
  assign regs_125_io_in = 64'h0; // @[RegFile.scala 75:16:@36169.4]
  assign regs_125_io_reset = reset; // @[RegFile.scala 78:19:@36173.4]
  assign regs_125_io_enable = 1'h1; // @[RegFile.scala 74:20:@36167.4]
  assign regs_126_clock = clock; // @[:@36176.4]
  assign regs_126_reset = io_reset; // @[:@36177.4 RegFile.scala 76:16:@36184.4]
  assign regs_126_io_in = 64'h0; // @[RegFile.scala 75:16:@36183.4]
  assign regs_126_io_reset = reset; // @[RegFile.scala 78:19:@36187.4]
  assign regs_126_io_enable = 1'h1; // @[RegFile.scala 74:20:@36181.4]
  assign regs_127_clock = clock; // @[:@36190.4]
  assign regs_127_reset = io_reset; // @[:@36191.4 RegFile.scala 76:16:@36198.4]
  assign regs_127_io_in = 64'h0; // @[RegFile.scala 75:16:@36197.4]
  assign regs_127_io_reset = reset; // @[RegFile.scala 78:19:@36201.4]
  assign regs_127_io_enable = 1'h1; // @[RegFile.scala 74:20:@36195.4]
  assign regs_128_clock = clock; // @[:@36204.4]
  assign regs_128_reset = io_reset; // @[:@36205.4 RegFile.scala 76:16:@36212.4]
  assign regs_128_io_in = 64'h0; // @[RegFile.scala 75:16:@36211.4]
  assign regs_128_io_reset = reset; // @[RegFile.scala 78:19:@36215.4]
  assign regs_128_io_enable = 1'h1; // @[RegFile.scala 74:20:@36209.4]
  assign regs_129_clock = clock; // @[:@36218.4]
  assign regs_129_reset = io_reset; // @[:@36219.4 RegFile.scala 76:16:@36226.4]
  assign regs_129_io_in = 64'h0; // @[RegFile.scala 75:16:@36225.4]
  assign regs_129_io_reset = reset; // @[RegFile.scala 78:19:@36229.4]
  assign regs_129_io_enable = 1'h1; // @[RegFile.scala 74:20:@36223.4]
  assign regs_130_clock = clock; // @[:@36232.4]
  assign regs_130_reset = io_reset; // @[:@36233.4 RegFile.scala 76:16:@36240.4]
  assign regs_130_io_in = 64'h0; // @[RegFile.scala 75:16:@36239.4]
  assign regs_130_io_reset = reset; // @[RegFile.scala 78:19:@36243.4]
  assign regs_130_io_enable = 1'h1; // @[RegFile.scala 74:20:@36237.4]
  assign regs_131_clock = clock; // @[:@36246.4]
  assign regs_131_reset = io_reset; // @[:@36247.4 RegFile.scala 76:16:@36254.4]
  assign regs_131_io_in = 64'h0; // @[RegFile.scala 75:16:@36253.4]
  assign regs_131_io_reset = reset; // @[RegFile.scala 78:19:@36257.4]
  assign regs_131_io_enable = 1'h1; // @[RegFile.scala 74:20:@36251.4]
  assign regs_132_clock = clock; // @[:@36260.4]
  assign regs_132_reset = io_reset; // @[:@36261.4 RegFile.scala 76:16:@36268.4]
  assign regs_132_io_in = 64'h0; // @[RegFile.scala 75:16:@36267.4]
  assign regs_132_io_reset = reset; // @[RegFile.scala 78:19:@36271.4]
  assign regs_132_io_enable = 1'h1; // @[RegFile.scala 74:20:@36265.4]
  assign regs_133_clock = clock; // @[:@36274.4]
  assign regs_133_reset = io_reset; // @[:@36275.4 RegFile.scala 76:16:@36282.4]
  assign regs_133_io_in = 64'h0; // @[RegFile.scala 75:16:@36281.4]
  assign regs_133_io_reset = reset; // @[RegFile.scala 78:19:@36285.4]
  assign regs_133_io_enable = 1'h1; // @[RegFile.scala 74:20:@36279.4]
  assign regs_134_clock = clock; // @[:@36288.4]
  assign regs_134_reset = io_reset; // @[:@36289.4 RegFile.scala 76:16:@36296.4]
  assign regs_134_io_in = 64'h0; // @[RegFile.scala 75:16:@36295.4]
  assign regs_134_io_reset = reset; // @[RegFile.scala 78:19:@36299.4]
  assign regs_134_io_enable = 1'h1; // @[RegFile.scala 74:20:@36293.4]
  assign regs_135_clock = clock; // @[:@36302.4]
  assign regs_135_reset = io_reset; // @[:@36303.4 RegFile.scala 76:16:@36310.4]
  assign regs_135_io_in = 64'h0; // @[RegFile.scala 75:16:@36309.4]
  assign regs_135_io_reset = reset; // @[RegFile.scala 78:19:@36313.4]
  assign regs_135_io_enable = 1'h1; // @[RegFile.scala 74:20:@36307.4]
  assign regs_136_clock = clock; // @[:@36316.4]
  assign regs_136_reset = io_reset; // @[:@36317.4 RegFile.scala 76:16:@36324.4]
  assign regs_136_io_in = 64'h0; // @[RegFile.scala 75:16:@36323.4]
  assign regs_136_io_reset = reset; // @[RegFile.scala 78:19:@36327.4]
  assign regs_136_io_enable = 1'h1; // @[RegFile.scala 74:20:@36321.4]
  assign regs_137_clock = clock; // @[:@36330.4]
  assign regs_137_reset = io_reset; // @[:@36331.4 RegFile.scala 76:16:@36338.4]
  assign regs_137_io_in = 64'h0; // @[RegFile.scala 75:16:@36337.4]
  assign regs_137_io_reset = reset; // @[RegFile.scala 78:19:@36341.4]
  assign regs_137_io_enable = 1'h1; // @[RegFile.scala 74:20:@36335.4]
  assign regs_138_clock = clock; // @[:@36344.4]
  assign regs_138_reset = io_reset; // @[:@36345.4 RegFile.scala 76:16:@36352.4]
  assign regs_138_io_in = 64'h0; // @[RegFile.scala 75:16:@36351.4]
  assign regs_138_io_reset = reset; // @[RegFile.scala 78:19:@36355.4]
  assign regs_138_io_enable = 1'h1; // @[RegFile.scala 74:20:@36349.4]
  assign regs_139_clock = clock; // @[:@36358.4]
  assign regs_139_reset = io_reset; // @[:@36359.4 RegFile.scala 76:16:@36366.4]
  assign regs_139_io_in = 64'h0; // @[RegFile.scala 75:16:@36365.4]
  assign regs_139_io_reset = reset; // @[RegFile.scala 78:19:@36369.4]
  assign regs_139_io_enable = 1'h1; // @[RegFile.scala 74:20:@36363.4]
  assign regs_140_clock = clock; // @[:@36372.4]
  assign regs_140_reset = io_reset; // @[:@36373.4 RegFile.scala 76:16:@36380.4]
  assign regs_140_io_in = 64'h0; // @[RegFile.scala 75:16:@36379.4]
  assign regs_140_io_reset = reset; // @[RegFile.scala 78:19:@36383.4]
  assign regs_140_io_enable = 1'h1; // @[RegFile.scala 74:20:@36377.4]
  assign regs_141_clock = clock; // @[:@36386.4]
  assign regs_141_reset = io_reset; // @[:@36387.4 RegFile.scala 76:16:@36394.4]
  assign regs_141_io_in = 64'h0; // @[RegFile.scala 75:16:@36393.4]
  assign regs_141_io_reset = reset; // @[RegFile.scala 78:19:@36397.4]
  assign regs_141_io_enable = 1'h1; // @[RegFile.scala 74:20:@36391.4]
  assign regs_142_clock = clock; // @[:@36400.4]
  assign regs_142_reset = io_reset; // @[:@36401.4 RegFile.scala 76:16:@36408.4]
  assign regs_142_io_in = 64'h0; // @[RegFile.scala 75:16:@36407.4]
  assign regs_142_io_reset = reset; // @[RegFile.scala 78:19:@36411.4]
  assign regs_142_io_enable = 1'h1; // @[RegFile.scala 74:20:@36405.4]
  assign regs_143_clock = clock; // @[:@36414.4]
  assign regs_143_reset = io_reset; // @[:@36415.4 RegFile.scala 76:16:@36422.4]
  assign regs_143_io_in = 64'h0; // @[RegFile.scala 75:16:@36421.4]
  assign regs_143_io_reset = reset; // @[RegFile.scala 78:19:@36425.4]
  assign regs_143_io_enable = 1'h1; // @[RegFile.scala 74:20:@36419.4]
  assign regs_144_clock = clock; // @[:@36428.4]
  assign regs_144_reset = io_reset; // @[:@36429.4 RegFile.scala 76:16:@36436.4]
  assign regs_144_io_in = 64'h0; // @[RegFile.scala 75:16:@36435.4]
  assign regs_144_io_reset = reset; // @[RegFile.scala 78:19:@36439.4]
  assign regs_144_io_enable = 1'h1; // @[RegFile.scala 74:20:@36433.4]
  assign regs_145_clock = clock; // @[:@36442.4]
  assign regs_145_reset = io_reset; // @[:@36443.4 RegFile.scala 76:16:@36450.4]
  assign regs_145_io_in = 64'h0; // @[RegFile.scala 75:16:@36449.4]
  assign regs_145_io_reset = reset; // @[RegFile.scala 78:19:@36453.4]
  assign regs_145_io_enable = 1'h1; // @[RegFile.scala 74:20:@36447.4]
  assign regs_146_clock = clock; // @[:@36456.4]
  assign regs_146_reset = io_reset; // @[:@36457.4 RegFile.scala 76:16:@36464.4]
  assign regs_146_io_in = 64'h0; // @[RegFile.scala 75:16:@36463.4]
  assign regs_146_io_reset = reset; // @[RegFile.scala 78:19:@36467.4]
  assign regs_146_io_enable = 1'h1; // @[RegFile.scala 74:20:@36461.4]
  assign regs_147_clock = clock; // @[:@36470.4]
  assign regs_147_reset = io_reset; // @[:@36471.4 RegFile.scala 76:16:@36478.4]
  assign regs_147_io_in = 64'h0; // @[RegFile.scala 75:16:@36477.4]
  assign regs_147_io_reset = reset; // @[RegFile.scala 78:19:@36481.4]
  assign regs_147_io_enable = 1'h1; // @[RegFile.scala 74:20:@36475.4]
  assign regs_148_clock = clock; // @[:@36484.4]
  assign regs_148_reset = io_reset; // @[:@36485.4 RegFile.scala 76:16:@36492.4]
  assign regs_148_io_in = 64'h0; // @[RegFile.scala 75:16:@36491.4]
  assign regs_148_io_reset = reset; // @[RegFile.scala 78:19:@36495.4]
  assign regs_148_io_enable = 1'h1; // @[RegFile.scala 74:20:@36489.4]
  assign regs_149_clock = clock; // @[:@36498.4]
  assign regs_149_reset = io_reset; // @[:@36499.4 RegFile.scala 76:16:@36506.4]
  assign regs_149_io_in = 64'h0; // @[RegFile.scala 75:16:@36505.4]
  assign regs_149_io_reset = reset; // @[RegFile.scala 78:19:@36509.4]
  assign regs_149_io_enable = 1'h1; // @[RegFile.scala 74:20:@36503.4]
  assign regs_150_clock = clock; // @[:@36512.4]
  assign regs_150_reset = io_reset; // @[:@36513.4 RegFile.scala 76:16:@36520.4]
  assign regs_150_io_in = 64'h0; // @[RegFile.scala 75:16:@36519.4]
  assign regs_150_io_reset = reset; // @[RegFile.scala 78:19:@36523.4]
  assign regs_150_io_enable = 1'h1; // @[RegFile.scala 74:20:@36517.4]
  assign regs_151_clock = clock; // @[:@36526.4]
  assign regs_151_reset = io_reset; // @[:@36527.4 RegFile.scala 76:16:@36534.4]
  assign regs_151_io_in = 64'h0; // @[RegFile.scala 75:16:@36533.4]
  assign regs_151_io_reset = reset; // @[RegFile.scala 78:19:@36537.4]
  assign regs_151_io_enable = 1'h1; // @[RegFile.scala 74:20:@36531.4]
  assign regs_152_clock = clock; // @[:@36540.4]
  assign regs_152_reset = io_reset; // @[:@36541.4 RegFile.scala 76:16:@36548.4]
  assign regs_152_io_in = 64'h0; // @[RegFile.scala 75:16:@36547.4]
  assign regs_152_io_reset = reset; // @[RegFile.scala 78:19:@36551.4]
  assign regs_152_io_enable = 1'h1; // @[RegFile.scala 74:20:@36545.4]
  assign regs_153_clock = clock; // @[:@36554.4]
  assign regs_153_reset = io_reset; // @[:@36555.4 RegFile.scala 76:16:@36562.4]
  assign regs_153_io_in = 64'h0; // @[RegFile.scala 75:16:@36561.4]
  assign regs_153_io_reset = reset; // @[RegFile.scala 78:19:@36565.4]
  assign regs_153_io_enable = 1'h1; // @[RegFile.scala 74:20:@36559.4]
  assign regs_154_clock = clock; // @[:@36568.4]
  assign regs_154_reset = io_reset; // @[:@36569.4 RegFile.scala 76:16:@36576.4]
  assign regs_154_io_in = 64'h0; // @[RegFile.scala 75:16:@36575.4]
  assign regs_154_io_reset = reset; // @[RegFile.scala 78:19:@36579.4]
  assign regs_154_io_enable = 1'h1; // @[RegFile.scala 74:20:@36573.4]
  assign regs_155_clock = clock; // @[:@36582.4]
  assign regs_155_reset = io_reset; // @[:@36583.4 RegFile.scala 76:16:@36590.4]
  assign regs_155_io_in = 64'h0; // @[RegFile.scala 75:16:@36589.4]
  assign regs_155_io_reset = reset; // @[RegFile.scala 78:19:@36593.4]
  assign regs_155_io_enable = 1'h1; // @[RegFile.scala 74:20:@36587.4]
  assign regs_156_clock = clock; // @[:@36596.4]
  assign regs_156_reset = io_reset; // @[:@36597.4 RegFile.scala 76:16:@36604.4]
  assign regs_156_io_in = 64'h0; // @[RegFile.scala 75:16:@36603.4]
  assign regs_156_io_reset = reset; // @[RegFile.scala 78:19:@36607.4]
  assign regs_156_io_enable = 1'h1; // @[RegFile.scala 74:20:@36601.4]
  assign regs_157_clock = clock; // @[:@36610.4]
  assign regs_157_reset = io_reset; // @[:@36611.4 RegFile.scala 76:16:@36618.4]
  assign regs_157_io_in = 64'h0; // @[RegFile.scala 75:16:@36617.4]
  assign regs_157_io_reset = reset; // @[RegFile.scala 78:19:@36621.4]
  assign regs_157_io_enable = 1'h1; // @[RegFile.scala 74:20:@36615.4]
  assign regs_158_clock = clock; // @[:@36624.4]
  assign regs_158_reset = io_reset; // @[:@36625.4 RegFile.scala 76:16:@36632.4]
  assign regs_158_io_in = 64'h0; // @[RegFile.scala 75:16:@36631.4]
  assign regs_158_io_reset = reset; // @[RegFile.scala 78:19:@36635.4]
  assign regs_158_io_enable = 1'h1; // @[RegFile.scala 74:20:@36629.4]
  assign regs_159_clock = clock; // @[:@36638.4]
  assign regs_159_reset = io_reset; // @[:@36639.4 RegFile.scala 76:16:@36646.4]
  assign regs_159_io_in = 64'h0; // @[RegFile.scala 75:16:@36645.4]
  assign regs_159_io_reset = reset; // @[RegFile.scala 78:19:@36649.4]
  assign regs_159_io_enable = 1'h1; // @[RegFile.scala 74:20:@36643.4]
  assign regs_160_clock = clock; // @[:@36652.4]
  assign regs_160_reset = io_reset; // @[:@36653.4 RegFile.scala 76:16:@36660.4]
  assign regs_160_io_in = 64'h0; // @[RegFile.scala 75:16:@36659.4]
  assign regs_160_io_reset = reset; // @[RegFile.scala 78:19:@36663.4]
  assign regs_160_io_enable = 1'h1; // @[RegFile.scala 74:20:@36657.4]
  assign regs_161_clock = clock; // @[:@36666.4]
  assign regs_161_reset = io_reset; // @[:@36667.4 RegFile.scala 76:16:@36674.4]
  assign regs_161_io_in = 64'h0; // @[RegFile.scala 75:16:@36673.4]
  assign regs_161_io_reset = reset; // @[RegFile.scala 78:19:@36677.4]
  assign regs_161_io_enable = 1'h1; // @[RegFile.scala 74:20:@36671.4]
  assign regs_162_clock = clock; // @[:@36680.4]
  assign regs_162_reset = io_reset; // @[:@36681.4 RegFile.scala 76:16:@36688.4]
  assign regs_162_io_in = 64'h0; // @[RegFile.scala 75:16:@36687.4]
  assign regs_162_io_reset = reset; // @[RegFile.scala 78:19:@36691.4]
  assign regs_162_io_enable = 1'h1; // @[RegFile.scala 74:20:@36685.4]
  assign regs_163_clock = clock; // @[:@36694.4]
  assign regs_163_reset = io_reset; // @[:@36695.4 RegFile.scala 76:16:@36702.4]
  assign regs_163_io_in = 64'h0; // @[RegFile.scala 75:16:@36701.4]
  assign regs_163_io_reset = reset; // @[RegFile.scala 78:19:@36705.4]
  assign regs_163_io_enable = 1'h1; // @[RegFile.scala 74:20:@36699.4]
  assign regs_164_clock = clock; // @[:@36708.4]
  assign regs_164_reset = io_reset; // @[:@36709.4 RegFile.scala 76:16:@36716.4]
  assign regs_164_io_in = 64'h0; // @[RegFile.scala 75:16:@36715.4]
  assign regs_164_io_reset = reset; // @[RegFile.scala 78:19:@36719.4]
  assign regs_164_io_enable = 1'h1; // @[RegFile.scala 74:20:@36713.4]
  assign regs_165_clock = clock; // @[:@36722.4]
  assign regs_165_reset = io_reset; // @[:@36723.4 RegFile.scala 76:16:@36730.4]
  assign regs_165_io_in = 64'h0; // @[RegFile.scala 75:16:@36729.4]
  assign regs_165_io_reset = reset; // @[RegFile.scala 78:19:@36733.4]
  assign regs_165_io_enable = 1'h1; // @[RegFile.scala 74:20:@36727.4]
  assign regs_166_clock = clock; // @[:@36736.4]
  assign regs_166_reset = io_reset; // @[:@36737.4 RegFile.scala 76:16:@36744.4]
  assign regs_166_io_in = 64'h0; // @[RegFile.scala 75:16:@36743.4]
  assign regs_166_io_reset = reset; // @[RegFile.scala 78:19:@36747.4]
  assign regs_166_io_enable = 1'h1; // @[RegFile.scala 74:20:@36741.4]
  assign regs_167_clock = clock; // @[:@36750.4]
  assign regs_167_reset = io_reset; // @[:@36751.4 RegFile.scala 76:16:@36758.4]
  assign regs_167_io_in = 64'h0; // @[RegFile.scala 75:16:@36757.4]
  assign regs_167_io_reset = reset; // @[RegFile.scala 78:19:@36761.4]
  assign regs_167_io_enable = 1'h1; // @[RegFile.scala 74:20:@36755.4]
  assign regs_168_clock = clock; // @[:@36764.4]
  assign regs_168_reset = io_reset; // @[:@36765.4 RegFile.scala 76:16:@36772.4]
  assign regs_168_io_in = 64'h0; // @[RegFile.scala 75:16:@36771.4]
  assign regs_168_io_reset = reset; // @[RegFile.scala 78:19:@36775.4]
  assign regs_168_io_enable = 1'h1; // @[RegFile.scala 74:20:@36769.4]
  assign regs_169_clock = clock; // @[:@36778.4]
  assign regs_169_reset = io_reset; // @[:@36779.4 RegFile.scala 76:16:@36786.4]
  assign regs_169_io_in = 64'h0; // @[RegFile.scala 75:16:@36785.4]
  assign regs_169_io_reset = reset; // @[RegFile.scala 78:19:@36789.4]
  assign regs_169_io_enable = 1'h1; // @[RegFile.scala 74:20:@36783.4]
  assign regs_170_clock = clock; // @[:@36792.4]
  assign regs_170_reset = io_reset; // @[:@36793.4 RegFile.scala 76:16:@36800.4]
  assign regs_170_io_in = 64'h0; // @[RegFile.scala 75:16:@36799.4]
  assign regs_170_io_reset = reset; // @[RegFile.scala 78:19:@36803.4]
  assign regs_170_io_enable = 1'h1; // @[RegFile.scala 74:20:@36797.4]
  assign regs_171_clock = clock; // @[:@36806.4]
  assign regs_171_reset = io_reset; // @[:@36807.4 RegFile.scala 76:16:@36814.4]
  assign regs_171_io_in = 64'h0; // @[RegFile.scala 75:16:@36813.4]
  assign regs_171_io_reset = reset; // @[RegFile.scala 78:19:@36817.4]
  assign regs_171_io_enable = 1'h1; // @[RegFile.scala 74:20:@36811.4]
  assign regs_172_clock = clock; // @[:@36820.4]
  assign regs_172_reset = io_reset; // @[:@36821.4 RegFile.scala 76:16:@36828.4]
  assign regs_172_io_in = 64'h0; // @[RegFile.scala 75:16:@36827.4]
  assign regs_172_io_reset = reset; // @[RegFile.scala 78:19:@36831.4]
  assign regs_172_io_enable = 1'h1; // @[RegFile.scala 74:20:@36825.4]
  assign regs_173_clock = clock; // @[:@36834.4]
  assign regs_173_reset = io_reset; // @[:@36835.4 RegFile.scala 76:16:@36842.4]
  assign regs_173_io_in = 64'h0; // @[RegFile.scala 75:16:@36841.4]
  assign regs_173_io_reset = reset; // @[RegFile.scala 78:19:@36845.4]
  assign regs_173_io_enable = 1'h1; // @[RegFile.scala 74:20:@36839.4]
  assign regs_174_clock = clock; // @[:@36848.4]
  assign regs_174_reset = io_reset; // @[:@36849.4 RegFile.scala 76:16:@36856.4]
  assign regs_174_io_in = 64'h0; // @[RegFile.scala 75:16:@36855.4]
  assign regs_174_io_reset = reset; // @[RegFile.scala 78:19:@36859.4]
  assign regs_174_io_enable = 1'h1; // @[RegFile.scala 74:20:@36853.4]
  assign regs_175_clock = clock; // @[:@36862.4]
  assign regs_175_reset = io_reset; // @[:@36863.4 RegFile.scala 76:16:@36870.4]
  assign regs_175_io_in = 64'h0; // @[RegFile.scala 75:16:@36869.4]
  assign regs_175_io_reset = reset; // @[RegFile.scala 78:19:@36873.4]
  assign regs_175_io_enable = 1'h1; // @[RegFile.scala 74:20:@36867.4]
  assign regs_176_clock = clock; // @[:@36876.4]
  assign regs_176_reset = io_reset; // @[:@36877.4 RegFile.scala 76:16:@36884.4]
  assign regs_176_io_in = 64'h0; // @[RegFile.scala 75:16:@36883.4]
  assign regs_176_io_reset = reset; // @[RegFile.scala 78:19:@36887.4]
  assign regs_176_io_enable = 1'h1; // @[RegFile.scala 74:20:@36881.4]
  assign regs_177_clock = clock; // @[:@36890.4]
  assign regs_177_reset = io_reset; // @[:@36891.4 RegFile.scala 76:16:@36898.4]
  assign regs_177_io_in = 64'h0; // @[RegFile.scala 75:16:@36897.4]
  assign regs_177_io_reset = reset; // @[RegFile.scala 78:19:@36901.4]
  assign regs_177_io_enable = 1'h1; // @[RegFile.scala 74:20:@36895.4]
  assign regs_178_clock = clock; // @[:@36904.4]
  assign regs_178_reset = io_reset; // @[:@36905.4 RegFile.scala 76:16:@36912.4]
  assign regs_178_io_in = 64'h0; // @[RegFile.scala 75:16:@36911.4]
  assign regs_178_io_reset = reset; // @[RegFile.scala 78:19:@36915.4]
  assign regs_178_io_enable = 1'h1; // @[RegFile.scala 74:20:@36909.4]
  assign regs_179_clock = clock; // @[:@36918.4]
  assign regs_179_reset = io_reset; // @[:@36919.4 RegFile.scala 76:16:@36926.4]
  assign regs_179_io_in = 64'h0; // @[RegFile.scala 75:16:@36925.4]
  assign regs_179_io_reset = reset; // @[RegFile.scala 78:19:@36929.4]
  assign regs_179_io_enable = 1'h1; // @[RegFile.scala 74:20:@36923.4]
  assign regs_180_clock = clock; // @[:@36932.4]
  assign regs_180_reset = io_reset; // @[:@36933.4 RegFile.scala 76:16:@36940.4]
  assign regs_180_io_in = 64'h0; // @[RegFile.scala 75:16:@36939.4]
  assign regs_180_io_reset = reset; // @[RegFile.scala 78:19:@36943.4]
  assign regs_180_io_enable = 1'h1; // @[RegFile.scala 74:20:@36937.4]
  assign regs_181_clock = clock; // @[:@36946.4]
  assign regs_181_reset = io_reset; // @[:@36947.4 RegFile.scala 76:16:@36954.4]
  assign regs_181_io_in = 64'h0; // @[RegFile.scala 75:16:@36953.4]
  assign regs_181_io_reset = reset; // @[RegFile.scala 78:19:@36957.4]
  assign regs_181_io_enable = 1'h1; // @[RegFile.scala 74:20:@36951.4]
  assign regs_182_clock = clock; // @[:@36960.4]
  assign regs_182_reset = io_reset; // @[:@36961.4 RegFile.scala 76:16:@36968.4]
  assign regs_182_io_in = 64'h0; // @[RegFile.scala 75:16:@36967.4]
  assign regs_182_io_reset = reset; // @[RegFile.scala 78:19:@36971.4]
  assign regs_182_io_enable = 1'h1; // @[RegFile.scala 74:20:@36965.4]
  assign regs_183_clock = clock; // @[:@36974.4]
  assign regs_183_reset = io_reset; // @[:@36975.4 RegFile.scala 76:16:@36982.4]
  assign regs_183_io_in = 64'h0; // @[RegFile.scala 75:16:@36981.4]
  assign regs_183_io_reset = reset; // @[RegFile.scala 78:19:@36985.4]
  assign regs_183_io_enable = 1'h1; // @[RegFile.scala 74:20:@36979.4]
  assign regs_184_clock = clock; // @[:@36988.4]
  assign regs_184_reset = io_reset; // @[:@36989.4 RegFile.scala 76:16:@36996.4]
  assign regs_184_io_in = 64'h0; // @[RegFile.scala 75:16:@36995.4]
  assign regs_184_io_reset = reset; // @[RegFile.scala 78:19:@36999.4]
  assign regs_184_io_enable = 1'h1; // @[RegFile.scala 74:20:@36993.4]
  assign regs_185_clock = clock; // @[:@37002.4]
  assign regs_185_reset = io_reset; // @[:@37003.4 RegFile.scala 76:16:@37010.4]
  assign regs_185_io_in = 64'h0; // @[RegFile.scala 75:16:@37009.4]
  assign regs_185_io_reset = reset; // @[RegFile.scala 78:19:@37013.4]
  assign regs_185_io_enable = 1'h1; // @[RegFile.scala 74:20:@37007.4]
  assign regs_186_clock = clock; // @[:@37016.4]
  assign regs_186_reset = io_reset; // @[:@37017.4 RegFile.scala 76:16:@37024.4]
  assign regs_186_io_in = 64'h0; // @[RegFile.scala 75:16:@37023.4]
  assign regs_186_io_reset = reset; // @[RegFile.scala 78:19:@37027.4]
  assign regs_186_io_enable = 1'h1; // @[RegFile.scala 74:20:@37021.4]
  assign regs_187_clock = clock; // @[:@37030.4]
  assign regs_187_reset = io_reset; // @[:@37031.4 RegFile.scala 76:16:@37038.4]
  assign regs_187_io_in = 64'h0; // @[RegFile.scala 75:16:@37037.4]
  assign regs_187_io_reset = reset; // @[RegFile.scala 78:19:@37041.4]
  assign regs_187_io_enable = 1'h1; // @[RegFile.scala 74:20:@37035.4]
  assign regs_188_clock = clock; // @[:@37044.4]
  assign regs_188_reset = io_reset; // @[:@37045.4 RegFile.scala 76:16:@37052.4]
  assign regs_188_io_in = 64'h0; // @[RegFile.scala 75:16:@37051.4]
  assign regs_188_io_reset = reset; // @[RegFile.scala 78:19:@37055.4]
  assign regs_188_io_enable = 1'h1; // @[RegFile.scala 74:20:@37049.4]
  assign regs_189_clock = clock; // @[:@37058.4]
  assign regs_189_reset = io_reset; // @[:@37059.4 RegFile.scala 76:16:@37066.4]
  assign regs_189_io_in = 64'h0; // @[RegFile.scala 75:16:@37065.4]
  assign regs_189_io_reset = reset; // @[RegFile.scala 78:19:@37069.4]
  assign regs_189_io_enable = 1'h1; // @[RegFile.scala 74:20:@37063.4]
  assign regs_190_clock = clock; // @[:@37072.4]
  assign regs_190_reset = io_reset; // @[:@37073.4 RegFile.scala 76:16:@37080.4]
  assign regs_190_io_in = 64'h0; // @[RegFile.scala 75:16:@37079.4]
  assign regs_190_io_reset = reset; // @[RegFile.scala 78:19:@37083.4]
  assign regs_190_io_enable = 1'h1; // @[RegFile.scala 74:20:@37077.4]
  assign regs_191_clock = clock; // @[:@37086.4]
  assign regs_191_reset = io_reset; // @[:@37087.4 RegFile.scala 76:16:@37094.4]
  assign regs_191_io_in = 64'h0; // @[RegFile.scala 75:16:@37093.4]
  assign regs_191_io_reset = reset; // @[RegFile.scala 78:19:@37097.4]
  assign regs_191_io_enable = 1'h1; // @[RegFile.scala 74:20:@37091.4]
  assign regs_192_clock = clock; // @[:@37100.4]
  assign regs_192_reset = io_reset; // @[:@37101.4 RegFile.scala 76:16:@37108.4]
  assign regs_192_io_in = 64'h0; // @[RegFile.scala 75:16:@37107.4]
  assign regs_192_io_reset = reset; // @[RegFile.scala 78:19:@37111.4]
  assign regs_192_io_enable = 1'h1; // @[RegFile.scala 74:20:@37105.4]
  assign regs_193_clock = clock; // @[:@37114.4]
  assign regs_193_reset = io_reset; // @[:@37115.4 RegFile.scala 76:16:@37122.4]
  assign regs_193_io_in = 64'h0; // @[RegFile.scala 75:16:@37121.4]
  assign regs_193_io_reset = reset; // @[RegFile.scala 78:19:@37125.4]
  assign regs_193_io_enable = 1'h1; // @[RegFile.scala 74:20:@37119.4]
  assign regs_194_clock = clock; // @[:@37128.4]
  assign regs_194_reset = io_reset; // @[:@37129.4 RegFile.scala 76:16:@37136.4]
  assign regs_194_io_in = 64'h0; // @[RegFile.scala 75:16:@37135.4]
  assign regs_194_io_reset = reset; // @[RegFile.scala 78:19:@37139.4]
  assign regs_194_io_enable = 1'h1; // @[RegFile.scala 74:20:@37133.4]
  assign regs_195_clock = clock; // @[:@37142.4]
  assign regs_195_reset = io_reset; // @[:@37143.4 RegFile.scala 76:16:@37150.4]
  assign regs_195_io_in = 64'h0; // @[RegFile.scala 75:16:@37149.4]
  assign regs_195_io_reset = reset; // @[RegFile.scala 78:19:@37153.4]
  assign regs_195_io_enable = 1'h1; // @[RegFile.scala 74:20:@37147.4]
  assign regs_196_clock = clock; // @[:@37156.4]
  assign regs_196_reset = io_reset; // @[:@37157.4 RegFile.scala 76:16:@37164.4]
  assign regs_196_io_in = 64'h0; // @[RegFile.scala 75:16:@37163.4]
  assign regs_196_io_reset = reset; // @[RegFile.scala 78:19:@37167.4]
  assign regs_196_io_enable = 1'h1; // @[RegFile.scala 74:20:@37161.4]
  assign regs_197_clock = clock; // @[:@37170.4]
  assign regs_197_reset = io_reset; // @[:@37171.4 RegFile.scala 76:16:@37178.4]
  assign regs_197_io_in = 64'h0; // @[RegFile.scala 75:16:@37177.4]
  assign regs_197_io_reset = reset; // @[RegFile.scala 78:19:@37181.4]
  assign regs_197_io_enable = 1'h1; // @[RegFile.scala 74:20:@37175.4]
  assign regs_198_clock = clock; // @[:@37184.4]
  assign regs_198_reset = io_reset; // @[:@37185.4 RegFile.scala 76:16:@37192.4]
  assign regs_198_io_in = 64'h0; // @[RegFile.scala 75:16:@37191.4]
  assign regs_198_io_reset = reset; // @[RegFile.scala 78:19:@37195.4]
  assign regs_198_io_enable = 1'h1; // @[RegFile.scala 74:20:@37189.4]
  assign regs_199_clock = clock; // @[:@37198.4]
  assign regs_199_reset = io_reset; // @[:@37199.4 RegFile.scala 76:16:@37206.4]
  assign regs_199_io_in = 64'h0; // @[RegFile.scala 75:16:@37205.4]
  assign regs_199_io_reset = reset; // @[RegFile.scala 78:19:@37209.4]
  assign regs_199_io_enable = 1'h1; // @[RegFile.scala 74:20:@37203.4]
  assign regs_200_clock = clock; // @[:@37212.4]
  assign regs_200_reset = io_reset; // @[:@37213.4 RegFile.scala 76:16:@37220.4]
  assign regs_200_io_in = 64'h0; // @[RegFile.scala 75:16:@37219.4]
  assign regs_200_io_reset = reset; // @[RegFile.scala 78:19:@37223.4]
  assign regs_200_io_enable = 1'h1; // @[RegFile.scala 74:20:@37217.4]
  assign regs_201_clock = clock; // @[:@37226.4]
  assign regs_201_reset = io_reset; // @[:@37227.4 RegFile.scala 76:16:@37234.4]
  assign regs_201_io_in = 64'h0; // @[RegFile.scala 75:16:@37233.4]
  assign regs_201_io_reset = reset; // @[RegFile.scala 78:19:@37237.4]
  assign regs_201_io_enable = 1'h1; // @[RegFile.scala 74:20:@37231.4]
  assign regs_202_clock = clock; // @[:@37240.4]
  assign regs_202_reset = io_reset; // @[:@37241.4 RegFile.scala 76:16:@37248.4]
  assign regs_202_io_in = 64'h0; // @[RegFile.scala 75:16:@37247.4]
  assign regs_202_io_reset = reset; // @[RegFile.scala 78:19:@37251.4]
  assign regs_202_io_enable = 1'h1; // @[RegFile.scala 74:20:@37245.4]
  assign regs_203_clock = clock; // @[:@37254.4]
  assign regs_203_reset = io_reset; // @[:@37255.4 RegFile.scala 76:16:@37262.4]
  assign regs_203_io_in = 64'h0; // @[RegFile.scala 75:16:@37261.4]
  assign regs_203_io_reset = reset; // @[RegFile.scala 78:19:@37265.4]
  assign regs_203_io_enable = 1'h1; // @[RegFile.scala 74:20:@37259.4]
  assign regs_204_clock = clock; // @[:@37268.4]
  assign regs_204_reset = io_reset; // @[:@37269.4 RegFile.scala 76:16:@37276.4]
  assign regs_204_io_in = 64'h0; // @[RegFile.scala 75:16:@37275.4]
  assign regs_204_io_reset = reset; // @[RegFile.scala 78:19:@37279.4]
  assign regs_204_io_enable = 1'h1; // @[RegFile.scala 74:20:@37273.4]
  assign regs_205_clock = clock; // @[:@37282.4]
  assign regs_205_reset = io_reset; // @[:@37283.4 RegFile.scala 76:16:@37290.4]
  assign regs_205_io_in = 64'h0; // @[RegFile.scala 75:16:@37289.4]
  assign regs_205_io_reset = reset; // @[RegFile.scala 78:19:@37293.4]
  assign regs_205_io_enable = 1'h1; // @[RegFile.scala 74:20:@37287.4]
  assign regs_206_clock = clock; // @[:@37296.4]
  assign regs_206_reset = io_reset; // @[:@37297.4 RegFile.scala 76:16:@37304.4]
  assign regs_206_io_in = 64'h0; // @[RegFile.scala 75:16:@37303.4]
  assign regs_206_io_reset = reset; // @[RegFile.scala 78:19:@37307.4]
  assign regs_206_io_enable = 1'h1; // @[RegFile.scala 74:20:@37301.4]
  assign regs_207_clock = clock; // @[:@37310.4]
  assign regs_207_reset = io_reset; // @[:@37311.4 RegFile.scala 76:16:@37318.4]
  assign regs_207_io_in = 64'h0; // @[RegFile.scala 75:16:@37317.4]
  assign regs_207_io_reset = reset; // @[RegFile.scala 78:19:@37321.4]
  assign regs_207_io_enable = 1'h1; // @[RegFile.scala 74:20:@37315.4]
  assign regs_208_clock = clock; // @[:@37324.4]
  assign regs_208_reset = io_reset; // @[:@37325.4 RegFile.scala 76:16:@37332.4]
  assign regs_208_io_in = 64'h0; // @[RegFile.scala 75:16:@37331.4]
  assign regs_208_io_reset = reset; // @[RegFile.scala 78:19:@37335.4]
  assign regs_208_io_enable = 1'h1; // @[RegFile.scala 74:20:@37329.4]
  assign regs_209_clock = clock; // @[:@37338.4]
  assign regs_209_reset = io_reset; // @[:@37339.4 RegFile.scala 76:16:@37346.4]
  assign regs_209_io_in = 64'h0; // @[RegFile.scala 75:16:@37345.4]
  assign regs_209_io_reset = reset; // @[RegFile.scala 78:19:@37349.4]
  assign regs_209_io_enable = 1'h1; // @[RegFile.scala 74:20:@37343.4]
  assign regs_210_clock = clock; // @[:@37352.4]
  assign regs_210_reset = io_reset; // @[:@37353.4 RegFile.scala 76:16:@37360.4]
  assign regs_210_io_in = 64'h0; // @[RegFile.scala 75:16:@37359.4]
  assign regs_210_io_reset = reset; // @[RegFile.scala 78:19:@37363.4]
  assign regs_210_io_enable = 1'h1; // @[RegFile.scala 74:20:@37357.4]
  assign regs_211_clock = clock; // @[:@37366.4]
  assign regs_211_reset = io_reset; // @[:@37367.4 RegFile.scala 76:16:@37374.4]
  assign regs_211_io_in = 64'h0; // @[RegFile.scala 75:16:@37373.4]
  assign regs_211_io_reset = reset; // @[RegFile.scala 78:19:@37377.4]
  assign regs_211_io_enable = 1'h1; // @[RegFile.scala 74:20:@37371.4]
  assign regs_212_clock = clock; // @[:@37380.4]
  assign regs_212_reset = io_reset; // @[:@37381.4 RegFile.scala 76:16:@37388.4]
  assign regs_212_io_in = 64'h0; // @[RegFile.scala 75:16:@37387.4]
  assign regs_212_io_reset = reset; // @[RegFile.scala 78:19:@37391.4]
  assign regs_212_io_enable = 1'h1; // @[RegFile.scala 74:20:@37385.4]
  assign regs_213_clock = clock; // @[:@37394.4]
  assign regs_213_reset = io_reset; // @[:@37395.4 RegFile.scala 76:16:@37402.4]
  assign regs_213_io_in = 64'h0; // @[RegFile.scala 75:16:@37401.4]
  assign regs_213_io_reset = reset; // @[RegFile.scala 78:19:@37405.4]
  assign regs_213_io_enable = 1'h1; // @[RegFile.scala 74:20:@37399.4]
  assign regs_214_clock = clock; // @[:@37408.4]
  assign regs_214_reset = io_reset; // @[:@37409.4 RegFile.scala 76:16:@37416.4]
  assign regs_214_io_in = 64'h0; // @[RegFile.scala 75:16:@37415.4]
  assign regs_214_io_reset = reset; // @[RegFile.scala 78:19:@37419.4]
  assign regs_214_io_enable = 1'h1; // @[RegFile.scala 74:20:@37413.4]
  assign regs_215_clock = clock; // @[:@37422.4]
  assign regs_215_reset = io_reset; // @[:@37423.4 RegFile.scala 76:16:@37430.4]
  assign regs_215_io_in = 64'h0; // @[RegFile.scala 75:16:@37429.4]
  assign regs_215_io_reset = reset; // @[RegFile.scala 78:19:@37433.4]
  assign regs_215_io_enable = 1'h1; // @[RegFile.scala 74:20:@37427.4]
  assign regs_216_clock = clock; // @[:@37436.4]
  assign regs_216_reset = io_reset; // @[:@37437.4 RegFile.scala 76:16:@37444.4]
  assign regs_216_io_in = 64'h0; // @[RegFile.scala 75:16:@37443.4]
  assign regs_216_io_reset = reset; // @[RegFile.scala 78:19:@37447.4]
  assign regs_216_io_enable = 1'h1; // @[RegFile.scala 74:20:@37441.4]
  assign regs_217_clock = clock; // @[:@37450.4]
  assign regs_217_reset = io_reset; // @[:@37451.4 RegFile.scala 76:16:@37458.4]
  assign regs_217_io_in = 64'h0; // @[RegFile.scala 75:16:@37457.4]
  assign regs_217_io_reset = reset; // @[RegFile.scala 78:19:@37461.4]
  assign regs_217_io_enable = 1'h1; // @[RegFile.scala 74:20:@37455.4]
  assign regs_218_clock = clock; // @[:@37464.4]
  assign regs_218_reset = io_reset; // @[:@37465.4 RegFile.scala 76:16:@37472.4]
  assign regs_218_io_in = 64'h0; // @[RegFile.scala 75:16:@37471.4]
  assign regs_218_io_reset = reset; // @[RegFile.scala 78:19:@37475.4]
  assign regs_218_io_enable = 1'h1; // @[RegFile.scala 74:20:@37469.4]
  assign regs_219_clock = clock; // @[:@37478.4]
  assign regs_219_reset = io_reset; // @[:@37479.4 RegFile.scala 76:16:@37486.4]
  assign regs_219_io_in = 64'h0; // @[RegFile.scala 75:16:@37485.4]
  assign regs_219_io_reset = reset; // @[RegFile.scala 78:19:@37489.4]
  assign regs_219_io_enable = 1'h1; // @[RegFile.scala 74:20:@37483.4]
  assign regs_220_clock = clock; // @[:@37492.4]
  assign regs_220_reset = io_reset; // @[:@37493.4 RegFile.scala 76:16:@37500.4]
  assign regs_220_io_in = 64'h0; // @[RegFile.scala 75:16:@37499.4]
  assign regs_220_io_reset = reset; // @[RegFile.scala 78:19:@37503.4]
  assign regs_220_io_enable = 1'h1; // @[RegFile.scala 74:20:@37497.4]
  assign regs_221_clock = clock; // @[:@37506.4]
  assign regs_221_reset = io_reset; // @[:@37507.4 RegFile.scala 76:16:@37514.4]
  assign regs_221_io_in = 64'h0; // @[RegFile.scala 75:16:@37513.4]
  assign regs_221_io_reset = reset; // @[RegFile.scala 78:19:@37517.4]
  assign regs_221_io_enable = 1'h1; // @[RegFile.scala 74:20:@37511.4]
  assign regs_222_clock = clock; // @[:@37520.4]
  assign regs_222_reset = io_reset; // @[:@37521.4 RegFile.scala 76:16:@37528.4]
  assign regs_222_io_in = 64'h0; // @[RegFile.scala 75:16:@37527.4]
  assign regs_222_io_reset = reset; // @[RegFile.scala 78:19:@37531.4]
  assign regs_222_io_enable = 1'h1; // @[RegFile.scala 74:20:@37525.4]
  assign regs_223_clock = clock; // @[:@37534.4]
  assign regs_223_reset = io_reset; // @[:@37535.4 RegFile.scala 76:16:@37542.4]
  assign regs_223_io_in = 64'h0; // @[RegFile.scala 75:16:@37541.4]
  assign regs_223_io_reset = reset; // @[RegFile.scala 78:19:@37545.4]
  assign regs_223_io_enable = 1'h1; // @[RegFile.scala 74:20:@37539.4]
  assign regs_224_clock = clock; // @[:@37548.4]
  assign regs_224_reset = io_reset; // @[:@37549.4 RegFile.scala 76:16:@37556.4]
  assign regs_224_io_in = 64'h0; // @[RegFile.scala 75:16:@37555.4]
  assign regs_224_io_reset = reset; // @[RegFile.scala 78:19:@37559.4]
  assign regs_224_io_enable = 1'h1; // @[RegFile.scala 74:20:@37553.4]
  assign regs_225_clock = clock; // @[:@37562.4]
  assign regs_225_reset = io_reset; // @[:@37563.4 RegFile.scala 76:16:@37570.4]
  assign regs_225_io_in = 64'h0; // @[RegFile.scala 75:16:@37569.4]
  assign regs_225_io_reset = reset; // @[RegFile.scala 78:19:@37573.4]
  assign regs_225_io_enable = 1'h1; // @[RegFile.scala 74:20:@37567.4]
  assign regs_226_clock = clock; // @[:@37576.4]
  assign regs_226_reset = io_reset; // @[:@37577.4 RegFile.scala 76:16:@37584.4]
  assign regs_226_io_in = 64'h0; // @[RegFile.scala 75:16:@37583.4]
  assign regs_226_io_reset = reset; // @[RegFile.scala 78:19:@37587.4]
  assign regs_226_io_enable = 1'h1; // @[RegFile.scala 74:20:@37581.4]
  assign regs_227_clock = clock; // @[:@37590.4]
  assign regs_227_reset = io_reset; // @[:@37591.4 RegFile.scala 76:16:@37598.4]
  assign regs_227_io_in = 64'h0; // @[RegFile.scala 75:16:@37597.4]
  assign regs_227_io_reset = reset; // @[RegFile.scala 78:19:@37601.4]
  assign regs_227_io_enable = 1'h1; // @[RegFile.scala 74:20:@37595.4]
  assign regs_228_clock = clock; // @[:@37604.4]
  assign regs_228_reset = io_reset; // @[:@37605.4 RegFile.scala 76:16:@37612.4]
  assign regs_228_io_in = 64'h0; // @[RegFile.scala 75:16:@37611.4]
  assign regs_228_io_reset = reset; // @[RegFile.scala 78:19:@37615.4]
  assign regs_228_io_enable = 1'h1; // @[RegFile.scala 74:20:@37609.4]
  assign regs_229_clock = clock; // @[:@37618.4]
  assign regs_229_reset = io_reset; // @[:@37619.4 RegFile.scala 76:16:@37626.4]
  assign regs_229_io_in = 64'h0; // @[RegFile.scala 75:16:@37625.4]
  assign regs_229_io_reset = reset; // @[RegFile.scala 78:19:@37629.4]
  assign regs_229_io_enable = 1'h1; // @[RegFile.scala 74:20:@37623.4]
  assign regs_230_clock = clock; // @[:@37632.4]
  assign regs_230_reset = io_reset; // @[:@37633.4 RegFile.scala 76:16:@37640.4]
  assign regs_230_io_in = 64'h0; // @[RegFile.scala 75:16:@37639.4]
  assign regs_230_io_reset = reset; // @[RegFile.scala 78:19:@37643.4]
  assign regs_230_io_enable = 1'h1; // @[RegFile.scala 74:20:@37637.4]
  assign regs_231_clock = clock; // @[:@37646.4]
  assign regs_231_reset = io_reset; // @[:@37647.4 RegFile.scala 76:16:@37654.4]
  assign regs_231_io_in = 64'h0; // @[RegFile.scala 75:16:@37653.4]
  assign regs_231_io_reset = reset; // @[RegFile.scala 78:19:@37657.4]
  assign regs_231_io_enable = 1'h1; // @[RegFile.scala 74:20:@37651.4]
  assign regs_232_clock = clock; // @[:@37660.4]
  assign regs_232_reset = io_reset; // @[:@37661.4 RegFile.scala 76:16:@37668.4]
  assign regs_232_io_in = 64'h0; // @[RegFile.scala 75:16:@37667.4]
  assign regs_232_io_reset = reset; // @[RegFile.scala 78:19:@37671.4]
  assign regs_232_io_enable = 1'h1; // @[RegFile.scala 74:20:@37665.4]
  assign regs_233_clock = clock; // @[:@37674.4]
  assign regs_233_reset = io_reset; // @[:@37675.4 RegFile.scala 76:16:@37682.4]
  assign regs_233_io_in = 64'h0; // @[RegFile.scala 75:16:@37681.4]
  assign regs_233_io_reset = reset; // @[RegFile.scala 78:19:@37685.4]
  assign regs_233_io_enable = 1'h1; // @[RegFile.scala 74:20:@37679.4]
  assign regs_234_clock = clock; // @[:@37688.4]
  assign regs_234_reset = io_reset; // @[:@37689.4 RegFile.scala 76:16:@37696.4]
  assign regs_234_io_in = 64'h0; // @[RegFile.scala 75:16:@37695.4]
  assign regs_234_io_reset = reset; // @[RegFile.scala 78:19:@37699.4]
  assign regs_234_io_enable = 1'h1; // @[RegFile.scala 74:20:@37693.4]
  assign regs_235_clock = clock; // @[:@37702.4]
  assign regs_235_reset = io_reset; // @[:@37703.4 RegFile.scala 76:16:@37710.4]
  assign regs_235_io_in = 64'h0; // @[RegFile.scala 75:16:@37709.4]
  assign regs_235_io_reset = reset; // @[RegFile.scala 78:19:@37713.4]
  assign regs_235_io_enable = 1'h1; // @[RegFile.scala 74:20:@37707.4]
  assign regs_236_clock = clock; // @[:@37716.4]
  assign regs_236_reset = io_reset; // @[:@37717.4 RegFile.scala 76:16:@37724.4]
  assign regs_236_io_in = 64'h0; // @[RegFile.scala 75:16:@37723.4]
  assign regs_236_io_reset = reset; // @[RegFile.scala 78:19:@37727.4]
  assign regs_236_io_enable = 1'h1; // @[RegFile.scala 74:20:@37721.4]
  assign regs_237_clock = clock; // @[:@37730.4]
  assign regs_237_reset = io_reset; // @[:@37731.4 RegFile.scala 76:16:@37738.4]
  assign regs_237_io_in = 64'h0; // @[RegFile.scala 75:16:@37737.4]
  assign regs_237_io_reset = reset; // @[RegFile.scala 78:19:@37741.4]
  assign regs_237_io_enable = 1'h1; // @[RegFile.scala 74:20:@37735.4]
  assign regs_238_clock = clock; // @[:@37744.4]
  assign regs_238_reset = io_reset; // @[:@37745.4 RegFile.scala 76:16:@37752.4]
  assign regs_238_io_in = 64'h0; // @[RegFile.scala 75:16:@37751.4]
  assign regs_238_io_reset = reset; // @[RegFile.scala 78:19:@37755.4]
  assign regs_238_io_enable = 1'h1; // @[RegFile.scala 74:20:@37749.4]
  assign regs_239_clock = clock; // @[:@37758.4]
  assign regs_239_reset = io_reset; // @[:@37759.4 RegFile.scala 76:16:@37766.4]
  assign regs_239_io_in = 64'h0; // @[RegFile.scala 75:16:@37765.4]
  assign regs_239_io_reset = reset; // @[RegFile.scala 78:19:@37769.4]
  assign regs_239_io_enable = 1'h1; // @[RegFile.scala 74:20:@37763.4]
  assign regs_240_clock = clock; // @[:@37772.4]
  assign regs_240_reset = io_reset; // @[:@37773.4 RegFile.scala 76:16:@37780.4]
  assign regs_240_io_in = 64'h0; // @[RegFile.scala 75:16:@37779.4]
  assign regs_240_io_reset = reset; // @[RegFile.scala 78:19:@37783.4]
  assign regs_240_io_enable = 1'h1; // @[RegFile.scala 74:20:@37777.4]
  assign regs_241_clock = clock; // @[:@37786.4]
  assign regs_241_reset = io_reset; // @[:@37787.4 RegFile.scala 76:16:@37794.4]
  assign regs_241_io_in = 64'h0; // @[RegFile.scala 75:16:@37793.4]
  assign regs_241_io_reset = reset; // @[RegFile.scala 78:19:@37797.4]
  assign regs_241_io_enable = 1'h1; // @[RegFile.scala 74:20:@37791.4]
  assign regs_242_clock = clock; // @[:@37800.4]
  assign regs_242_reset = io_reset; // @[:@37801.4 RegFile.scala 76:16:@37808.4]
  assign regs_242_io_in = 64'h0; // @[RegFile.scala 75:16:@37807.4]
  assign regs_242_io_reset = reset; // @[RegFile.scala 78:19:@37811.4]
  assign regs_242_io_enable = 1'h1; // @[RegFile.scala 74:20:@37805.4]
  assign regs_243_clock = clock; // @[:@37814.4]
  assign regs_243_reset = io_reset; // @[:@37815.4 RegFile.scala 76:16:@37822.4]
  assign regs_243_io_in = 64'h0; // @[RegFile.scala 75:16:@37821.4]
  assign regs_243_io_reset = reset; // @[RegFile.scala 78:19:@37825.4]
  assign regs_243_io_enable = 1'h1; // @[RegFile.scala 74:20:@37819.4]
  assign regs_244_clock = clock; // @[:@37828.4]
  assign regs_244_reset = io_reset; // @[:@37829.4 RegFile.scala 76:16:@37836.4]
  assign regs_244_io_in = 64'h0; // @[RegFile.scala 75:16:@37835.4]
  assign regs_244_io_reset = reset; // @[RegFile.scala 78:19:@37839.4]
  assign regs_244_io_enable = 1'h1; // @[RegFile.scala 74:20:@37833.4]
  assign regs_245_clock = clock; // @[:@37842.4]
  assign regs_245_reset = io_reset; // @[:@37843.4 RegFile.scala 76:16:@37850.4]
  assign regs_245_io_in = 64'h0; // @[RegFile.scala 75:16:@37849.4]
  assign regs_245_io_reset = reset; // @[RegFile.scala 78:19:@37853.4]
  assign regs_245_io_enable = 1'h1; // @[RegFile.scala 74:20:@37847.4]
  assign regs_246_clock = clock; // @[:@37856.4]
  assign regs_246_reset = io_reset; // @[:@37857.4 RegFile.scala 76:16:@37864.4]
  assign regs_246_io_in = 64'h0; // @[RegFile.scala 75:16:@37863.4]
  assign regs_246_io_reset = reset; // @[RegFile.scala 78:19:@37867.4]
  assign regs_246_io_enable = 1'h1; // @[RegFile.scala 74:20:@37861.4]
  assign regs_247_clock = clock; // @[:@37870.4]
  assign regs_247_reset = io_reset; // @[:@37871.4 RegFile.scala 76:16:@37878.4]
  assign regs_247_io_in = 64'h0; // @[RegFile.scala 75:16:@37877.4]
  assign regs_247_io_reset = reset; // @[RegFile.scala 78:19:@37881.4]
  assign regs_247_io_enable = 1'h1; // @[RegFile.scala 74:20:@37875.4]
  assign regs_248_clock = clock; // @[:@37884.4]
  assign regs_248_reset = io_reset; // @[:@37885.4 RegFile.scala 76:16:@37892.4]
  assign regs_248_io_in = 64'h0; // @[RegFile.scala 75:16:@37891.4]
  assign regs_248_io_reset = reset; // @[RegFile.scala 78:19:@37895.4]
  assign regs_248_io_enable = 1'h1; // @[RegFile.scala 74:20:@37889.4]
  assign regs_249_clock = clock; // @[:@37898.4]
  assign regs_249_reset = io_reset; // @[:@37899.4 RegFile.scala 76:16:@37906.4]
  assign regs_249_io_in = 64'h0; // @[RegFile.scala 75:16:@37905.4]
  assign regs_249_io_reset = reset; // @[RegFile.scala 78:19:@37909.4]
  assign regs_249_io_enable = 1'h1; // @[RegFile.scala 74:20:@37903.4]
  assign regs_250_clock = clock; // @[:@37912.4]
  assign regs_250_reset = io_reset; // @[:@37913.4 RegFile.scala 76:16:@37920.4]
  assign regs_250_io_in = 64'h0; // @[RegFile.scala 75:16:@37919.4]
  assign regs_250_io_reset = reset; // @[RegFile.scala 78:19:@37923.4]
  assign regs_250_io_enable = 1'h1; // @[RegFile.scala 74:20:@37917.4]
  assign regs_251_clock = clock; // @[:@37926.4]
  assign regs_251_reset = io_reset; // @[:@37927.4 RegFile.scala 76:16:@37934.4]
  assign regs_251_io_in = 64'h0; // @[RegFile.scala 75:16:@37933.4]
  assign regs_251_io_reset = reset; // @[RegFile.scala 78:19:@37937.4]
  assign regs_251_io_enable = 1'h1; // @[RegFile.scala 74:20:@37931.4]
  assign regs_252_clock = clock; // @[:@37940.4]
  assign regs_252_reset = io_reset; // @[:@37941.4 RegFile.scala 76:16:@37948.4]
  assign regs_252_io_in = 64'h0; // @[RegFile.scala 75:16:@37947.4]
  assign regs_252_io_reset = reset; // @[RegFile.scala 78:19:@37951.4]
  assign regs_252_io_enable = 1'h1; // @[RegFile.scala 74:20:@37945.4]
  assign regs_253_clock = clock; // @[:@37954.4]
  assign regs_253_reset = io_reset; // @[:@37955.4 RegFile.scala 76:16:@37962.4]
  assign regs_253_io_in = 64'h0; // @[RegFile.scala 75:16:@37961.4]
  assign regs_253_io_reset = reset; // @[RegFile.scala 78:19:@37965.4]
  assign regs_253_io_enable = 1'h1; // @[RegFile.scala 74:20:@37959.4]
  assign regs_254_clock = clock; // @[:@37968.4]
  assign regs_254_reset = io_reset; // @[:@37969.4 RegFile.scala 76:16:@37976.4]
  assign regs_254_io_in = 64'h0; // @[RegFile.scala 75:16:@37975.4]
  assign regs_254_io_reset = reset; // @[RegFile.scala 78:19:@37979.4]
  assign regs_254_io_enable = 1'h1; // @[RegFile.scala 74:20:@37973.4]
  assign regs_255_clock = clock; // @[:@37982.4]
  assign regs_255_reset = io_reset; // @[:@37983.4 RegFile.scala 76:16:@37990.4]
  assign regs_255_io_in = 64'h0; // @[RegFile.scala 75:16:@37989.4]
  assign regs_255_io_reset = reset; // @[RegFile.scala 78:19:@37993.4]
  assign regs_255_io_enable = 1'h1; // @[RegFile.scala 74:20:@37987.4]
  assign regs_256_clock = clock; // @[:@37996.4]
  assign regs_256_reset = io_reset; // @[:@37997.4 RegFile.scala 76:16:@38004.4]
  assign regs_256_io_in = 64'h0; // @[RegFile.scala 75:16:@38003.4]
  assign regs_256_io_reset = reset; // @[RegFile.scala 78:19:@38007.4]
  assign regs_256_io_enable = 1'h1; // @[RegFile.scala 74:20:@38001.4]
  assign regs_257_clock = clock; // @[:@38010.4]
  assign regs_257_reset = io_reset; // @[:@38011.4 RegFile.scala 76:16:@38018.4]
  assign regs_257_io_in = 64'h0; // @[RegFile.scala 75:16:@38017.4]
  assign regs_257_io_reset = reset; // @[RegFile.scala 78:19:@38021.4]
  assign regs_257_io_enable = 1'h1; // @[RegFile.scala 74:20:@38015.4]
  assign regs_258_clock = clock; // @[:@38024.4]
  assign regs_258_reset = io_reset; // @[:@38025.4 RegFile.scala 76:16:@38032.4]
  assign regs_258_io_in = 64'h0; // @[RegFile.scala 75:16:@38031.4]
  assign regs_258_io_reset = reset; // @[RegFile.scala 78:19:@38035.4]
  assign regs_258_io_enable = 1'h1; // @[RegFile.scala 74:20:@38029.4]
  assign regs_259_clock = clock; // @[:@38038.4]
  assign regs_259_reset = io_reset; // @[:@38039.4 RegFile.scala 76:16:@38046.4]
  assign regs_259_io_in = 64'h0; // @[RegFile.scala 75:16:@38045.4]
  assign regs_259_io_reset = reset; // @[RegFile.scala 78:19:@38049.4]
  assign regs_259_io_enable = 1'h1; // @[RegFile.scala 74:20:@38043.4]
  assign regs_260_clock = clock; // @[:@38052.4]
  assign regs_260_reset = io_reset; // @[:@38053.4 RegFile.scala 76:16:@38060.4]
  assign regs_260_io_in = 64'h0; // @[RegFile.scala 75:16:@38059.4]
  assign regs_260_io_reset = reset; // @[RegFile.scala 78:19:@38063.4]
  assign regs_260_io_enable = 1'h1; // @[RegFile.scala 74:20:@38057.4]
  assign regs_261_clock = clock; // @[:@38066.4]
  assign regs_261_reset = io_reset; // @[:@38067.4 RegFile.scala 76:16:@38074.4]
  assign regs_261_io_in = 64'h0; // @[RegFile.scala 75:16:@38073.4]
  assign regs_261_io_reset = reset; // @[RegFile.scala 78:19:@38077.4]
  assign regs_261_io_enable = 1'h1; // @[RegFile.scala 74:20:@38071.4]
  assign regs_262_clock = clock; // @[:@38080.4]
  assign regs_262_reset = io_reset; // @[:@38081.4 RegFile.scala 76:16:@38088.4]
  assign regs_262_io_in = 64'h0; // @[RegFile.scala 75:16:@38087.4]
  assign regs_262_io_reset = reset; // @[RegFile.scala 78:19:@38091.4]
  assign regs_262_io_enable = 1'h1; // @[RegFile.scala 74:20:@38085.4]
  assign regs_263_clock = clock; // @[:@38094.4]
  assign regs_263_reset = io_reset; // @[:@38095.4 RegFile.scala 76:16:@38102.4]
  assign regs_263_io_in = 64'h0; // @[RegFile.scala 75:16:@38101.4]
  assign regs_263_io_reset = reset; // @[RegFile.scala 78:19:@38105.4]
  assign regs_263_io_enable = 1'h1; // @[RegFile.scala 74:20:@38099.4]
  assign regs_264_clock = clock; // @[:@38108.4]
  assign regs_264_reset = io_reset; // @[:@38109.4 RegFile.scala 76:16:@38116.4]
  assign regs_264_io_in = 64'h0; // @[RegFile.scala 75:16:@38115.4]
  assign regs_264_io_reset = reset; // @[RegFile.scala 78:19:@38119.4]
  assign regs_264_io_enable = 1'h1; // @[RegFile.scala 74:20:@38113.4]
  assign regs_265_clock = clock; // @[:@38122.4]
  assign regs_265_reset = io_reset; // @[:@38123.4 RegFile.scala 76:16:@38130.4]
  assign regs_265_io_in = 64'h0; // @[RegFile.scala 75:16:@38129.4]
  assign regs_265_io_reset = reset; // @[RegFile.scala 78:19:@38133.4]
  assign regs_265_io_enable = 1'h1; // @[RegFile.scala 74:20:@38127.4]
  assign regs_266_clock = clock; // @[:@38136.4]
  assign regs_266_reset = io_reset; // @[:@38137.4 RegFile.scala 76:16:@38144.4]
  assign regs_266_io_in = 64'h0; // @[RegFile.scala 75:16:@38143.4]
  assign regs_266_io_reset = reset; // @[RegFile.scala 78:19:@38147.4]
  assign regs_266_io_enable = 1'h1; // @[RegFile.scala 74:20:@38141.4]
  assign regs_267_clock = clock; // @[:@38150.4]
  assign regs_267_reset = io_reset; // @[:@38151.4 RegFile.scala 76:16:@38158.4]
  assign regs_267_io_in = 64'h0; // @[RegFile.scala 75:16:@38157.4]
  assign regs_267_io_reset = reset; // @[RegFile.scala 78:19:@38161.4]
  assign regs_267_io_enable = 1'h1; // @[RegFile.scala 74:20:@38155.4]
  assign regs_268_clock = clock; // @[:@38164.4]
  assign regs_268_reset = io_reset; // @[:@38165.4 RegFile.scala 76:16:@38172.4]
  assign regs_268_io_in = 64'h0; // @[RegFile.scala 75:16:@38171.4]
  assign regs_268_io_reset = reset; // @[RegFile.scala 78:19:@38175.4]
  assign regs_268_io_enable = 1'h1; // @[RegFile.scala 74:20:@38169.4]
  assign regs_269_clock = clock; // @[:@38178.4]
  assign regs_269_reset = io_reset; // @[:@38179.4 RegFile.scala 76:16:@38186.4]
  assign regs_269_io_in = 64'h0; // @[RegFile.scala 75:16:@38185.4]
  assign regs_269_io_reset = reset; // @[RegFile.scala 78:19:@38189.4]
  assign regs_269_io_enable = 1'h1; // @[RegFile.scala 74:20:@38183.4]
  assign regs_270_clock = clock; // @[:@38192.4]
  assign regs_270_reset = io_reset; // @[:@38193.4 RegFile.scala 76:16:@38200.4]
  assign regs_270_io_in = 64'h0; // @[RegFile.scala 75:16:@38199.4]
  assign regs_270_io_reset = reset; // @[RegFile.scala 78:19:@38203.4]
  assign regs_270_io_enable = 1'h1; // @[RegFile.scala 74:20:@38197.4]
  assign regs_271_clock = clock; // @[:@38206.4]
  assign regs_271_reset = io_reset; // @[:@38207.4 RegFile.scala 76:16:@38214.4]
  assign regs_271_io_in = 64'h0; // @[RegFile.scala 75:16:@38213.4]
  assign regs_271_io_reset = reset; // @[RegFile.scala 78:19:@38217.4]
  assign regs_271_io_enable = 1'h1; // @[RegFile.scala 74:20:@38211.4]
  assign regs_272_clock = clock; // @[:@38220.4]
  assign regs_272_reset = io_reset; // @[:@38221.4 RegFile.scala 76:16:@38228.4]
  assign regs_272_io_in = 64'h0; // @[RegFile.scala 75:16:@38227.4]
  assign regs_272_io_reset = reset; // @[RegFile.scala 78:19:@38231.4]
  assign regs_272_io_enable = 1'h1; // @[RegFile.scala 74:20:@38225.4]
  assign regs_273_clock = clock; // @[:@38234.4]
  assign regs_273_reset = io_reset; // @[:@38235.4 RegFile.scala 76:16:@38242.4]
  assign regs_273_io_in = 64'h0; // @[RegFile.scala 75:16:@38241.4]
  assign regs_273_io_reset = reset; // @[RegFile.scala 78:19:@38245.4]
  assign regs_273_io_enable = 1'h1; // @[RegFile.scala 74:20:@38239.4]
  assign regs_274_clock = clock; // @[:@38248.4]
  assign regs_274_reset = io_reset; // @[:@38249.4 RegFile.scala 76:16:@38256.4]
  assign regs_274_io_in = 64'h0; // @[RegFile.scala 75:16:@38255.4]
  assign regs_274_io_reset = reset; // @[RegFile.scala 78:19:@38259.4]
  assign regs_274_io_enable = 1'h1; // @[RegFile.scala 74:20:@38253.4]
  assign regs_275_clock = clock; // @[:@38262.4]
  assign regs_275_reset = io_reset; // @[:@38263.4 RegFile.scala 76:16:@38270.4]
  assign regs_275_io_in = 64'h0; // @[RegFile.scala 75:16:@38269.4]
  assign regs_275_io_reset = reset; // @[RegFile.scala 78:19:@38273.4]
  assign regs_275_io_enable = 1'h1; // @[RegFile.scala 74:20:@38267.4]
  assign regs_276_clock = clock; // @[:@38276.4]
  assign regs_276_reset = io_reset; // @[:@38277.4 RegFile.scala 76:16:@38284.4]
  assign regs_276_io_in = 64'h0; // @[RegFile.scala 75:16:@38283.4]
  assign regs_276_io_reset = reset; // @[RegFile.scala 78:19:@38287.4]
  assign regs_276_io_enable = 1'h1; // @[RegFile.scala 74:20:@38281.4]
  assign regs_277_clock = clock; // @[:@38290.4]
  assign regs_277_reset = io_reset; // @[:@38291.4 RegFile.scala 76:16:@38298.4]
  assign regs_277_io_in = 64'h0; // @[RegFile.scala 75:16:@38297.4]
  assign regs_277_io_reset = reset; // @[RegFile.scala 78:19:@38301.4]
  assign regs_277_io_enable = 1'h1; // @[RegFile.scala 74:20:@38295.4]
  assign regs_278_clock = clock; // @[:@38304.4]
  assign regs_278_reset = io_reset; // @[:@38305.4 RegFile.scala 76:16:@38312.4]
  assign regs_278_io_in = 64'h0; // @[RegFile.scala 75:16:@38311.4]
  assign regs_278_io_reset = reset; // @[RegFile.scala 78:19:@38315.4]
  assign regs_278_io_enable = 1'h1; // @[RegFile.scala 74:20:@38309.4]
  assign regs_279_clock = clock; // @[:@38318.4]
  assign regs_279_reset = io_reset; // @[:@38319.4 RegFile.scala 76:16:@38326.4]
  assign regs_279_io_in = 64'h0; // @[RegFile.scala 75:16:@38325.4]
  assign regs_279_io_reset = reset; // @[RegFile.scala 78:19:@38329.4]
  assign regs_279_io_enable = 1'h1; // @[RegFile.scala 74:20:@38323.4]
  assign regs_280_clock = clock; // @[:@38332.4]
  assign regs_280_reset = io_reset; // @[:@38333.4 RegFile.scala 76:16:@38340.4]
  assign regs_280_io_in = 64'h0; // @[RegFile.scala 75:16:@38339.4]
  assign regs_280_io_reset = reset; // @[RegFile.scala 78:19:@38343.4]
  assign regs_280_io_enable = 1'h1; // @[RegFile.scala 74:20:@38337.4]
  assign regs_281_clock = clock; // @[:@38346.4]
  assign regs_281_reset = io_reset; // @[:@38347.4 RegFile.scala 76:16:@38354.4]
  assign regs_281_io_in = 64'h0; // @[RegFile.scala 75:16:@38353.4]
  assign regs_281_io_reset = reset; // @[RegFile.scala 78:19:@38357.4]
  assign regs_281_io_enable = 1'h1; // @[RegFile.scala 74:20:@38351.4]
  assign regs_282_clock = clock; // @[:@38360.4]
  assign regs_282_reset = io_reset; // @[:@38361.4 RegFile.scala 76:16:@38368.4]
  assign regs_282_io_in = 64'h0; // @[RegFile.scala 75:16:@38367.4]
  assign regs_282_io_reset = reset; // @[RegFile.scala 78:19:@38371.4]
  assign regs_282_io_enable = 1'h1; // @[RegFile.scala 74:20:@38365.4]
  assign regs_283_clock = clock; // @[:@38374.4]
  assign regs_283_reset = io_reset; // @[:@38375.4 RegFile.scala 76:16:@38382.4]
  assign regs_283_io_in = 64'h0; // @[RegFile.scala 75:16:@38381.4]
  assign regs_283_io_reset = reset; // @[RegFile.scala 78:19:@38385.4]
  assign regs_283_io_enable = 1'h1; // @[RegFile.scala 74:20:@38379.4]
  assign regs_284_clock = clock; // @[:@38388.4]
  assign regs_284_reset = io_reset; // @[:@38389.4 RegFile.scala 76:16:@38396.4]
  assign regs_284_io_in = 64'h0; // @[RegFile.scala 75:16:@38395.4]
  assign regs_284_io_reset = reset; // @[RegFile.scala 78:19:@38399.4]
  assign regs_284_io_enable = 1'h1; // @[RegFile.scala 74:20:@38393.4]
  assign regs_285_clock = clock; // @[:@38402.4]
  assign regs_285_reset = io_reset; // @[:@38403.4 RegFile.scala 76:16:@38410.4]
  assign regs_285_io_in = 64'h0; // @[RegFile.scala 75:16:@38409.4]
  assign regs_285_io_reset = reset; // @[RegFile.scala 78:19:@38413.4]
  assign regs_285_io_enable = 1'h1; // @[RegFile.scala 74:20:@38407.4]
  assign regs_286_clock = clock; // @[:@38416.4]
  assign regs_286_reset = io_reset; // @[:@38417.4 RegFile.scala 76:16:@38424.4]
  assign regs_286_io_in = 64'h0; // @[RegFile.scala 75:16:@38423.4]
  assign regs_286_io_reset = reset; // @[RegFile.scala 78:19:@38427.4]
  assign regs_286_io_enable = 1'h1; // @[RegFile.scala 74:20:@38421.4]
  assign regs_287_clock = clock; // @[:@38430.4]
  assign regs_287_reset = io_reset; // @[:@38431.4 RegFile.scala 76:16:@38438.4]
  assign regs_287_io_in = 64'h0; // @[RegFile.scala 75:16:@38437.4]
  assign regs_287_io_reset = reset; // @[RegFile.scala 78:19:@38441.4]
  assign regs_287_io_enable = 1'h1; // @[RegFile.scala 74:20:@38435.4]
  assign regs_288_clock = clock; // @[:@38444.4]
  assign regs_288_reset = io_reset; // @[:@38445.4 RegFile.scala 76:16:@38452.4]
  assign regs_288_io_in = 64'h0; // @[RegFile.scala 75:16:@38451.4]
  assign regs_288_io_reset = reset; // @[RegFile.scala 78:19:@38455.4]
  assign regs_288_io_enable = 1'h1; // @[RegFile.scala 74:20:@38449.4]
  assign regs_289_clock = clock; // @[:@38458.4]
  assign regs_289_reset = io_reset; // @[:@38459.4 RegFile.scala 76:16:@38466.4]
  assign regs_289_io_in = 64'h0; // @[RegFile.scala 75:16:@38465.4]
  assign regs_289_io_reset = reset; // @[RegFile.scala 78:19:@38469.4]
  assign regs_289_io_enable = 1'h1; // @[RegFile.scala 74:20:@38463.4]
  assign regs_290_clock = clock; // @[:@38472.4]
  assign regs_290_reset = io_reset; // @[:@38473.4 RegFile.scala 76:16:@38480.4]
  assign regs_290_io_in = 64'h0; // @[RegFile.scala 75:16:@38479.4]
  assign regs_290_io_reset = reset; // @[RegFile.scala 78:19:@38483.4]
  assign regs_290_io_enable = 1'h1; // @[RegFile.scala 74:20:@38477.4]
  assign regs_291_clock = clock; // @[:@38486.4]
  assign regs_291_reset = io_reset; // @[:@38487.4 RegFile.scala 76:16:@38494.4]
  assign regs_291_io_in = 64'h0; // @[RegFile.scala 75:16:@38493.4]
  assign regs_291_io_reset = reset; // @[RegFile.scala 78:19:@38497.4]
  assign regs_291_io_enable = 1'h1; // @[RegFile.scala 74:20:@38491.4]
  assign regs_292_clock = clock; // @[:@38500.4]
  assign regs_292_reset = io_reset; // @[:@38501.4 RegFile.scala 76:16:@38508.4]
  assign regs_292_io_in = 64'h0; // @[RegFile.scala 75:16:@38507.4]
  assign regs_292_io_reset = reset; // @[RegFile.scala 78:19:@38511.4]
  assign regs_292_io_enable = 1'h1; // @[RegFile.scala 74:20:@38505.4]
  assign regs_293_clock = clock; // @[:@38514.4]
  assign regs_293_reset = io_reset; // @[:@38515.4 RegFile.scala 76:16:@38522.4]
  assign regs_293_io_in = 64'h0; // @[RegFile.scala 75:16:@38521.4]
  assign regs_293_io_reset = reset; // @[RegFile.scala 78:19:@38525.4]
  assign regs_293_io_enable = 1'h1; // @[RegFile.scala 74:20:@38519.4]
  assign regs_294_clock = clock; // @[:@38528.4]
  assign regs_294_reset = io_reset; // @[:@38529.4 RegFile.scala 76:16:@38536.4]
  assign regs_294_io_in = 64'h0; // @[RegFile.scala 75:16:@38535.4]
  assign regs_294_io_reset = reset; // @[RegFile.scala 78:19:@38539.4]
  assign regs_294_io_enable = 1'h1; // @[RegFile.scala 74:20:@38533.4]
  assign regs_295_clock = clock; // @[:@38542.4]
  assign regs_295_reset = io_reset; // @[:@38543.4 RegFile.scala 76:16:@38550.4]
  assign regs_295_io_in = 64'h0; // @[RegFile.scala 75:16:@38549.4]
  assign regs_295_io_reset = reset; // @[RegFile.scala 78:19:@38553.4]
  assign regs_295_io_enable = 1'h1; // @[RegFile.scala 74:20:@38547.4]
  assign regs_296_clock = clock; // @[:@38556.4]
  assign regs_296_reset = io_reset; // @[:@38557.4 RegFile.scala 76:16:@38564.4]
  assign regs_296_io_in = 64'h0; // @[RegFile.scala 75:16:@38563.4]
  assign regs_296_io_reset = reset; // @[RegFile.scala 78:19:@38567.4]
  assign regs_296_io_enable = 1'h1; // @[RegFile.scala 74:20:@38561.4]
  assign regs_297_clock = clock; // @[:@38570.4]
  assign regs_297_reset = io_reset; // @[:@38571.4 RegFile.scala 76:16:@38578.4]
  assign regs_297_io_in = 64'h0; // @[RegFile.scala 75:16:@38577.4]
  assign regs_297_io_reset = reset; // @[RegFile.scala 78:19:@38581.4]
  assign regs_297_io_enable = 1'h1; // @[RegFile.scala 74:20:@38575.4]
  assign regs_298_clock = clock; // @[:@38584.4]
  assign regs_298_reset = io_reset; // @[:@38585.4 RegFile.scala 76:16:@38592.4]
  assign regs_298_io_in = 64'h0; // @[RegFile.scala 75:16:@38591.4]
  assign regs_298_io_reset = reset; // @[RegFile.scala 78:19:@38595.4]
  assign regs_298_io_enable = 1'h1; // @[RegFile.scala 74:20:@38589.4]
  assign regs_299_clock = clock; // @[:@38598.4]
  assign regs_299_reset = io_reset; // @[:@38599.4 RegFile.scala 76:16:@38606.4]
  assign regs_299_io_in = 64'h0; // @[RegFile.scala 75:16:@38605.4]
  assign regs_299_io_reset = reset; // @[RegFile.scala 78:19:@38609.4]
  assign regs_299_io_enable = 1'h1; // @[RegFile.scala 74:20:@38603.4]
  assign regs_300_clock = clock; // @[:@38612.4]
  assign regs_300_reset = io_reset; // @[:@38613.4 RegFile.scala 76:16:@38620.4]
  assign regs_300_io_in = 64'h0; // @[RegFile.scala 75:16:@38619.4]
  assign regs_300_io_reset = reset; // @[RegFile.scala 78:19:@38623.4]
  assign regs_300_io_enable = 1'h1; // @[RegFile.scala 74:20:@38617.4]
  assign regs_301_clock = clock; // @[:@38626.4]
  assign regs_301_reset = io_reset; // @[:@38627.4 RegFile.scala 76:16:@38634.4]
  assign regs_301_io_in = 64'h0; // @[RegFile.scala 75:16:@38633.4]
  assign regs_301_io_reset = reset; // @[RegFile.scala 78:19:@38637.4]
  assign regs_301_io_enable = 1'h1; // @[RegFile.scala 74:20:@38631.4]
  assign regs_302_clock = clock; // @[:@38640.4]
  assign regs_302_reset = io_reset; // @[:@38641.4 RegFile.scala 76:16:@38648.4]
  assign regs_302_io_in = 64'h0; // @[RegFile.scala 75:16:@38647.4]
  assign regs_302_io_reset = reset; // @[RegFile.scala 78:19:@38651.4]
  assign regs_302_io_enable = 1'h1; // @[RegFile.scala 74:20:@38645.4]
  assign regs_303_clock = clock; // @[:@38654.4]
  assign regs_303_reset = io_reset; // @[:@38655.4 RegFile.scala 76:16:@38662.4]
  assign regs_303_io_in = 64'h0; // @[RegFile.scala 75:16:@38661.4]
  assign regs_303_io_reset = reset; // @[RegFile.scala 78:19:@38665.4]
  assign regs_303_io_enable = 1'h1; // @[RegFile.scala 74:20:@38659.4]
  assign regs_304_clock = clock; // @[:@38668.4]
  assign regs_304_reset = io_reset; // @[:@38669.4 RegFile.scala 76:16:@38676.4]
  assign regs_304_io_in = 64'h0; // @[RegFile.scala 75:16:@38675.4]
  assign regs_304_io_reset = reset; // @[RegFile.scala 78:19:@38679.4]
  assign regs_304_io_enable = 1'h1; // @[RegFile.scala 74:20:@38673.4]
  assign regs_305_clock = clock; // @[:@38682.4]
  assign regs_305_reset = io_reset; // @[:@38683.4 RegFile.scala 76:16:@38690.4]
  assign regs_305_io_in = 64'h0; // @[RegFile.scala 75:16:@38689.4]
  assign regs_305_io_reset = reset; // @[RegFile.scala 78:19:@38693.4]
  assign regs_305_io_enable = 1'h1; // @[RegFile.scala 74:20:@38687.4]
  assign regs_306_clock = clock; // @[:@38696.4]
  assign regs_306_reset = io_reset; // @[:@38697.4 RegFile.scala 76:16:@38704.4]
  assign regs_306_io_in = 64'h0; // @[RegFile.scala 75:16:@38703.4]
  assign regs_306_io_reset = reset; // @[RegFile.scala 78:19:@38707.4]
  assign regs_306_io_enable = 1'h1; // @[RegFile.scala 74:20:@38701.4]
  assign regs_307_clock = clock; // @[:@38710.4]
  assign regs_307_reset = io_reset; // @[:@38711.4 RegFile.scala 76:16:@38718.4]
  assign regs_307_io_in = 64'h0; // @[RegFile.scala 75:16:@38717.4]
  assign regs_307_io_reset = reset; // @[RegFile.scala 78:19:@38721.4]
  assign regs_307_io_enable = 1'h1; // @[RegFile.scala 74:20:@38715.4]
  assign regs_308_clock = clock; // @[:@38724.4]
  assign regs_308_reset = io_reset; // @[:@38725.4 RegFile.scala 76:16:@38732.4]
  assign regs_308_io_in = 64'h0; // @[RegFile.scala 75:16:@38731.4]
  assign regs_308_io_reset = reset; // @[RegFile.scala 78:19:@38735.4]
  assign regs_308_io_enable = 1'h1; // @[RegFile.scala 74:20:@38729.4]
  assign regs_309_clock = clock; // @[:@38738.4]
  assign regs_309_reset = io_reset; // @[:@38739.4 RegFile.scala 76:16:@38746.4]
  assign regs_309_io_in = 64'h0; // @[RegFile.scala 75:16:@38745.4]
  assign regs_309_io_reset = reset; // @[RegFile.scala 78:19:@38749.4]
  assign regs_309_io_enable = 1'h1; // @[RegFile.scala 74:20:@38743.4]
  assign regs_310_clock = clock; // @[:@38752.4]
  assign regs_310_reset = io_reset; // @[:@38753.4 RegFile.scala 76:16:@38760.4]
  assign regs_310_io_in = 64'h0; // @[RegFile.scala 75:16:@38759.4]
  assign regs_310_io_reset = reset; // @[RegFile.scala 78:19:@38763.4]
  assign regs_310_io_enable = 1'h1; // @[RegFile.scala 74:20:@38757.4]
  assign regs_311_clock = clock; // @[:@38766.4]
  assign regs_311_reset = io_reset; // @[:@38767.4 RegFile.scala 76:16:@38774.4]
  assign regs_311_io_in = 64'h0; // @[RegFile.scala 75:16:@38773.4]
  assign regs_311_io_reset = reset; // @[RegFile.scala 78:19:@38777.4]
  assign regs_311_io_enable = 1'h1; // @[RegFile.scala 74:20:@38771.4]
  assign regs_312_clock = clock; // @[:@38780.4]
  assign regs_312_reset = io_reset; // @[:@38781.4 RegFile.scala 76:16:@38788.4]
  assign regs_312_io_in = 64'h0; // @[RegFile.scala 75:16:@38787.4]
  assign regs_312_io_reset = reset; // @[RegFile.scala 78:19:@38791.4]
  assign regs_312_io_enable = 1'h1; // @[RegFile.scala 74:20:@38785.4]
  assign regs_313_clock = clock; // @[:@38794.4]
  assign regs_313_reset = io_reset; // @[:@38795.4 RegFile.scala 76:16:@38802.4]
  assign regs_313_io_in = 64'h0; // @[RegFile.scala 75:16:@38801.4]
  assign regs_313_io_reset = reset; // @[RegFile.scala 78:19:@38805.4]
  assign regs_313_io_enable = 1'h1; // @[RegFile.scala 74:20:@38799.4]
  assign regs_314_clock = clock; // @[:@38808.4]
  assign regs_314_reset = io_reset; // @[:@38809.4 RegFile.scala 76:16:@38816.4]
  assign regs_314_io_in = 64'h0; // @[RegFile.scala 75:16:@38815.4]
  assign regs_314_io_reset = reset; // @[RegFile.scala 78:19:@38819.4]
  assign regs_314_io_enable = 1'h1; // @[RegFile.scala 74:20:@38813.4]
  assign regs_315_clock = clock; // @[:@38822.4]
  assign regs_315_reset = io_reset; // @[:@38823.4 RegFile.scala 76:16:@38830.4]
  assign regs_315_io_in = 64'h0; // @[RegFile.scala 75:16:@38829.4]
  assign regs_315_io_reset = reset; // @[RegFile.scala 78:19:@38833.4]
  assign regs_315_io_enable = 1'h1; // @[RegFile.scala 74:20:@38827.4]
  assign regs_316_clock = clock; // @[:@38836.4]
  assign regs_316_reset = io_reset; // @[:@38837.4 RegFile.scala 76:16:@38844.4]
  assign regs_316_io_in = 64'h0; // @[RegFile.scala 75:16:@38843.4]
  assign regs_316_io_reset = reset; // @[RegFile.scala 78:19:@38847.4]
  assign regs_316_io_enable = 1'h1; // @[RegFile.scala 74:20:@38841.4]
  assign regs_317_clock = clock; // @[:@38850.4]
  assign regs_317_reset = io_reset; // @[:@38851.4 RegFile.scala 76:16:@38858.4]
  assign regs_317_io_in = 64'h0; // @[RegFile.scala 75:16:@38857.4]
  assign regs_317_io_reset = reset; // @[RegFile.scala 78:19:@38861.4]
  assign regs_317_io_enable = 1'h1; // @[RegFile.scala 74:20:@38855.4]
  assign regs_318_clock = clock; // @[:@38864.4]
  assign regs_318_reset = io_reset; // @[:@38865.4 RegFile.scala 76:16:@38872.4]
  assign regs_318_io_in = 64'h0; // @[RegFile.scala 75:16:@38871.4]
  assign regs_318_io_reset = reset; // @[RegFile.scala 78:19:@38875.4]
  assign regs_318_io_enable = 1'h1; // @[RegFile.scala 74:20:@38869.4]
  assign regs_319_clock = clock; // @[:@38878.4]
  assign regs_319_reset = io_reset; // @[:@38879.4 RegFile.scala 76:16:@38886.4]
  assign regs_319_io_in = 64'h0; // @[RegFile.scala 75:16:@38885.4]
  assign regs_319_io_reset = reset; // @[RegFile.scala 78:19:@38889.4]
  assign regs_319_io_enable = 1'h1; // @[RegFile.scala 74:20:@38883.4]
  assign regs_320_clock = clock; // @[:@38892.4]
  assign regs_320_reset = io_reset; // @[:@38893.4 RegFile.scala 76:16:@38900.4]
  assign regs_320_io_in = 64'h0; // @[RegFile.scala 75:16:@38899.4]
  assign regs_320_io_reset = reset; // @[RegFile.scala 78:19:@38903.4]
  assign regs_320_io_enable = 1'h1; // @[RegFile.scala 74:20:@38897.4]
  assign regs_321_clock = clock; // @[:@38906.4]
  assign regs_321_reset = io_reset; // @[:@38907.4 RegFile.scala 76:16:@38914.4]
  assign regs_321_io_in = 64'h0; // @[RegFile.scala 75:16:@38913.4]
  assign regs_321_io_reset = reset; // @[RegFile.scala 78:19:@38917.4]
  assign regs_321_io_enable = 1'h1; // @[RegFile.scala 74:20:@38911.4]
  assign regs_322_clock = clock; // @[:@38920.4]
  assign regs_322_reset = io_reset; // @[:@38921.4 RegFile.scala 76:16:@38928.4]
  assign regs_322_io_in = 64'h0; // @[RegFile.scala 75:16:@38927.4]
  assign regs_322_io_reset = reset; // @[RegFile.scala 78:19:@38931.4]
  assign regs_322_io_enable = 1'h1; // @[RegFile.scala 74:20:@38925.4]
  assign regs_323_clock = clock; // @[:@38934.4]
  assign regs_323_reset = io_reset; // @[:@38935.4 RegFile.scala 76:16:@38942.4]
  assign regs_323_io_in = 64'h0; // @[RegFile.scala 75:16:@38941.4]
  assign regs_323_io_reset = reset; // @[RegFile.scala 78:19:@38945.4]
  assign regs_323_io_enable = 1'h1; // @[RegFile.scala 74:20:@38939.4]
  assign regs_324_clock = clock; // @[:@38948.4]
  assign regs_324_reset = io_reset; // @[:@38949.4 RegFile.scala 76:16:@38956.4]
  assign regs_324_io_in = 64'h0; // @[RegFile.scala 75:16:@38955.4]
  assign regs_324_io_reset = reset; // @[RegFile.scala 78:19:@38959.4]
  assign regs_324_io_enable = 1'h1; // @[RegFile.scala 74:20:@38953.4]
  assign regs_325_clock = clock; // @[:@38962.4]
  assign regs_325_reset = io_reset; // @[:@38963.4 RegFile.scala 76:16:@38970.4]
  assign regs_325_io_in = 64'h0; // @[RegFile.scala 75:16:@38969.4]
  assign regs_325_io_reset = reset; // @[RegFile.scala 78:19:@38973.4]
  assign regs_325_io_enable = 1'h1; // @[RegFile.scala 74:20:@38967.4]
  assign regs_326_clock = clock; // @[:@38976.4]
  assign regs_326_reset = io_reset; // @[:@38977.4 RegFile.scala 76:16:@38984.4]
  assign regs_326_io_in = 64'h0; // @[RegFile.scala 75:16:@38983.4]
  assign regs_326_io_reset = reset; // @[RegFile.scala 78:19:@38987.4]
  assign regs_326_io_enable = 1'h1; // @[RegFile.scala 74:20:@38981.4]
  assign regs_327_clock = clock; // @[:@38990.4]
  assign regs_327_reset = io_reset; // @[:@38991.4 RegFile.scala 76:16:@38998.4]
  assign regs_327_io_in = 64'h0; // @[RegFile.scala 75:16:@38997.4]
  assign regs_327_io_reset = reset; // @[RegFile.scala 78:19:@39001.4]
  assign regs_327_io_enable = 1'h1; // @[RegFile.scala 74:20:@38995.4]
  assign regs_328_clock = clock; // @[:@39004.4]
  assign regs_328_reset = io_reset; // @[:@39005.4 RegFile.scala 76:16:@39012.4]
  assign regs_328_io_in = 64'h0; // @[RegFile.scala 75:16:@39011.4]
  assign regs_328_io_reset = reset; // @[RegFile.scala 78:19:@39015.4]
  assign regs_328_io_enable = 1'h1; // @[RegFile.scala 74:20:@39009.4]
  assign regs_329_clock = clock; // @[:@39018.4]
  assign regs_329_reset = io_reset; // @[:@39019.4 RegFile.scala 76:16:@39026.4]
  assign regs_329_io_in = 64'h0; // @[RegFile.scala 75:16:@39025.4]
  assign regs_329_io_reset = reset; // @[RegFile.scala 78:19:@39029.4]
  assign regs_329_io_enable = 1'h1; // @[RegFile.scala 74:20:@39023.4]
  assign regs_330_clock = clock; // @[:@39032.4]
  assign regs_330_reset = io_reset; // @[:@39033.4 RegFile.scala 76:16:@39040.4]
  assign regs_330_io_in = 64'h0; // @[RegFile.scala 75:16:@39039.4]
  assign regs_330_io_reset = reset; // @[RegFile.scala 78:19:@39043.4]
  assign regs_330_io_enable = 1'h1; // @[RegFile.scala 74:20:@39037.4]
  assign regs_331_clock = clock; // @[:@39046.4]
  assign regs_331_reset = io_reset; // @[:@39047.4 RegFile.scala 76:16:@39054.4]
  assign regs_331_io_in = 64'h0; // @[RegFile.scala 75:16:@39053.4]
  assign regs_331_io_reset = reset; // @[RegFile.scala 78:19:@39057.4]
  assign regs_331_io_enable = 1'h1; // @[RegFile.scala 74:20:@39051.4]
  assign regs_332_clock = clock; // @[:@39060.4]
  assign regs_332_reset = io_reset; // @[:@39061.4 RegFile.scala 76:16:@39068.4]
  assign regs_332_io_in = 64'h0; // @[RegFile.scala 75:16:@39067.4]
  assign regs_332_io_reset = reset; // @[RegFile.scala 78:19:@39071.4]
  assign regs_332_io_enable = 1'h1; // @[RegFile.scala 74:20:@39065.4]
  assign regs_333_clock = clock; // @[:@39074.4]
  assign regs_333_reset = io_reset; // @[:@39075.4 RegFile.scala 76:16:@39082.4]
  assign regs_333_io_in = 64'h0; // @[RegFile.scala 75:16:@39081.4]
  assign regs_333_io_reset = reset; // @[RegFile.scala 78:19:@39085.4]
  assign regs_333_io_enable = 1'h1; // @[RegFile.scala 74:20:@39079.4]
  assign regs_334_clock = clock; // @[:@39088.4]
  assign regs_334_reset = io_reset; // @[:@39089.4 RegFile.scala 76:16:@39096.4]
  assign regs_334_io_in = 64'h0; // @[RegFile.scala 75:16:@39095.4]
  assign regs_334_io_reset = reset; // @[RegFile.scala 78:19:@39099.4]
  assign regs_334_io_enable = 1'h1; // @[RegFile.scala 74:20:@39093.4]
  assign regs_335_clock = clock; // @[:@39102.4]
  assign regs_335_reset = io_reset; // @[:@39103.4 RegFile.scala 76:16:@39110.4]
  assign regs_335_io_in = 64'h0; // @[RegFile.scala 75:16:@39109.4]
  assign regs_335_io_reset = reset; // @[RegFile.scala 78:19:@39113.4]
  assign regs_335_io_enable = 1'h1; // @[RegFile.scala 74:20:@39107.4]
  assign regs_336_clock = clock; // @[:@39116.4]
  assign regs_336_reset = io_reset; // @[:@39117.4 RegFile.scala 76:16:@39124.4]
  assign regs_336_io_in = 64'h0; // @[RegFile.scala 75:16:@39123.4]
  assign regs_336_io_reset = reset; // @[RegFile.scala 78:19:@39127.4]
  assign regs_336_io_enable = 1'h1; // @[RegFile.scala 74:20:@39121.4]
  assign regs_337_clock = clock; // @[:@39130.4]
  assign regs_337_reset = io_reset; // @[:@39131.4 RegFile.scala 76:16:@39138.4]
  assign regs_337_io_in = 64'h0; // @[RegFile.scala 75:16:@39137.4]
  assign regs_337_io_reset = reset; // @[RegFile.scala 78:19:@39141.4]
  assign regs_337_io_enable = 1'h1; // @[RegFile.scala 74:20:@39135.4]
  assign regs_338_clock = clock; // @[:@39144.4]
  assign regs_338_reset = io_reset; // @[:@39145.4 RegFile.scala 76:16:@39152.4]
  assign regs_338_io_in = 64'h0; // @[RegFile.scala 75:16:@39151.4]
  assign regs_338_io_reset = reset; // @[RegFile.scala 78:19:@39155.4]
  assign regs_338_io_enable = 1'h1; // @[RegFile.scala 74:20:@39149.4]
  assign regs_339_clock = clock; // @[:@39158.4]
  assign regs_339_reset = io_reset; // @[:@39159.4 RegFile.scala 76:16:@39166.4]
  assign regs_339_io_in = 64'h0; // @[RegFile.scala 75:16:@39165.4]
  assign regs_339_io_reset = reset; // @[RegFile.scala 78:19:@39169.4]
  assign regs_339_io_enable = 1'h1; // @[RegFile.scala 74:20:@39163.4]
  assign regs_340_clock = clock; // @[:@39172.4]
  assign regs_340_reset = io_reset; // @[:@39173.4 RegFile.scala 76:16:@39180.4]
  assign regs_340_io_in = 64'h0; // @[RegFile.scala 75:16:@39179.4]
  assign regs_340_io_reset = reset; // @[RegFile.scala 78:19:@39183.4]
  assign regs_340_io_enable = 1'h1; // @[RegFile.scala 74:20:@39177.4]
  assign regs_341_clock = clock; // @[:@39186.4]
  assign regs_341_reset = io_reset; // @[:@39187.4 RegFile.scala 76:16:@39194.4]
  assign regs_341_io_in = 64'h0; // @[RegFile.scala 75:16:@39193.4]
  assign regs_341_io_reset = reset; // @[RegFile.scala 78:19:@39197.4]
  assign regs_341_io_enable = 1'h1; // @[RegFile.scala 74:20:@39191.4]
  assign regs_342_clock = clock; // @[:@39200.4]
  assign regs_342_reset = io_reset; // @[:@39201.4 RegFile.scala 76:16:@39208.4]
  assign regs_342_io_in = 64'h0; // @[RegFile.scala 75:16:@39207.4]
  assign regs_342_io_reset = reset; // @[RegFile.scala 78:19:@39211.4]
  assign regs_342_io_enable = 1'h1; // @[RegFile.scala 74:20:@39205.4]
  assign regs_343_clock = clock; // @[:@39214.4]
  assign regs_343_reset = io_reset; // @[:@39215.4 RegFile.scala 76:16:@39222.4]
  assign regs_343_io_in = 64'h0; // @[RegFile.scala 75:16:@39221.4]
  assign regs_343_io_reset = reset; // @[RegFile.scala 78:19:@39225.4]
  assign regs_343_io_enable = 1'h1; // @[RegFile.scala 74:20:@39219.4]
  assign regs_344_clock = clock; // @[:@39228.4]
  assign regs_344_reset = io_reset; // @[:@39229.4 RegFile.scala 76:16:@39236.4]
  assign regs_344_io_in = 64'h0; // @[RegFile.scala 75:16:@39235.4]
  assign regs_344_io_reset = reset; // @[RegFile.scala 78:19:@39239.4]
  assign regs_344_io_enable = 1'h1; // @[RegFile.scala 74:20:@39233.4]
  assign regs_345_clock = clock; // @[:@39242.4]
  assign regs_345_reset = io_reset; // @[:@39243.4 RegFile.scala 76:16:@39250.4]
  assign regs_345_io_in = 64'h0; // @[RegFile.scala 75:16:@39249.4]
  assign regs_345_io_reset = reset; // @[RegFile.scala 78:19:@39253.4]
  assign regs_345_io_enable = 1'h1; // @[RegFile.scala 74:20:@39247.4]
  assign regs_346_clock = clock; // @[:@39256.4]
  assign regs_346_reset = io_reset; // @[:@39257.4 RegFile.scala 76:16:@39264.4]
  assign regs_346_io_in = 64'h0; // @[RegFile.scala 75:16:@39263.4]
  assign regs_346_io_reset = reset; // @[RegFile.scala 78:19:@39267.4]
  assign regs_346_io_enable = 1'h1; // @[RegFile.scala 74:20:@39261.4]
  assign regs_347_clock = clock; // @[:@39270.4]
  assign regs_347_reset = io_reset; // @[:@39271.4 RegFile.scala 76:16:@39278.4]
  assign regs_347_io_in = 64'h0; // @[RegFile.scala 75:16:@39277.4]
  assign regs_347_io_reset = reset; // @[RegFile.scala 78:19:@39281.4]
  assign regs_347_io_enable = 1'h1; // @[RegFile.scala 74:20:@39275.4]
  assign regs_348_clock = clock; // @[:@39284.4]
  assign regs_348_reset = io_reset; // @[:@39285.4 RegFile.scala 76:16:@39292.4]
  assign regs_348_io_in = 64'h0; // @[RegFile.scala 75:16:@39291.4]
  assign regs_348_io_reset = reset; // @[RegFile.scala 78:19:@39295.4]
  assign regs_348_io_enable = 1'h1; // @[RegFile.scala 74:20:@39289.4]
  assign regs_349_clock = clock; // @[:@39298.4]
  assign regs_349_reset = io_reset; // @[:@39299.4 RegFile.scala 76:16:@39306.4]
  assign regs_349_io_in = 64'h0; // @[RegFile.scala 75:16:@39305.4]
  assign regs_349_io_reset = reset; // @[RegFile.scala 78:19:@39309.4]
  assign regs_349_io_enable = 1'h1; // @[RegFile.scala 74:20:@39303.4]
  assign regs_350_clock = clock; // @[:@39312.4]
  assign regs_350_reset = io_reset; // @[:@39313.4 RegFile.scala 76:16:@39320.4]
  assign regs_350_io_in = 64'h0; // @[RegFile.scala 75:16:@39319.4]
  assign regs_350_io_reset = reset; // @[RegFile.scala 78:19:@39323.4]
  assign regs_350_io_enable = 1'h1; // @[RegFile.scala 74:20:@39317.4]
  assign regs_351_clock = clock; // @[:@39326.4]
  assign regs_351_reset = io_reset; // @[:@39327.4 RegFile.scala 76:16:@39334.4]
  assign regs_351_io_in = 64'h0; // @[RegFile.scala 75:16:@39333.4]
  assign regs_351_io_reset = reset; // @[RegFile.scala 78:19:@39337.4]
  assign regs_351_io_enable = 1'h1; // @[RegFile.scala 74:20:@39331.4]
  assign regs_352_clock = clock; // @[:@39340.4]
  assign regs_352_reset = io_reset; // @[:@39341.4 RegFile.scala 76:16:@39348.4]
  assign regs_352_io_in = 64'h0; // @[RegFile.scala 75:16:@39347.4]
  assign regs_352_io_reset = reset; // @[RegFile.scala 78:19:@39351.4]
  assign regs_352_io_enable = 1'h1; // @[RegFile.scala 74:20:@39345.4]
  assign regs_353_clock = clock; // @[:@39354.4]
  assign regs_353_reset = io_reset; // @[:@39355.4 RegFile.scala 76:16:@39362.4]
  assign regs_353_io_in = 64'h0; // @[RegFile.scala 75:16:@39361.4]
  assign regs_353_io_reset = reset; // @[RegFile.scala 78:19:@39365.4]
  assign regs_353_io_enable = 1'h1; // @[RegFile.scala 74:20:@39359.4]
  assign regs_354_clock = clock; // @[:@39368.4]
  assign regs_354_reset = io_reset; // @[:@39369.4 RegFile.scala 76:16:@39376.4]
  assign regs_354_io_in = 64'h0; // @[RegFile.scala 75:16:@39375.4]
  assign regs_354_io_reset = reset; // @[RegFile.scala 78:19:@39379.4]
  assign regs_354_io_enable = 1'h1; // @[RegFile.scala 74:20:@39373.4]
  assign regs_355_clock = clock; // @[:@39382.4]
  assign regs_355_reset = io_reset; // @[:@39383.4 RegFile.scala 76:16:@39390.4]
  assign regs_355_io_in = 64'h0; // @[RegFile.scala 75:16:@39389.4]
  assign regs_355_io_reset = reset; // @[RegFile.scala 78:19:@39393.4]
  assign regs_355_io_enable = 1'h1; // @[RegFile.scala 74:20:@39387.4]
  assign regs_356_clock = clock; // @[:@39396.4]
  assign regs_356_reset = io_reset; // @[:@39397.4 RegFile.scala 76:16:@39404.4]
  assign regs_356_io_in = 64'h0; // @[RegFile.scala 75:16:@39403.4]
  assign regs_356_io_reset = reset; // @[RegFile.scala 78:19:@39407.4]
  assign regs_356_io_enable = 1'h1; // @[RegFile.scala 74:20:@39401.4]
  assign regs_357_clock = clock; // @[:@39410.4]
  assign regs_357_reset = io_reset; // @[:@39411.4 RegFile.scala 76:16:@39418.4]
  assign regs_357_io_in = 64'h0; // @[RegFile.scala 75:16:@39417.4]
  assign regs_357_io_reset = reset; // @[RegFile.scala 78:19:@39421.4]
  assign regs_357_io_enable = 1'h1; // @[RegFile.scala 74:20:@39415.4]
  assign regs_358_clock = clock; // @[:@39424.4]
  assign regs_358_reset = io_reset; // @[:@39425.4 RegFile.scala 76:16:@39432.4]
  assign regs_358_io_in = 64'h0; // @[RegFile.scala 75:16:@39431.4]
  assign regs_358_io_reset = reset; // @[RegFile.scala 78:19:@39435.4]
  assign regs_358_io_enable = 1'h1; // @[RegFile.scala 74:20:@39429.4]
  assign regs_359_clock = clock; // @[:@39438.4]
  assign regs_359_reset = io_reset; // @[:@39439.4 RegFile.scala 76:16:@39446.4]
  assign regs_359_io_in = 64'h0; // @[RegFile.scala 75:16:@39445.4]
  assign regs_359_io_reset = reset; // @[RegFile.scala 78:19:@39449.4]
  assign regs_359_io_enable = 1'h1; // @[RegFile.scala 74:20:@39443.4]
  assign regs_360_clock = clock; // @[:@39452.4]
  assign regs_360_reset = io_reset; // @[:@39453.4 RegFile.scala 76:16:@39460.4]
  assign regs_360_io_in = 64'h0; // @[RegFile.scala 75:16:@39459.4]
  assign regs_360_io_reset = reset; // @[RegFile.scala 78:19:@39463.4]
  assign regs_360_io_enable = 1'h1; // @[RegFile.scala 74:20:@39457.4]
  assign regs_361_clock = clock; // @[:@39466.4]
  assign regs_361_reset = io_reset; // @[:@39467.4 RegFile.scala 76:16:@39474.4]
  assign regs_361_io_in = 64'h0; // @[RegFile.scala 75:16:@39473.4]
  assign regs_361_io_reset = reset; // @[RegFile.scala 78:19:@39477.4]
  assign regs_361_io_enable = 1'h1; // @[RegFile.scala 74:20:@39471.4]
  assign regs_362_clock = clock; // @[:@39480.4]
  assign regs_362_reset = io_reset; // @[:@39481.4 RegFile.scala 76:16:@39488.4]
  assign regs_362_io_in = 64'h0; // @[RegFile.scala 75:16:@39487.4]
  assign regs_362_io_reset = reset; // @[RegFile.scala 78:19:@39491.4]
  assign regs_362_io_enable = 1'h1; // @[RegFile.scala 74:20:@39485.4]
  assign regs_363_clock = clock; // @[:@39494.4]
  assign regs_363_reset = io_reset; // @[:@39495.4 RegFile.scala 76:16:@39502.4]
  assign regs_363_io_in = 64'h0; // @[RegFile.scala 75:16:@39501.4]
  assign regs_363_io_reset = reset; // @[RegFile.scala 78:19:@39505.4]
  assign regs_363_io_enable = 1'h1; // @[RegFile.scala 74:20:@39499.4]
  assign regs_364_clock = clock; // @[:@39508.4]
  assign regs_364_reset = io_reset; // @[:@39509.4 RegFile.scala 76:16:@39516.4]
  assign regs_364_io_in = 64'h0; // @[RegFile.scala 75:16:@39515.4]
  assign regs_364_io_reset = reset; // @[RegFile.scala 78:19:@39519.4]
  assign regs_364_io_enable = 1'h1; // @[RegFile.scala 74:20:@39513.4]
  assign regs_365_clock = clock; // @[:@39522.4]
  assign regs_365_reset = io_reset; // @[:@39523.4 RegFile.scala 76:16:@39530.4]
  assign regs_365_io_in = 64'h0; // @[RegFile.scala 75:16:@39529.4]
  assign regs_365_io_reset = reset; // @[RegFile.scala 78:19:@39533.4]
  assign regs_365_io_enable = 1'h1; // @[RegFile.scala 74:20:@39527.4]
  assign regs_366_clock = clock; // @[:@39536.4]
  assign regs_366_reset = io_reset; // @[:@39537.4 RegFile.scala 76:16:@39544.4]
  assign regs_366_io_in = 64'h0; // @[RegFile.scala 75:16:@39543.4]
  assign regs_366_io_reset = reset; // @[RegFile.scala 78:19:@39547.4]
  assign regs_366_io_enable = 1'h1; // @[RegFile.scala 74:20:@39541.4]
  assign regs_367_clock = clock; // @[:@39550.4]
  assign regs_367_reset = io_reset; // @[:@39551.4 RegFile.scala 76:16:@39558.4]
  assign regs_367_io_in = 64'h0; // @[RegFile.scala 75:16:@39557.4]
  assign regs_367_io_reset = reset; // @[RegFile.scala 78:19:@39561.4]
  assign regs_367_io_enable = 1'h1; // @[RegFile.scala 74:20:@39555.4]
  assign regs_368_clock = clock; // @[:@39564.4]
  assign regs_368_reset = io_reset; // @[:@39565.4 RegFile.scala 76:16:@39572.4]
  assign regs_368_io_in = 64'h0; // @[RegFile.scala 75:16:@39571.4]
  assign regs_368_io_reset = reset; // @[RegFile.scala 78:19:@39575.4]
  assign regs_368_io_enable = 1'h1; // @[RegFile.scala 74:20:@39569.4]
  assign regs_369_clock = clock; // @[:@39578.4]
  assign regs_369_reset = io_reset; // @[:@39579.4 RegFile.scala 76:16:@39586.4]
  assign regs_369_io_in = 64'h0; // @[RegFile.scala 75:16:@39585.4]
  assign regs_369_io_reset = reset; // @[RegFile.scala 78:19:@39589.4]
  assign regs_369_io_enable = 1'h1; // @[RegFile.scala 74:20:@39583.4]
  assign regs_370_clock = clock; // @[:@39592.4]
  assign regs_370_reset = io_reset; // @[:@39593.4 RegFile.scala 76:16:@39600.4]
  assign regs_370_io_in = 64'h0; // @[RegFile.scala 75:16:@39599.4]
  assign regs_370_io_reset = reset; // @[RegFile.scala 78:19:@39603.4]
  assign regs_370_io_enable = 1'h1; // @[RegFile.scala 74:20:@39597.4]
  assign regs_371_clock = clock; // @[:@39606.4]
  assign regs_371_reset = io_reset; // @[:@39607.4 RegFile.scala 76:16:@39614.4]
  assign regs_371_io_in = 64'h0; // @[RegFile.scala 75:16:@39613.4]
  assign regs_371_io_reset = reset; // @[RegFile.scala 78:19:@39617.4]
  assign regs_371_io_enable = 1'h1; // @[RegFile.scala 74:20:@39611.4]
  assign regs_372_clock = clock; // @[:@39620.4]
  assign regs_372_reset = io_reset; // @[:@39621.4 RegFile.scala 76:16:@39628.4]
  assign regs_372_io_in = 64'h0; // @[RegFile.scala 75:16:@39627.4]
  assign regs_372_io_reset = reset; // @[RegFile.scala 78:19:@39631.4]
  assign regs_372_io_enable = 1'h1; // @[RegFile.scala 74:20:@39625.4]
  assign regs_373_clock = clock; // @[:@39634.4]
  assign regs_373_reset = io_reset; // @[:@39635.4 RegFile.scala 76:16:@39642.4]
  assign regs_373_io_in = 64'h0; // @[RegFile.scala 75:16:@39641.4]
  assign regs_373_io_reset = reset; // @[RegFile.scala 78:19:@39645.4]
  assign regs_373_io_enable = 1'h1; // @[RegFile.scala 74:20:@39639.4]
  assign regs_374_clock = clock; // @[:@39648.4]
  assign regs_374_reset = io_reset; // @[:@39649.4 RegFile.scala 76:16:@39656.4]
  assign regs_374_io_in = 64'h0; // @[RegFile.scala 75:16:@39655.4]
  assign regs_374_io_reset = reset; // @[RegFile.scala 78:19:@39659.4]
  assign regs_374_io_enable = 1'h1; // @[RegFile.scala 74:20:@39653.4]
  assign regs_375_clock = clock; // @[:@39662.4]
  assign regs_375_reset = io_reset; // @[:@39663.4 RegFile.scala 76:16:@39670.4]
  assign regs_375_io_in = 64'h0; // @[RegFile.scala 75:16:@39669.4]
  assign regs_375_io_reset = reset; // @[RegFile.scala 78:19:@39673.4]
  assign regs_375_io_enable = 1'h1; // @[RegFile.scala 74:20:@39667.4]
  assign regs_376_clock = clock; // @[:@39676.4]
  assign regs_376_reset = io_reset; // @[:@39677.4 RegFile.scala 76:16:@39684.4]
  assign regs_376_io_in = 64'h0; // @[RegFile.scala 75:16:@39683.4]
  assign regs_376_io_reset = reset; // @[RegFile.scala 78:19:@39687.4]
  assign regs_376_io_enable = 1'h1; // @[RegFile.scala 74:20:@39681.4]
  assign regs_377_clock = clock; // @[:@39690.4]
  assign regs_377_reset = io_reset; // @[:@39691.4 RegFile.scala 76:16:@39698.4]
  assign regs_377_io_in = 64'h0; // @[RegFile.scala 75:16:@39697.4]
  assign regs_377_io_reset = reset; // @[RegFile.scala 78:19:@39701.4]
  assign regs_377_io_enable = 1'h1; // @[RegFile.scala 74:20:@39695.4]
  assign regs_378_clock = clock; // @[:@39704.4]
  assign regs_378_reset = io_reset; // @[:@39705.4 RegFile.scala 76:16:@39712.4]
  assign regs_378_io_in = 64'h0; // @[RegFile.scala 75:16:@39711.4]
  assign regs_378_io_reset = reset; // @[RegFile.scala 78:19:@39715.4]
  assign regs_378_io_enable = 1'h1; // @[RegFile.scala 74:20:@39709.4]
  assign regs_379_clock = clock; // @[:@39718.4]
  assign regs_379_reset = io_reset; // @[:@39719.4 RegFile.scala 76:16:@39726.4]
  assign regs_379_io_in = 64'h0; // @[RegFile.scala 75:16:@39725.4]
  assign regs_379_io_reset = reset; // @[RegFile.scala 78:19:@39729.4]
  assign regs_379_io_enable = 1'h1; // @[RegFile.scala 74:20:@39723.4]
  assign regs_380_clock = clock; // @[:@39732.4]
  assign regs_380_reset = io_reset; // @[:@39733.4 RegFile.scala 76:16:@39740.4]
  assign regs_380_io_in = 64'h0; // @[RegFile.scala 75:16:@39739.4]
  assign regs_380_io_reset = reset; // @[RegFile.scala 78:19:@39743.4]
  assign regs_380_io_enable = 1'h1; // @[RegFile.scala 74:20:@39737.4]
  assign regs_381_clock = clock; // @[:@39746.4]
  assign regs_381_reset = io_reset; // @[:@39747.4 RegFile.scala 76:16:@39754.4]
  assign regs_381_io_in = 64'h0; // @[RegFile.scala 75:16:@39753.4]
  assign regs_381_io_reset = reset; // @[RegFile.scala 78:19:@39757.4]
  assign regs_381_io_enable = 1'h1; // @[RegFile.scala 74:20:@39751.4]
  assign regs_382_clock = clock; // @[:@39760.4]
  assign regs_382_reset = io_reset; // @[:@39761.4 RegFile.scala 76:16:@39768.4]
  assign regs_382_io_in = 64'h0; // @[RegFile.scala 75:16:@39767.4]
  assign regs_382_io_reset = reset; // @[RegFile.scala 78:19:@39771.4]
  assign regs_382_io_enable = 1'h1; // @[RegFile.scala 74:20:@39765.4]
  assign regs_383_clock = clock; // @[:@39774.4]
  assign regs_383_reset = io_reset; // @[:@39775.4 RegFile.scala 76:16:@39782.4]
  assign regs_383_io_in = 64'h0; // @[RegFile.scala 75:16:@39781.4]
  assign regs_383_io_reset = reset; // @[RegFile.scala 78:19:@39785.4]
  assign regs_383_io_enable = 1'h1; // @[RegFile.scala 74:20:@39779.4]
  assign regs_384_clock = clock; // @[:@39788.4]
  assign regs_384_reset = io_reset; // @[:@39789.4 RegFile.scala 76:16:@39796.4]
  assign regs_384_io_in = 64'h0; // @[RegFile.scala 75:16:@39795.4]
  assign regs_384_io_reset = reset; // @[RegFile.scala 78:19:@39799.4]
  assign regs_384_io_enable = 1'h1; // @[RegFile.scala 74:20:@39793.4]
  assign regs_385_clock = clock; // @[:@39802.4]
  assign regs_385_reset = io_reset; // @[:@39803.4 RegFile.scala 76:16:@39810.4]
  assign regs_385_io_in = 64'h0; // @[RegFile.scala 75:16:@39809.4]
  assign regs_385_io_reset = reset; // @[RegFile.scala 78:19:@39813.4]
  assign regs_385_io_enable = 1'h1; // @[RegFile.scala 74:20:@39807.4]
  assign regs_386_clock = clock; // @[:@39816.4]
  assign regs_386_reset = io_reset; // @[:@39817.4 RegFile.scala 76:16:@39824.4]
  assign regs_386_io_in = 64'h0; // @[RegFile.scala 75:16:@39823.4]
  assign regs_386_io_reset = reset; // @[RegFile.scala 78:19:@39827.4]
  assign regs_386_io_enable = 1'h1; // @[RegFile.scala 74:20:@39821.4]
  assign regs_387_clock = clock; // @[:@39830.4]
  assign regs_387_reset = io_reset; // @[:@39831.4 RegFile.scala 76:16:@39838.4]
  assign regs_387_io_in = 64'h0; // @[RegFile.scala 75:16:@39837.4]
  assign regs_387_io_reset = reset; // @[RegFile.scala 78:19:@39841.4]
  assign regs_387_io_enable = 1'h1; // @[RegFile.scala 74:20:@39835.4]
  assign regs_388_clock = clock; // @[:@39844.4]
  assign regs_388_reset = io_reset; // @[:@39845.4 RegFile.scala 76:16:@39852.4]
  assign regs_388_io_in = 64'h0; // @[RegFile.scala 75:16:@39851.4]
  assign regs_388_io_reset = reset; // @[RegFile.scala 78:19:@39855.4]
  assign regs_388_io_enable = 1'h1; // @[RegFile.scala 74:20:@39849.4]
  assign regs_389_clock = clock; // @[:@39858.4]
  assign regs_389_reset = io_reset; // @[:@39859.4 RegFile.scala 76:16:@39866.4]
  assign regs_389_io_in = 64'h0; // @[RegFile.scala 75:16:@39865.4]
  assign regs_389_io_reset = reset; // @[RegFile.scala 78:19:@39869.4]
  assign regs_389_io_enable = 1'h1; // @[RegFile.scala 74:20:@39863.4]
  assign regs_390_clock = clock; // @[:@39872.4]
  assign regs_390_reset = io_reset; // @[:@39873.4 RegFile.scala 76:16:@39880.4]
  assign regs_390_io_in = 64'h0; // @[RegFile.scala 75:16:@39879.4]
  assign regs_390_io_reset = reset; // @[RegFile.scala 78:19:@39883.4]
  assign regs_390_io_enable = 1'h1; // @[RegFile.scala 74:20:@39877.4]
  assign regs_391_clock = clock; // @[:@39886.4]
  assign regs_391_reset = io_reset; // @[:@39887.4 RegFile.scala 76:16:@39894.4]
  assign regs_391_io_in = 64'h0; // @[RegFile.scala 75:16:@39893.4]
  assign regs_391_io_reset = reset; // @[RegFile.scala 78:19:@39897.4]
  assign regs_391_io_enable = 1'h1; // @[RegFile.scala 74:20:@39891.4]
  assign regs_392_clock = clock; // @[:@39900.4]
  assign regs_392_reset = io_reset; // @[:@39901.4 RegFile.scala 76:16:@39908.4]
  assign regs_392_io_in = 64'h0; // @[RegFile.scala 75:16:@39907.4]
  assign regs_392_io_reset = reset; // @[RegFile.scala 78:19:@39911.4]
  assign regs_392_io_enable = 1'h1; // @[RegFile.scala 74:20:@39905.4]
  assign regs_393_clock = clock; // @[:@39914.4]
  assign regs_393_reset = io_reset; // @[:@39915.4 RegFile.scala 76:16:@39922.4]
  assign regs_393_io_in = 64'h0; // @[RegFile.scala 75:16:@39921.4]
  assign regs_393_io_reset = reset; // @[RegFile.scala 78:19:@39925.4]
  assign regs_393_io_enable = 1'h1; // @[RegFile.scala 74:20:@39919.4]
  assign regs_394_clock = clock; // @[:@39928.4]
  assign regs_394_reset = io_reset; // @[:@39929.4 RegFile.scala 76:16:@39936.4]
  assign regs_394_io_in = 64'h0; // @[RegFile.scala 75:16:@39935.4]
  assign regs_394_io_reset = reset; // @[RegFile.scala 78:19:@39939.4]
  assign regs_394_io_enable = 1'h1; // @[RegFile.scala 74:20:@39933.4]
  assign regs_395_clock = clock; // @[:@39942.4]
  assign regs_395_reset = io_reset; // @[:@39943.4 RegFile.scala 76:16:@39950.4]
  assign regs_395_io_in = 64'h0; // @[RegFile.scala 75:16:@39949.4]
  assign regs_395_io_reset = reset; // @[RegFile.scala 78:19:@39953.4]
  assign regs_395_io_enable = 1'h1; // @[RegFile.scala 74:20:@39947.4]
  assign regs_396_clock = clock; // @[:@39956.4]
  assign regs_396_reset = io_reset; // @[:@39957.4 RegFile.scala 76:16:@39964.4]
  assign regs_396_io_in = 64'h0; // @[RegFile.scala 75:16:@39963.4]
  assign regs_396_io_reset = reset; // @[RegFile.scala 78:19:@39967.4]
  assign regs_396_io_enable = 1'h1; // @[RegFile.scala 74:20:@39961.4]
  assign regs_397_clock = clock; // @[:@39970.4]
  assign regs_397_reset = io_reset; // @[:@39971.4 RegFile.scala 76:16:@39978.4]
  assign regs_397_io_in = 64'h0; // @[RegFile.scala 75:16:@39977.4]
  assign regs_397_io_reset = reset; // @[RegFile.scala 78:19:@39981.4]
  assign regs_397_io_enable = 1'h1; // @[RegFile.scala 74:20:@39975.4]
  assign regs_398_clock = clock; // @[:@39984.4]
  assign regs_398_reset = io_reset; // @[:@39985.4 RegFile.scala 76:16:@39992.4]
  assign regs_398_io_in = 64'h0; // @[RegFile.scala 75:16:@39991.4]
  assign regs_398_io_reset = reset; // @[RegFile.scala 78:19:@39995.4]
  assign regs_398_io_enable = 1'h1; // @[RegFile.scala 74:20:@39989.4]
  assign regs_399_clock = clock; // @[:@39998.4]
  assign regs_399_reset = io_reset; // @[:@39999.4 RegFile.scala 76:16:@40006.4]
  assign regs_399_io_in = 64'h0; // @[RegFile.scala 75:16:@40005.4]
  assign regs_399_io_reset = reset; // @[RegFile.scala 78:19:@40009.4]
  assign regs_399_io_enable = 1'h1; // @[RegFile.scala 74:20:@40003.4]
  assign regs_400_clock = clock; // @[:@40012.4]
  assign regs_400_reset = io_reset; // @[:@40013.4 RegFile.scala 76:16:@40020.4]
  assign regs_400_io_in = 64'h0; // @[RegFile.scala 75:16:@40019.4]
  assign regs_400_io_reset = reset; // @[RegFile.scala 78:19:@40023.4]
  assign regs_400_io_enable = 1'h1; // @[RegFile.scala 74:20:@40017.4]
  assign regs_401_clock = clock; // @[:@40026.4]
  assign regs_401_reset = io_reset; // @[:@40027.4 RegFile.scala 76:16:@40034.4]
  assign regs_401_io_in = 64'h0; // @[RegFile.scala 75:16:@40033.4]
  assign regs_401_io_reset = reset; // @[RegFile.scala 78:19:@40037.4]
  assign regs_401_io_enable = 1'h1; // @[RegFile.scala 74:20:@40031.4]
  assign regs_402_clock = clock; // @[:@40040.4]
  assign regs_402_reset = io_reset; // @[:@40041.4 RegFile.scala 76:16:@40048.4]
  assign regs_402_io_in = 64'h0; // @[RegFile.scala 75:16:@40047.4]
  assign regs_402_io_reset = reset; // @[RegFile.scala 78:19:@40051.4]
  assign regs_402_io_enable = 1'h1; // @[RegFile.scala 74:20:@40045.4]
  assign regs_403_clock = clock; // @[:@40054.4]
  assign regs_403_reset = io_reset; // @[:@40055.4 RegFile.scala 76:16:@40062.4]
  assign regs_403_io_in = 64'h0; // @[RegFile.scala 75:16:@40061.4]
  assign regs_403_io_reset = reset; // @[RegFile.scala 78:19:@40065.4]
  assign regs_403_io_enable = 1'h1; // @[RegFile.scala 74:20:@40059.4]
  assign regs_404_clock = clock; // @[:@40068.4]
  assign regs_404_reset = io_reset; // @[:@40069.4 RegFile.scala 76:16:@40076.4]
  assign regs_404_io_in = 64'h0; // @[RegFile.scala 75:16:@40075.4]
  assign regs_404_io_reset = reset; // @[RegFile.scala 78:19:@40079.4]
  assign regs_404_io_enable = 1'h1; // @[RegFile.scala 74:20:@40073.4]
  assign regs_405_clock = clock; // @[:@40082.4]
  assign regs_405_reset = io_reset; // @[:@40083.4 RegFile.scala 76:16:@40090.4]
  assign regs_405_io_in = 64'h0; // @[RegFile.scala 75:16:@40089.4]
  assign regs_405_io_reset = reset; // @[RegFile.scala 78:19:@40093.4]
  assign regs_405_io_enable = 1'h1; // @[RegFile.scala 74:20:@40087.4]
  assign regs_406_clock = clock; // @[:@40096.4]
  assign regs_406_reset = io_reset; // @[:@40097.4 RegFile.scala 76:16:@40104.4]
  assign regs_406_io_in = 64'h0; // @[RegFile.scala 75:16:@40103.4]
  assign regs_406_io_reset = reset; // @[RegFile.scala 78:19:@40107.4]
  assign regs_406_io_enable = 1'h1; // @[RegFile.scala 74:20:@40101.4]
  assign regs_407_clock = clock; // @[:@40110.4]
  assign regs_407_reset = io_reset; // @[:@40111.4 RegFile.scala 76:16:@40118.4]
  assign regs_407_io_in = 64'h0; // @[RegFile.scala 75:16:@40117.4]
  assign regs_407_io_reset = reset; // @[RegFile.scala 78:19:@40121.4]
  assign regs_407_io_enable = 1'h1; // @[RegFile.scala 74:20:@40115.4]
  assign regs_408_clock = clock; // @[:@40124.4]
  assign regs_408_reset = io_reset; // @[:@40125.4 RegFile.scala 76:16:@40132.4]
  assign regs_408_io_in = 64'h0; // @[RegFile.scala 75:16:@40131.4]
  assign regs_408_io_reset = reset; // @[RegFile.scala 78:19:@40135.4]
  assign regs_408_io_enable = 1'h1; // @[RegFile.scala 74:20:@40129.4]
  assign regs_409_clock = clock; // @[:@40138.4]
  assign regs_409_reset = io_reset; // @[:@40139.4 RegFile.scala 76:16:@40146.4]
  assign regs_409_io_in = 64'h0; // @[RegFile.scala 75:16:@40145.4]
  assign regs_409_io_reset = reset; // @[RegFile.scala 78:19:@40149.4]
  assign regs_409_io_enable = 1'h1; // @[RegFile.scala 74:20:@40143.4]
  assign regs_410_clock = clock; // @[:@40152.4]
  assign regs_410_reset = io_reset; // @[:@40153.4 RegFile.scala 76:16:@40160.4]
  assign regs_410_io_in = 64'h0; // @[RegFile.scala 75:16:@40159.4]
  assign regs_410_io_reset = reset; // @[RegFile.scala 78:19:@40163.4]
  assign regs_410_io_enable = 1'h1; // @[RegFile.scala 74:20:@40157.4]
  assign regs_411_clock = clock; // @[:@40166.4]
  assign regs_411_reset = io_reset; // @[:@40167.4 RegFile.scala 76:16:@40174.4]
  assign regs_411_io_in = 64'h0; // @[RegFile.scala 75:16:@40173.4]
  assign regs_411_io_reset = reset; // @[RegFile.scala 78:19:@40177.4]
  assign regs_411_io_enable = 1'h1; // @[RegFile.scala 74:20:@40171.4]
  assign regs_412_clock = clock; // @[:@40180.4]
  assign regs_412_reset = io_reset; // @[:@40181.4 RegFile.scala 76:16:@40188.4]
  assign regs_412_io_in = 64'h0; // @[RegFile.scala 75:16:@40187.4]
  assign regs_412_io_reset = reset; // @[RegFile.scala 78:19:@40191.4]
  assign regs_412_io_enable = 1'h1; // @[RegFile.scala 74:20:@40185.4]
  assign regs_413_clock = clock; // @[:@40194.4]
  assign regs_413_reset = io_reset; // @[:@40195.4 RegFile.scala 76:16:@40202.4]
  assign regs_413_io_in = 64'h0; // @[RegFile.scala 75:16:@40201.4]
  assign regs_413_io_reset = reset; // @[RegFile.scala 78:19:@40205.4]
  assign regs_413_io_enable = 1'h1; // @[RegFile.scala 74:20:@40199.4]
  assign regs_414_clock = clock; // @[:@40208.4]
  assign regs_414_reset = io_reset; // @[:@40209.4 RegFile.scala 76:16:@40216.4]
  assign regs_414_io_in = 64'h0; // @[RegFile.scala 75:16:@40215.4]
  assign regs_414_io_reset = reset; // @[RegFile.scala 78:19:@40219.4]
  assign regs_414_io_enable = 1'h1; // @[RegFile.scala 74:20:@40213.4]
  assign regs_415_clock = clock; // @[:@40222.4]
  assign regs_415_reset = io_reset; // @[:@40223.4 RegFile.scala 76:16:@40230.4]
  assign regs_415_io_in = 64'h0; // @[RegFile.scala 75:16:@40229.4]
  assign regs_415_io_reset = reset; // @[RegFile.scala 78:19:@40233.4]
  assign regs_415_io_enable = 1'h1; // @[RegFile.scala 74:20:@40227.4]
  assign regs_416_clock = clock; // @[:@40236.4]
  assign regs_416_reset = io_reset; // @[:@40237.4 RegFile.scala 76:16:@40244.4]
  assign regs_416_io_in = 64'h0; // @[RegFile.scala 75:16:@40243.4]
  assign regs_416_io_reset = reset; // @[RegFile.scala 78:19:@40247.4]
  assign regs_416_io_enable = 1'h1; // @[RegFile.scala 74:20:@40241.4]
  assign regs_417_clock = clock; // @[:@40250.4]
  assign regs_417_reset = io_reset; // @[:@40251.4 RegFile.scala 76:16:@40258.4]
  assign regs_417_io_in = 64'h0; // @[RegFile.scala 75:16:@40257.4]
  assign regs_417_io_reset = reset; // @[RegFile.scala 78:19:@40261.4]
  assign regs_417_io_enable = 1'h1; // @[RegFile.scala 74:20:@40255.4]
  assign regs_418_clock = clock; // @[:@40264.4]
  assign regs_418_reset = io_reset; // @[:@40265.4 RegFile.scala 76:16:@40272.4]
  assign regs_418_io_in = 64'h0; // @[RegFile.scala 75:16:@40271.4]
  assign regs_418_io_reset = reset; // @[RegFile.scala 78:19:@40275.4]
  assign regs_418_io_enable = 1'h1; // @[RegFile.scala 74:20:@40269.4]
  assign regs_419_clock = clock; // @[:@40278.4]
  assign regs_419_reset = io_reset; // @[:@40279.4 RegFile.scala 76:16:@40286.4]
  assign regs_419_io_in = 64'h0; // @[RegFile.scala 75:16:@40285.4]
  assign regs_419_io_reset = reset; // @[RegFile.scala 78:19:@40289.4]
  assign regs_419_io_enable = 1'h1; // @[RegFile.scala 74:20:@40283.4]
  assign regs_420_clock = clock; // @[:@40292.4]
  assign regs_420_reset = io_reset; // @[:@40293.4 RegFile.scala 76:16:@40300.4]
  assign regs_420_io_in = 64'h0; // @[RegFile.scala 75:16:@40299.4]
  assign regs_420_io_reset = reset; // @[RegFile.scala 78:19:@40303.4]
  assign regs_420_io_enable = 1'h1; // @[RegFile.scala 74:20:@40297.4]
  assign regs_421_clock = clock; // @[:@40306.4]
  assign regs_421_reset = io_reset; // @[:@40307.4 RegFile.scala 76:16:@40314.4]
  assign regs_421_io_in = 64'h0; // @[RegFile.scala 75:16:@40313.4]
  assign regs_421_io_reset = reset; // @[RegFile.scala 78:19:@40317.4]
  assign regs_421_io_enable = 1'h1; // @[RegFile.scala 74:20:@40311.4]
  assign regs_422_clock = clock; // @[:@40320.4]
  assign regs_422_reset = io_reset; // @[:@40321.4 RegFile.scala 76:16:@40328.4]
  assign regs_422_io_in = 64'h0; // @[RegFile.scala 75:16:@40327.4]
  assign regs_422_io_reset = reset; // @[RegFile.scala 78:19:@40331.4]
  assign regs_422_io_enable = 1'h1; // @[RegFile.scala 74:20:@40325.4]
  assign regs_423_clock = clock; // @[:@40334.4]
  assign regs_423_reset = io_reset; // @[:@40335.4 RegFile.scala 76:16:@40342.4]
  assign regs_423_io_in = 64'h0; // @[RegFile.scala 75:16:@40341.4]
  assign regs_423_io_reset = reset; // @[RegFile.scala 78:19:@40345.4]
  assign regs_423_io_enable = 1'h1; // @[RegFile.scala 74:20:@40339.4]
  assign regs_424_clock = clock; // @[:@40348.4]
  assign regs_424_reset = io_reset; // @[:@40349.4 RegFile.scala 76:16:@40356.4]
  assign regs_424_io_in = 64'h0; // @[RegFile.scala 75:16:@40355.4]
  assign regs_424_io_reset = reset; // @[RegFile.scala 78:19:@40359.4]
  assign regs_424_io_enable = 1'h1; // @[RegFile.scala 74:20:@40353.4]
  assign regs_425_clock = clock; // @[:@40362.4]
  assign regs_425_reset = io_reset; // @[:@40363.4 RegFile.scala 76:16:@40370.4]
  assign regs_425_io_in = 64'h0; // @[RegFile.scala 75:16:@40369.4]
  assign regs_425_io_reset = reset; // @[RegFile.scala 78:19:@40373.4]
  assign regs_425_io_enable = 1'h1; // @[RegFile.scala 74:20:@40367.4]
  assign regs_426_clock = clock; // @[:@40376.4]
  assign regs_426_reset = io_reset; // @[:@40377.4 RegFile.scala 76:16:@40384.4]
  assign regs_426_io_in = 64'h0; // @[RegFile.scala 75:16:@40383.4]
  assign regs_426_io_reset = reset; // @[RegFile.scala 78:19:@40387.4]
  assign regs_426_io_enable = 1'h1; // @[RegFile.scala 74:20:@40381.4]
  assign regs_427_clock = clock; // @[:@40390.4]
  assign regs_427_reset = io_reset; // @[:@40391.4 RegFile.scala 76:16:@40398.4]
  assign regs_427_io_in = 64'h0; // @[RegFile.scala 75:16:@40397.4]
  assign regs_427_io_reset = reset; // @[RegFile.scala 78:19:@40401.4]
  assign regs_427_io_enable = 1'h1; // @[RegFile.scala 74:20:@40395.4]
  assign regs_428_clock = clock; // @[:@40404.4]
  assign regs_428_reset = io_reset; // @[:@40405.4 RegFile.scala 76:16:@40412.4]
  assign regs_428_io_in = 64'h0; // @[RegFile.scala 75:16:@40411.4]
  assign regs_428_io_reset = reset; // @[RegFile.scala 78:19:@40415.4]
  assign regs_428_io_enable = 1'h1; // @[RegFile.scala 74:20:@40409.4]
  assign regs_429_clock = clock; // @[:@40418.4]
  assign regs_429_reset = io_reset; // @[:@40419.4 RegFile.scala 76:16:@40426.4]
  assign regs_429_io_in = 64'h0; // @[RegFile.scala 75:16:@40425.4]
  assign regs_429_io_reset = reset; // @[RegFile.scala 78:19:@40429.4]
  assign regs_429_io_enable = 1'h1; // @[RegFile.scala 74:20:@40423.4]
  assign regs_430_clock = clock; // @[:@40432.4]
  assign regs_430_reset = io_reset; // @[:@40433.4 RegFile.scala 76:16:@40440.4]
  assign regs_430_io_in = 64'h0; // @[RegFile.scala 75:16:@40439.4]
  assign regs_430_io_reset = reset; // @[RegFile.scala 78:19:@40443.4]
  assign regs_430_io_enable = 1'h1; // @[RegFile.scala 74:20:@40437.4]
  assign regs_431_clock = clock; // @[:@40446.4]
  assign regs_431_reset = io_reset; // @[:@40447.4 RegFile.scala 76:16:@40454.4]
  assign regs_431_io_in = 64'h0; // @[RegFile.scala 75:16:@40453.4]
  assign regs_431_io_reset = reset; // @[RegFile.scala 78:19:@40457.4]
  assign regs_431_io_enable = 1'h1; // @[RegFile.scala 74:20:@40451.4]
  assign regs_432_clock = clock; // @[:@40460.4]
  assign regs_432_reset = io_reset; // @[:@40461.4 RegFile.scala 76:16:@40468.4]
  assign regs_432_io_in = 64'h0; // @[RegFile.scala 75:16:@40467.4]
  assign regs_432_io_reset = reset; // @[RegFile.scala 78:19:@40471.4]
  assign regs_432_io_enable = 1'h1; // @[RegFile.scala 74:20:@40465.4]
  assign regs_433_clock = clock; // @[:@40474.4]
  assign regs_433_reset = io_reset; // @[:@40475.4 RegFile.scala 76:16:@40482.4]
  assign regs_433_io_in = 64'h0; // @[RegFile.scala 75:16:@40481.4]
  assign regs_433_io_reset = reset; // @[RegFile.scala 78:19:@40485.4]
  assign regs_433_io_enable = 1'h1; // @[RegFile.scala 74:20:@40479.4]
  assign regs_434_clock = clock; // @[:@40488.4]
  assign regs_434_reset = io_reset; // @[:@40489.4 RegFile.scala 76:16:@40496.4]
  assign regs_434_io_in = 64'h0; // @[RegFile.scala 75:16:@40495.4]
  assign regs_434_io_reset = reset; // @[RegFile.scala 78:19:@40499.4]
  assign regs_434_io_enable = 1'h1; // @[RegFile.scala 74:20:@40493.4]
  assign regs_435_clock = clock; // @[:@40502.4]
  assign regs_435_reset = io_reset; // @[:@40503.4 RegFile.scala 76:16:@40510.4]
  assign regs_435_io_in = 64'h0; // @[RegFile.scala 75:16:@40509.4]
  assign regs_435_io_reset = reset; // @[RegFile.scala 78:19:@40513.4]
  assign regs_435_io_enable = 1'h1; // @[RegFile.scala 74:20:@40507.4]
  assign regs_436_clock = clock; // @[:@40516.4]
  assign regs_436_reset = io_reset; // @[:@40517.4 RegFile.scala 76:16:@40524.4]
  assign regs_436_io_in = 64'h0; // @[RegFile.scala 75:16:@40523.4]
  assign regs_436_io_reset = reset; // @[RegFile.scala 78:19:@40527.4]
  assign regs_436_io_enable = 1'h1; // @[RegFile.scala 74:20:@40521.4]
  assign regs_437_clock = clock; // @[:@40530.4]
  assign regs_437_reset = io_reset; // @[:@40531.4 RegFile.scala 76:16:@40538.4]
  assign regs_437_io_in = 64'h0; // @[RegFile.scala 75:16:@40537.4]
  assign regs_437_io_reset = reset; // @[RegFile.scala 78:19:@40541.4]
  assign regs_437_io_enable = 1'h1; // @[RegFile.scala 74:20:@40535.4]
  assign regs_438_clock = clock; // @[:@40544.4]
  assign regs_438_reset = io_reset; // @[:@40545.4 RegFile.scala 76:16:@40552.4]
  assign regs_438_io_in = 64'h0; // @[RegFile.scala 75:16:@40551.4]
  assign regs_438_io_reset = reset; // @[RegFile.scala 78:19:@40555.4]
  assign regs_438_io_enable = 1'h1; // @[RegFile.scala 74:20:@40549.4]
  assign regs_439_clock = clock; // @[:@40558.4]
  assign regs_439_reset = io_reset; // @[:@40559.4 RegFile.scala 76:16:@40566.4]
  assign regs_439_io_in = 64'h0; // @[RegFile.scala 75:16:@40565.4]
  assign regs_439_io_reset = reset; // @[RegFile.scala 78:19:@40569.4]
  assign regs_439_io_enable = 1'h1; // @[RegFile.scala 74:20:@40563.4]
  assign regs_440_clock = clock; // @[:@40572.4]
  assign regs_440_reset = io_reset; // @[:@40573.4 RegFile.scala 76:16:@40580.4]
  assign regs_440_io_in = 64'h0; // @[RegFile.scala 75:16:@40579.4]
  assign regs_440_io_reset = reset; // @[RegFile.scala 78:19:@40583.4]
  assign regs_440_io_enable = 1'h1; // @[RegFile.scala 74:20:@40577.4]
  assign regs_441_clock = clock; // @[:@40586.4]
  assign regs_441_reset = io_reset; // @[:@40587.4 RegFile.scala 76:16:@40594.4]
  assign regs_441_io_in = 64'h0; // @[RegFile.scala 75:16:@40593.4]
  assign regs_441_io_reset = reset; // @[RegFile.scala 78:19:@40597.4]
  assign regs_441_io_enable = 1'h1; // @[RegFile.scala 74:20:@40591.4]
  assign regs_442_clock = clock; // @[:@40600.4]
  assign regs_442_reset = io_reset; // @[:@40601.4 RegFile.scala 76:16:@40608.4]
  assign regs_442_io_in = 64'h0; // @[RegFile.scala 75:16:@40607.4]
  assign regs_442_io_reset = reset; // @[RegFile.scala 78:19:@40611.4]
  assign regs_442_io_enable = 1'h1; // @[RegFile.scala 74:20:@40605.4]
  assign regs_443_clock = clock; // @[:@40614.4]
  assign regs_443_reset = io_reset; // @[:@40615.4 RegFile.scala 76:16:@40622.4]
  assign regs_443_io_in = 64'h0; // @[RegFile.scala 75:16:@40621.4]
  assign regs_443_io_reset = reset; // @[RegFile.scala 78:19:@40625.4]
  assign regs_443_io_enable = 1'h1; // @[RegFile.scala 74:20:@40619.4]
  assign regs_444_clock = clock; // @[:@40628.4]
  assign regs_444_reset = io_reset; // @[:@40629.4 RegFile.scala 76:16:@40636.4]
  assign regs_444_io_in = 64'h0; // @[RegFile.scala 75:16:@40635.4]
  assign regs_444_io_reset = reset; // @[RegFile.scala 78:19:@40639.4]
  assign regs_444_io_enable = 1'h1; // @[RegFile.scala 74:20:@40633.4]
  assign regs_445_clock = clock; // @[:@40642.4]
  assign regs_445_reset = io_reset; // @[:@40643.4 RegFile.scala 76:16:@40650.4]
  assign regs_445_io_in = 64'h0; // @[RegFile.scala 75:16:@40649.4]
  assign regs_445_io_reset = reset; // @[RegFile.scala 78:19:@40653.4]
  assign regs_445_io_enable = 1'h1; // @[RegFile.scala 74:20:@40647.4]
  assign regs_446_clock = clock; // @[:@40656.4]
  assign regs_446_reset = io_reset; // @[:@40657.4 RegFile.scala 76:16:@40664.4]
  assign regs_446_io_in = 64'h0; // @[RegFile.scala 75:16:@40663.4]
  assign regs_446_io_reset = reset; // @[RegFile.scala 78:19:@40667.4]
  assign regs_446_io_enable = 1'h1; // @[RegFile.scala 74:20:@40661.4]
  assign regs_447_clock = clock; // @[:@40670.4]
  assign regs_447_reset = io_reset; // @[:@40671.4 RegFile.scala 76:16:@40678.4]
  assign regs_447_io_in = 64'h0; // @[RegFile.scala 75:16:@40677.4]
  assign regs_447_io_reset = reset; // @[RegFile.scala 78:19:@40681.4]
  assign regs_447_io_enable = 1'h1; // @[RegFile.scala 74:20:@40675.4]
  assign regs_448_clock = clock; // @[:@40684.4]
  assign regs_448_reset = io_reset; // @[:@40685.4 RegFile.scala 76:16:@40692.4]
  assign regs_448_io_in = 64'h0; // @[RegFile.scala 75:16:@40691.4]
  assign regs_448_io_reset = reset; // @[RegFile.scala 78:19:@40695.4]
  assign regs_448_io_enable = 1'h1; // @[RegFile.scala 74:20:@40689.4]
  assign regs_449_clock = clock; // @[:@40698.4]
  assign regs_449_reset = io_reset; // @[:@40699.4 RegFile.scala 76:16:@40706.4]
  assign regs_449_io_in = 64'h0; // @[RegFile.scala 75:16:@40705.4]
  assign regs_449_io_reset = reset; // @[RegFile.scala 78:19:@40709.4]
  assign regs_449_io_enable = 1'h1; // @[RegFile.scala 74:20:@40703.4]
  assign regs_450_clock = clock; // @[:@40712.4]
  assign regs_450_reset = io_reset; // @[:@40713.4 RegFile.scala 76:16:@40720.4]
  assign regs_450_io_in = 64'h0; // @[RegFile.scala 75:16:@40719.4]
  assign regs_450_io_reset = reset; // @[RegFile.scala 78:19:@40723.4]
  assign regs_450_io_enable = 1'h1; // @[RegFile.scala 74:20:@40717.4]
  assign regs_451_clock = clock; // @[:@40726.4]
  assign regs_451_reset = io_reset; // @[:@40727.4 RegFile.scala 76:16:@40734.4]
  assign regs_451_io_in = 64'h0; // @[RegFile.scala 75:16:@40733.4]
  assign regs_451_io_reset = reset; // @[RegFile.scala 78:19:@40737.4]
  assign regs_451_io_enable = 1'h1; // @[RegFile.scala 74:20:@40731.4]
  assign regs_452_clock = clock; // @[:@40740.4]
  assign regs_452_reset = io_reset; // @[:@40741.4 RegFile.scala 76:16:@40748.4]
  assign regs_452_io_in = 64'h0; // @[RegFile.scala 75:16:@40747.4]
  assign regs_452_io_reset = reset; // @[RegFile.scala 78:19:@40751.4]
  assign regs_452_io_enable = 1'h1; // @[RegFile.scala 74:20:@40745.4]
  assign regs_453_clock = clock; // @[:@40754.4]
  assign regs_453_reset = io_reset; // @[:@40755.4 RegFile.scala 76:16:@40762.4]
  assign regs_453_io_in = 64'h0; // @[RegFile.scala 75:16:@40761.4]
  assign regs_453_io_reset = reset; // @[RegFile.scala 78:19:@40765.4]
  assign regs_453_io_enable = 1'h1; // @[RegFile.scala 74:20:@40759.4]
  assign regs_454_clock = clock; // @[:@40768.4]
  assign regs_454_reset = io_reset; // @[:@40769.4 RegFile.scala 76:16:@40776.4]
  assign regs_454_io_in = 64'h0; // @[RegFile.scala 75:16:@40775.4]
  assign regs_454_io_reset = reset; // @[RegFile.scala 78:19:@40779.4]
  assign regs_454_io_enable = 1'h1; // @[RegFile.scala 74:20:@40773.4]
  assign regs_455_clock = clock; // @[:@40782.4]
  assign regs_455_reset = io_reset; // @[:@40783.4 RegFile.scala 76:16:@40790.4]
  assign regs_455_io_in = 64'h0; // @[RegFile.scala 75:16:@40789.4]
  assign regs_455_io_reset = reset; // @[RegFile.scala 78:19:@40793.4]
  assign regs_455_io_enable = 1'h1; // @[RegFile.scala 74:20:@40787.4]
  assign regs_456_clock = clock; // @[:@40796.4]
  assign regs_456_reset = io_reset; // @[:@40797.4 RegFile.scala 76:16:@40804.4]
  assign regs_456_io_in = 64'h0; // @[RegFile.scala 75:16:@40803.4]
  assign regs_456_io_reset = reset; // @[RegFile.scala 78:19:@40807.4]
  assign regs_456_io_enable = 1'h1; // @[RegFile.scala 74:20:@40801.4]
  assign regs_457_clock = clock; // @[:@40810.4]
  assign regs_457_reset = io_reset; // @[:@40811.4 RegFile.scala 76:16:@40818.4]
  assign regs_457_io_in = 64'h0; // @[RegFile.scala 75:16:@40817.4]
  assign regs_457_io_reset = reset; // @[RegFile.scala 78:19:@40821.4]
  assign regs_457_io_enable = 1'h1; // @[RegFile.scala 74:20:@40815.4]
  assign regs_458_clock = clock; // @[:@40824.4]
  assign regs_458_reset = io_reset; // @[:@40825.4 RegFile.scala 76:16:@40832.4]
  assign regs_458_io_in = 64'h0; // @[RegFile.scala 75:16:@40831.4]
  assign regs_458_io_reset = reset; // @[RegFile.scala 78:19:@40835.4]
  assign regs_458_io_enable = 1'h1; // @[RegFile.scala 74:20:@40829.4]
  assign regs_459_clock = clock; // @[:@40838.4]
  assign regs_459_reset = io_reset; // @[:@40839.4 RegFile.scala 76:16:@40846.4]
  assign regs_459_io_in = 64'h0; // @[RegFile.scala 75:16:@40845.4]
  assign regs_459_io_reset = reset; // @[RegFile.scala 78:19:@40849.4]
  assign regs_459_io_enable = 1'h1; // @[RegFile.scala 74:20:@40843.4]
  assign regs_460_clock = clock; // @[:@40852.4]
  assign regs_460_reset = io_reset; // @[:@40853.4 RegFile.scala 76:16:@40860.4]
  assign regs_460_io_in = 64'h0; // @[RegFile.scala 75:16:@40859.4]
  assign regs_460_io_reset = reset; // @[RegFile.scala 78:19:@40863.4]
  assign regs_460_io_enable = 1'h1; // @[RegFile.scala 74:20:@40857.4]
  assign regs_461_clock = clock; // @[:@40866.4]
  assign regs_461_reset = io_reset; // @[:@40867.4 RegFile.scala 76:16:@40874.4]
  assign regs_461_io_in = 64'h0; // @[RegFile.scala 75:16:@40873.4]
  assign regs_461_io_reset = reset; // @[RegFile.scala 78:19:@40877.4]
  assign regs_461_io_enable = 1'h1; // @[RegFile.scala 74:20:@40871.4]
  assign regs_462_clock = clock; // @[:@40880.4]
  assign regs_462_reset = io_reset; // @[:@40881.4 RegFile.scala 76:16:@40888.4]
  assign regs_462_io_in = 64'h0; // @[RegFile.scala 75:16:@40887.4]
  assign regs_462_io_reset = reset; // @[RegFile.scala 78:19:@40891.4]
  assign regs_462_io_enable = 1'h1; // @[RegFile.scala 74:20:@40885.4]
  assign regs_463_clock = clock; // @[:@40894.4]
  assign regs_463_reset = io_reset; // @[:@40895.4 RegFile.scala 76:16:@40902.4]
  assign regs_463_io_in = 64'h0; // @[RegFile.scala 75:16:@40901.4]
  assign regs_463_io_reset = reset; // @[RegFile.scala 78:19:@40905.4]
  assign regs_463_io_enable = 1'h1; // @[RegFile.scala 74:20:@40899.4]
  assign regs_464_clock = clock; // @[:@40908.4]
  assign regs_464_reset = io_reset; // @[:@40909.4 RegFile.scala 76:16:@40916.4]
  assign regs_464_io_in = 64'h0; // @[RegFile.scala 75:16:@40915.4]
  assign regs_464_io_reset = reset; // @[RegFile.scala 78:19:@40919.4]
  assign regs_464_io_enable = 1'h1; // @[RegFile.scala 74:20:@40913.4]
  assign regs_465_clock = clock; // @[:@40922.4]
  assign regs_465_reset = io_reset; // @[:@40923.4 RegFile.scala 76:16:@40930.4]
  assign regs_465_io_in = 64'h0; // @[RegFile.scala 75:16:@40929.4]
  assign regs_465_io_reset = reset; // @[RegFile.scala 78:19:@40933.4]
  assign regs_465_io_enable = 1'h1; // @[RegFile.scala 74:20:@40927.4]
  assign regs_466_clock = clock; // @[:@40936.4]
  assign regs_466_reset = io_reset; // @[:@40937.4 RegFile.scala 76:16:@40944.4]
  assign regs_466_io_in = 64'h0; // @[RegFile.scala 75:16:@40943.4]
  assign regs_466_io_reset = reset; // @[RegFile.scala 78:19:@40947.4]
  assign regs_466_io_enable = 1'h1; // @[RegFile.scala 74:20:@40941.4]
  assign regs_467_clock = clock; // @[:@40950.4]
  assign regs_467_reset = io_reset; // @[:@40951.4 RegFile.scala 76:16:@40958.4]
  assign regs_467_io_in = 64'h0; // @[RegFile.scala 75:16:@40957.4]
  assign regs_467_io_reset = reset; // @[RegFile.scala 78:19:@40961.4]
  assign regs_467_io_enable = 1'h1; // @[RegFile.scala 74:20:@40955.4]
  assign regs_468_clock = clock; // @[:@40964.4]
  assign regs_468_reset = io_reset; // @[:@40965.4 RegFile.scala 76:16:@40972.4]
  assign regs_468_io_in = 64'h0; // @[RegFile.scala 75:16:@40971.4]
  assign regs_468_io_reset = reset; // @[RegFile.scala 78:19:@40975.4]
  assign regs_468_io_enable = 1'h1; // @[RegFile.scala 74:20:@40969.4]
  assign regs_469_clock = clock; // @[:@40978.4]
  assign regs_469_reset = io_reset; // @[:@40979.4 RegFile.scala 76:16:@40986.4]
  assign regs_469_io_in = 64'h0; // @[RegFile.scala 75:16:@40985.4]
  assign regs_469_io_reset = reset; // @[RegFile.scala 78:19:@40989.4]
  assign regs_469_io_enable = 1'h1; // @[RegFile.scala 74:20:@40983.4]
  assign regs_470_clock = clock; // @[:@40992.4]
  assign regs_470_reset = io_reset; // @[:@40993.4 RegFile.scala 76:16:@41000.4]
  assign regs_470_io_in = 64'h0; // @[RegFile.scala 75:16:@40999.4]
  assign regs_470_io_reset = reset; // @[RegFile.scala 78:19:@41003.4]
  assign regs_470_io_enable = 1'h1; // @[RegFile.scala 74:20:@40997.4]
  assign regs_471_clock = clock; // @[:@41006.4]
  assign regs_471_reset = io_reset; // @[:@41007.4 RegFile.scala 76:16:@41014.4]
  assign regs_471_io_in = 64'h0; // @[RegFile.scala 75:16:@41013.4]
  assign regs_471_io_reset = reset; // @[RegFile.scala 78:19:@41017.4]
  assign regs_471_io_enable = 1'h1; // @[RegFile.scala 74:20:@41011.4]
  assign regs_472_clock = clock; // @[:@41020.4]
  assign regs_472_reset = io_reset; // @[:@41021.4 RegFile.scala 76:16:@41028.4]
  assign regs_472_io_in = 64'h0; // @[RegFile.scala 75:16:@41027.4]
  assign regs_472_io_reset = reset; // @[RegFile.scala 78:19:@41031.4]
  assign regs_472_io_enable = 1'h1; // @[RegFile.scala 74:20:@41025.4]
  assign regs_473_clock = clock; // @[:@41034.4]
  assign regs_473_reset = io_reset; // @[:@41035.4 RegFile.scala 76:16:@41042.4]
  assign regs_473_io_in = 64'h0; // @[RegFile.scala 75:16:@41041.4]
  assign regs_473_io_reset = reset; // @[RegFile.scala 78:19:@41045.4]
  assign regs_473_io_enable = 1'h1; // @[RegFile.scala 74:20:@41039.4]
  assign regs_474_clock = clock; // @[:@41048.4]
  assign regs_474_reset = io_reset; // @[:@41049.4 RegFile.scala 76:16:@41056.4]
  assign regs_474_io_in = 64'h0; // @[RegFile.scala 75:16:@41055.4]
  assign regs_474_io_reset = reset; // @[RegFile.scala 78:19:@41059.4]
  assign regs_474_io_enable = 1'h1; // @[RegFile.scala 74:20:@41053.4]
  assign regs_475_clock = clock; // @[:@41062.4]
  assign regs_475_reset = io_reset; // @[:@41063.4 RegFile.scala 76:16:@41070.4]
  assign regs_475_io_in = 64'h0; // @[RegFile.scala 75:16:@41069.4]
  assign regs_475_io_reset = reset; // @[RegFile.scala 78:19:@41073.4]
  assign regs_475_io_enable = 1'h1; // @[RegFile.scala 74:20:@41067.4]
  assign regs_476_clock = clock; // @[:@41076.4]
  assign regs_476_reset = io_reset; // @[:@41077.4 RegFile.scala 76:16:@41084.4]
  assign regs_476_io_in = 64'h0; // @[RegFile.scala 75:16:@41083.4]
  assign regs_476_io_reset = reset; // @[RegFile.scala 78:19:@41087.4]
  assign regs_476_io_enable = 1'h1; // @[RegFile.scala 74:20:@41081.4]
  assign regs_477_clock = clock; // @[:@41090.4]
  assign regs_477_reset = io_reset; // @[:@41091.4 RegFile.scala 76:16:@41098.4]
  assign regs_477_io_in = 64'h0; // @[RegFile.scala 75:16:@41097.4]
  assign regs_477_io_reset = reset; // @[RegFile.scala 78:19:@41101.4]
  assign regs_477_io_enable = 1'h1; // @[RegFile.scala 74:20:@41095.4]
  assign regs_478_clock = clock; // @[:@41104.4]
  assign regs_478_reset = io_reset; // @[:@41105.4 RegFile.scala 76:16:@41112.4]
  assign regs_478_io_in = 64'h0; // @[RegFile.scala 75:16:@41111.4]
  assign regs_478_io_reset = reset; // @[RegFile.scala 78:19:@41115.4]
  assign regs_478_io_enable = 1'h1; // @[RegFile.scala 74:20:@41109.4]
  assign regs_479_clock = clock; // @[:@41118.4]
  assign regs_479_reset = io_reset; // @[:@41119.4 RegFile.scala 76:16:@41126.4]
  assign regs_479_io_in = 64'h0; // @[RegFile.scala 75:16:@41125.4]
  assign regs_479_io_reset = reset; // @[RegFile.scala 78:19:@41129.4]
  assign regs_479_io_enable = 1'h1; // @[RegFile.scala 74:20:@41123.4]
  assign regs_480_clock = clock; // @[:@41132.4]
  assign regs_480_reset = io_reset; // @[:@41133.4 RegFile.scala 76:16:@41140.4]
  assign regs_480_io_in = 64'h0; // @[RegFile.scala 75:16:@41139.4]
  assign regs_480_io_reset = reset; // @[RegFile.scala 78:19:@41143.4]
  assign regs_480_io_enable = 1'h1; // @[RegFile.scala 74:20:@41137.4]
  assign regs_481_clock = clock; // @[:@41146.4]
  assign regs_481_reset = io_reset; // @[:@41147.4 RegFile.scala 76:16:@41154.4]
  assign regs_481_io_in = 64'h0; // @[RegFile.scala 75:16:@41153.4]
  assign regs_481_io_reset = reset; // @[RegFile.scala 78:19:@41157.4]
  assign regs_481_io_enable = 1'h1; // @[RegFile.scala 74:20:@41151.4]
  assign regs_482_clock = clock; // @[:@41160.4]
  assign regs_482_reset = io_reset; // @[:@41161.4 RegFile.scala 76:16:@41168.4]
  assign regs_482_io_in = 64'h0; // @[RegFile.scala 75:16:@41167.4]
  assign regs_482_io_reset = reset; // @[RegFile.scala 78:19:@41171.4]
  assign regs_482_io_enable = 1'h1; // @[RegFile.scala 74:20:@41165.4]
  assign regs_483_clock = clock; // @[:@41174.4]
  assign regs_483_reset = io_reset; // @[:@41175.4 RegFile.scala 76:16:@41182.4]
  assign regs_483_io_in = 64'h0; // @[RegFile.scala 75:16:@41181.4]
  assign regs_483_io_reset = reset; // @[RegFile.scala 78:19:@41185.4]
  assign regs_483_io_enable = 1'h1; // @[RegFile.scala 74:20:@41179.4]
  assign regs_484_clock = clock; // @[:@41188.4]
  assign regs_484_reset = io_reset; // @[:@41189.4 RegFile.scala 76:16:@41196.4]
  assign regs_484_io_in = 64'h0; // @[RegFile.scala 75:16:@41195.4]
  assign regs_484_io_reset = reset; // @[RegFile.scala 78:19:@41199.4]
  assign regs_484_io_enable = 1'h1; // @[RegFile.scala 74:20:@41193.4]
  assign regs_485_clock = clock; // @[:@41202.4]
  assign regs_485_reset = io_reset; // @[:@41203.4 RegFile.scala 76:16:@41210.4]
  assign regs_485_io_in = 64'h0; // @[RegFile.scala 75:16:@41209.4]
  assign regs_485_io_reset = reset; // @[RegFile.scala 78:19:@41213.4]
  assign regs_485_io_enable = 1'h1; // @[RegFile.scala 74:20:@41207.4]
  assign regs_486_clock = clock; // @[:@41216.4]
  assign regs_486_reset = io_reset; // @[:@41217.4 RegFile.scala 76:16:@41224.4]
  assign regs_486_io_in = 64'h0; // @[RegFile.scala 75:16:@41223.4]
  assign regs_486_io_reset = reset; // @[RegFile.scala 78:19:@41227.4]
  assign regs_486_io_enable = 1'h1; // @[RegFile.scala 74:20:@41221.4]
  assign regs_487_clock = clock; // @[:@41230.4]
  assign regs_487_reset = io_reset; // @[:@41231.4 RegFile.scala 76:16:@41238.4]
  assign regs_487_io_in = 64'h0; // @[RegFile.scala 75:16:@41237.4]
  assign regs_487_io_reset = reset; // @[RegFile.scala 78:19:@41241.4]
  assign regs_487_io_enable = 1'h1; // @[RegFile.scala 74:20:@41235.4]
  assign regs_488_clock = clock; // @[:@41244.4]
  assign regs_488_reset = io_reset; // @[:@41245.4 RegFile.scala 76:16:@41252.4]
  assign regs_488_io_in = 64'h0; // @[RegFile.scala 75:16:@41251.4]
  assign regs_488_io_reset = reset; // @[RegFile.scala 78:19:@41255.4]
  assign regs_488_io_enable = 1'h1; // @[RegFile.scala 74:20:@41249.4]
  assign regs_489_clock = clock; // @[:@41258.4]
  assign regs_489_reset = io_reset; // @[:@41259.4 RegFile.scala 76:16:@41266.4]
  assign regs_489_io_in = 64'h0; // @[RegFile.scala 75:16:@41265.4]
  assign regs_489_io_reset = reset; // @[RegFile.scala 78:19:@41269.4]
  assign regs_489_io_enable = 1'h1; // @[RegFile.scala 74:20:@41263.4]
  assign regs_490_clock = clock; // @[:@41272.4]
  assign regs_490_reset = io_reset; // @[:@41273.4 RegFile.scala 76:16:@41280.4]
  assign regs_490_io_in = 64'h0; // @[RegFile.scala 75:16:@41279.4]
  assign regs_490_io_reset = reset; // @[RegFile.scala 78:19:@41283.4]
  assign regs_490_io_enable = 1'h1; // @[RegFile.scala 74:20:@41277.4]
  assign regs_491_clock = clock; // @[:@41286.4]
  assign regs_491_reset = io_reset; // @[:@41287.4 RegFile.scala 76:16:@41294.4]
  assign regs_491_io_in = 64'h0; // @[RegFile.scala 75:16:@41293.4]
  assign regs_491_io_reset = reset; // @[RegFile.scala 78:19:@41297.4]
  assign regs_491_io_enable = 1'h1; // @[RegFile.scala 74:20:@41291.4]
  assign regs_492_clock = clock; // @[:@41300.4]
  assign regs_492_reset = io_reset; // @[:@41301.4 RegFile.scala 76:16:@41308.4]
  assign regs_492_io_in = 64'h0; // @[RegFile.scala 75:16:@41307.4]
  assign regs_492_io_reset = reset; // @[RegFile.scala 78:19:@41311.4]
  assign regs_492_io_enable = 1'h1; // @[RegFile.scala 74:20:@41305.4]
  assign regs_493_clock = clock; // @[:@41314.4]
  assign regs_493_reset = io_reset; // @[:@41315.4 RegFile.scala 76:16:@41322.4]
  assign regs_493_io_in = 64'h0; // @[RegFile.scala 75:16:@41321.4]
  assign regs_493_io_reset = reset; // @[RegFile.scala 78:19:@41325.4]
  assign regs_493_io_enable = 1'h1; // @[RegFile.scala 74:20:@41319.4]
  assign regs_494_clock = clock; // @[:@41328.4]
  assign regs_494_reset = io_reset; // @[:@41329.4 RegFile.scala 76:16:@41336.4]
  assign regs_494_io_in = 64'h0; // @[RegFile.scala 75:16:@41335.4]
  assign regs_494_io_reset = reset; // @[RegFile.scala 78:19:@41339.4]
  assign regs_494_io_enable = 1'h1; // @[RegFile.scala 74:20:@41333.4]
  assign regs_495_clock = clock; // @[:@41342.4]
  assign regs_495_reset = io_reset; // @[:@41343.4 RegFile.scala 76:16:@41350.4]
  assign regs_495_io_in = 64'h0; // @[RegFile.scala 75:16:@41349.4]
  assign regs_495_io_reset = reset; // @[RegFile.scala 78:19:@41353.4]
  assign regs_495_io_enable = 1'h1; // @[RegFile.scala 74:20:@41347.4]
  assign regs_496_clock = clock; // @[:@41356.4]
  assign regs_496_reset = io_reset; // @[:@41357.4 RegFile.scala 76:16:@41364.4]
  assign regs_496_io_in = 64'h0; // @[RegFile.scala 75:16:@41363.4]
  assign regs_496_io_reset = reset; // @[RegFile.scala 78:19:@41367.4]
  assign regs_496_io_enable = 1'h1; // @[RegFile.scala 74:20:@41361.4]
  assign regs_497_clock = clock; // @[:@41370.4]
  assign regs_497_reset = io_reset; // @[:@41371.4 RegFile.scala 76:16:@41378.4]
  assign regs_497_io_in = 64'h0; // @[RegFile.scala 75:16:@41377.4]
  assign regs_497_io_reset = reset; // @[RegFile.scala 78:19:@41381.4]
  assign regs_497_io_enable = 1'h1; // @[RegFile.scala 74:20:@41375.4]
  assign regs_498_clock = clock; // @[:@41384.4]
  assign regs_498_reset = io_reset; // @[:@41385.4 RegFile.scala 76:16:@41392.4]
  assign regs_498_io_in = 64'h0; // @[RegFile.scala 75:16:@41391.4]
  assign regs_498_io_reset = reset; // @[RegFile.scala 78:19:@41395.4]
  assign regs_498_io_enable = 1'h1; // @[RegFile.scala 74:20:@41389.4]
  assign regs_499_clock = clock; // @[:@41398.4]
  assign regs_499_reset = io_reset; // @[:@41399.4 RegFile.scala 76:16:@41406.4]
  assign regs_499_io_in = 64'h0; // @[RegFile.scala 75:16:@41405.4]
  assign regs_499_io_reset = reset; // @[RegFile.scala 78:19:@41409.4]
  assign regs_499_io_enable = 1'h1; // @[RegFile.scala 74:20:@41403.4]
  assign regs_500_clock = clock; // @[:@41412.4]
  assign regs_500_reset = io_reset; // @[:@41413.4 RegFile.scala 76:16:@41420.4]
  assign regs_500_io_in = 64'h0; // @[RegFile.scala 75:16:@41419.4]
  assign regs_500_io_reset = reset; // @[RegFile.scala 78:19:@41423.4]
  assign regs_500_io_enable = 1'h1; // @[RegFile.scala 74:20:@41417.4]
  assign regs_501_clock = clock; // @[:@41426.4]
  assign regs_501_reset = io_reset; // @[:@41427.4 RegFile.scala 76:16:@41434.4]
  assign regs_501_io_in = 64'h0; // @[RegFile.scala 75:16:@41433.4]
  assign regs_501_io_reset = reset; // @[RegFile.scala 78:19:@41437.4]
  assign regs_501_io_enable = 1'h1; // @[RegFile.scala 74:20:@41431.4]
  assign regs_502_clock = clock; // @[:@41440.4]
  assign regs_502_reset = io_reset; // @[:@41441.4 RegFile.scala 76:16:@41448.4]
  assign regs_502_io_in = 64'h0; // @[RegFile.scala 75:16:@41447.4]
  assign regs_502_io_reset = reset; // @[RegFile.scala 78:19:@41451.4]
  assign regs_502_io_enable = 1'h1; // @[RegFile.scala 74:20:@41445.4]
  assign rport_io_ins_0 = regs_0_io_out; // @[RegFile.scala 97:16:@41960.4]
  assign rport_io_ins_1 = regs_1_io_out; // @[RegFile.scala 97:16:@41961.4]
  assign rport_io_ins_2 = regs_2_io_out; // @[RegFile.scala 97:16:@41962.4]
  assign rport_io_ins_3 = regs_3_io_out; // @[RegFile.scala 97:16:@41963.4]
  assign rport_io_ins_4 = regs_4_io_out; // @[RegFile.scala 97:16:@41964.4]
  assign rport_io_ins_5 = regs_5_io_out; // @[RegFile.scala 97:16:@41965.4]
  assign rport_io_ins_6 = regs_6_io_out; // @[RegFile.scala 97:16:@41966.4]
  assign rport_io_ins_7 = regs_7_io_out; // @[RegFile.scala 97:16:@41967.4]
  assign rport_io_ins_8 = regs_8_io_out; // @[RegFile.scala 97:16:@41968.4]
  assign rport_io_ins_9 = regs_9_io_out; // @[RegFile.scala 97:16:@41969.4]
  assign rport_io_ins_10 = regs_10_io_out; // @[RegFile.scala 97:16:@41970.4]
  assign rport_io_ins_11 = regs_11_io_out; // @[RegFile.scala 97:16:@41971.4]
  assign rport_io_ins_12 = regs_12_io_out; // @[RegFile.scala 97:16:@41972.4]
  assign rport_io_ins_13 = regs_13_io_out; // @[RegFile.scala 97:16:@41973.4]
  assign rport_io_ins_14 = regs_14_io_out; // @[RegFile.scala 97:16:@41974.4]
  assign rport_io_ins_15 = regs_15_io_out; // @[RegFile.scala 97:16:@41975.4]
  assign rport_io_ins_16 = regs_16_io_out; // @[RegFile.scala 97:16:@41976.4]
  assign rport_io_ins_17 = regs_17_io_out; // @[RegFile.scala 97:16:@41977.4]
  assign rport_io_ins_18 = regs_18_io_out; // @[RegFile.scala 97:16:@41978.4]
  assign rport_io_ins_19 = regs_19_io_out; // @[RegFile.scala 97:16:@41979.4]
  assign rport_io_ins_20 = regs_20_io_out; // @[RegFile.scala 97:16:@41980.4]
  assign rport_io_ins_21 = regs_21_io_out; // @[RegFile.scala 97:16:@41981.4]
  assign rport_io_ins_22 = regs_22_io_out; // @[RegFile.scala 97:16:@41982.4]
  assign rport_io_ins_23 = regs_23_io_out; // @[RegFile.scala 97:16:@41983.4]
  assign rport_io_ins_24 = regs_24_io_out; // @[RegFile.scala 97:16:@41984.4]
  assign rport_io_ins_25 = regs_25_io_out; // @[RegFile.scala 97:16:@41985.4]
  assign rport_io_ins_26 = regs_26_io_out; // @[RegFile.scala 97:16:@41986.4]
  assign rport_io_ins_27 = regs_27_io_out; // @[RegFile.scala 97:16:@41987.4]
  assign rport_io_ins_28 = regs_28_io_out; // @[RegFile.scala 97:16:@41988.4]
  assign rport_io_ins_29 = regs_29_io_out; // @[RegFile.scala 97:16:@41989.4]
  assign rport_io_ins_30 = regs_30_io_out; // @[RegFile.scala 97:16:@41990.4]
  assign rport_io_ins_31 = regs_31_io_out; // @[RegFile.scala 97:16:@41991.4]
  assign rport_io_ins_32 = regs_32_io_out; // @[RegFile.scala 97:16:@41992.4]
  assign rport_io_ins_33 = regs_33_io_out; // @[RegFile.scala 97:16:@41993.4]
  assign rport_io_ins_34 = regs_34_io_out; // @[RegFile.scala 97:16:@41994.4]
  assign rport_io_ins_35 = regs_35_io_out; // @[RegFile.scala 97:16:@41995.4]
  assign rport_io_ins_36 = regs_36_io_out; // @[RegFile.scala 97:16:@41996.4]
  assign rport_io_ins_37 = regs_37_io_out; // @[RegFile.scala 97:16:@41997.4]
  assign rport_io_ins_38 = regs_38_io_out; // @[RegFile.scala 97:16:@41998.4]
  assign rport_io_ins_39 = regs_39_io_out; // @[RegFile.scala 97:16:@41999.4]
  assign rport_io_ins_40 = regs_40_io_out; // @[RegFile.scala 97:16:@42000.4]
  assign rport_io_ins_41 = regs_41_io_out; // @[RegFile.scala 97:16:@42001.4]
  assign rport_io_ins_42 = regs_42_io_out; // @[RegFile.scala 97:16:@42002.4]
  assign rport_io_ins_43 = regs_43_io_out; // @[RegFile.scala 97:16:@42003.4]
  assign rport_io_ins_44 = regs_44_io_out; // @[RegFile.scala 97:16:@42004.4]
  assign rport_io_ins_45 = regs_45_io_out; // @[RegFile.scala 97:16:@42005.4]
  assign rport_io_ins_46 = regs_46_io_out; // @[RegFile.scala 97:16:@42006.4]
  assign rport_io_ins_47 = regs_47_io_out; // @[RegFile.scala 97:16:@42007.4]
  assign rport_io_ins_48 = regs_48_io_out; // @[RegFile.scala 97:16:@42008.4]
  assign rport_io_ins_49 = regs_49_io_out; // @[RegFile.scala 97:16:@42009.4]
  assign rport_io_ins_50 = regs_50_io_out; // @[RegFile.scala 97:16:@42010.4]
  assign rport_io_ins_51 = regs_51_io_out; // @[RegFile.scala 97:16:@42011.4]
  assign rport_io_ins_52 = regs_52_io_out; // @[RegFile.scala 97:16:@42012.4]
  assign rport_io_ins_53 = regs_53_io_out; // @[RegFile.scala 97:16:@42013.4]
  assign rport_io_ins_54 = regs_54_io_out; // @[RegFile.scala 97:16:@42014.4]
  assign rport_io_ins_55 = regs_55_io_out; // @[RegFile.scala 97:16:@42015.4]
  assign rport_io_ins_56 = regs_56_io_out; // @[RegFile.scala 97:16:@42016.4]
  assign rport_io_ins_57 = regs_57_io_out; // @[RegFile.scala 97:16:@42017.4]
  assign rport_io_ins_58 = regs_58_io_out; // @[RegFile.scala 97:16:@42018.4]
  assign rport_io_ins_59 = regs_59_io_out; // @[RegFile.scala 97:16:@42019.4]
  assign rport_io_ins_60 = regs_60_io_out; // @[RegFile.scala 97:16:@42020.4]
  assign rport_io_ins_61 = regs_61_io_out; // @[RegFile.scala 97:16:@42021.4]
  assign rport_io_ins_62 = regs_62_io_out; // @[RegFile.scala 97:16:@42022.4]
  assign rport_io_ins_63 = regs_63_io_out; // @[RegFile.scala 97:16:@42023.4]
  assign rport_io_ins_64 = regs_64_io_out; // @[RegFile.scala 97:16:@42024.4]
  assign rport_io_ins_65 = regs_65_io_out; // @[RegFile.scala 97:16:@42025.4]
  assign rport_io_ins_66 = regs_66_io_out; // @[RegFile.scala 97:16:@42026.4]
  assign rport_io_ins_67 = regs_67_io_out; // @[RegFile.scala 97:16:@42027.4]
  assign rport_io_ins_68 = regs_68_io_out; // @[RegFile.scala 97:16:@42028.4]
  assign rport_io_ins_69 = regs_69_io_out; // @[RegFile.scala 97:16:@42029.4]
  assign rport_io_ins_70 = regs_70_io_out; // @[RegFile.scala 97:16:@42030.4]
  assign rport_io_ins_71 = regs_71_io_out; // @[RegFile.scala 97:16:@42031.4]
  assign rport_io_ins_72 = regs_72_io_out; // @[RegFile.scala 97:16:@42032.4]
  assign rport_io_ins_73 = regs_73_io_out; // @[RegFile.scala 97:16:@42033.4]
  assign rport_io_ins_74 = regs_74_io_out; // @[RegFile.scala 97:16:@42034.4]
  assign rport_io_ins_75 = regs_75_io_out; // @[RegFile.scala 97:16:@42035.4]
  assign rport_io_ins_76 = regs_76_io_out; // @[RegFile.scala 97:16:@42036.4]
  assign rport_io_ins_77 = regs_77_io_out; // @[RegFile.scala 97:16:@42037.4]
  assign rport_io_ins_78 = regs_78_io_out; // @[RegFile.scala 97:16:@42038.4]
  assign rport_io_ins_79 = regs_79_io_out; // @[RegFile.scala 97:16:@42039.4]
  assign rport_io_ins_80 = regs_80_io_out; // @[RegFile.scala 97:16:@42040.4]
  assign rport_io_ins_81 = regs_81_io_out; // @[RegFile.scala 97:16:@42041.4]
  assign rport_io_ins_82 = regs_82_io_out; // @[RegFile.scala 97:16:@42042.4]
  assign rport_io_ins_83 = regs_83_io_out; // @[RegFile.scala 97:16:@42043.4]
  assign rport_io_ins_84 = regs_84_io_out; // @[RegFile.scala 97:16:@42044.4]
  assign rport_io_ins_85 = regs_85_io_out; // @[RegFile.scala 97:16:@42045.4]
  assign rport_io_ins_86 = regs_86_io_out; // @[RegFile.scala 97:16:@42046.4]
  assign rport_io_ins_87 = regs_87_io_out; // @[RegFile.scala 97:16:@42047.4]
  assign rport_io_ins_88 = regs_88_io_out; // @[RegFile.scala 97:16:@42048.4]
  assign rport_io_ins_89 = regs_89_io_out; // @[RegFile.scala 97:16:@42049.4]
  assign rport_io_ins_90 = regs_90_io_out; // @[RegFile.scala 97:16:@42050.4]
  assign rport_io_ins_91 = regs_91_io_out; // @[RegFile.scala 97:16:@42051.4]
  assign rport_io_ins_92 = regs_92_io_out; // @[RegFile.scala 97:16:@42052.4]
  assign rport_io_ins_93 = regs_93_io_out; // @[RegFile.scala 97:16:@42053.4]
  assign rport_io_ins_94 = regs_94_io_out; // @[RegFile.scala 97:16:@42054.4]
  assign rport_io_ins_95 = regs_95_io_out; // @[RegFile.scala 97:16:@42055.4]
  assign rport_io_ins_96 = regs_96_io_out; // @[RegFile.scala 97:16:@42056.4]
  assign rport_io_ins_97 = regs_97_io_out; // @[RegFile.scala 97:16:@42057.4]
  assign rport_io_ins_98 = regs_98_io_out; // @[RegFile.scala 97:16:@42058.4]
  assign rport_io_ins_99 = regs_99_io_out; // @[RegFile.scala 97:16:@42059.4]
  assign rport_io_ins_100 = regs_100_io_out; // @[RegFile.scala 97:16:@42060.4]
  assign rport_io_ins_101 = regs_101_io_out; // @[RegFile.scala 97:16:@42061.4]
  assign rport_io_ins_102 = regs_102_io_out; // @[RegFile.scala 97:16:@42062.4]
  assign rport_io_ins_103 = regs_103_io_out; // @[RegFile.scala 97:16:@42063.4]
  assign rport_io_ins_104 = regs_104_io_out; // @[RegFile.scala 97:16:@42064.4]
  assign rport_io_ins_105 = regs_105_io_out; // @[RegFile.scala 97:16:@42065.4]
  assign rport_io_ins_106 = regs_106_io_out; // @[RegFile.scala 97:16:@42066.4]
  assign rport_io_ins_107 = regs_107_io_out; // @[RegFile.scala 97:16:@42067.4]
  assign rport_io_ins_108 = regs_108_io_out; // @[RegFile.scala 97:16:@42068.4]
  assign rport_io_ins_109 = regs_109_io_out; // @[RegFile.scala 97:16:@42069.4]
  assign rport_io_ins_110 = regs_110_io_out; // @[RegFile.scala 97:16:@42070.4]
  assign rport_io_ins_111 = regs_111_io_out; // @[RegFile.scala 97:16:@42071.4]
  assign rport_io_ins_112 = regs_112_io_out; // @[RegFile.scala 97:16:@42072.4]
  assign rport_io_ins_113 = regs_113_io_out; // @[RegFile.scala 97:16:@42073.4]
  assign rport_io_ins_114 = regs_114_io_out; // @[RegFile.scala 97:16:@42074.4]
  assign rport_io_ins_115 = regs_115_io_out; // @[RegFile.scala 97:16:@42075.4]
  assign rport_io_ins_116 = regs_116_io_out; // @[RegFile.scala 97:16:@42076.4]
  assign rport_io_ins_117 = regs_117_io_out; // @[RegFile.scala 97:16:@42077.4]
  assign rport_io_ins_118 = regs_118_io_out; // @[RegFile.scala 97:16:@42078.4]
  assign rport_io_ins_119 = regs_119_io_out; // @[RegFile.scala 97:16:@42079.4]
  assign rport_io_ins_120 = regs_120_io_out; // @[RegFile.scala 97:16:@42080.4]
  assign rport_io_ins_121 = regs_121_io_out; // @[RegFile.scala 97:16:@42081.4]
  assign rport_io_ins_122 = regs_122_io_out; // @[RegFile.scala 97:16:@42082.4]
  assign rport_io_ins_123 = regs_123_io_out; // @[RegFile.scala 97:16:@42083.4]
  assign rport_io_ins_124 = regs_124_io_out; // @[RegFile.scala 97:16:@42084.4]
  assign rport_io_ins_125 = regs_125_io_out; // @[RegFile.scala 97:16:@42085.4]
  assign rport_io_ins_126 = regs_126_io_out; // @[RegFile.scala 97:16:@42086.4]
  assign rport_io_ins_127 = regs_127_io_out; // @[RegFile.scala 97:16:@42087.4]
  assign rport_io_ins_128 = regs_128_io_out; // @[RegFile.scala 97:16:@42088.4]
  assign rport_io_ins_129 = regs_129_io_out; // @[RegFile.scala 97:16:@42089.4]
  assign rport_io_ins_130 = regs_130_io_out; // @[RegFile.scala 97:16:@42090.4]
  assign rport_io_ins_131 = regs_131_io_out; // @[RegFile.scala 97:16:@42091.4]
  assign rport_io_ins_132 = regs_132_io_out; // @[RegFile.scala 97:16:@42092.4]
  assign rport_io_ins_133 = regs_133_io_out; // @[RegFile.scala 97:16:@42093.4]
  assign rport_io_ins_134 = regs_134_io_out; // @[RegFile.scala 97:16:@42094.4]
  assign rport_io_ins_135 = regs_135_io_out; // @[RegFile.scala 97:16:@42095.4]
  assign rport_io_ins_136 = regs_136_io_out; // @[RegFile.scala 97:16:@42096.4]
  assign rport_io_ins_137 = regs_137_io_out; // @[RegFile.scala 97:16:@42097.4]
  assign rport_io_ins_138 = regs_138_io_out; // @[RegFile.scala 97:16:@42098.4]
  assign rport_io_ins_139 = regs_139_io_out; // @[RegFile.scala 97:16:@42099.4]
  assign rport_io_ins_140 = regs_140_io_out; // @[RegFile.scala 97:16:@42100.4]
  assign rport_io_ins_141 = regs_141_io_out; // @[RegFile.scala 97:16:@42101.4]
  assign rport_io_ins_142 = regs_142_io_out; // @[RegFile.scala 97:16:@42102.4]
  assign rport_io_ins_143 = regs_143_io_out; // @[RegFile.scala 97:16:@42103.4]
  assign rport_io_ins_144 = regs_144_io_out; // @[RegFile.scala 97:16:@42104.4]
  assign rport_io_ins_145 = regs_145_io_out; // @[RegFile.scala 97:16:@42105.4]
  assign rport_io_ins_146 = regs_146_io_out; // @[RegFile.scala 97:16:@42106.4]
  assign rport_io_ins_147 = regs_147_io_out; // @[RegFile.scala 97:16:@42107.4]
  assign rport_io_ins_148 = regs_148_io_out; // @[RegFile.scala 97:16:@42108.4]
  assign rport_io_ins_149 = regs_149_io_out; // @[RegFile.scala 97:16:@42109.4]
  assign rport_io_ins_150 = regs_150_io_out; // @[RegFile.scala 97:16:@42110.4]
  assign rport_io_ins_151 = regs_151_io_out; // @[RegFile.scala 97:16:@42111.4]
  assign rport_io_ins_152 = regs_152_io_out; // @[RegFile.scala 97:16:@42112.4]
  assign rport_io_ins_153 = regs_153_io_out; // @[RegFile.scala 97:16:@42113.4]
  assign rport_io_ins_154 = regs_154_io_out; // @[RegFile.scala 97:16:@42114.4]
  assign rport_io_ins_155 = regs_155_io_out; // @[RegFile.scala 97:16:@42115.4]
  assign rport_io_ins_156 = regs_156_io_out; // @[RegFile.scala 97:16:@42116.4]
  assign rport_io_ins_157 = regs_157_io_out; // @[RegFile.scala 97:16:@42117.4]
  assign rport_io_ins_158 = regs_158_io_out; // @[RegFile.scala 97:16:@42118.4]
  assign rport_io_ins_159 = regs_159_io_out; // @[RegFile.scala 97:16:@42119.4]
  assign rport_io_ins_160 = regs_160_io_out; // @[RegFile.scala 97:16:@42120.4]
  assign rport_io_ins_161 = regs_161_io_out; // @[RegFile.scala 97:16:@42121.4]
  assign rport_io_ins_162 = regs_162_io_out; // @[RegFile.scala 97:16:@42122.4]
  assign rport_io_ins_163 = regs_163_io_out; // @[RegFile.scala 97:16:@42123.4]
  assign rport_io_ins_164 = regs_164_io_out; // @[RegFile.scala 97:16:@42124.4]
  assign rport_io_ins_165 = regs_165_io_out; // @[RegFile.scala 97:16:@42125.4]
  assign rport_io_ins_166 = regs_166_io_out; // @[RegFile.scala 97:16:@42126.4]
  assign rport_io_ins_167 = regs_167_io_out; // @[RegFile.scala 97:16:@42127.4]
  assign rport_io_ins_168 = regs_168_io_out; // @[RegFile.scala 97:16:@42128.4]
  assign rport_io_ins_169 = regs_169_io_out; // @[RegFile.scala 97:16:@42129.4]
  assign rport_io_ins_170 = regs_170_io_out; // @[RegFile.scala 97:16:@42130.4]
  assign rport_io_ins_171 = regs_171_io_out; // @[RegFile.scala 97:16:@42131.4]
  assign rport_io_ins_172 = regs_172_io_out; // @[RegFile.scala 97:16:@42132.4]
  assign rport_io_ins_173 = regs_173_io_out; // @[RegFile.scala 97:16:@42133.4]
  assign rport_io_ins_174 = regs_174_io_out; // @[RegFile.scala 97:16:@42134.4]
  assign rport_io_ins_175 = regs_175_io_out; // @[RegFile.scala 97:16:@42135.4]
  assign rport_io_ins_176 = regs_176_io_out; // @[RegFile.scala 97:16:@42136.4]
  assign rport_io_ins_177 = regs_177_io_out; // @[RegFile.scala 97:16:@42137.4]
  assign rport_io_ins_178 = regs_178_io_out; // @[RegFile.scala 97:16:@42138.4]
  assign rport_io_ins_179 = regs_179_io_out; // @[RegFile.scala 97:16:@42139.4]
  assign rport_io_ins_180 = regs_180_io_out; // @[RegFile.scala 97:16:@42140.4]
  assign rport_io_ins_181 = regs_181_io_out; // @[RegFile.scala 97:16:@42141.4]
  assign rport_io_ins_182 = regs_182_io_out; // @[RegFile.scala 97:16:@42142.4]
  assign rport_io_ins_183 = regs_183_io_out; // @[RegFile.scala 97:16:@42143.4]
  assign rport_io_ins_184 = regs_184_io_out; // @[RegFile.scala 97:16:@42144.4]
  assign rport_io_ins_185 = regs_185_io_out; // @[RegFile.scala 97:16:@42145.4]
  assign rport_io_ins_186 = regs_186_io_out; // @[RegFile.scala 97:16:@42146.4]
  assign rport_io_ins_187 = regs_187_io_out; // @[RegFile.scala 97:16:@42147.4]
  assign rport_io_ins_188 = regs_188_io_out; // @[RegFile.scala 97:16:@42148.4]
  assign rport_io_ins_189 = regs_189_io_out; // @[RegFile.scala 97:16:@42149.4]
  assign rport_io_ins_190 = regs_190_io_out; // @[RegFile.scala 97:16:@42150.4]
  assign rport_io_ins_191 = regs_191_io_out; // @[RegFile.scala 97:16:@42151.4]
  assign rport_io_ins_192 = regs_192_io_out; // @[RegFile.scala 97:16:@42152.4]
  assign rport_io_ins_193 = regs_193_io_out; // @[RegFile.scala 97:16:@42153.4]
  assign rport_io_ins_194 = regs_194_io_out; // @[RegFile.scala 97:16:@42154.4]
  assign rport_io_ins_195 = regs_195_io_out; // @[RegFile.scala 97:16:@42155.4]
  assign rport_io_ins_196 = regs_196_io_out; // @[RegFile.scala 97:16:@42156.4]
  assign rport_io_ins_197 = regs_197_io_out; // @[RegFile.scala 97:16:@42157.4]
  assign rport_io_ins_198 = regs_198_io_out; // @[RegFile.scala 97:16:@42158.4]
  assign rport_io_ins_199 = regs_199_io_out; // @[RegFile.scala 97:16:@42159.4]
  assign rport_io_ins_200 = regs_200_io_out; // @[RegFile.scala 97:16:@42160.4]
  assign rport_io_ins_201 = regs_201_io_out; // @[RegFile.scala 97:16:@42161.4]
  assign rport_io_ins_202 = regs_202_io_out; // @[RegFile.scala 97:16:@42162.4]
  assign rport_io_ins_203 = regs_203_io_out; // @[RegFile.scala 97:16:@42163.4]
  assign rport_io_ins_204 = regs_204_io_out; // @[RegFile.scala 97:16:@42164.4]
  assign rport_io_ins_205 = regs_205_io_out; // @[RegFile.scala 97:16:@42165.4]
  assign rport_io_ins_206 = regs_206_io_out; // @[RegFile.scala 97:16:@42166.4]
  assign rport_io_ins_207 = regs_207_io_out; // @[RegFile.scala 97:16:@42167.4]
  assign rport_io_ins_208 = regs_208_io_out; // @[RegFile.scala 97:16:@42168.4]
  assign rport_io_ins_209 = regs_209_io_out; // @[RegFile.scala 97:16:@42169.4]
  assign rport_io_ins_210 = regs_210_io_out; // @[RegFile.scala 97:16:@42170.4]
  assign rport_io_ins_211 = regs_211_io_out; // @[RegFile.scala 97:16:@42171.4]
  assign rport_io_ins_212 = regs_212_io_out; // @[RegFile.scala 97:16:@42172.4]
  assign rport_io_ins_213 = regs_213_io_out; // @[RegFile.scala 97:16:@42173.4]
  assign rport_io_ins_214 = regs_214_io_out; // @[RegFile.scala 97:16:@42174.4]
  assign rport_io_ins_215 = regs_215_io_out; // @[RegFile.scala 97:16:@42175.4]
  assign rport_io_ins_216 = regs_216_io_out; // @[RegFile.scala 97:16:@42176.4]
  assign rport_io_ins_217 = regs_217_io_out; // @[RegFile.scala 97:16:@42177.4]
  assign rport_io_ins_218 = regs_218_io_out; // @[RegFile.scala 97:16:@42178.4]
  assign rport_io_ins_219 = regs_219_io_out; // @[RegFile.scala 97:16:@42179.4]
  assign rport_io_ins_220 = regs_220_io_out; // @[RegFile.scala 97:16:@42180.4]
  assign rport_io_ins_221 = regs_221_io_out; // @[RegFile.scala 97:16:@42181.4]
  assign rport_io_ins_222 = regs_222_io_out; // @[RegFile.scala 97:16:@42182.4]
  assign rport_io_ins_223 = regs_223_io_out; // @[RegFile.scala 97:16:@42183.4]
  assign rport_io_ins_224 = regs_224_io_out; // @[RegFile.scala 97:16:@42184.4]
  assign rport_io_ins_225 = regs_225_io_out; // @[RegFile.scala 97:16:@42185.4]
  assign rport_io_ins_226 = regs_226_io_out; // @[RegFile.scala 97:16:@42186.4]
  assign rport_io_ins_227 = regs_227_io_out; // @[RegFile.scala 97:16:@42187.4]
  assign rport_io_ins_228 = regs_228_io_out; // @[RegFile.scala 97:16:@42188.4]
  assign rport_io_ins_229 = regs_229_io_out; // @[RegFile.scala 97:16:@42189.4]
  assign rport_io_ins_230 = regs_230_io_out; // @[RegFile.scala 97:16:@42190.4]
  assign rport_io_ins_231 = regs_231_io_out; // @[RegFile.scala 97:16:@42191.4]
  assign rport_io_ins_232 = regs_232_io_out; // @[RegFile.scala 97:16:@42192.4]
  assign rport_io_ins_233 = regs_233_io_out; // @[RegFile.scala 97:16:@42193.4]
  assign rport_io_ins_234 = regs_234_io_out; // @[RegFile.scala 97:16:@42194.4]
  assign rport_io_ins_235 = regs_235_io_out; // @[RegFile.scala 97:16:@42195.4]
  assign rport_io_ins_236 = regs_236_io_out; // @[RegFile.scala 97:16:@42196.4]
  assign rport_io_ins_237 = regs_237_io_out; // @[RegFile.scala 97:16:@42197.4]
  assign rport_io_ins_238 = regs_238_io_out; // @[RegFile.scala 97:16:@42198.4]
  assign rport_io_ins_239 = regs_239_io_out; // @[RegFile.scala 97:16:@42199.4]
  assign rport_io_ins_240 = regs_240_io_out; // @[RegFile.scala 97:16:@42200.4]
  assign rport_io_ins_241 = regs_241_io_out; // @[RegFile.scala 97:16:@42201.4]
  assign rport_io_ins_242 = regs_242_io_out; // @[RegFile.scala 97:16:@42202.4]
  assign rport_io_ins_243 = regs_243_io_out; // @[RegFile.scala 97:16:@42203.4]
  assign rport_io_ins_244 = regs_244_io_out; // @[RegFile.scala 97:16:@42204.4]
  assign rport_io_ins_245 = regs_245_io_out; // @[RegFile.scala 97:16:@42205.4]
  assign rport_io_ins_246 = regs_246_io_out; // @[RegFile.scala 97:16:@42206.4]
  assign rport_io_ins_247 = regs_247_io_out; // @[RegFile.scala 97:16:@42207.4]
  assign rport_io_ins_248 = regs_248_io_out; // @[RegFile.scala 97:16:@42208.4]
  assign rport_io_ins_249 = regs_249_io_out; // @[RegFile.scala 97:16:@42209.4]
  assign rport_io_ins_250 = regs_250_io_out; // @[RegFile.scala 97:16:@42210.4]
  assign rport_io_ins_251 = regs_251_io_out; // @[RegFile.scala 97:16:@42211.4]
  assign rport_io_ins_252 = regs_252_io_out; // @[RegFile.scala 97:16:@42212.4]
  assign rport_io_ins_253 = regs_253_io_out; // @[RegFile.scala 97:16:@42213.4]
  assign rport_io_ins_254 = regs_254_io_out; // @[RegFile.scala 97:16:@42214.4]
  assign rport_io_ins_255 = regs_255_io_out; // @[RegFile.scala 97:16:@42215.4]
  assign rport_io_ins_256 = regs_256_io_out; // @[RegFile.scala 97:16:@42216.4]
  assign rport_io_ins_257 = regs_257_io_out; // @[RegFile.scala 97:16:@42217.4]
  assign rport_io_ins_258 = regs_258_io_out; // @[RegFile.scala 97:16:@42218.4]
  assign rport_io_ins_259 = regs_259_io_out; // @[RegFile.scala 97:16:@42219.4]
  assign rport_io_ins_260 = regs_260_io_out; // @[RegFile.scala 97:16:@42220.4]
  assign rport_io_ins_261 = regs_261_io_out; // @[RegFile.scala 97:16:@42221.4]
  assign rport_io_ins_262 = regs_262_io_out; // @[RegFile.scala 97:16:@42222.4]
  assign rport_io_ins_263 = regs_263_io_out; // @[RegFile.scala 97:16:@42223.4]
  assign rport_io_ins_264 = regs_264_io_out; // @[RegFile.scala 97:16:@42224.4]
  assign rport_io_ins_265 = regs_265_io_out; // @[RegFile.scala 97:16:@42225.4]
  assign rport_io_ins_266 = regs_266_io_out; // @[RegFile.scala 97:16:@42226.4]
  assign rport_io_ins_267 = regs_267_io_out; // @[RegFile.scala 97:16:@42227.4]
  assign rport_io_ins_268 = regs_268_io_out; // @[RegFile.scala 97:16:@42228.4]
  assign rport_io_ins_269 = regs_269_io_out; // @[RegFile.scala 97:16:@42229.4]
  assign rport_io_ins_270 = regs_270_io_out; // @[RegFile.scala 97:16:@42230.4]
  assign rport_io_ins_271 = regs_271_io_out; // @[RegFile.scala 97:16:@42231.4]
  assign rport_io_ins_272 = regs_272_io_out; // @[RegFile.scala 97:16:@42232.4]
  assign rport_io_ins_273 = regs_273_io_out; // @[RegFile.scala 97:16:@42233.4]
  assign rport_io_ins_274 = regs_274_io_out; // @[RegFile.scala 97:16:@42234.4]
  assign rport_io_ins_275 = regs_275_io_out; // @[RegFile.scala 97:16:@42235.4]
  assign rport_io_ins_276 = regs_276_io_out; // @[RegFile.scala 97:16:@42236.4]
  assign rport_io_ins_277 = regs_277_io_out; // @[RegFile.scala 97:16:@42237.4]
  assign rport_io_ins_278 = regs_278_io_out; // @[RegFile.scala 97:16:@42238.4]
  assign rport_io_ins_279 = regs_279_io_out; // @[RegFile.scala 97:16:@42239.4]
  assign rport_io_ins_280 = regs_280_io_out; // @[RegFile.scala 97:16:@42240.4]
  assign rport_io_ins_281 = regs_281_io_out; // @[RegFile.scala 97:16:@42241.4]
  assign rport_io_ins_282 = regs_282_io_out; // @[RegFile.scala 97:16:@42242.4]
  assign rport_io_ins_283 = regs_283_io_out; // @[RegFile.scala 97:16:@42243.4]
  assign rport_io_ins_284 = regs_284_io_out; // @[RegFile.scala 97:16:@42244.4]
  assign rport_io_ins_285 = regs_285_io_out; // @[RegFile.scala 97:16:@42245.4]
  assign rport_io_ins_286 = regs_286_io_out; // @[RegFile.scala 97:16:@42246.4]
  assign rport_io_ins_287 = regs_287_io_out; // @[RegFile.scala 97:16:@42247.4]
  assign rport_io_ins_288 = regs_288_io_out; // @[RegFile.scala 97:16:@42248.4]
  assign rport_io_ins_289 = regs_289_io_out; // @[RegFile.scala 97:16:@42249.4]
  assign rport_io_ins_290 = regs_290_io_out; // @[RegFile.scala 97:16:@42250.4]
  assign rport_io_ins_291 = regs_291_io_out; // @[RegFile.scala 97:16:@42251.4]
  assign rport_io_ins_292 = regs_292_io_out; // @[RegFile.scala 97:16:@42252.4]
  assign rport_io_ins_293 = regs_293_io_out; // @[RegFile.scala 97:16:@42253.4]
  assign rport_io_ins_294 = regs_294_io_out; // @[RegFile.scala 97:16:@42254.4]
  assign rport_io_ins_295 = regs_295_io_out; // @[RegFile.scala 97:16:@42255.4]
  assign rport_io_ins_296 = regs_296_io_out; // @[RegFile.scala 97:16:@42256.4]
  assign rport_io_ins_297 = regs_297_io_out; // @[RegFile.scala 97:16:@42257.4]
  assign rport_io_ins_298 = regs_298_io_out; // @[RegFile.scala 97:16:@42258.4]
  assign rport_io_ins_299 = regs_299_io_out; // @[RegFile.scala 97:16:@42259.4]
  assign rport_io_ins_300 = regs_300_io_out; // @[RegFile.scala 97:16:@42260.4]
  assign rport_io_ins_301 = regs_301_io_out; // @[RegFile.scala 97:16:@42261.4]
  assign rport_io_ins_302 = regs_302_io_out; // @[RegFile.scala 97:16:@42262.4]
  assign rport_io_ins_303 = regs_303_io_out; // @[RegFile.scala 97:16:@42263.4]
  assign rport_io_ins_304 = regs_304_io_out; // @[RegFile.scala 97:16:@42264.4]
  assign rport_io_ins_305 = regs_305_io_out; // @[RegFile.scala 97:16:@42265.4]
  assign rport_io_ins_306 = regs_306_io_out; // @[RegFile.scala 97:16:@42266.4]
  assign rport_io_ins_307 = regs_307_io_out; // @[RegFile.scala 97:16:@42267.4]
  assign rport_io_ins_308 = regs_308_io_out; // @[RegFile.scala 97:16:@42268.4]
  assign rport_io_ins_309 = regs_309_io_out; // @[RegFile.scala 97:16:@42269.4]
  assign rport_io_ins_310 = regs_310_io_out; // @[RegFile.scala 97:16:@42270.4]
  assign rport_io_ins_311 = regs_311_io_out; // @[RegFile.scala 97:16:@42271.4]
  assign rport_io_ins_312 = regs_312_io_out; // @[RegFile.scala 97:16:@42272.4]
  assign rport_io_ins_313 = regs_313_io_out; // @[RegFile.scala 97:16:@42273.4]
  assign rport_io_ins_314 = regs_314_io_out; // @[RegFile.scala 97:16:@42274.4]
  assign rport_io_ins_315 = regs_315_io_out; // @[RegFile.scala 97:16:@42275.4]
  assign rport_io_ins_316 = regs_316_io_out; // @[RegFile.scala 97:16:@42276.4]
  assign rport_io_ins_317 = regs_317_io_out; // @[RegFile.scala 97:16:@42277.4]
  assign rport_io_ins_318 = regs_318_io_out; // @[RegFile.scala 97:16:@42278.4]
  assign rport_io_ins_319 = regs_319_io_out; // @[RegFile.scala 97:16:@42279.4]
  assign rport_io_ins_320 = regs_320_io_out; // @[RegFile.scala 97:16:@42280.4]
  assign rport_io_ins_321 = regs_321_io_out; // @[RegFile.scala 97:16:@42281.4]
  assign rport_io_ins_322 = regs_322_io_out; // @[RegFile.scala 97:16:@42282.4]
  assign rport_io_ins_323 = regs_323_io_out; // @[RegFile.scala 97:16:@42283.4]
  assign rport_io_ins_324 = regs_324_io_out; // @[RegFile.scala 97:16:@42284.4]
  assign rport_io_ins_325 = regs_325_io_out; // @[RegFile.scala 97:16:@42285.4]
  assign rport_io_ins_326 = regs_326_io_out; // @[RegFile.scala 97:16:@42286.4]
  assign rport_io_ins_327 = regs_327_io_out; // @[RegFile.scala 97:16:@42287.4]
  assign rport_io_ins_328 = regs_328_io_out; // @[RegFile.scala 97:16:@42288.4]
  assign rport_io_ins_329 = regs_329_io_out; // @[RegFile.scala 97:16:@42289.4]
  assign rport_io_ins_330 = regs_330_io_out; // @[RegFile.scala 97:16:@42290.4]
  assign rport_io_ins_331 = regs_331_io_out; // @[RegFile.scala 97:16:@42291.4]
  assign rport_io_ins_332 = regs_332_io_out; // @[RegFile.scala 97:16:@42292.4]
  assign rport_io_ins_333 = regs_333_io_out; // @[RegFile.scala 97:16:@42293.4]
  assign rport_io_ins_334 = regs_334_io_out; // @[RegFile.scala 97:16:@42294.4]
  assign rport_io_ins_335 = regs_335_io_out; // @[RegFile.scala 97:16:@42295.4]
  assign rport_io_ins_336 = regs_336_io_out; // @[RegFile.scala 97:16:@42296.4]
  assign rport_io_ins_337 = regs_337_io_out; // @[RegFile.scala 97:16:@42297.4]
  assign rport_io_ins_338 = regs_338_io_out; // @[RegFile.scala 97:16:@42298.4]
  assign rport_io_ins_339 = regs_339_io_out; // @[RegFile.scala 97:16:@42299.4]
  assign rport_io_ins_340 = regs_340_io_out; // @[RegFile.scala 97:16:@42300.4]
  assign rport_io_ins_341 = regs_341_io_out; // @[RegFile.scala 97:16:@42301.4]
  assign rport_io_ins_342 = regs_342_io_out; // @[RegFile.scala 97:16:@42302.4]
  assign rport_io_ins_343 = regs_343_io_out; // @[RegFile.scala 97:16:@42303.4]
  assign rport_io_ins_344 = regs_344_io_out; // @[RegFile.scala 97:16:@42304.4]
  assign rport_io_ins_345 = regs_345_io_out; // @[RegFile.scala 97:16:@42305.4]
  assign rport_io_ins_346 = regs_346_io_out; // @[RegFile.scala 97:16:@42306.4]
  assign rport_io_ins_347 = regs_347_io_out; // @[RegFile.scala 97:16:@42307.4]
  assign rport_io_ins_348 = regs_348_io_out; // @[RegFile.scala 97:16:@42308.4]
  assign rport_io_ins_349 = regs_349_io_out; // @[RegFile.scala 97:16:@42309.4]
  assign rport_io_ins_350 = regs_350_io_out; // @[RegFile.scala 97:16:@42310.4]
  assign rport_io_ins_351 = regs_351_io_out; // @[RegFile.scala 97:16:@42311.4]
  assign rport_io_ins_352 = regs_352_io_out; // @[RegFile.scala 97:16:@42312.4]
  assign rport_io_ins_353 = regs_353_io_out; // @[RegFile.scala 97:16:@42313.4]
  assign rport_io_ins_354 = regs_354_io_out; // @[RegFile.scala 97:16:@42314.4]
  assign rport_io_ins_355 = regs_355_io_out; // @[RegFile.scala 97:16:@42315.4]
  assign rport_io_ins_356 = regs_356_io_out; // @[RegFile.scala 97:16:@42316.4]
  assign rport_io_ins_357 = regs_357_io_out; // @[RegFile.scala 97:16:@42317.4]
  assign rport_io_ins_358 = regs_358_io_out; // @[RegFile.scala 97:16:@42318.4]
  assign rport_io_ins_359 = regs_359_io_out; // @[RegFile.scala 97:16:@42319.4]
  assign rport_io_ins_360 = regs_360_io_out; // @[RegFile.scala 97:16:@42320.4]
  assign rport_io_ins_361 = regs_361_io_out; // @[RegFile.scala 97:16:@42321.4]
  assign rport_io_ins_362 = regs_362_io_out; // @[RegFile.scala 97:16:@42322.4]
  assign rport_io_ins_363 = regs_363_io_out; // @[RegFile.scala 97:16:@42323.4]
  assign rport_io_ins_364 = regs_364_io_out; // @[RegFile.scala 97:16:@42324.4]
  assign rport_io_ins_365 = regs_365_io_out; // @[RegFile.scala 97:16:@42325.4]
  assign rport_io_ins_366 = regs_366_io_out; // @[RegFile.scala 97:16:@42326.4]
  assign rport_io_ins_367 = regs_367_io_out; // @[RegFile.scala 97:16:@42327.4]
  assign rport_io_ins_368 = regs_368_io_out; // @[RegFile.scala 97:16:@42328.4]
  assign rport_io_ins_369 = regs_369_io_out; // @[RegFile.scala 97:16:@42329.4]
  assign rport_io_ins_370 = regs_370_io_out; // @[RegFile.scala 97:16:@42330.4]
  assign rport_io_ins_371 = regs_371_io_out; // @[RegFile.scala 97:16:@42331.4]
  assign rport_io_ins_372 = regs_372_io_out; // @[RegFile.scala 97:16:@42332.4]
  assign rport_io_ins_373 = regs_373_io_out; // @[RegFile.scala 97:16:@42333.4]
  assign rport_io_ins_374 = regs_374_io_out; // @[RegFile.scala 97:16:@42334.4]
  assign rport_io_ins_375 = regs_375_io_out; // @[RegFile.scala 97:16:@42335.4]
  assign rport_io_ins_376 = regs_376_io_out; // @[RegFile.scala 97:16:@42336.4]
  assign rport_io_ins_377 = regs_377_io_out; // @[RegFile.scala 97:16:@42337.4]
  assign rport_io_ins_378 = regs_378_io_out; // @[RegFile.scala 97:16:@42338.4]
  assign rport_io_ins_379 = regs_379_io_out; // @[RegFile.scala 97:16:@42339.4]
  assign rport_io_ins_380 = regs_380_io_out; // @[RegFile.scala 97:16:@42340.4]
  assign rport_io_ins_381 = regs_381_io_out; // @[RegFile.scala 97:16:@42341.4]
  assign rport_io_ins_382 = regs_382_io_out; // @[RegFile.scala 97:16:@42342.4]
  assign rport_io_ins_383 = regs_383_io_out; // @[RegFile.scala 97:16:@42343.4]
  assign rport_io_ins_384 = regs_384_io_out; // @[RegFile.scala 97:16:@42344.4]
  assign rport_io_ins_385 = regs_385_io_out; // @[RegFile.scala 97:16:@42345.4]
  assign rport_io_ins_386 = regs_386_io_out; // @[RegFile.scala 97:16:@42346.4]
  assign rport_io_ins_387 = regs_387_io_out; // @[RegFile.scala 97:16:@42347.4]
  assign rport_io_ins_388 = regs_388_io_out; // @[RegFile.scala 97:16:@42348.4]
  assign rport_io_ins_389 = regs_389_io_out; // @[RegFile.scala 97:16:@42349.4]
  assign rport_io_ins_390 = regs_390_io_out; // @[RegFile.scala 97:16:@42350.4]
  assign rport_io_ins_391 = regs_391_io_out; // @[RegFile.scala 97:16:@42351.4]
  assign rport_io_ins_392 = regs_392_io_out; // @[RegFile.scala 97:16:@42352.4]
  assign rport_io_ins_393 = regs_393_io_out; // @[RegFile.scala 97:16:@42353.4]
  assign rport_io_ins_394 = regs_394_io_out; // @[RegFile.scala 97:16:@42354.4]
  assign rport_io_ins_395 = regs_395_io_out; // @[RegFile.scala 97:16:@42355.4]
  assign rport_io_ins_396 = regs_396_io_out; // @[RegFile.scala 97:16:@42356.4]
  assign rport_io_ins_397 = regs_397_io_out; // @[RegFile.scala 97:16:@42357.4]
  assign rport_io_ins_398 = regs_398_io_out; // @[RegFile.scala 97:16:@42358.4]
  assign rport_io_ins_399 = regs_399_io_out; // @[RegFile.scala 97:16:@42359.4]
  assign rport_io_ins_400 = regs_400_io_out; // @[RegFile.scala 97:16:@42360.4]
  assign rport_io_ins_401 = regs_401_io_out; // @[RegFile.scala 97:16:@42361.4]
  assign rport_io_ins_402 = regs_402_io_out; // @[RegFile.scala 97:16:@42362.4]
  assign rport_io_ins_403 = regs_403_io_out; // @[RegFile.scala 97:16:@42363.4]
  assign rport_io_ins_404 = regs_404_io_out; // @[RegFile.scala 97:16:@42364.4]
  assign rport_io_ins_405 = regs_405_io_out; // @[RegFile.scala 97:16:@42365.4]
  assign rport_io_ins_406 = regs_406_io_out; // @[RegFile.scala 97:16:@42366.4]
  assign rport_io_ins_407 = regs_407_io_out; // @[RegFile.scala 97:16:@42367.4]
  assign rport_io_ins_408 = regs_408_io_out; // @[RegFile.scala 97:16:@42368.4]
  assign rport_io_ins_409 = regs_409_io_out; // @[RegFile.scala 97:16:@42369.4]
  assign rport_io_ins_410 = regs_410_io_out; // @[RegFile.scala 97:16:@42370.4]
  assign rport_io_ins_411 = regs_411_io_out; // @[RegFile.scala 97:16:@42371.4]
  assign rport_io_ins_412 = regs_412_io_out; // @[RegFile.scala 97:16:@42372.4]
  assign rport_io_ins_413 = regs_413_io_out; // @[RegFile.scala 97:16:@42373.4]
  assign rport_io_ins_414 = regs_414_io_out; // @[RegFile.scala 97:16:@42374.4]
  assign rport_io_ins_415 = regs_415_io_out; // @[RegFile.scala 97:16:@42375.4]
  assign rport_io_ins_416 = regs_416_io_out; // @[RegFile.scala 97:16:@42376.4]
  assign rport_io_ins_417 = regs_417_io_out; // @[RegFile.scala 97:16:@42377.4]
  assign rport_io_ins_418 = regs_418_io_out; // @[RegFile.scala 97:16:@42378.4]
  assign rport_io_ins_419 = regs_419_io_out; // @[RegFile.scala 97:16:@42379.4]
  assign rport_io_ins_420 = regs_420_io_out; // @[RegFile.scala 97:16:@42380.4]
  assign rport_io_ins_421 = regs_421_io_out; // @[RegFile.scala 97:16:@42381.4]
  assign rport_io_ins_422 = regs_422_io_out; // @[RegFile.scala 97:16:@42382.4]
  assign rport_io_ins_423 = regs_423_io_out; // @[RegFile.scala 97:16:@42383.4]
  assign rport_io_ins_424 = regs_424_io_out; // @[RegFile.scala 97:16:@42384.4]
  assign rport_io_ins_425 = regs_425_io_out; // @[RegFile.scala 97:16:@42385.4]
  assign rport_io_ins_426 = regs_426_io_out; // @[RegFile.scala 97:16:@42386.4]
  assign rport_io_ins_427 = regs_427_io_out; // @[RegFile.scala 97:16:@42387.4]
  assign rport_io_ins_428 = regs_428_io_out; // @[RegFile.scala 97:16:@42388.4]
  assign rport_io_ins_429 = regs_429_io_out; // @[RegFile.scala 97:16:@42389.4]
  assign rport_io_ins_430 = regs_430_io_out; // @[RegFile.scala 97:16:@42390.4]
  assign rport_io_ins_431 = regs_431_io_out; // @[RegFile.scala 97:16:@42391.4]
  assign rport_io_ins_432 = regs_432_io_out; // @[RegFile.scala 97:16:@42392.4]
  assign rport_io_ins_433 = regs_433_io_out; // @[RegFile.scala 97:16:@42393.4]
  assign rport_io_ins_434 = regs_434_io_out; // @[RegFile.scala 97:16:@42394.4]
  assign rport_io_ins_435 = regs_435_io_out; // @[RegFile.scala 97:16:@42395.4]
  assign rport_io_ins_436 = regs_436_io_out; // @[RegFile.scala 97:16:@42396.4]
  assign rport_io_ins_437 = regs_437_io_out; // @[RegFile.scala 97:16:@42397.4]
  assign rport_io_ins_438 = regs_438_io_out; // @[RegFile.scala 97:16:@42398.4]
  assign rport_io_ins_439 = regs_439_io_out; // @[RegFile.scala 97:16:@42399.4]
  assign rport_io_ins_440 = regs_440_io_out; // @[RegFile.scala 97:16:@42400.4]
  assign rport_io_ins_441 = regs_441_io_out; // @[RegFile.scala 97:16:@42401.4]
  assign rport_io_ins_442 = regs_442_io_out; // @[RegFile.scala 97:16:@42402.4]
  assign rport_io_ins_443 = regs_443_io_out; // @[RegFile.scala 97:16:@42403.4]
  assign rport_io_ins_444 = regs_444_io_out; // @[RegFile.scala 97:16:@42404.4]
  assign rport_io_ins_445 = regs_445_io_out; // @[RegFile.scala 97:16:@42405.4]
  assign rport_io_ins_446 = regs_446_io_out; // @[RegFile.scala 97:16:@42406.4]
  assign rport_io_ins_447 = regs_447_io_out; // @[RegFile.scala 97:16:@42407.4]
  assign rport_io_ins_448 = regs_448_io_out; // @[RegFile.scala 97:16:@42408.4]
  assign rport_io_ins_449 = regs_449_io_out; // @[RegFile.scala 97:16:@42409.4]
  assign rport_io_ins_450 = regs_450_io_out; // @[RegFile.scala 97:16:@42410.4]
  assign rport_io_ins_451 = regs_451_io_out; // @[RegFile.scala 97:16:@42411.4]
  assign rport_io_ins_452 = regs_452_io_out; // @[RegFile.scala 97:16:@42412.4]
  assign rport_io_ins_453 = regs_453_io_out; // @[RegFile.scala 97:16:@42413.4]
  assign rport_io_ins_454 = regs_454_io_out; // @[RegFile.scala 97:16:@42414.4]
  assign rport_io_ins_455 = regs_455_io_out; // @[RegFile.scala 97:16:@42415.4]
  assign rport_io_ins_456 = regs_456_io_out; // @[RegFile.scala 97:16:@42416.4]
  assign rport_io_ins_457 = regs_457_io_out; // @[RegFile.scala 97:16:@42417.4]
  assign rport_io_ins_458 = regs_458_io_out; // @[RegFile.scala 97:16:@42418.4]
  assign rport_io_ins_459 = regs_459_io_out; // @[RegFile.scala 97:16:@42419.4]
  assign rport_io_ins_460 = regs_460_io_out; // @[RegFile.scala 97:16:@42420.4]
  assign rport_io_ins_461 = regs_461_io_out; // @[RegFile.scala 97:16:@42421.4]
  assign rport_io_ins_462 = regs_462_io_out; // @[RegFile.scala 97:16:@42422.4]
  assign rport_io_ins_463 = regs_463_io_out; // @[RegFile.scala 97:16:@42423.4]
  assign rport_io_ins_464 = regs_464_io_out; // @[RegFile.scala 97:16:@42424.4]
  assign rport_io_ins_465 = regs_465_io_out; // @[RegFile.scala 97:16:@42425.4]
  assign rport_io_ins_466 = regs_466_io_out; // @[RegFile.scala 97:16:@42426.4]
  assign rport_io_ins_467 = regs_467_io_out; // @[RegFile.scala 97:16:@42427.4]
  assign rport_io_ins_468 = regs_468_io_out; // @[RegFile.scala 97:16:@42428.4]
  assign rport_io_ins_469 = regs_469_io_out; // @[RegFile.scala 97:16:@42429.4]
  assign rport_io_ins_470 = regs_470_io_out; // @[RegFile.scala 97:16:@42430.4]
  assign rport_io_ins_471 = regs_471_io_out; // @[RegFile.scala 97:16:@42431.4]
  assign rport_io_ins_472 = regs_472_io_out; // @[RegFile.scala 97:16:@42432.4]
  assign rport_io_ins_473 = regs_473_io_out; // @[RegFile.scala 97:16:@42433.4]
  assign rport_io_ins_474 = regs_474_io_out; // @[RegFile.scala 97:16:@42434.4]
  assign rport_io_ins_475 = regs_475_io_out; // @[RegFile.scala 97:16:@42435.4]
  assign rport_io_ins_476 = regs_476_io_out; // @[RegFile.scala 97:16:@42436.4]
  assign rport_io_ins_477 = regs_477_io_out; // @[RegFile.scala 97:16:@42437.4]
  assign rport_io_ins_478 = regs_478_io_out; // @[RegFile.scala 97:16:@42438.4]
  assign rport_io_ins_479 = regs_479_io_out; // @[RegFile.scala 97:16:@42439.4]
  assign rport_io_ins_480 = regs_480_io_out; // @[RegFile.scala 97:16:@42440.4]
  assign rport_io_ins_481 = regs_481_io_out; // @[RegFile.scala 97:16:@42441.4]
  assign rport_io_ins_482 = regs_482_io_out; // @[RegFile.scala 97:16:@42442.4]
  assign rport_io_ins_483 = regs_483_io_out; // @[RegFile.scala 97:16:@42443.4]
  assign rport_io_ins_484 = regs_484_io_out; // @[RegFile.scala 97:16:@42444.4]
  assign rport_io_ins_485 = regs_485_io_out; // @[RegFile.scala 97:16:@42445.4]
  assign rport_io_ins_486 = regs_486_io_out; // @[RegFile.scala 97:16:@42446.4]
  assign rport_io_ins_487 = regs_487_io_out; // @[RegFile.scala 97:16:@42447.4]
  assign rport_io_ins_488 = regs_488_io_out; // @[RegFile.scala 97:16:@42448.4]
  assign rport_io_ins_489 = regs_489_io_out; // @[RegFile.scala 97:16:@42449.4]
  assign rport_io_ins_490 = regs_490_io_out; // @[RegFile.scala 97:16:@42450.4]
  assign rport_io_ins_491 = regs_491_io_out; // @[RegFile.scala 97:16:@42451.4]
  assign rport_io_ins_492 = regs_492_io_out; // @[RegFile.scala 97:16:@42452.4]
  assign rport_io_ins_493 = regs_493_io_out; // @[RegFile.scala 97:16:@42453.4]
  assign rport_io_ins_494 = regs_494_io_out; // @[RegFile.scala 97:16:@42454.4]
  assign rport_io_ins_495 = regs_495_io_out; // @[RegFile.scala 97:16:@42455.4]
  assign rport_io_ins_496 = regs_496_io_out; // @[RegFile.scala 97:16:@42456.4]
  assign rport_io_ins_497 = regs_497_io_out; // @[RegFile.scala 97:16:@42457.4]
  assign rport_io_ins_498 = regs_498_io_out; // @[RegFile.scala 97:16:@42458.4]
  assign rport_io_ins_499 = regs_499_io_out; // @[RegFile.scala 97:16:@42459.4]
  assign rport_io_ins_500 = regs_500_io_out; // @[RegFile.scala 97:16:@42460.4]
  assign rport_io_ins_501 = regs_501_io_out; // @[RegFile.scala 97:16:@42461.4]
  assign rport_io_ins_502 = regs_502_io_out; // @[RegFile.scala 97:16:@42462.4]
  assign rport_io_sel = io_raddr[8:0]; // @[RegFile.scala 106:18:@42463.4]
endmodule
module RetimeWrapper_521( // @[:@42485.2]
  input         clock, // @[:@42486.4]
  input         reset, // @[:@42487.4]
  input  [39:0] io_in, // @[:@42488.4]
  output [39:0] io_out // @[:@42488.4]
);
  wire [39:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@42490.4]
  wire [39:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@42490.4]
  wire [39:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@42490.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@42490.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@42490.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@42490.4]
  RetimeShiftRegister #(.WIDTH(40), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@42490.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@42503.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@42502.4]
  assign sr_init = 40'h0; // @[RetimeShiftRegister.scala 19:16:@42501.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@42500.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@42499.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@42497.4]
endmodule
module FringeFF_503( // @[:@42505.2]
  input         clock, // @[:@42506.4]
  input         reset, // @[:@42507.4]
  input  [39:0] io_in, // @[:@42508.4]
  output [39:0] io_out, // @[:@42508.4]
  input         io_enable // @[:@42508.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@42511.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@42511.4]
  wire [39:0] RetimeWrapper_io_in; // @[package.scala 93:22:@42511.4]
  wire [39:0] RetimeWrapper_io_out; // @[package.scala 93:22:@42511.4]
  wire [39:0] _T_18; // @[package.scala 96:25:@42516.4 package.scala 96:25:@42517.4]
  RetimeWrapper_521 RetimeWrapper ( // @[package.scala 93:22:@42511.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@42516.4 package.scala 96:25:@42517.4]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@42528.4]
  assign RetimeWrapper_clock = clock; // @[:@42512.4]
  assign RetimeWrapper_reset = reset; // @[:@42513.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _T_18; // @[package.scala 94:16:@42514.4]
endmodule
module FringeCounter( // @[:@42530.2]
  input   clock, // @[:@42531.4]
  input   reset, // @[:@42532.4]
  input   io_enable, // @[:@42533.4]
  output  io_done // @[:@42533.4]
);
  wire  reg$_clock; // @[FringeCounter.scala 24:19:@42535.4]
  wire  reg$_reset; // @[FringeCounter.scala 24:19:@42535.4]
  wire [39:0] reg$_io_in; // @[FringeCounter.scala 24:19:@42535.4]
  wire [39:0] reg$_io_out; // @[FringeCounter.scala 24:19:@42535.4]
  wire  reg$_io_enable; // @[FringeCounter.scala 24:19:@42535.4]
  wire [40:0] count; // @[Cat.scala 30:58:@42542.4]
  wire [41:0] _T_25; // @[FringeCounter.scala 31:22:@42543.4]
  wire [40:0] newval; // @[FringeCounter.scala 31:22:@42544.4]
  wire  isMax; // @[FringeCounter.scala 32:22:@42545.4]
  wire [40:0] next; // @[FringeCounter.scala 33:17:@42547.4]
  FringeFF_503 reg$ ( // @[FringeCounter.scala 24:19:@42535.4]
    .clock(reg$_clock),
    .reset(reg$_reset),
    .io_in(reg$_io_in),
    .io_out(reg$_io_out),
    .io_enable(reg$_io_enable)
  );
  assign count = {1'h0,reg$_io_out}; // @[Cat.scala 30:58:@42542.4]
  assign _T_25 = count + 41'h1; // @[FringeCounter.scala 31:22:@42543.4]
  assign newval = count + 41'h1; // @[FringeCounter.scala 31:22:@42544.4]
  assign isMax = newval >= 41'h2cb417800; // @[FringeCounter.scala 32:22:@42545.4]
  assign next = isMax ? count : newval; // @[FringeCounter.scala 33:17:@42547.4]
  assign io_done = io_enable & isMax; // @[FringeCounter.scala 43:11:@42558.4]
  assign reg$_clock = clock; // @[:@42536.4]
  assign reg$_reset = reset; // @[:@42537.4]
  assign reg$_io_in = next[39:0]; // @[FringeCounter.scala 35:15:@42549.6 FringeCounter.scala 37:15:@42552.6]
  assign reg$_io_enable = io_enable; // @[FringeCounter.scala 27:17:@42540.4]
endmodule
module FringeFF_504( // @[:@42592.2]
  input   clock, // @[:@42593.4]
  input   reset, // @[:@42594.4]
  input   io_in, // @[:@42595.4]
  input   io_reset, // @[:@42595.4]
  output  io_out, // @[:@42595.4]
  input   io_enable // @[:@42595.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@42598.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@42598.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@42598.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@42598.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@42598.4]
  wire  _T_18; // @[package.scala 96:25:@42603.4 package.scala 96:25:@42604.4]
  wire  _GEN_0; // @[FringeFF.scala 21:27:@42609.6]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@42598.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@42603.4 package.scala 96:25:@42604.4]
  assign _GEN_0 = io_reset ? 1'h0 : _T_18; // @[FringeFF.scala 21:27:@42609.6]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@42615.4]
  assign RetimeWrapper_clock = clock; // @[:@42599.4]
  assign RetimeWrapper_reset = reset; // @[:@42600.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@42602.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _GEN_0; // @[package.scala 94:16:@42601.4]
endmodule
module Depulser( // @[:@42617.2]
  input   clock, // @[:@42618.4]
  input   reset, // @[:@42619.4]
  input   io_in, // @[:@42620.4]
  input   io_rst, // @[:@42620.4]
  output  io_out // @[:@42620.4]
);
  wire  r_clock; // @[Depulser.scala 14:17:@42622.4]
  wire  r_reset; // @[Depulser.scala 14:17:@42622.4]
  wire  r_io_in; // @[Depulser.scala 14:17:@42622.4]
  wire  r_io_reset; // @[Depulser.scala 14:17:@42622.4]
  wire  r_io_out; // @[Depulser.scala 14:17:@42622.4]
  wire  r_io_enable; // @[Depulser.scala 14:17:@42622.4]
  FringeFF_504 r ( // @[Depulser.scala 14:17:@42622.4]
    .clock(r_clock),
    .reset(r_reset),
    .io_in(r_io_in),
    .io_reset(r_io_reset),
    .io_out(r_io_out),
    .io_enable(r_io_enable)
  );
  assign io_out = r_io_out; // @[Depulser.scala 19:10:@42631.4]
  assign r_clock = clock; // @[:@42623.4]
  assign r_reset = reset; // @[:@42624.4]
  assign r_io_in = io_rst ? 1'h0 : io_in; // @[Depulser.scala 15:11:@42626.4]
  assign r_io_reset = io_rst; // @[Depulser.scala 18:14:@42630.4]
  assign r_io_enable = io_in | io_rst; // @[Depulser.scala 17:15:@42629.4]
endmodule
module Fringe( // @[:@42633.2]
  input         clock, // @[:@42634.4]
  input         reset, // @[:@42635.4]
  input  [31:0] io_raddr, // @[:@42636.4]
  input         io_wen, // @[:@42636.4]
  input  [31:0] io_waddr, // @[:@42636.4]
  input  [63:0] io_wdata, // @[:@42636.4]
  output [63:0] io_rdata, // @[:@42636.4]
  output        io_enable, // @[:@42636.4]
  input         io_done, // @[:@42636.4]
  output        io_reset, // @[:@42636.4]
  output [63:0] io_argIns_0, // @[:@42636.4]
  input         io_argOuts_0_valid, // @[:@42636.4]
  input  [63:0] io_argOuts_0_bits, // @[:@42636.4]
  output [63:0] io_argEchos_0, // @[:@42636.4]
  input         io_heap_0_req_valid, // @[:@42636.4]
  input         io_heap_0_req_bits_allocDealloc, // @[:@42636.4]
  input  [63:0] io_heap_0_req_bits_sizeAddr, // @[:@42636.4]
  output        io_heap_0_resp_valid, // @[:@42636.4]
  output        io_heap_0_resp_bits_allocDealloc, // @[:@42636.4]
  output [63:0] io_heap_0_resp_bits_sizeAddr // @[:@42636.4]
);
  wire  heap_io_accel_0_req_valid; // @[Fringe.scala 107:20:@44337.4]
  wire  heap_io_accel_0_req_bits_allocDealloc; // @[Fringe.scala 107:20:@44337.4]
  wire [63:0] heap_io_accel_0_req_bits_sizeAddr; // @[Fringe.scala 107:20:@44337.4]
  wire  heap_io_accel_0_resp_valid; // @[Fringe.scala 107:20:@44337.4]
  wire  heap_io_accel_0_resp_bits_allocDealloc; // @[Fringe.scala 107:20:@44337.4]
  wire [63:0] heap_io_accel_0_resp_bits_sizeAddr; // @[Fringe.scala 107:20:@44337.4]
  wire  heap_io_host_0_req_valid; // @[Fringe.scala 107:20:@44337.4]
  wire  heap_io_host_0_req_bits_allocDealloc; // @[Fringe.scala 107:20:@44337.4]
  wire [63:0] heap_io_host_0_req_bits_sizeAddr; // @[Fringe.scala 107:20:@44337.4]
  wire  heap_io_host_0_resp_valid; // @[Fringe.scala 107:20:@44337.4]
  wire  heap_io_host_0_resp_bits_allocDealloc; // @[Fringe.scala 107:20:@44337.4]
  wire [63:0] heap_io_host_0_resp_bits_sizeAddr; // @[Fringe.scala 107:20:@44337.4]
  wire  regs_clock; // @[Fringe.scala 116:20:@44346.4]
  wire  regs_reset; // @[Fringe.scala 116:20:@44346.4]
  wire [9:0] regs_io_raddr; // @[Fringe.scala 116:20:@44346.4]
  wire  regs_io_wen; // @[Fringe.scala 116:20:@44346.4]
  wire [9:0] regs_io_waddr; // @[Fringe.scala 116:20:@44346.4]
  wire [63:0] regs_io_wdata; // @[Fringe.scala 116:20:@44346.4]
  wire [63:0] regs_io_rdata; // @[Fringe.scala 116:20:@44346.4]
  wire  regs_io_reset; // @[Fringe.scala 116:20:@44346.4]
  wire [63:0] regs_io_argIns_0; // @[Fringe.scala 116:20:@44346.4]
  wire [63:0] regs_io_argIns_1; // @[Fringe.scala 116:20:@44346.4]
  wire [63:0] regs_io_argIns_2; // @[Fringe.scala 116:20:@44346.4]
  wire  regs_io_argOuts_0_valid; // @[Fringe.scala 116:20:@44346.4]
  wire [63:0] regs_io_argOuts_0_bits; // @[Fringe.scala 116:20:@44346.4]
  wire  regs_io_argOuts_1_valid; // @[Fringe.scala 116:20:@44346.4]
  wire [63:0] regs_io_argOuts_1_bits; // @[Fringe.scala 116:20:@44346.4]
  wire [63:0] regs_io_argEchos_1; // @[Fringe.scala 116:20:@44346.4]
  wire  timeoutCtr_clock; // @[Fringe.scala 143:26:@46399.4]
  wire  timeoutCtr_reset; // @[Fringe.scala 143:26:@46399.4]
  wire  timeoutCtr_io_enable; // @[Fringe.scala 143:26:@46399.4]
  wire  timeoutCtr_io_done; // @[Fringe.scala 143:26:@46399.4]
  wire  depulser_clock; // @[Fringe.scala 153:24:@46417.4]
  wire  depulser_reset; // @[Fringe.scala 153:24:@46417.4]
  wire  depulser_io_in; // @[Fringe.scala 153:24:@46417.4]
  wire  depulser_io_rst; // @[Fringe.scala 153:24:@46417.4]
  wire  depulser_io_out; // @[Fringe.scala 153:24:@46417.4]
  reg [63:0] _T_921; // @[Reg.scala 11:16:@46370.4]
  reg [63:0] _RAND_0;
  wire [63:0] _T_925; // @[:@46376.4 :@46377.4]
  wire  curStatus_done; // @[Fringe.scala 133:45:@46378.4]
  wire  curStatus_timeout; // @[Fringe.scala 133:45:@46380.4]
  wire [2:0] curStatus_allocDealloc; // @[Fringe.scala 133:45:@46382.4]
  wire [58:0] curStatus_sizeAddr; // @[Fringe.scala 133:45:@46384.4]
  wire  _T_930; // @[Fringe.scala 134:28:@46386.4]
  wire  _T_934; // @[Fringe.scala 134:42:@46388.4]
  wire  _T_935; // @[Fringe.scala 135:27:@46390.4]
  wire [63:0] _T_945; // @[Fringe.scala 156:22:@46425.4]
  reg  _T_952; // @[package.scala 152:20:@46428.4]
  reg [31:0] _RAND_1;
  wire  _T_953; // @[package.scala 153:13:@46430.4]
  wire  _T_954; // @[package.scala 153:8:@46431.4]
  wire  _T_957; // @[Fringe.scala 160:55:@46435.4]
  wire  status_bits_done; // @[Fringe.scala 160:26:@46436.4]
  wire  _T_960; // @[Fringe.scala 161:58:@46439.4]
  wire  status_bits_timeout; // @[Fringe.scala 161:29:@46440.4]
  wire [1:0] _T_964; // @[Fringe.scala 162:57:@46442.4]
  wire [1:0] _T_966; // @[Fringe.scala 162:34:@46443.4]
  wire [63:0] _T_968; // @[Fringe.scala 163:30:@46445.4]
  wire [1:0] _T_969; // @[Fringe.scala 171:37:@46448.4]
  wire [58:0] status_bits_sizeAddr; // @[Fringe.scala 158:20:@46427.4 Fringe.scala 163:24:@46446.4]
  wire [2:0] status_bits_allocDealloc; // @[Fringe.scala 158:20:@46427.4 Fringe.scala 162:28:@46444.4]
  wire [61:0] _T_970; // @[Fringe.scala 171:37:@46449.4]
  wire  alloc; // @[Fringe.scala 202:38:@47830.4]
  wire  dealloc; // @[Fringe.scala 203:40:@47831.4]
  wire  _T_1474; // @[Fringe.scala 204:37:@47832.4]
  reg  _T_1477; // @[package.scala 152:20:@47833.4]
  reg [31:0] _RAND_2;
  wire  _T_1478; // @[package.scala 153:13:@47835.4]
  DRAMHeap heap ( // @[Fringe.scala 107:20:@44337.4]
    .io_accel_0_req_valid(heap_io_accel_0_req_valid),
    .io_accel_0_req_bits_allocDealloc(heap_io_accel_0_req_bits_allocDealloc),
    .io_accel_0_req_bits_sizeAddr(heap_io_accel_0_req_bits_sizeAddr),
    .io_accel_0_resp_valid(heap_io_accel_0_resp_valid),
    .io_accel_0_resp_bits_allocDealloc(heap_io_accel_0_resp_bits_allocDealloc),
    .io_accel_0_resp_bits_sizeAddr(heap_io_accel_0_resp_bits_sizeAddr),
    .io_host_0_req_valid(heap_io_host_0_req_valid),
    .io_host_0_req_bits_allocDealloc(heap_io_host_0_req_bits_allocDealloc),
    .io_host_0_req_bits_sizeAddr(heap_io_host_0_req_bits_sizeAddr),
    .io_host_0_resp_valid(heap_io_host_0_resp_valid),
    .io_host_0_resp_bits_allocDealloc(heap_io_host_0_resp_bits_allocDealloc),
    .io_host_0_resp_bits_sizeAddr(heap_io_host_0_resp_bits_sizeAddr)
  );
  RegFile regs ( // @[Fringe.scala 116:20:@44346.4]
    .clock(regs_clock),
    .reset(regs_reset),
    .io_raddr(regs_io_raddr),
    .io_wen(regs_io_wen),
    .io_waddr(regs_io_waddr),
    .io_wdata(regs_io_wdata),
    .io_rdata(regs_io_rdata),
    .io_reset(regs_io_reset),
    .io_argIns_0(regs_io_argIns_0),
    .io_argIns_1(regs_io_argIns_1),
    .io_argIns_2(regs_io_argIns_2),
    .io_argOuts_0_valid(regs_io_argOuts_0_valid),
    .io_argOuts_0_bits(regs_io_argOuts_0_bits),
    .io_argOuts_1_valid(regs_io_argOuts_1_valid),
    .io_argOuts_1_bits(regs_io_argOuts_1_bits),
    .io_argEchos_1(regs_io_argEchos_1)
  );
  FringeCounter timeoutCtr ( // @[Fringe.scala 143:26:@46399.4]
    .clock(timeoutCtr_clock),
    .reset(timeoutCtr_reset),
    .io_enable(timeoutCtr_io_enable),
    .io_done(timeoutCtr_io_done)
  );
  Depulser depulser ( // @[Fringe.scala 153:24:@46417.4]
    .clock(depulser_clock),
    .reset(depulser_reset),
    .io_in(depulser_io_in),
    .io_rst(depulser_io_rst),
    .io_out(depulser_io_out)
  );
  assign _T_925 = regs_io_argIns_1; // @[:@46376.4 :@46377.4]
  assign curStatus_done = _T_925[0]; // @[Fringe.scala 133:45:@46378.4]
  assign curStatus_timeout = _T_925[1]; // @[Fringe.scala 133:45:@46380.4]
  assign curStatus_allocDealloc = _T_925[4:2]; // @[Fringe.scala 133:45:@46382.4]
  assign curStatus_sizeAddr = _T_925[63:5]; // @[Fringe.scala 133:45:@46384.4]
  assign _T_930 = regs_io_argIns_0[0]; // @[Fringe.scala 134:28:@46386.4]
  assign _T_934 = curStatus_done == 1'h0; // @[Fringe.scala 134:42:@46388.4]
  assign _T_935 = regs_io_argIns_0[1]; // @[Fringe.scala 135:27:@46390.4]
  assign _T_945 = ~ regs_io_argIns_0; // @[Fringe.scala 156:22:@46425.4]
  assign _T_953 = _T_952 ^ heap_io_host_0_req_valid; // @[package.scala 153:13:@46430.4]
  assign _T_954 = heap_io_host_0_req_valid & _T_953; // @[package.scala 153:8:@46431.4]
  assign _T_957 = _T_930 & depulser_io_out; // @[Fringe.scala 160:55:@46435.4]
  assign status_bits_done = depulser_io_out ? _T_957 : curStatus_done; // @[Fringe.scala 160:26:@46436.4]
  assign _T_960 = _T_930 & timeoutCtr_io_done; // @[Fringe.scala 161:58:@46439.4]
  assign status_bits_timeout = depulser_io_out ? _T_960 : curStatus_timeout; // @[Fringe.scala 161:29:@46440.4]
  assign _T_964 = heap_io_host_0_req_bits_allocDealloc ? 2'h1 : 2'h2; // @[Fringe.scala 162:57:@46442.4]
  assign _T_966 = heap_io_host_0_req_valid ? _T_964 : 2'h0; // @[Fringe.scala 162:34:@46443.4]
  assign _T_968 = heap_io_host_0_req_valid ? heap_io_host_0_req_bits_sizeAddr : 64'h0; // @[Fringe.scala 163:30:@46445.4]
  assign _T_969 = {status_bits_timeout,status_bits_done}; // @[Fringe.scala 171:37:@46448.4]
  assign status_bits_sizeAddr = _T_968[58:0]; // @[Fringe.scala 158:20:@46427.4 Fringe.scala 163:24:@46446.4]
  assign status_bits_allocDealloc = {{1'd0}, _T_966}; // @[Fringe.scala 158:20:@46427.4 Fringe.scala 162:28:@46444.4]
  assign _T_970 = {status_bits_sizeAddr,status_bits_allocDealloc}; // @[Fringe.scala 171:37:@46449.4]
  assign alloc = curStatus_allocDealloc == 3'h3; // @[Fringe.scala 202:38:@47830.4]
  assign dealloc = curStatus_allocDealloc == 3'h4; // @[Fringe.scala 203:40:@47831.4]
  assign _T_1474 = alloc | dealloc; // @[Fringe.scala 204:37:@47832.4]
  assign _T_1478 = _T_1477 ^ _T_1474; // @[package.scala 153:13:@47835.4]
  assign io_rdata = _T_921; // @[Fringe.scala 128:14:@46374.4]
  assign io_enable = _T_930 & _T_934; // @[Fringe.scala 136:13:@46394.4]
  assign io_reset = _T_935 | reset; // @[Fringe.scala 137:12:@46395.4]
  assign io_argIns_0 = regs_io_argIns_2; // @[Fringe.scala 151:51:@46416.4]
  assign io_argEchos_0 = regs_io_argEchos_1; // @[Fringe.scala 174:24:@46452.4]
  assign io_heap_0_resp_valid = heap_io_accel_0_resp_valid; // @[Fringe.scala 108:17:@44342.4]
  assign io_heap_0_resp_bits_allocDealloc = heap_io_accel_0_resp_bits_allocDealloc; // @[Fringe.scala 108:17:@44341.4]
  assign io_heap_0_resp_bits_sizeAddr = heap_io_accel_0_resp_bits_sizeAddr; // @[Fringe.scala 108:17:@44340.4]
  assign heap_io_accel_0_req_valid = io_heap_0_req_valid; // @[Fringe.scala 108:17:@44345.4]
  assign heap_io_accel_0_req_bits_allocDealloc = io_heap_0_req_bits_allocDealloc; // @[Fringe.scala 108:17:@44344.4]
  assign heap_io_accel_0_req_bits_sizeAddr = io_heap_0_req_bits_sizeAddr; // @[Fringe.scala 108:17:@44343.4]
  assign heap_io_host_0_resp_valid = _T_1474 & _T_1478; // @[Fringe.scala 204:22:@47837.4]
  assign heap_io_host_0_resp_bits_allocDealloc = curStatus_allocDealloc == 3'h3; // @[Fringe.scala 205:34:@47838.4]
  assign heap_io_host_0_resp_bits_sizeAddr = {{5'd0}, curStatus_sizeAddr}; // @[Fringe.scala 206:30:@47839.4]
  assign regs_clock = clock; // @[:@44347.4]
  assign regs_reset = reset; // @[:@44348.4 Fringe.scala 139:14:@46398.4]
  assign regs_io_raddr = io_raddr[9:0]; // @[Fringe.scala 118:17:@46366.4]
  assign regs_io_wen = io_wen; // @[Fringe.scala 120:15:@46368.4]
  assign regs_io_waddr = io_waddr[9:0]; // @[Fringe.scala 119:17:@46367.4]
  assign regs_io_wdata = io_wdata; // @[Fringe.scala 121:17:@46369.4]
  assign regs_io_reset = _T_935 | reset; // @[Fringe.scala 138:17:@46396.4]
  assign regs_io_argOuts_0_valid = depulser_io_out | _T_954; // @[Fringe.scala 170:23:@46447.4]
  assign regs_io_argOuts_0_bits = {_T_970,_T_969}; // @[Fringe.scala 171:22:@46451.4]
  assign regs_io_argOuts_1_valid = io_argOuts_0_valid; // @[Fringe.scala 176:23:@46454.4]
  assign regs_io_argOuts_1_bits = io_argOuts_0_bits; // @[Fringe.scala 175:22:@46453.4]
  assign timeoutCtr_clock = clock; // @[:@46400.4]
  assign timeoutCtr_reset = reset; // @[:@46401.4]
  assign timeoutCtr_io_enable = _T_930 & _T_934; // @[Fringe.scala 149:24:@46415.4]
  assign depulser_clock = clock; // @[:@46418.4]
  assign depulser_reset = reset; // @[:@46419.4]
  assign depulser_io_in = io_done | timeoutCtr_io_done; // @[Fringe.scala 155:18:@46424.4]
  assign depulser_io_rst = _T_945[0]; // @[Fringe.scala 156:19:@46426.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  _T_921 = _RAND_0[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_952 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_1477 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    _T_921 <= regs_io_rdata;
    if (reset) begin
      _T_952 <= 1'h0;
    end else begin
      _T_952 <= heap_io_host_0_req_valid;
    end
    if (reset) begin
      _T_1477 <= 1'h0;
    end else begin
      _T_1477 <= _T_1474;
    end
  end
endmodule
module SpatialIP( // @[:@47841.2]
  input         clock, // @[:@47842.4]
  input         reset, // @[:@47843.4]
  input  [31:0] io_raddr, // @[:@47844.4]
  input         io_wen, // @[:@47844.4]
  input  [31:0] io_waddr, // @[:@47844.4]
  input  [63:0] io_wdata, // @[:@47844.4]
  output [63:0] io_rdata, // @[:@47844.4]
  input         io_dram_0_cmd_ready, // @[:@47844.4]
  output        io_dram_0_cmd_valid, // @[:@47844.4]
  output [63:0] io_dram_0_cmd_bits_addr, // @[:@47844.4]
  output [31:0] io_dram_0_cmd_bits_size, // @[:@47844.4]
  output [63:0] io_dram_0_cmd_bits_rawAddr, // @[:@47844.4]
  output        io_dram_0_cmd_bits_isWr, // @[:@47844.4]
  output [31:0] io_dram_0_cmd_bits_tag, // @[:@47844.4]
  input         io_dram_0_wdata_ready, // @[:@47844.4]
  output        io_dram_0_wdata_valid, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_0, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_1, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_2, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_3, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_4, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_5, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_6, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_7, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_8, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_9, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_10, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_11, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_12, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_13, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_14, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_15, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_16, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_17, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_18, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_19, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_20, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_21, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_22, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_23, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_24, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_25, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_26, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_27, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_28, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_29, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_30, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_31, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_32, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_33, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_34, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_35, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_36, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_37, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_38, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_39, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_40, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_41, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_42, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_43, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_44, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_45, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_46, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_47, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_48, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_49, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_50, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_51, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_52, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_53, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_54, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_55, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_56, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_57, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_58, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_59, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_60, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_61, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_62, // @[:@47844.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_63, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_0, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_1, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_2, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_3, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_4, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_5, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_6, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_7, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_8, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_9, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_10, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_11, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_12, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_13, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_14, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_15, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_16, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_17, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_18, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_19, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_20, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_21, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_22, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_23, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_24, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_25, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_26, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_27, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_28, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_29, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_30, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_31, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_32, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_33, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_34, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_35, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_36, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_37, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_38, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_39, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_40, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_41, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_42, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_43, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_44, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_45, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_46, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_47, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_48, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_49, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_50, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_51, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_52, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_53, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_54, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_55, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_56, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_57, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_58, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_59, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_60, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_61, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_62, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wstrb_63, // @[:@47844.4]
  output        io_dram_0_wdata_bits_wlast, // @[:@47844.4]
  output        io_dram_0_rresp_ready, // @[:@47844.4]
  input         io_dram_0_rresp_valid, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_0, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_1, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_2, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_3, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_4, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_5, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_6, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_7, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_8, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_9, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_10, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_11, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_12, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_13, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_14, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_15, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_16, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_17, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_18, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_19, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_20, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_21, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_22, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_23, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_24, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_25, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_26, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_27, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_28, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_29, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_30, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_31, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_32, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_33, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_34, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_35, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_36, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_37, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_38, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_39, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_40, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_41, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_42, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_43, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_44, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_45, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_46, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_47, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_48, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_49, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_50, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_51, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_52, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_53, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_54, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_55, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_56, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_57, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_58, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_59, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_60, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_61, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_62, // @[:@47844.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_63, // @[:@47844.4]
  input  [31:0] io_dram_0_rresp_bits_tag, // @[:@47844.4]
  output        io_dram_0_wresp_ready, // @[:@47844.4]
  input         io_dram_0_wresp_valid, // @[:@47844.4]
  input  [31:0] io_dram_0_wresp_bits_tag // @[:@47844.4]
);
  wire  accel_clock; // @[Instantiator.scala 53:44:@47846.4]
  wire  accel_reset; // @[Instantiator.scala 53:44:@47846.4]
  wire  accel_io_enable; // @[Instantiator.scala 53:44:@47846.4]
  wire  accel_io_done; // @[Instantiator.scala 53:44:@47846.4]
  wire  accel_io_reset; // @[Instantiator.scala 53:44:@47846.4]
  wire  accel_io_memStreams_loads_0_cmd_ready; // @[Instantiator.scala 53:44:@47846.4]
  wire  accel_io_memStreams_loads_0_cmd_valid; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_loads_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@47846.4]
  wire [31:0] accel_io_memStreams_loads_0_cmd_bits_size; // @[Instantiator.scala 53:44:@47846.4]
  wire  accel_io_memStreams_loads_0_data_ready; // @[Instantiator.scala 53:44:@47846.4]
  wire  accel_io_memStreams_loads_0_data_valid; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_0; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_1; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_2; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_3; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_4; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_5; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_6; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_7; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_8; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_9; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_10; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_11; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_12; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_13; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_14; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_15; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_16; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_17; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_18; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_19; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_20; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_21; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_22; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_23; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_24; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_25; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_26; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_27; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_28; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_29; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_30; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_31; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_32; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_33; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_34; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_35; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_36; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_37; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_38; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_39; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_40; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_41; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_42; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_43; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_44; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_45; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_46; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_47; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_48; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_49; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_50; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_51; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_52; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_53; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_54; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_55; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_56; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_57; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_58; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_59; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_60; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_61; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_62; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_loads_0_data_bits_rdata_63; // @[Instantiator.scala 53:44:@47846.4]
  wire  accel_io_memStreams_stores_0_cmd_ready; // @[Instantiator.scala 53:44:@47846.4]
  wire  accel_io_memStreams_stores_0_cmd_valid; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_stores_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@47846.4]
  wire [31:0] accel_io_memStreams_stores_0_cmd_bits_size; // @[Instantiator.scala 53:44:@47846.4]
  wire  accel_io_memStreams_stores_0_data_ready; // @[Instantiator.scala 53:44:@47846.4]
  wire  accel_io_memStreams_stores_0_data_valid; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_1; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_2; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_3; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_4; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_5; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_6; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_7; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_8; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_9; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_10; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_11; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_12; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_13; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_14; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_15; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_16; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_17; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_18; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_19; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_20; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_21; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_22; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_23; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_24; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_25; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_26; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_27; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_28; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_29; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_30; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_31; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_32; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_33; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_34; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_35; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_36; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_37; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_38; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_39; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_40; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_41; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_42; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_43; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_44; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_45; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_46; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_47; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_48; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_49; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_50; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_51; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_52; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_53; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_54; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_55; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_56; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_57; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_58; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_59; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_60; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_61; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_62; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_63; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_stores_0_data_bits_wstrb; // @[Instantiator.scala 53:44:@47846.4]
  wire  accel_io_memStreams_stores_0_wresp_ready; // @[Instantiator.scala 53:44:@47846.4]
  wire  accel_io_memStreams_stores_0_wresp_valid; // @[Instantiator.scala 53:44:@47846.4]
  wire  accel_io_memStreams_stores_0_wresp_bits; // @[Instantiator.scala 53:44:@47846.4]
  wire  accel_io_memStreams_gathers_0_cmd_ready; // @[Instantiator.scala 53:44:@47846.4]
  wire  accel_io_memStreams_gathers_0_cmd_valid; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_0; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_1; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_2; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_3; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_4; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_5; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_6; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_7; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_8; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_9; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_10; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_11; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_12; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_13; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_14; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_15; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_16; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_17; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_18; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_19; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_20; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_21; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_22; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_23; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_24; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_25; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_26; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_27; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_28; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_29; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_30; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_31; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_32; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_33; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_34; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_35; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_36; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_37; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_38; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_39; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_40; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_41; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_42; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_43; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_44; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_45; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_46; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_47; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_48; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_49; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_50; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_51; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_52; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_53; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_54; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_55; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_56; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_57; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_58; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_59; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_60; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_61; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_62; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_63; // @[Instantiator.scala 53:44:@47846.4]
  wire  accel_io_memStreams_gathers_0_data_ready; // @[Instantiator.scala 53:44:@47846.4]
  wire  accel_io_memStreams_gathers_0_data_valid; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_0; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_1; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_2; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_3; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_4; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_5; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_6; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_7; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_8; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_9; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_10; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_11; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_12; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_13; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_14; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_15; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_16; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_17; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_18; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_19; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_20; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_21; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_22; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_23; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_24; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_25; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_26; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_27; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_28; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_29; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_30; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_31; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_32; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_33; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_34; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_35; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_36; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_37; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_38; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_39; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_40; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_41; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_42; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_43; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_44; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_45; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_46; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_47; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_48; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_49; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_50; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_51; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_52; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_53; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_54; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_55; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_56; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_57; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_58; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_59; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_60; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_61; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_62; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_63; // @[Instantiator.scala 53:44:@47846.4]
  wire  accel_io_memStreams_scatters_0_cmd_ready; // @[Instantiator.scala 53:44:@47846.4]
  wire  accel_io_memStreams_scatters_0_cmd_valid; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_16; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_17; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_18; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_19; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_20; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_21; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_22; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_23; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_24; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_25; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_26; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_27; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_28; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_29; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_30; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_31; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_32; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_33; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_34; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_35; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_36; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_37; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_38; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_39; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_40; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_41; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_42; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_43; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_44; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_45; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_46; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_47; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_48; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_49; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_50; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_51; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_52; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_53; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_54; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_55; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_56; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_57; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_58; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_59; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_60; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_61; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_62; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_63; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_0; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_1; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_2; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_3; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_4; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_5; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_6; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_7; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_8; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_9; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_10; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_11; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_12; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_13; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_14; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_15; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_16; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_17; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_18; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_19; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_20; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_21; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_22; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_23; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_24; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_25; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_26; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_27; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_28; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_29; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_30; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_31; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_32; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_33; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_34; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_35; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_36; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_37; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_38; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_39; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_40; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_41; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_42; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_43; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_44; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_45; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_46; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_47; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_48; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_49; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_50; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_51; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_52; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_53; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_54; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_55; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_56; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_57; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_58; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_59; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_60; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_61; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_62; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_63; // @[Instantiator.scala 53:44:@47846.4]
  wire  accel_io_memStreams_scatters_0_wresp_ready; // @[Instantiator.scala 53:44:@47846.4]
  wire  accel_io_memStreams_scatters_0_wresp_valid; // @[Instantiator.scala 53:44:@47846.4]
  wire  accel_io_memStreams_scatters_0_wresp_bits; // @[Instantiator.scala 53:44:@47846.4]
  wire  accel_io_axiStreamsIn_0_TVALID; // @[Instantiator.scala 53:44:@47846.4]
  wire  accel_io_axiStreamsIn_0_TREADY; // @[Instantiator.scala 53:44:@47846.4]
  wire [255:0] accel_io_axiStreamsIn_0_TDATA; // @[Instantiator.scala 53:44:@47846.4]
  wire [31:0] accel_io_axiStreamsIn_0_TSTRB; // @[Instantiator.scala 53:44:@47846.4]
  wire [31:0] accel_io_axiStreamsIn_0_TKEEP; // @[Instantiator.scala 53:44:@47846.4]
  wire  accel_io_axiStreamsIn_0_TLAST; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_axiStreamsIn_0_TID; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_axiStreamsIn_0_TDEST; // @[Instantiator.scala 53:44:@47846.4]
  wire [31:0] accel_io_axiStreamsIn_0_TUSER; // @[Instantiator.scala 53:44:@47846.4]
  wire  accel_io_axiStreamsOut_0_TVALID; // @[Instantiator.scala 53:44:@47846.4]
  wire  accel_io_axiStreamsOut_0_TREADY; // @[Instantiator.scala 53:44:@47846.4]
  wire [255:0] accel_io_axiStreamsOut_0_TDATA; // @[Instantiator.scala 53:44:@47846.4]
  wire [31:0] accel_io_axiStreamsOut_0_TSTRB; // @[Instantiator.scala 53:44:@47846.4]
  wire [31:0] accel_io_axiStreamsOut_0_TKEEP; // @[Instantiator.scala 53:44:@47846.4]
  wire  accel_io_axiStreamsOut_0_TLAST; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_axiStreamsOut_0_TID; // @[Instantiator.scala 53:44:@47846.4]
  wire [7:0] accel_io_axiStreamsOut_0_TDEST; // @[Instantiator.scala 53:44:@47846.4]
  wire [31:0] accel_io_axiStreamsOut_0_TUSER; // @[Instantiator.scala 53:44:@47846.4]
  wire  accel_io_heap_0_req_valid; // @[Instantiator.scala 53:44:@47846.4]
  wire  accel_io_heap_0_req_bits_allocDealloc; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_heap_0_req_bits_sizeAddr; // @[Instantiator.scala 53:44:@47846.4]
  wire  accel_io_heap_0_resp_valid; // @[Instantiator.scala 53:44:@47846.4]
  wire  accel_io_heap_0_resp_bits_allocDealloc; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_heap_0_resp_bits_sizeAddr; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_argIns_0; // @[Instantiator.scala 53:44:@47846.4]
  wire  accel_io_argOuts_0_port_ready; // @[Instantiator.scala 53:44:@47846.4]
  wire  accel_io_argOuts_0_port_valid; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_argOuts_0_port_bits; // @[Instantiator.scala 53:44:@47846.4]
  wire [63:0] accel_io_argOuts_0_echo; // @[Instantiator.scala 53:44:@47846.4]
  wire  Fringe_clock; // @[SimTarget.scala 16:24:@48290.4]
  wire  Fringe_reset; // @[SimTarget.scala 16:24:@48290.4]
  wire [31:0] Fringe_io_raddr; // @[SimTarget.scala 16:24:@48290.4]
  wire  Fringe_io_wen; // @[SimTarget.scala 16:24:@48290.4]
  wire [31:0] Fringe_io_waddr; // @[SimTarget.scala 16:24:@48290.4]
  wire [63:0] Fringe_io_wdata; // @[SimTarget.scala 16:24:@48290.4]
  wire [63:0] Fringe_io_rdata; // @[SimTarget.scala 16:24:@48290.4]
  wire  Fringe_io_enable; // @[SimTarget.scala 16:24:@48290.4]
  wire  Fringe_io_done; // @[SimTarget.scala 16:24:@48290.4]
  wire  Fringe_io_reset; // @[SimTarget.scala 16:24:@48290.4]
  wire [63:0] Fringe_io_argIns_0; // @[SimTarget.scala 16:24:@48290.4]
  wire  Fringe_io_argOuts_0_valid; // @[SimTarget.scala 16:24:@48290.4]
  wire [63:0] Fringe_io_argOuts_0_bits; // @[SimTarget.scala 16:24:@48290.4]
  wire [63:0] Fringe_io_argEchos_0; // @[SimTarget.scala 16:24:@48290.4]
  wire  Fringe_io_heap_0_req_valid; // @[SimTarget.scala 16:24:@48290.4]
  wire  Fringe_io_heap_0_req_bits_allocDealloc; // @[SimTarget.scala 16:24:@48290.4]
  wire [63:0] Fringe_io_heap_0_req_bits_sizeAddr; // @[SimTarget.scala 16:24:@48290.4]
  wire  Fringe_io_heap_0_resp_valid; // @[SimTarget.scala 16:24:@48290.4]
  wire  Fringe_io_heap_0_resp_bits_allocDealloc; // @[SimTarget.scala 16:24:@48290.4]
  wire [63:0] Fringe_io_heap_0_resp_bits_sizeAddr; // @[SimTarget.scala 16:24:@48290.4]
  AccelUnit accel ( // @[Instantiator.scala 53:44:@47846.4]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_enable(accel_io_enable),
    .io_done(accel_io_done),
    .io_reset(accel_io_reset),
    .io_memStreams_loads_0_cmd_ready(accel_io_memStreams_loads_0_cmd_ready),
    .io_memStreams_loads_0_cmd_valid(accel_io_memStreams_loads_0_cmd_valid),
    .io_memStreams_loads_0_cmd_bits_addr(accel_io_memStreams_loads_0_cmd_bits_addr),
    .io_memStreams_loads_0_cmd_bits_size(accel_io_memStreams_loads_0_cmd_bits_size),
    .io_memStreams_loads_0_data_ready(accel_io_memStreams_loads_0_data_ready),
    .io_memStreams_loads_0_data_valid(accel_io_memStreams_loads_0_data_valid),
    .io_memStreams_loads_0_data_bits_rdata_0(accel_io_memStreams_loads_0_data_bits_rdata_0),
    .io_memStreams_loads_0_data_bits_rdata_1(accel_io_memStreams_loads_0_data_bits_rdata_1),
    .io_memStreams_loads_0_data_bits_rdata_2(accel_io_memStreams_loads_0_data_bits_rdata_2),
    .io_memStreams_loads_0_data_bits_rdata_3(accel_io_memStreams_loads_0_data_bits_rdata_3),
    .io_memStreams_loads_0_data_bits_rdata_4(accel_io_memStreams_loads_0_data_bits_rdata_4),
    .io_memStreams_loads_0_data_bits_rdata_5(accel_io_memStreams_loads_0_data_bits_rdata_5),
    .io_memStreams_loads_0_data_bits_rdata_6(accel_io_memStreams_loads_0_data_bits_rdata_6),
    .io_memStreams_loads_0_data_bits_rdata_7(accel_io_memStreams_loads_0_data_bits_rdata_7),
    .io_memStreams_loads_0_data_bits_rdata_8(accel_io_memStreams_loads_0_data_bits_rdata_8),
    .io_memStreams_loads_0_data_bits_rdata_9(accel_io_memStreams_loads_0_data_bits_rdata_9),
    .io_memStreams_loads_0_data_bits_rdata_10(accel_io_memStreams_loads_0_data_bits_rdata_10),
    .io_memStreams_loads_0_data_bits_rdata_11(accel_io_memStreams_loads_0_data_bits_rdata_11),
    .io_memStreams_loads_0_data_bits_rdata_12(accel_io_memStreams_loads_0_data_bits_rdata_12),
    .io_memStreams_loads_0_data_bits_rdata_13(accel_io_memStreams_loads_0_data_bits_rdata_13),
    .io_memStreams_loads_0_data_bits_rdata_14(accel_io_memStreams_loads_0_data_bits_rdata_14),
    .io_memStreams_loads_0_data_bits_rdata_15(accel_io_memStreams_loads_0_data_bits_rdata_15),
    .io_memStreams_loads_0_data_bits_rdata_16(accel_io_memStreams_loads_0_data_bits_rdata_16),
    .io_memStreams_loads_0_data_bits_rdata_17(accel_io_memStreams_loads_0_data_bits_rdata_17),
    .io_memStreams_loads_0_data_bits_rdata_18(accel_io_memStreams_loads_0_data_bits_rdata_18),
    .io_memStreams_loads_0_data_bits_rdata_19(accel_io_memStreams_loads_0_data_bits_rdata_19),
    .io_memStreams_loads_0_data_bits_rdata_20(accel_io_memStreams_loads_0_data_bits_rdata_20),
    .io_memStreams_loads_0_data_bits_rdata_21(accel_io_memStreams_loads_0_data_bits_rdata_21),
    .io_memStreams_loads_0_data_bits_rdata_22(accel_io_memStreams_loads_0_data_bits_rdata_22),
    .io_memStreams_loads_0_data_bits_rdata_23(accel_io_memStreams_loads_0_data_bits_rdata_23),
    .io_memStreams_loads_0_data_bits_rdata_24(accel_io_memStreams_loads_0_data_bits_rdata_24),
    .io_memStreams_loads_0_data_bits_rdata_25(accel_io_memStreams_loads_0_data_bits_rdata_25),
    .io_memStreams_loads_0_data_bits_rdata_26(accel_io_memStreams_loads_0_data_bits_rdata_26),
    .io_memStreams_loads_0_data_bits_rdata_27(accel_io_memStreams_loads_0_data_bits_rdata_27),
    .io_memStreams_loads_0_data_bits_rdata_28(accel_io_memStreams_loads_0_data_bits_rdata_28),
    .io_memStreams_loads_0_data_bits_rdata_29(accel_io_memStreams_loads_0_data_bits_rdata_29),
    .io_memStreams_loads_0_data_bits_rdata_30(accel_io_memStreams_loads_0_data_bits_rdata_30),
    .io_memStreams_loads_0_data_bits_rdata_31(accel_io_memStreams_loads_0_data_bits_rdata_31),
    .io_memStreams_loads_0_data_bits_rdata_32(accel_io_memStreams_loads_0_data_bits_rdata_32),
    .io_memStreams_loads_0_data_bits_rdata_33(accel_io_memStreams_loads_0_data_bits_rdata_33),
    .io_memStreams_loads_0_data_bits_rdata_34(accel_io_memStreams_loads_0_data_bits_rdata_34),
    .io_memStreams_loads_0_data_bits_rdata_35(accel_io_memStreams_loads_0_data_bits_rdata_35),
    .io_memStreams_loads_0_data_bits_rdata_36(accel_io_memStreams_loads_0_data_bits_rdata_36),
    .io_memStreams_loads_0_data_bits_rdata_37(accel_io_memStreams_loads_0_data_bits_rdata_37),
    .io_memStreams_loads_0_data_bits_rdata_38(accel_io_memStreams_loads_0_data_bits_rdata_38),
    .io_memStreams_loads_0_data_bits_rdata_39(accel_io_memStreams_loads_0_data_bits_rdata_39),
    .io_memStreams_loads_0_data_bits_rdata_40(accel_io_memStreams_loads_0_data_bits_rdata_40),
    .io_memStreams_loads_0_data_bits_rdata_41(accel_io_memStreams_loads_0_data_bits_rdata_41),
    .io_memStreams_loads_0_data_bits_rdata_42(accel_io_memStreams_loads_0_data_bits_rdata_42),
    .io_memStreams_loads_0_data_bits_rdata_43(accel_io_memStreams_loads_0_data_bits_rdata_43),
    .io_memStreams_loads_0_data_bits_rdata_44(accel_io_memStreams_loads_0_data_bits_rdata_44),
    .io_memStreams_loads_0_data_bits_rdata_45(accel_io_memStreams_loads_0_data_bits_rdata_45),
    .io_memStreams_loads_0_data_bits_rdata_46(accel_io_memStreams_loads_0_data_bits_rdata_46),
    .io_memStreams_loads_0_data_bits_rdata_47(accel_io_memStreams_loads_0_data_bits_rdata_47),
    .io_memStreams_loads_0_data_bits_rdata_48(accel_io_memStreams_loads_0_data_bits_rdata_48),
    .io_memStreams_loads_0_data_bits_rdata_49(accel_io_memStreams_loads_0_data_bits_rdata_49),
    .io_memStreams_loads_0_data_bits_rdata_50(accel_io_memStreams_loads_0_data_bits_rdata_50),
    .io_memStreams_loads_0_data_bits_rdata_51(accel_io_memStreams_loads_0_data_bits_rdata_51),
    .io_memStreams_loads_0_data_bits_rdata_52(accel_io_memStreams_loads_0_data_bits_rdata_52),
    .io_memStreams_loads_0_data_bits_rdata_53(accel_io_memStreams_loads_0_data_bits_rdata_53),
    .io_memStreams_loads_0_data_bits_rdata_54(accel_io_memStreams_loads_0_data_bits_rdata_54),
    .io_memStreams_loads_0_data_bits_rdata_55(accel_io_memStreams_loads_0_data_bits_rdata_55),
    .io_memStreams_loads_0_data_bits_rdata_56(accel_io_memStreams_loads_0_data_bits_rdata_56),
    .io_memStreams_loads_0_data_bits_rdata_57(accel_io_memStreams_loads_0_data_bits_rdata_57),
    .io_memStreams_loads_0_data_bits_rdata_58(accel_io_memStreams_loads_0_data_bits_rdata_58),
    .io_memStreams_loads_0_data_bits_rdata_59(accel_io_memStreams_loads_0_data_bits_rdata_59),
    .io_memStreams_loads_0_data_bits_rdata_60(accel_io_memStreams_loads_0_data_bits_rdata_60),
    .io_memStreams_loads_0_data_bits_rdata_61(accel_io_memStreams_loads_0_data_bits_rdata_61),
    .io_memStreams_loads_0_data_bits_rdata_62(accel_io_memStreams_loads_0_data_bits_rdata_62),
    .io_memStreams_loads_0_data_bits_rdata_63(accel_io_memStreams_loads_0_data_bits_rdata_63),
    .io_memStreams_stores_0_cmd_ready(accel_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(accel_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(accel_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(accel_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(accel_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(accel_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(accel_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wdata_1(accel_io_memStreams_stores_0_data_bits_wdata_1),
    .io_memStreams_stores_0_data_bits_wdata_2(accel_io_memStreams_stores_0_data_bits_wdata_2),
    .io_memStreams_stores_0_data_bits_wdata_3(accel_io_memStreams_stores_0_data_bits_wdata_3),
    .io_memStreams_stores_0_data_bits_wdata_4(accel_io_memStreams_stores_0_data_bits_wdata_4),
    .io_memStreams_stores_0_data_bits_wdata_5(accel_io_memStreams_stores_0_data_bits_wdata_5),
    .io_memStreams_stores_0_data_bits_wdata_6(accel_io_memStreams_stores_0_data_bits_wdata_6),
    .io_memStreams_stores_0_data_bits_wdata_7(accel_io_memStreams_stores_0_data_bits_wdata_7),
    .io_memStreams_stores_0_data_bits_wdata_8(accel_io_memStreams_stores_0_data_bits_wdata_8),
    .io_memStreams_stores_0_data_bits_wdata_9(accel_io_memStreams_stores_0_data_bits_wdata_9),
    .io_memStreams_stores_0_data_bits_wdata_10(accel_io_memStreams_stores_0_data_bits_wdata_10),
    .io_memStreams_stores_0_data_bits_wdata_11(accel_io_memStreams_stores_0_data_bits_wdata_11),
    .io_memStreams_stores_0_data_bits_wdata_12(accel_io_memStreams_stores_0_data_bits_wdata_12),
    .io_memStreams_stores_0_data_bits_wdata_13(accel_io_memStreams_stores_0_data_bits_wdata_13),
    .io_memStreams_stores_0_data_bits_wdata_14(accel_io_memStreams_stores_0_data_bits_wdata_14),
    .io_memStreams_stores_0_data_bits_wdata_15(accel_io_memStreams_stores_0_data_bits_wdata_15),
    .io_memStreams_stores_0_data_bits_wdata_16(accel_io_memStreams_stores_0_data_bits_wdata_16),
    .io_memStreams_stores_0_data_bits_wdata_17(accel_io_memStreams_stores_0_data_bits_wdata_17),
    .io_memStreams_stores_0_data_bits_wdata_18(accel_io_memStreams_stores_0_data_bits_wdata_18),
    .io_memStreams_stores_0_data_bits_wdata_19(accel_io_memStreams_stores_0_data_bits_wdata_19),
    .io_memStreams_stores_0_data_bits_wdata_20(accel_io_memStreams_stores_0_data_bits_wdata_20),
    .io_memStreams_stores_0_data_bits_wdata_21(accel_io_memStreams_stores_0_data_bits_wdata_21),
    .io_memStreams_stores_0_data_bits_wdata_22(accel_io_memStreams_stores_0_data_bits_wdata_22),
    .io_memStreams_stores_0_data_bits_wdata_23(accel_io_memStreams_stores_0_data_bits_wdata_23),
    .io_memStreams_stores_0_data_bits_wdata_24(accel_io_memStreams_stores_0_data_bits_wdata_24),
    .io_memStreams_stores_0_data_bits_wdata_25(accel_io_memStreams_stores_0_data_bits_wdata_25),
    .io_memStreams_stores_0_data_bits_wdata_26(accel_io_memStreams_stores_0_data_bits_wdata_26),
    .io_memStreams_stores_0_data_bits_wdata_27(accel_io_memStreams_stores_0_data_bits_wdata_27),
    .io_memStreams_stores_0_data_bits_wdata_28(accel_io_memStreams_stores_0_data_bits_wdata_28),
    .io_memStreams_stores_0_data_bits_wdata_29(accel_io_memStreams_stores_0_data_bits_wdata_29),
    .io_memStreams_stores_0_data_bits_wdata_30(accel_io_memStreams_stores_0_data_bits_wdata_30),
    .io_memStreams_stores_0_data_bits_wdata_31(accel_io_memStreams_stores_0_data_bits_wdata_31),
    .io_memStreams_stores_0_data_bits_wdata_32(accel_io_memStreams_stores_0_data_bits_wdata_32),
    .io_memStreams_stores_0_data_bits_wdata_33(accel_io_memStreams_stores_0_data_bits_wdata_33),
    .io_memStreams_stores_0_data_bits_wdata_34(accel_io_memStreams_stores_0_data_bits_wdata_34),
    .io_memStreams_stores_0_data_bits_wdata_35(accel_io_memStreams_stores_0_data_bits_wdata_35),
    .io_memStreams_stores_0_data_bits_wdata_36(accel_io_memStreams_stores_0_data_bits_wdata_36),
    .io_memStreams_stores_0_data_bits_wdata_37(accel_io_memStreams_stores_0_data_bits_wdata_37),
    .io_memStreams_stores_0_data_bits_wdata_38(accel_io_memStreams_stores_0_data_bits_wdata_38),
    .io_memStreams_stores_0_data_bits_wdata_39(accel_io_memStreams_stores_0_data_bits_wdata_39),
    .io_memStreams_stores_0_data_bits_wdata_40(accel_io_memStreams_stores_0_data_bits_wdata_40),
    .io_memStreams_stores_0_data_bits_wdata_41(accel_io_memStreams_stores_0_data_bits_wdata_41),
    .io_memStreams_stores_0_data_bits_wdata_42(accel_io_memStreams_stores_0_data_bits_wdata_42),
    .io_memStreams_stores_0_data_bits_wdata_43(accel_io_memStreams_stores_0_data_bits_wdata_43),
    .io_memStreams_stores_0_data_bits_wdata_44(accel_io_memStreams_stores_0_data_bits_wdata_44),
    .io_memStreams_stores_0_data_bits_wdata_45(accel_io_memStreams_stores_0_data_bits_wdata_45),
    .io_memStreams_stores_0_data_bits_wdata_46(accel_io_memStreams_stores_0_data_bits_wdata_46),
    .io_memStreams_stores_0_data_bits_wdata_47(accel_io_memStreams_stores_0_data_bits_wdata_47),
    .io_memStreams_stores_0_data_bits_wdata_48(accel_io_memStreams_stores_0_data_bits_wdata_48),
    .io_memStreams_stores_0_data_bits_wdata_49(accel_io_memStreams_stores_0_data_bits_wdata_49),
    .io_memStreams_stores_0_data_bits_wdata_50(accel_io_memStreams_stores_0_data_bits_wdata_50),
    .io_memStreams_stores_0_data_bits_wdata_51(accel_io_memStreams_stores_0_data_bits_wdata_51),
    .io_memStreams_stores_0_data_bits_wdata_52(accel_io_memStreams_stores_0_data_bits_wdata_52),
    .io_memStreams_stores_0_data_bits_wdata_53(accel_io_memStreams_stores_0_data_bits_wdata_53),
    .io_memStreams_stores_0_data_bits_wdata_54(accel_io_memStreams_stores_0_data_bits_wdata_54),
    .io_memStreams_stores_0_data_bits_wdata_55(accel_io_memStreams_stores_0_data_bits_wdata_55),
    .io_memStreams_stores_0_data_bits_wdata_56(accel_io_memStreams_stores_0_data_bits_wdata_56),
    .io_memStreams_stores_0_data_bits_wdata_57(accel_io_memStreams_stores_0_data_bits_wdata_57),
    .io_memStreams_stores_0_data_bits_wdata_58(accel_io_memStreams_stores_0_data_bits_wdata_58),
    .io_memStreams_stores_0_data_bits_wdata_59(accel_io_memStreams_stores_0_data_bits_wdata_59),
    .io_memStreams_stores_0_data_bits_wdata_60(accel_io_memStreams_stores_0_data_bits_wdata_60),
    .io_memStreams_stores_0_data_bits_wdata_61(accel_io_memStreams_stores_0_data_bits_wdata_61),
    .io_memStreams_stores_0_data_bits_wdata_62(accel_io_memStreams_stores_0_data_bits_wdata_62),
    .io_memStreams_stores_0_data_bits_wdata_63(accel_io_memStreams_stores_0_data_bits_wdata_63),
    .io_memStreams_stores_0_data_bits_wstrb(accel_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(accel_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(accel_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(accel_io_memStreams_stores_0_wresp_bits),
    .io_memStreams_gathers_0_cmd_ready(accel_io_memStreams_gathers_0_cmd_ready),
    .io_memStreams_gathers_0_cmd_valid(accel_io_memStreams_gathers_0_cmd_valid),
    .io_memStreams_gathers_0_cmd_bits_addr_0(accel_io_memStreams_gathers_0_cmd_bits_addr_0),
    .io_memStreams_gathers_0_cmd_bits_addr_1(accel_io_memStreams_gathers_0_cmd_bits_addr_1),
    .io_memStreams_gathers_0_cmd_bits_addr_2(accel_io_memStreams_gathers_0_cmd_bits_addr_2),
    .io_memStreams_gathers_0_cmd_bits_addr_3(accel_io_memStreams_gathers_0_cmd_bits_addr_3),
    .io_memStreams_gathers_0_cmd_bits_addr_4(accel_io_memStreams_gathers_0_cmd_bits_addr_4),
    .io_memStreams_gathers_0_cmd_bits_addr_5(accel_io_memStreams_gathers_0_cmd_bits_addr_5),
    .io_memStreams_gathers_0_cmd_bits_addr_6(accel_io_memStreams_gathers_0_cmd_bits_addr_6),
    .io_memStreams_gathers_0_cmd_bits_addr_7(accel_io_memStreams_gathers_0_cmd_bits_addr_7),
    .io_memStreams_gathers_0_cmd_bits_addr_8(accel_io_memStreams_gathers_0_cmd_bits_addr_8),
    .io_memStreams_gathers_0_cmd_bits_addr_9(accel_io_memStreams_gathers_0_cmd_bits_addr_9),
    .io_memStreams_gathers_0_cmd_bits_addr_10(accel_io_memStreams_gathers_0_cmd_bits_addr_10),
    .io_memStreams_gathers_0_cmd_bits_addr_11(accel_io_memStreams_gathers_0_cmd_bits_addr_11),
    .io_memStreams_gathers_0_cmd_bits_addr_12(accel_io_memStreams_gathers_0_cmd_bits_addr_12),
    .io_memStreams_gathers_0_cmd_bits_addr_13(accel_io_memStreams_gathers_0_cmd_bits_addr_13),
    .io_memStreams_gathers_0_cmd_bits_addr_14(accel_io_memStreams_gathers_0_cmd_bits_addr_14),
    .io_memStreams_gathers_0_cmd_bits_addr_15(accel_io_memStreams_gathers_0_cmd_bits_addr_15),
    .io_memStreams_gathers_0_cmd_bits_addr_16(accel_io_memStreams_gathers_0_cmd_bits_addr_16),
    .io_memStreams_gathers_0_cmd_bits_addr_17(accel_io_memStreams_gathers_0_cmd_bits_addr_17),
    .io_memStreams_gathers_0_cmd_bits_addr_18(accel_io_memStreams_gathers_0_cmd_bits_addr_18),
    .io_memStreams_gathers_0_cmd_bits_addr_19(accel_io_memStreams_gathers_0_cmd_bits_addr_19),
    .io_memStreams_gathers_0_cmd_bits_addr_20(accel_io_memStreams_gathers_0_cmd_bits_addr_20),
    .io_memStreams_gathers_0_cmd_bits_addr_21(accel_io_memStreams_gathers_0_cmd_bits_addr_21),
    .io_memStreams_gathers_0_cmd_bits_addr_22(accel_io_memStreams_gathers_0_cmd_bits_addr_22),
    .io_memStreams_gathers_0_cmd_bits_addr_23(accel_io_memStreams_gathers_0_cmd_bits_addr_23),
    .io_memStreams_gathers_0_cmd_bits_addr_24(accel_io_memStreams_gathers_0_cmd_bits_addr_24),
    .io_memStreams_gathers_0_cmd_bits_addr_25(accel_io_memStreams_gathers_0_cmd_bits_addr_25),
    .io_memStreams_gathers_0_cmd_bits_addr_26(accel_io_memStreams_gathers_0_cmd_bits_addr_26),
    .io_memStreams_gathers_0_cmd_bits_addr_27(accel_io_memStreams_gathers_0_cmd_bits_addr_27),
    .io_memStreams_gathers_0_cmd_bits_addr_28(accel_io_memStreams_gathers_0_cmd_bits_addr_28),
    .io_memStreams_gathers_0_cmd_bits_addr_29(accel_io_memStreams_gathers_0_cmd_bits_addr_29),
    .io_memStreams_gathers_0_cmd_bits_addr_30(accel_io_memStreams_gathers_0_cmd_bits_addr_30),
    .io_memStreams_gathers_0_cmd_bits_addr_31(accel_io_memStreams_gathers_0_cmd_bits_addr_31),
    .io_memStreams_gathers_0_cmd_bits_addr_32(accel_io_memStreams_gathers_0_cmd_bits_addr_32),
    .io_memStreams_gathers_0_cmd_bits_addr_33(accel_io_memStreams_gathers_0_cmd_bits_addr_33),
    .io_memStreams_gathers_0_cmd_bits_addr_34(accel_io_memStreams_gathers_0_cmd_bits_addr_34),
    .io_memStreams_gathers_0_cmd_bits_addr_35(accel_io_memStreams_gathers_0_cmd_bits_addr_35),
    .io_memStreams_gathers_0_cmd_bits_addr_36(accel_io_memStreams_gathers_0_cmd_bits_addr_36),
    .io_memStreams_gathers_0_cmd_bits_addr_37(accel_io_memStreams_gathers_0_cmd_bits_addr_37),
    .io_memStreams_gathers_0_cmd_bits_addr_38(accel_io_memStreams_gathers_0_cmd_bits_addr_38),
    .io_memStreams_gathers_0_cmd_bits_addr_39(accel_io_memStreams_gathers_0_cmd_bits_addr_39),
    .io_memStreams_gathers_0_cmd_bits_addr_40(accel_io_memStreams_gathers_0_cmd_bits_addr_40),
    .io_memStreams_gathers_0_cmd_bits_addr_41(accel_io_memStreams_gathers_0_cmd_bits_addr_41),
    .io_memStreams_gathers_0_cmd_bits_addr_42(accel_io_memStreams_gathers_0_cmd_bits_addr_42),
    .io_memStreams_gathers_0_cmd_bits_addr_43(accel_io_memStreams_gathers_0_cmd_bits_addr_43),
    .io_memStreams_gathers_0_cmd_bits_addr_44(accel_io_memStreams_gathers_0_cmd_bits_addr_44),
    .io_memStreams_gathers_0_cmd_bits_addr_45(accel_io_memStreams_gathers_0_cmd_bits_addr_45),
    .io_memStreams_gathers_0_cmd_bits_addr_46(accel_io_memStreams_gathers_0_cmd_bits_addr_46),
    .io_memStreams_gathers_0_cmd_bits_addr_47(accel_io_memStreams_gathers_0_cmd_bits_addr_47),
    .io_memStreams_gathers_0_cmd_bits_addr_48(accel_io_memStreams_gathers_0_cmd_bits_addr_48),
    .io_memStreams_gathers_0_cmd_bits_addr_49(accel_io_memStreams_gathers_0_cmd_bits_addr_49),
    .io_memStreams_gathers_0_cmd_bits_addr_50(accel_io_memStreams_gathers_0_cmd_bits_addr_50),
    .io_memStreams_gathers_0_cmd_bits_addr_51(accel_io_memStreams_gathers_0_cmd_bits_addr_51),
    .io_memStreams_gathers_0_cmd_bits_addr_52(accel_io_memStreams_gathers_0_cmd_bits_addr_52),
    .io_memStreams_gathers_0_cmd_bits_addr_53(accel_io_memStreams_gathers_0_cmd_bits_addr_53),
    .io_memStreams_gathers_0_cmd_bits_addr_54(accel_io_memStreams_gathers_0_cmd_bits_addr_54),
    .io_memStreams_gathers_0_cmd_bits_addr_55(accel_io_memStreams_gathers_0_cmd_bits_addr_55),
    .io_memStreams_gathers_0_cmd_bits_addr_56(accel_io_memStreams_gathers_0_cmd_bits_addr_56),
    .io_memStreams_gathers_0_cmd_bits_addr_57(accel_io_memStreams_gathers_0_cmd_bits_addr_57),
    .io_memStreams_gathers_0_cmd_bits_addr_58(accel_io_memStreams_gathers_0_cmd_bits_addr_58),
    .io_memStreams_gathers_0_cmd_bits_addr_59(accel_io_memStreams_gathers_0_cmd_bits_addr_59),
    .io_memStreams_gathers_0_cmd_bits_addr_60(accel_io_memStreams_gathers_0_cmd_bits_addr_60),
    .io_memStreams_gathers_0_cmd_bits_addr_61(accel_io_memStreams_gathers_0_cmd_bits_addr_61),
    .io_memStreams_gathers_0_cmd_bits_addr_62(accel_io_memStreams_gathers_0_cmd_bits_addr_62),
    .io_memStreams_gathers_0_cmd_bits_addr_63(accel_io_memStreams_gathers_0_cmd_bits_addr_63),
    .io_memStreams_gathers_0_data_ready(accel_io_memStreams_gathers_0_data_ready),
    .io_memStreams_gathers_0_data_valid(accel_io_memStreams_gathers_0_data_valid),
    .io_memStreams_gathers_0_data_bits_0(accel_io_memStreams_gathers_0_data_bits_0),
    .io_memStreams_gathers_0_data_bits_1(accel_io_memStreams_gathers_0_data_bits_1),
    .io_memStreams_gathers_0_data_bits_2(accel_io_memStreams_gathers_0_data_bits_2),
    .io_memStreams_gathers_0_data_bits_3(accel_io_memStreams_gathers_0_data_bits_3),
    .io_memStreams_gathers_0_data_bits_4(accel_io_memStreams_gathers_0_data_bits_4),
    .io_memStreams_gathers_0_data_bits_5(accel_io_memStreams_gathers_0_data_bits_5),
    .io_memStreams_gathers_0_data_bits_6(accel_io_memStreams_gathers_0_data_bits_6),
    .io_memStreams_gathers_0_data_bits_7(accel_io_memStreams_gathers_0_data_bits_7),
    .io_memStreams_gathers_0_data_bits_8(accel_io_memStreams_gathers_0_data_bits_8),
    .io_memStreams_gathers_0_data_bits_9(accel_io_memStreams_gathers_0_data_bits_9),
    .io_memStreams_gathers_0_data_bits_10(accel_io_memStreams_gathers_0_data_bits_10),
    .io_memStreams_gathers_0_data_bits_11(accel_io_memStreams_gathers_0_data_bits_11),
    .io_memStreams_gathers_0_data_bits_12(accel_io_memStreams_gathers_0_data_bits_12),
    .io_memStreams_gathers_0_data_bits_13(accel_io_memStreams_gathers_0_data_bits_13),
    .io_memStreams_gathers_0_data_bits_14(accel_io_memStreams_gathers_0_data_bits_14),
    .io_memStreams_gathers_0_data_bits_15(accel_io_memStreams_gathers_0_data_bits_15),
    .io_memStreams_gathers_0_data_bits_16(accel_io_memStreams_gathers_0_data_bits_16),
    .io_memStreams_gathers_0_data_bits_17(accel_io_memStreams_gathers_0_data_bits_17),
    .io_memStreams_gathers_0_data_bits_18(accel_io_memStreams_gathers_0_data_bits_18),
    .io_memStreams_gathers_0_data_bits_19(accel_io_memStreams_gathers_0_data_bits_19),
    .io_memStreams_gathers_0_data_bits_20(accel_io_memStreams_gathers_0_data_bits_20),
    .io_memStreams_gathers_0_data_bits_21(accel_io_memStreams_gathers_0_data_bits_21),
    .io_memStreams_gathers_0_data_bits_22(accel_io_memStreams_gathers_0_data_bits_22),
    .io_memStreams_gathers_0_data_bits_23(accel_io_memStreams_gathers_0_data_bits_23),
    .io_memStreams_gathers_0_data_bits_24(accel_io_memStreams_gathers_0_data_bits_24),
    .io_memStreams_gathers_0_data_bits_25(accel_io_memStreams_gathers_0_data_bits_25),
    .io_memStreams_gathers_0_data_bits_26(accel_io_memStreams_gathers_0_data_bits_26),
    .io_memStreams_gathers_0_data_bits_27(accel_io_memStreams_gathers_0_data_bits_27),
    .io_memStreams_gathers_0_data_bits_28(accel_io_memStreams_gathers_0_data_bits_28),
    .io_memStreams_gathers_0_data_bits_29(accel_io_memStreams_gathers_0_data_bits_29),
    .io_memStreams_gathers_0_data_bits_30(accel_io_memStreams_gathers_0_data_bits_30),
    .io_memStreams_gathers_0_data_bits_31(accel_io_memStreams_gathers_0_data_bits_31),
    .io_memStreams_gathers_0_data_bits_32(accel_io_memStreams_gathers_0_data_bits_32),
    .io_memStreams_gathers_0_data_bits_33(accel_io_memStreams_gathers_0_data_bits_33),
    .io_memStreams_gathers_0_data_bits_34(accel_io_memStreams_gathers_0_data_bits_34),
    .io_memStreams_gathers_0_data_bits_35(accel_io_memStreams_gathers_0_data_bits_35),
    .io_memStreams_gathers_0_data_bits_36(accel_io_memStreams_gathers_0_data_bits_36),
    .io_memStreams_gathers_0_data_bits_37(accel_io_memStreams_gathers_0_data_bits_37),
    .io_memStreams_gathers_0_data_bits_38(accel_io_memStreams_gathers_0_data_bits_38),
    .io_memStreams_gathers_0_data_bits_39(accel_io_memStreams_gathers_0_data_bits_39),
    .io_memStreams_gathers_0_data_bits_40(accel_io_memStreams_gathers_0_data_bits_40),
    .io_memStreams_gathers_0_data_bits_41(accel_io_memStreams_gathers_0_data_bits_41),
    .io_memStreams_gathers_0_data_bits_42(accel_io_memStreams_gathers_0_data_bits_42),
    .io_memStreams_gathers_0_data_bits_43(accel_io_memStreams_gathers_0_data_bits_43),
    .io_memStreams_gathers_0_data_bits_44(accel_io_memStreams_gathers_0_data_bits_44),
    .io_memStreams_gathers_0_data_bits_45(accel_io_memStreams_gathers_0_data_bits_45),
    .io_memStreams_gathers_0_data_bits_46(accel_io_memStreams_gathers_0_data_bits_46),
    .io_memStreams_gathers_0_data_bits_47(accel_io_memStreams_gathers_0_data_bits_47),
    .io_memStreams_gathers_0_data_bits_48(accel_io_memStreams_gathers_0_data_bits_48),
    .io_memStreams_gathers_0_data_bits_49(accel_io_memStreams_gathers_0_data_bits_49),
    .io_memStreams_gathers_0_data_bits_50(accel_io_memStreams_gathers_0_data_bits_50),
    .io_memStreams_gathers_0_data_bits_51(accel_io_memStreams_gathers_0_data_bits_51),
    .io_memStreams_gathers_0_data_bits_52(accel_io_memStreams_gathers_0_data_bits_52),
    .io_memStreams_gathers_0_data_bits_53(accel_io_memStreams_gathers_0_data_bits_53),
    .io_memStreams_gathers_0_data_bits_54(accel_io_memStreams_gathers_0_data_bits_54),
    .io_memStreams_gathers_0_data_bits_55(accel_io_memStreams_gathers_0_data_bits_55),
    .io_memStreams_gathers_0_data_bits_56(accel_io_memStreams_gathers_0_data_bits_56),
    .io_memStreams_gathers_0_data_bits_57(accel_io_memStreams_gathers_0_data_bits_57),
    .io_memStreams_gathers_0_data_bits_58(accel_io_memStreams_gathers_0_data_bits_58),
    .io_memStreams_gathers_0_data_bits_59(accel_io_memStreams_gathers_0_data_bits_59),
    .io_memStreams_gathers_0_data_bits_60(accel_io_memStreams_gathers_0_data_bits_60),
    .io_memStreams_gathers_0_data_bits_61(accel_io_memStreams_gathers_0_data_bits_61),
    .io_memStreams_gathers_0_data_bits_62(accel_io_memStreams_gathers_0_data_bits_62),
    .io_memStreams_gathers_0_data_bits_63(accel_io_memStreams_gathers_0_data_bits_63),
    .io_memStreams_scatters_0_cmd_ready(accel_io_memStreams_scatters_0_cmd_ready),
    .io_memStreams_scatters_0_cmd_valid(accel_io_memStreams_scatters_0_cmd_valid),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_0(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_1(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_2(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_3(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_4(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_5(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_6(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_7(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_8(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_9(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_10(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_11(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_12(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_13(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_14(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_15(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_16(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_16),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_17(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_17),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_18(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_18),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_19(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_19),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_20(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_20),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_21(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_21),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_22(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_22),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_23(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_23),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_24(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_24),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_25(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_25),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_26(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_26),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_27(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_27),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_28(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_28),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_29(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_29),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_30(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_30),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_31(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_31),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_32(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_32),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_33(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_33),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_34(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_34),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_35(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_35),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_36(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_36),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_37(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_37),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_38(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_38),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_39(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_39),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_40(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_40),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_41(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_41),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_42(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_42),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_43(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_43),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_44(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_44),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_45(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_45),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_46(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_46),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_47(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_47),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_48(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_48),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_49(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_49),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_50(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_50),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_51(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_51),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_52(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_52),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_53(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_53),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_54(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_54),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_55(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_55),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_56(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_56),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_57(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_57),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_58(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_58),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_59(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_59),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_60(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_60),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_61(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_61),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_62(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_62),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_63(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_63),
    .io_memStreams_scatters_0_cmd_bits_wdata_0(accel_io_memStreams_scatters_0_cmd_bits_wdata_0),
    .io_memStreams_scatters_0_cmd_bits_wdata_1(accel_io_memStreams_scatters_0_cmd_bits_wdata_1),
    .io_memStreams_scatters_0_cmd_bits_wdata_2(accel_io_memStreams_scatters_0_cmd_bits_wdata_2),
    .io_memStreams_scatters_0_cmd_bits_wdata_3(accel_io_memStreams_scatters_0_cmd_bits_wdata_3),
    .io_memStreams_scatters_0_cmd_bits_wdata_4(accel_io_memStreams_scatters_0_cmd_bits_wdata_4),
    .io_memStreams_scatters_0_cmd_bits_wdata_5(accel_io_memStreams_scatters_0_cmd_bits_wdata_5),
    .io_memStreams_scatters_0_cmd_bits_wdata_6(accel_io_memStreams_scatters_0_cmd_bits_wdata_6),
    .io_memStreams_scatters_0_cmd_bits_wdata_7(accel_io_memStreams_scatters_0_cmd_bits_wdata_7),
    .io_memStreams_scatters_0_cmd_bits_wdata_8(accel_io_memStreams_scatters_0_cmd_bits_wdata_8),
    .io_memStreams_scatters_0_cmd_bits_wdata_9(accel_io_memStreams_scatters_0_cmd_bits_wdata_9),
    .io_memStreams_scatters_0_cmd_bits_wdata_10(accel_io_memStreams_scatters_0_cmd_bits_wdata_10),
    .io_memStreams_scatters_0_cmd_bits_wdata_11(accel_io_memStreams_scatters_0_cmd_bits_wdata_11),
    .io_memStreams_scatters_0_cmd_bits_wdata_12(accel_io_memStreams_scatters_0_cmd_bits_wdata_12),
    .io_memStreams_scatters_0_cmd_bits_wdata_13(accel_io_memStreams_scatters_0_cmd_bits_wdata_13),
    .io_memStreams_scatters_0_cmd_bits_wdata_14(accel_io_memStreams_scatters_0_cmd_bits_wdata_14),
    .io_memStreams_scatters_0_cmd_bits_wdata_15(accel_io_memStreams_scatters_0_cmd_bits_wdata_15),
    .io_memStreams_scatters_0_cmd_bits_wdata_16(accel_io_memStreams_scatters_0_cmd_bits_wdata_16),
    .io_memStreams_scatters_0_cmd_bits_wdata_17(accel_io_memStreams_scatters_0_cmd_bits_wdata_17),
    .io_memStreams_scatters_0_cmd_bits_wdata_18(accel_io_memStreams_scatters_0_cmd_bits_wdata_18),
    .io_memStreams_scatters_0_cmd_bits_wdata_19(accel_io_memStreams_scatters_0_cmd_bits_wdata_19),
    .io_memStreams_scatters_0_cmd_bits_wdata_20(accel_io_memStreams_scatters_0_cmd_bits_wdata_20),
    .io_memStreams_scatters_0_cmd_bits_wdata_21(accel_io_memStreams_scatters_0_cmd_bits_wdata_21),
    .io_memStreams_scatters_0_cmd_bits_wdata_22(accel_io_memStreams_scatters_0_cmd_bits_wdata_22),
    .io_memStreams_scatters_0_cmd_bits_wdata_23(accel_io_memStreams_scatters_0_cmd_bits_wdata_23),
    .io_memStreams_scatters_0_cmd_bits_wdata_24(accel_io_memStreams_scatters_0_cmd_bits_wdata_24),
    .io_memStreams_scatters_0_cmd_bits_wdata_25(accel_io_memStreams_scatters_0_cmd_bits_wdata_25),
    .io_memStreams_scatters_0_cmd_bits_wdata_26(accel_io_memStreams_scatters_0_cmd_bits_wdata_26),
    .io_memStreams_scatters_0_cmd_bits_wdata_27(accel_io_memStreams_scatters_0_cmd_bits_wdata_27),
    .io_memStreams_scatters_0_cmd_bits_wdata_28(accel_io_memStreams_scatters_0_cmd_bits_wdata_28),
    .io_memStreams_scatters_0_cmd_bits_wdata_29(accel_io_memStreams_scatters_0_cmd_bits_wdata_29),
    .io_memStreams_scatters_0_cmd_bits_wdata_30(accel_io_memStreams_scatters_0_cmd_bits_wdata_30),
    .io_memStreams_scatters_0_cmd_bits_wdata_31(accel_io_memStreams_scatters_0_cmd_bits_wdata_31),
    .io_memStreams_scatters_0_cmd_bits_wdata_32(accel_io_memStreams_scatters_0_cmd_bits_wdata_32),
    .io_memStreams_scatters_0_cmd_bits_wdata_33(accel_io_memStreams_scatters_0_cmd_bits_wdata_33),
    .io_memStreams_scatters_0_cmd_bits_wdata_34(accel_io_memStreams_scatters_0_cmd_bits_wdata_34),
    .io_memStreams_scatters_0_cmd_bits_wdata_35(accel_io_memStreams_scatters_0_cmd_bits_wdata_35),
    .io_memStreams_scatters_0_cmd_bits_wdata_36(accel_io_memStreams_scatters_0_cmd_bits_wdata_36),
    .io_memStreams_scatters_0_cmd_bits_wdata_37(accel_io_memStreams_scatters_0_cmd_bits_wdata_37),
    .io_memStreams_scatters_0_cmd_bits_wdata_38(accel_io_memStreams_scatters_0_cmd_bits_wdata_38),
    .io_memStreams_scatters_0_cmd_bits_wdata_39(accel_io_memStreams_scatters_0_cmd_bits_wdata_39),
    .io_memStreams_scatters_0_cmd_bits_wdata_40(accel_io_memStreams_scatters_0_cmd_bits_wdata_40),
    .io_memStreams_scatters_0_cmd_bits_wdata_41(accel_io_memStreams_scatters_0_cmd_bits_wdata_41),
    .io_memStreams_scatters_0_cmd_bits_wdata_42(accel_io_memStreams_scatters_0_cmd_bits_wdata_42),
    .io_memStreams_scatters_0_cmd_bits_wdata_43(accel_io_memStreams_scatters_0_cmd_bits_wdata_43),
    .io_memStreams_scatters_0_cmd_bits_wdata_44(accel_io_memStreams_scatters_0_cmd_bits_wdata_44),
    .io_memStreams_scatters_0_cmd_bits_wdata_45(accel_io_memStreams_scatters_0_cmd_bits_wdata_45),
    .io_memStreams_scatters_0_cmd_bits_wdata_46(accel_io_memStreams_scatters_0_cmd_bits_wdata_46),
    .io_memStreams_scatters_0_cmd_bits_wdata_47(accel_io_memStreams_scatters_0_cmd_bits_wdata_47),
    .io_memStreams_scatters_0_cmd_bits_wdata_48(accel_io_memStreams_scatters_0_cmd_bits_wdata_48),
    .io_memStreams_scatters_0_cmd_bits_wdata_49(accel_io_memStreams_scatters_0_cmd_bits_wdata_49),
    .io_memStreams_scatters_0_cmd_bits_wdata_50(accel_io_memStreams_scatters_0_cmd_bits_wdata_50),
    .io_memStreams_scatters_0_cmd_bits_wdata_51(accel_io_memStreams_scatters_0_cmd_bits_wdata_51),
    .io_memStreams_scatters_0_cmd_bits_wdata_52(accel_io_memStreams_scatters_0_cmd_bits_wdata_52),
    .io_memStreams_scatters_0_cmd_bits_wdata_53(accel_io_memStreams_scatters_0_cmd_bits_wdata_53),
    .io_memStreams_scatters_0_cmd_bits_wdata_54(accel_io_memStreams_scatters_0_cmd_bits_wdata_54),
    .io_memStreams_scatters_0_cmd_bits_wdata_55(accel_io_memStreams_scatters_0_cmd_bits_wdata_55),
    .io_memStreams_scatters_0_cmd_bits_wdata_56(accel_io_memStreams_scatters_0_cmd_bits_wdata_56),
    .io_memStreams_scatters_0_cmd_bits_wdata_57(accel_io_memStreams_scatters_0_cmd_bits_wdata_57),
    .io_memStreams_scatters_0_cmd_bits_wdata_58(accel_io_memStreams_scatters_0_cmd_bits_wdata_58),
    .io_memStreams_scatters_0_cmd_bits_wdata_59(accel_io_memStreams_scatters_0_cmd_bits_wdata_59),
    .io_memStreams_scatters_0_cmd_bits_wdata_60(accel_io_memStreams_scatters_0_cmd_bits_wdata_60),
    .io_memStreams_scatters_0_cmd_bits_wdata_61(accel_io_memStreams_scatters_0_cmd_bits_wdata_61),
    .io_memStreams_scatters_0_cmd_bits_wdata_62(accel_io_memStreams_scatters_0_cmd_bits_wdata_62),
    .io_memStreams_scatters_0_cmd_bits_wdata_63(accel_io_memStreams_scatters_0_cmd_bits_wdata_63),
    .io_memStreams_scatters_0_wresp_ready(accel_io_memStreams_scatters_0_wresp_ready),
    .io_memStreams_scatters_0_wresp_valid(accel_io_memStreams_scatters_0_wresp_valid),
    .io_memStreams_scatters_0_wresp_bits(accel_io_memStreams_scatters_0_wresp_bits),
    .io_axiStreamsIn_0_TVALID(accel_io_axiStreamsIn_0_TVALID),
    .io_axiStreamsIn_0_TREADY(accel_io_axiStreamsIn_0_TREADY),
    .io_axiStreamsIn_0_TDATA(accel_io_axiStreamsIn_0_TDATA),
    .io_axiStreamsIn_0_TSTRB(accel_io_axiStreamsIn_0_TSTRB),
    .io_axiStreamsIn_0_TKEEP(accel_io_axiStreamsIn_0_TKEEP),
    .io_axiStreamsIn_0_TLAST(accel_io_axiStreamsIn_0_TLAST),
    .io_axiStreamsIn_0_TID(accel_io_axiStreamsIn_0_TID),
    .io_axiStreamsIn_0_TDEST(accel_io_axiStreamsIn_0_TDEST),
    .io_axiStreamsIn_0_TUSER(accel_io_axiStreamsIn_0_TUSER),
    .io_axiStreamsOut_0_TVALID(accel_io_axiStreamsOut_0_TVALID),
    .io_axiStreamsOut_0_TREADY(accel_io_axiStreamsOut_0_TREADY),
    .io_axiStreamsOut_0_TDATA(accel_io_axiStreamsOut_0_TDATA),
    .io_axiStreamsOut_0_TSTRB(accel_io_axiStreamsOut_0_TSTRB),
    .io_axiStreamsOut_0_TKEEP(accel_io_axiStreamsOut_0_TKEEP),
    .io_axiStreamsOut_0_TLAST(accel_io_axiStreamsOut_0_TLAST),
    .io_axiStreamsOut_0_TID(accel_io_axiStreamsOut_0_TID),
    .io_axiStreamsOut_0_TDEST(accel_io_axiStreamsOut_0_TDEST),
    .io_axiStreamsOut_0_TUSER(accel_io_axiStreamsOut_0_TUSER),
    .io_heap_0_req_valid(accel_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(accel_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(accel_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(accel_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(accel_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(accel_io_heap_0_resp_bits_sizeAddr),
    .io_argIns_0(accel_io_argIns_0),
    .io_argOuts_0_port_ready(accel_io_argOuts_0_port_ready),
    .io_argOuts_0_port_valid(accel_io_argOuts_0_port_valid),
    .io_argOuts_0_port_bits(accel_io_argOuts_0_port_bits),
    .io_argOuts_0_echo(accel_io_argOuts_0_echo)
  );
  Fringe Fringe ( // @[SimTarget.scala 16:24:@48290.4]
    .clock(Fringe_clock),
    .reset(Fringe_reset),
    .io_raddr(Fringe_io_raddr),
    .io_wen(Fringe_io_wen),
    .io_waddr(Fringe_io_waddr),
    .io_wdata(Fringe_io_wdata),
    .io_rdata(Fringe_io_rdata),
    .io_enable(Fringe_io_enable),
    .io_done(Fringe_io_done),
    .io_reset(Fringe_io_reset),
    .io_argIns_0(Fringe_io_argIns_0),
    .io_argOuts_0_valid(Fringe_io_argOuts_0_valid),
    .io_argOuts_0_bits(Fringe_io_argOuts_0_bits),
    .io_argEchos_0(Fringe_io_argEchos_0),
    .io_heap_0_req_valid(Fringe_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(Fringe_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(Fringe_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(Fringe_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(Fringe_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(Fringe_io_heap_0_resp_bits_sizeAddr)
  );
  assign io_rdata = Fringe_io_rdata; // @[SimTarget.scala 24:14:@49098.4]
  assign io_dram_0_cmd_valid = 1'h0; // @[SimTarget.scala 27:13:@49305.4]
  assign io_dram_0_cmd_bits_addr = 64'h0; // @[SimTarget.scala 27:13:@49304.4]
  assign io_dram_0_cmd_bits_size = 32'h0; // @[SimTarget.scala 27:13:@49303.4]
  assign io_dram_0_cmd_bits_rawAddr = 64'h0; // @[SimTarget.scala 27:13:@49302.4]
  assign io_dram_0_cmd_bits_isWr = 1'h0; // @[SimTarget.scala 27:13:@49301.4]
  assign io_dram_0_cmd_bits_tag = 32'h0; // @[SimTarget.scala 27:13:@49300.4]
  assign io_dram_0_wdata_valid = 1'h0; // @[SimTarget.scala 27:13:@49298.4]
  assign io_dram_0_wdata_bits_wdata_0 = 8'h0; // @[SimTarget.scala 27:13:@49234.4]
  assign io_dram_0_wdata_bits_wdata_1 = 8'h0; // @[SimTarget.scala 27:13:@49235.4]
  assign io_dram_0_wdata_bits_wdata_2 = 8'h0; // @[SimTarget.scala 27:13:@49236.4]
  assign io_dram_0_wdata_bits_wdata_3 = 8'h0; // @[SimTarget.scala 27:13:@49237.4]
  assign io_dram_0_wdata_bits_wdata_4 = 8'h0; // @[SimTarget.scala 27:13:@49238.4]
  assign io_dram_0_wdata_bits_wdata_5 = 8'h0; // @[SimTarget.scala 27:13:@49239.4]
  assign io_dram_0_wdata_bits_wdata_6 = 8'h0; // @[SimTarget.scala 27:13:@49240.4]
  assign io_dram_0_wdata_bits_wdata_7 = 8'h0; // @[SimTarget.scala 27:13:@49241.4]
  assign io_dram_0_wdata_bits_wdata_8 = 8'h0; // @[SimTarget.scala 27:13:@49242.4]
  assign io_dram_0_wdata_bits_wdata_9 = 8'h0; // @[SimTarget.scala 27:13:@49243.4]
  assign io_dram_0_wdata_bits_wdata_10 = 8'h0; // @[SimTarget.scala 27:13:@49244.4]
  assign io_dram_0_wdata_bits_wdata_11 = 8'h0; // @[SimTarget.scala 27:13:@49245.4]
  assign io_dram_0_wdata_bits_wdata_12 = 8'h0; // @[SimTarget.scala 27:13:@49246.4]
  assign io_dram_0_wdata_bits_wdata_13 = 8'h0; // @[SimTarget.scala 27:13:@49247.4]
  assign io_dram_0_wdata_bits_wdata_14 = 8'h0; // @[SimTarget.scala 27:13:@49248.4]
  assign io_dram_0_wdata_bits_wdata_15 = 8'h0; // @[SimTarget.scala 27:13:@49249.4]
  assign io_dram_0_wdata_bits_wdata_16 = 8'h0; // @[SimTarget.scala 27:13:@49250.4]
  assign io_dram_0_wdata_bits_wdata_17 = 8'h0; // @[SimTarget.scala 27:13:@49251.4]
  assign io_dram_0_wdata_bits_wdata_18 = 8'h0; // @[SimTarget.scala 27:13:@49252.4]
  assign io_dram_0_wdata_bits_wdata_19 = 8'h0; // @[SimTarget.scala 27:13:@49253.4]
  assign io_dram_0_wdata_bits_wdata_20 = 8'h0; // @[SimTarget.scala 27:13:@49254.4]
  assign io_dram_0_wdata_bits_wdata_21 = 8'h0; // @[SimTarget.scala 27:13:@49255.4]
  assign io_dram_0_wdata_bits_wdata_22 = 8'h0; // @[SimTarget.scala 27:13:@49256.4]
  assign io_dram_0_wdata_bits_wdata_23 = 8'h0; // @[SimTarget.scala 27:13:@49257.4]
  assign io_dram_0_wdata_bits_wdata_24 = 8'h0; // @[SimTarget.scala 27:13:@49258.4]
  assign io_dram_0_wdata_bits_wdata_25 = 8'h0; // @[SimTarget.scala 27:13:@49259.4]
  assign io_dram_0_wdata_bits_wdata_26 = 8'h0; // @[SimTarget.scala 27:13:@49260.4]
  assign io_dram_0_wdata_bits_wdata_27 = 8'h0; // @[SimTarget.scala 27:13:@49261.4]
  assign io_dram_0_wdata_bits_wdata_28 = 8'h0; // @[SimTarget.scala 27:13:@49262.4]
  assign io_dram_0_wdata_bits_wdata_29 = 8'h0; // @[SimTarget.scala 27:13:@49263.4]
  assign io_dram_0_wdata_bits_wdata_30 = 8'h0; // @[SimTarget.scala 27:13:@49264.4]
  assign io_dram_0_wdata_bits_wdata_31 = 8'h0; // @[SimTarget.scala 27:13:@49265.4]
  assign io_dram_0_wdata_bits_wdata_32 = 8'h0; // @[SimTarget.scala 27:13:@49266.4]
  assign io_dram_0_wdata_bits_wdata_33 = 8'h0; // @[SimTarget.scala 27:13:@49267.4]
  assign io_dram_0_wdata_bits_wdata_34 = 8'h0; // @[SimTarget.scala 27:13:@49268.4]
  assign io_dram_0_wdata_bits_wdata_35 = 8'h0; // @[SimTarget.scala 27:13:@49269.4]
  assign io_dram_0_wdata_bits_wdata_36 = 8'h0; // @[SimTarget.scala 27:13:@49270.4]
  assign io_dram_0_wdata_bits_wdata_37 = 8'h0; // @[SimTarget.scala 27:13:@49271.4]
  assign io_dram_0_wdata_bits_wdata_38 = 8'h0; // @[SimTarget.scala 27:13:@49272.4]
  assign io_dram_0_wdata_bits_wdata_39 = 8'h0; // @[SimTarget.scala 27:13:@49273.4]
  assign io_dram_0_wdata_bits_wdata_40 = 8'h0; // @[SimTarget.scala 27:13:@49274.4]
  assign io_dram_0_wdata_bits_wdata_41 = 8'h0; // @[SimTarget.scala 27:13:@49275.4]
  assign io_dram_0_wdata_bits_wdata_42 = 8'h0; // @[SimTarget.scala 27:13:@49276.4]
  assign io_dram_0_wdata_bits_wdata_43 = 8'h0; // @[SimTarget.scala 27:13:@49277.4]
  assign io_dram_0_wdata_bits_wdata_44 = 8'h0; // @[SimTarget.scala 27:13:@49278.4]
  assign io_dram_0_wdata_bits_wdata_45 = 8'h0; // @[SimTarget.scala 27:13:@49279.4]
  assign io_dram_0_wdata_bits_wdata_46 = 8'h0; // @[SimTarget.scala 27:13:@49280.4]
  assign io_dram_0_wdata_bits_wdata_47 = 8'h0; // @[SimTarget.scala 27:13:@49281.4]
  assign io_dram_0_wdata_bits_wdata_48 = 8'h0; // @[SimTarget.scala 27:13:@49282.4]
  assign io_dram_0_wdata_bits_wdata_49 = 8'h0; // @[SimTarget.scala 27:13:@49283.4]
  assign io_dram_0_wdata_bits_wdata_50 = 8'h0; // @[SimTarget.scala 27:13:@49284.4]
  assign io_dram_0_wdata_bits_wdata_51 = 8'h0; // @[SimTarget.scala 27:13:@49285.4]
  assign io_dram_0_wdata_bits_wdata_52 = 8'h0; // @[SimTarget.scala 27:13:@49286.4]
  assign io_dram_0_wdata_bits_wdata_53 = 8'h0; // @[SimTarget.scala 27:13:@49287.4]
  assign io_dram_0_wdata_bits_wdata_54 = 8'h0; // @[SimTarget.scala 27:13:@49288.4]
  assign io_dram_0_wdata_bits_wdata_55 = 8'h0; // @[SimTarget.scala 27:13:@49289.4]
  assign io_dram_0_wdata_bits_wdata_56 = 8'h0; // @[SimTarget.scala 27:13:@49290.4]
  assign io_dram_0_wdata_bits_wdata_57 = 8'h0; // @[SimTarget.scala 27:13:@49291.4]
  assign io_dram_0_wdata_bits_wdata_58 = 8'h0; // @[SimTarget.scala 27:13:@49292.4]
  assign io_dram_0_wdata_bits_wdata_59 = 8'h0; // @[SimTarget.scala 27:13:@49293.4]
  assign io_dram_0_wdata_bits_wdata_60 = 8'h0; // @[SimTarget.scala 27:13:@49294.4]
  assign io_dram_0_wdata_bits_wdata_61 = 8'h0; // @[SimTarget.scala 27:13:@49295.4]
  assign io_dram_0_wdata_bits_wdata_62 = 8'h0; // @[SimTarget.scala 27:13:@49296.4]
  assign io_dram_0_wdata_bits_wdata_63 = 8'h0; // @[SimTarget.scala 27:13:@49297.4]
  assign io_dram_0_wdata_bits_wstrb_0 = 1'h0; // @[SimTarget.scala 27:13:@49170.4]
  assign io_dram_0_wdata_bits_wstrb_1 = 1'h0; // @[SimTarget.scala 27:13:@49171.4]
  assign io_dram_0_wdata_bits_wstrb_2 = 1'h0; // @[SimTarget.scala 27:13:@49172.4]
  assign io_dram_0_wdata_bits_wstrb_3 = 1'h0; // @[SimTarget.scala 27:13:@49173.4]
  assign io_dram_0_wdata_bits_wstrb_4 = 1'h0; // @[SimTarget.scala 27:13:@49174.4]
  assign io_dram_0_wdata_bits_wstrb_5 = 1'h0; // @[SimTarget.scala 27:13:@49175.4]
  assign io_dram_0_wdata_bits_wstrb_6 = 1'h0; // @[SimTarget.scala 27:13:@49176.4]
  assign io_dram_0_wdata_bits_wstrb_7 = 1'h0; // @[SimTarget.scala 27:13:@49177.4]
  assign io_dram_0_wdata_bits_wstrb_8 = 1'h0; // @[SimTarget.scala 27:13:@49178.4]
  assign io_dram_0_wdata_bits_wstrb_9 = 1'h0; // @[SimTarget.scala 27:13:@49179.4]
  assign io_dram_0_wdata_bits_wstrb_10 = 1'h0; // @[SimTarget.scala 27:13:@49180.4]
  assign io_dram_0_wdata_bits_wstrb_11 = 1'h0; // @[SimTarget.scala 27:13:@49181.4]
  assign io_dram_0_wdata_bits_wstrb_12 = 1'h0; // @[SimTarget.scala 27:13:@49182.4]
  assign io_dram_0_wdata_bits_wstrb_13 = 1'h0; // @[SimTarget.scala 27:13:@49183.4]
  assign io_dram_0_wdata_bits_wstrb_14 = 1'h0; // @[SimTarget.scala 27:13:@49184.4]
  assign io_dram_0_wdata_bits_wstrb_15 = 1'h0; // @[SimTarget.scala 27:13:@49185.4]
  assign io_dram_0_wdata_bits_wstrb_16 = 1'h0; // @[SimTarget.scala 27:13:@49186.4]
  assign io_dram_0_wdata_bits_wstrb_17 = 1'h0; // @[SimTarget.scala 27:13:@49187.4]
  assign io_dram_0_wdata_bits_wstrb_18 = 1'h0; // @[SimTarget.scala 27:13:@49188.4]
  assign io_dram_0_wdata_bits_wstrb_19 = 1'h0; // @[SimTarget.scala 27:13:@49189.4]
  assign io_dram_0_wdata_bits_wstrb_20 = 1'h0; // @[SimTarget.scala 27:13:@49190.4]
  assign io_dram_0_wdata_bits_wstrb_21 = 1'h0; // @[SimTarget.scala 27:13:@49191.4]
  assign io_dram_0_wdata_bits_wstrb_22 = 1'h0; // @[SimTarget.scala 27:13:@49192.4]
  assign io_dram_0_wdata_bits_wstrb_23 = 1'h0; // @[SimTarget.scala 27:13:@49193.4]
  assign io_dram_0_wdata_bits_wstrb_24 = 1'h0; // @[SimTarget.scala 27:13:@49194.4]
  assign io_dram_0_wdata_bits_wstrb_25 = 1'h0; // @[SimTarget.scala 27:13:@49195.4]
  assign io_dram_0_wdata_bits_wstrb_26 = 1'h0; // @[SimTarget.scala 27:13:@49196.4]
  assign io_dram_0_wdata_bits_wstrb_27 = 1'h0; // @[SimTarget.scala 27:13:@49197.4]
  assign io_dram_0_wdata_bits_wstrb_28 = 1'h0; // @[SimTarget.scala 27:13:@49198.4]
  assign io_dram_0_wdata_bits_wstrb_29 = 1'h0; // @[SimTarget.scala 27:13:@49199.4]
  assign io_dram_0_wdata_bits_wstrb_30 = 1'h0; // @[SimTarget.scala 27:13:@49200.4]
  assign io_dram_0_wdata_bits_wstrb_31 = 1'h0; // @[SimTarget.scala 27:13:@49201.4]
  assign io_dram_0_wdata_bits_wstrb_32 = 1'h0; // @[SimTarget.scala 27:13:@49202.4]
  assign io_dram_0_wdata_bits_wstrb_33 = 1'h0; // @[SimTarget.scala 27:13:@49203.4]
  assign io_dram_0_wdata_bits_wstrb_34 = 1'h0; // @[SimTarget.scala 27:13:@49204.4]
  assign io_dram_0_wdata_bits_wstrb_35 = 1'h0; // @[SimTarget.scala 27:13:@49205.4]
  assign io_dram_0_wdata_bits_wstrb_36 = 1'h0; // @[SimTarget.scala 27:13:@49206.4]
  assign io_dram_0_wdata_bits_wstrb_37 = 1'h0; // @[SimTarget.scala 27:13:@49207.4]
  assign io_dram_0_wdata_bits_wstrb_38 = 1'h0; // @[SimTarget.scala 27:13:@49208.4]
  assign io_dram_0_wdata_bits_wstrb_39 = 1'h0; // @[SimTarget.scala 27:13:@49209.4]
  assign io_dram_0_wdata_bits_wstrb_40 = 1'h0; // @[SimTarget.scala 27:13:@49210.4]
  assign io_dram_0_wdata_bits_wstrb_41 = 1'h0; // @[SimTarget.scala 27:13:@49211.4]
  assign io_dram_0_wdata_bits_wstrb_42 = 1'h0; // @[SimTarget.scala 27:13:@49212.4]
  assign io_dram_0_wdata_bits_wstrb_43 = 1'h0; // @[SimTarget.scala 27:13:@49213.4]
  assign io_dram_0_wdata_bits_wstrb_44 = 1'h0; // @[SimTarget.scala 27:13:@49214.4]
  assign io_dram_0_wdata_bits_wstrb_45 = 1'h0; // @[SimTarget.scala 27:13:@49215.4]
  assign io_dram_0_wdata_bits_wstrb_46 = 1'h0; // @[SimTarget.scala 27:13:@49216.4]
  assign io_dram_0_wdata_bits_wstrb_47 = 1'h0; // @[SimTarget.scala 27:13:@49217.4]
  assign io_dram_0_wdata_bits_wstrb_48 = 1'h0; // @[SimTarget.scala 27:13:@49218.4]
  assign io_dram_0_wdata_bits_wstrb_49 = 1'h0; // @[SimTarget.scala 27:13:@49219.4]
  assign io_dram_0_wdata_bits_wstrb_50 = 1'h0; // @[SimTarget.scala 27:13:@49220.4]
  assign io_dram_0_wdata_bits_wstrb_51 = 1'h0; // @[SimTarget.scala 27:13:@49221.4]
  assign io_dram_0_wdata_bits_wstrb_52 = 1'h0; // @[SimTarget.scala 27:13:@49222.4]
  assign io_dram_0_wdata_bits_wstrb_53 = 1'h0; // @[SimTarget.scala 27:13:@49223.4]
  assign io_dram_0_wdata_bits_wstrb_54 = 1'h0; // @[SimTarget.scala 27:13:@49224.4]
  assign io_dram_0_wdata_bits_wstrb_55 = 1'h0; // @[SimTarget.scala 27:13:@49225.4]
  assign io_dram_0_wdata_bits_wstrb_56 = 1'h0; // @[SimTarget.scala 27:13:@49226.4]
  assign io_dram_0_wdata_bits_wstrb_57 = 1'h0; // @[SimTarget.scala 27:13:@49227.4]
  assign io_dram_0_wdata_bits_wstrb_58 = 1'h0; // @[SimTarget.scala 27:13:@49228.4]
  assign io_dram_0_wdata_bits_wstrb_59 = 1'h0; // @[SimTarget.scala 27:13:@49229.4]
  assign io_dram_0_wdata_bits_wstrb_60 = 1'h0; // @[SimTarget.scala 27:13:@49230.4]
  assign io_dram_0_wdata_bits_wstrb_61 = 1'h0; // @[SimTarget.scala 27:13:@49231.4]
  assign io_dram_0_wdata_bits_wstrb_62 = 1'h0; // @[SimTarget.scala 27:13:@49232.4]
  assign io_dram_0_wdata_bits_wstrb_63 = 1'h0; // @[SimTarget.scala 27:13:@49233.4]
  assign io_dram_0_wdata_bits_wlast = 1'h0; // @[SimTarget.scala 27:13:@49169.4]
  assign io_dram_0_rresp_ready = 1'h0; // @[SimTarget.scala 27:13:@49168.4]
  assign io_dram_0_wresp_ready = 1'h0; // @[SimTarget.scala 27:13:@49101.4]
  assign accel_clock = clock; // @[:@47847.4]
  assign accel_reset = reset; // @[:@47848.4]
  assign accel_io_enable = Fringe_io_enable; // @[SimTarget.scala 45:21:@49727.4]
  assign accel_io_reset = Fringe_io_reset; // @[SimTarget.scala 47:20:@49729.4]
  assign accel_io_memStreams_loads_0_cmd_ready = 1'h0; // @[SimTarget.scala 43:26:@49720.4]
  assign accel_io_memStreams_loads_0_data_valid = 1'h0; // @[SimTarget.scala 43:26:@49715.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_0 = 8'h0; // @[SimTarget.scala 43:26:@49651.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_1 = 8'h0; // @[SimTarget.scala 43:26:@49652.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_2 = 8'h0; // @[SimTarget.scala 43:26:@49653.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_3 = 8'h0; // @[SimTarget.scala 43:26:@49654.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_4 = 8'h0; // @[SimTarget.scala 43:26:@49655.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_5 = 8'h0; // @[SimTarget.scala 43:26:@49656.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_6 = 8'h0; // @[SimTarget.scala 43:26:@49657.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_7 = 8'h0; // @[SimTarget.scala 43:26:@49658.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_8 = 8'h0; // @[SimTarget.scala 43:26:@49659.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_9 = 8'h0; // @[SimTarget.scala 43:26:@49660.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_10 = 8'h0; // @[SimTarget.scala 43:26:@49661.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_11 = 8'h0; // @[SimTarget.scala 43:26:@49662.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_12 = 8'h0; // @[SimTarget.scala 43:26:@49663.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_13 = 8'h0; // @[SimTarget.scala 43:26:@49664.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_14 = 8'h0; // @[SimTarget.scala 43:26:@49665.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_15 = 8'h0; // @[SimTarget.scala 43:26:@49666.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_16 = 8'h0; // @[SimTarget.scala 43:26:@49667.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_17 = 8'h0; // @[SimTarget.scala 43:26:@49668.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_18 = 8'h0; // @[SimTarget.scala 43:26:@49669.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_19 = 8'h0; // @[SimTarget.scala 43:26:@49670.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_20 = 8'h0; // @[SimTarget.scala 43:26:@49671.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_21 = 8'h0; // @[SimTarget.scala 43:26:@49672.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_22 = 8'h0; // @[SimTarget.scala 43:26:@49673.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_23 = 8'h0; // @[SimTarget.scala 43:26:@49674.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_24 = 8'h0; // @[SimTarget.scala 43:26:@49675.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_25 = 8'h0; // @[SimTarget.scala 43:26:@49676.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_26 = 8'h0; // @[SimTarget.scala 43:26:@49677.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_27 = 8'h0; // @[SimTarget.scala 43:26:@49678.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_28 = 8'h0; // @[SimTarget.scala 43:26:@49679.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_29 = 8'h0; // @[SimTarget.scala 43:26:@49680.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_30 = 8'h0; // @[SimTarget.scala 43:26:@49681.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_31 = 8'h0; // @[SimTarget.scala 43:26:@49682.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_32 = 8'h0; // @[SimTarget.scala 43:26:@49683.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_33 = 8'h0; // @[SimTarget.scala 43:26:@49684.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_34 = 8'h0; // @[SimTarget.scala 43:26:@49685.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_35 = 8'h0; // @[SimTarget.scala 43:26:@49686.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_36 = 8'h0; // @[SimTarget.scala 43:26:@49687.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_37 = 8'h0; // @[SimTarget.scala 43:26:@49688.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_38 = 8'h0; // @[SimTarget.scala 43:26:@49689.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_39 = 8'h0; // @[SimTarget.scala 43:26:@49690.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_40 = 8'h0; // @[SimTarget.scala 43:26:@49691.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_41 = 8'h0; // @[SimTarget.scala 43:26:@49692.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_42 = 8'h0; // @[SimTarget.scala 43:26:@49693.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_43 = 8'h0; // @[SimTarget.scala 43:26:@49694.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_44 = 8'h0; // @[SimTarget.scala 43:26:@49695.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_45 = 8'h0; // @[SimTarget.scala 43:26:@49696.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_46 = 8'h0; // @[SimTarget.scala 43:26:@49697.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_47 = 8'h0; // @[SimTarget.scala 43:26:@49698.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_48 = 8'h0; // @[SimTarget.scala 43:26:@49699.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_49 = 8'h0; // @[SimTarget.scala 43:26:@49700.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_50 = 8'h0; // @[SimTarget.scala 43:26:@49701.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_51 = 8'h0; // @[SimTarget.scala 43:26:@49702.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_52 = 8'h0; // @[SimTarget.scala 43:26:@49703.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_53 = 8'h0; // @[SimTarget.scala 43:26:@49704.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_54 = 8'h0; // @[SimTarget.scala 43:26:@49705.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_55 = 8'h0; // @[SimTarget.scala 43:26:@49706.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_56 = 8'h0; // @[SimTarget.scala 43:26:@49707.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_57 = 8'h0; // @[SimTarget.scala 43:26:@49708.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_58 = 8'h0; // @[SimTarget.scala 43:26:@49709.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_59 = 8'h0; // @[SimTarget.scala 43:26:@49710.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_60 = 8'h0; // @[SimTarget.scala 43:26:@49711.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_61 = 8'h0; // @[SimTarget.scala 43:26:@49712.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_62 = 8'h0; // @[SimTarget.scala 43:26:@49713.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_63 = 8'h0; // @[SimTarget.scala 43:26:@49714.4]
  assign accel_io_memStreams_stores_0_cmd_ready = 1'h0; // @[SimTarget.scala 43:26:@49650.4]
  assign accel_io_memStreams_stores_0_data_ready = 1'h0; // @[SimTarget.scala 43:26:@49646.4]
  assign accel_io_memStreams_stores_0_wresp_valid = 1'h0; // @[SimTarget.scala 43:26:@49578.4]
  assign accel_io_memStreams_stores_0_wresp_bits = 1'h0; // @[SimTarget.scala 43:26:@49577.4]
  assign accel_io_memStreams_gathers_0_cmd_ready = 1'h0; // @[SimTarget.scala 43:26:@49576.4]
  assign accel_io_memStreams_gathers_0_data_valid = 1'h0; // @[SimTarget.scala 43:26:@49509.4]
  assign accel_io_memStreams_gathers_0_data_bits_0 = 8'h0; // @[SimTarget.scala 43:26:@49445.4]
  assign accel_io_memStreams_gathers_0_data_bits_1 = 8'h0; // @[SimTarget.scala 43:26:@49446.4]
  assign accel_io_memStreams_gathers_0_data_bits_2 = 8'h0; // @[SimTarget.scala 43:26:@49447.4]
  assign accel_io_memStreams_gathers_0_data_bits_3 = 8'h0; // @[SimTarget.scala 43:26:@49448.4]
  assign accel_io_memStreams_gathers_0_data_bits_4 = 8'h0; // @[SimTarget.scala 43:26:@49449.4]
  assign accel_io_memStreams_gathers_0_data_bits_5 = 8'h0; // @[SimTarget.scala 43:26:@49450.4]
  assign accel_io_memStreams_gathers_0_data_bits_6 = 8'h0; // @[SimTarget.scala 43:26:@49451.4]
  assign accel_io_memStreams_gathers_0_data_bits_7 = 8'h0; // @[SimTarget.scala 43:26:@49452.4]
  assign accel_io_memStreams_gathers_0_data_bits_8 = 8'h0; // @[SimTarget.scala 43:26:@49453.4]
  assign accel_io_memStreams_gathers_0_data_bits_9 = 8'h0; // @[SimTarget.scala 43:26:@49454.4]
  assign accel_io_memStreams_gathers_0_data_bits_10 = 8'h0; // @[SimTarget.scala 43:26:@49455.4]
  assign accel_io_memStreams_gathers_0_data_bits_11 = 8'h0; // @[SimTarget.scala 43:26:@49456.4]
  assign accel_io_memStreams_gathers_0_data_bits_12 = 8'h0; // @[SimTarget.scala 43:26:@49457.4]
  assign accel_io_memStreams_gathers_0_data_bits_13 = 8'h0; // @[SimTarget.scala 43:26:@49458.4]
  assign accel_io_memStreams_gathers_0_data_bits_14 = 8'h0; // @[SimTarget.scala 43:26:@49459.4]
  assign accel_io_memStreams_gathers_0_data_bits_15 = 8'h0; // @[SimTarget.scala 43:26:@49460.4]
  assign accel_io_memStreams_gathers_0_data_bits_16 = 8'h0; // @[SimTarget.scala 43:26:@49461.4]
  assign accel_io_memStreams_gathers_0_data_bits_17 = 8'h0; // @[SimTarget.scala 43:26:@49462.4]
  assign accel_io_memStreams_gathers_0_data_bits_18 = 8'h0; // @[SimTarget.scala 43:26:@49463.4]
  assign accel_io_memStreams_gathers_0_data_bits_19 = 8'h0; // @[SimTarget.scala 43:26:@49464.4]
  assign accel_io_memStreams_gathers_0_data_bits_20 = 8'h0; // @[SimTarget.scala 43:26:@49465.4]
  assign accel_io_memStreams_gathers_0_data_bits_21 = 8'h0; // @[SimTarget.scala 43:26:@49466.4]
  assign accel_io_memStreams_gathers_0_data_bits_22 = 8'h0; // @[SimTarget.scala 43:26:@49467.4]
  assign accel_io_memStreams_gathers_0_data_bits_23 = 8'h0; // @[SimTarget.scala 43:26:@49468.4]
  assign accel_io_memStreams_gathers_0_data_bits_24 = 8'h0; // @[SimTarget.scala 43:26:@49469.4]
  assign accel_io_memStreams_gathers_0_data_bits_25 = 8'h0; // @[SimTarget.scala 43:26:@49470.4]
  assign accel_io_memStreams_gathers_0_data_bits_26 = 8'h0; // @[SimTarget.scala 43:26:@49471.4]
  assign accel_io_memStreams_gathers_0_data_bits_27 = 8'h0; // @[SimTarget.scala 43:26:@49472.4]
  assign accel_io_memStreams_gathers_0_data_bits_28 = 8'h0; // @[SimTarget.scala 43:26:@49473.4]
  assign accel_io_memStreams_gathers_0_data_bits_29 = 8'h0; // @[SimTarget.scala 43:26:@49474.4]
  assign accel_io_memStreams_gathers_0_data_bits_30 = 8'h0; // @[SimTarget.scala 43:26:@49475.4]
  assign accel_io_memStreams_gathers_0_data_bits_31 = 8'h0; // @[SimTarget.scala 43:26:@49476.4]
  assign accel_io_memStreams_gathers_0_data_bits_32 = 8'h0; // @[SimTarget.scala 43:26:@49477.4]
  assign accel_io_memStreams_gathers_0_data_bits_33 = 8'h0; // @[SimTarget.scala 43:26:@49478.4]
  assign accel_io_memStreams_gathers_0_data_bits_34 = 8'h0; // @[SimTarget.scala 43:26:@49479.4]
  assign accel_io_memStreams_gathers_0_data_bits_35 = 8'h0; // @[SimTarget.scala 43:26:@49480.4]
  assign accel_io_memStreams_gathers_0_data_bits_36 = 8'h0; // @[SimTarget.scala 43:26:@49481.4]
  assign accel_io_memStreams_gathers_0_data_bits_37 = 8'h0; // @[SimTarget.scala 43:26:@49482.4]
  assign accel_io_memStreams_gathers_0_data_bits_38 = 8'h0; // @[SimTarget.scala 43:26:@49483.4]
  assign accel_io_memStreams_gathers_0_data_bits_39 = 8'h0; // @[SimTarget.scala 43:26:@49484.4]
  assign accel_io_memStreams_gathers_0_data_bits_40 = 8'h0; // @[SimTarget.scala 43:26:@49485.4]
  assign accel_io_memStreams_gathers_0_data_bits_41 = 8'h0; // @[SimTarget.scala 43:26:@49486.4]
  assign accel_io_memStreams_gathers_0_data_bits_42 = 8'h0; // @[SimTarget.scala 43:26:@49487.4]
  assign accel_io_memStreams_gathers_0_data_bits_43 = 8'h0; // @[SimTarget.scala 43:26:@49488.4]
  assign accel_io_memStreams_gathers_0_data_bits_44 = 8'h0; // @[SimTarget.scala 43:26:@49489.4]
  assign accel_io_memStreams_gathers_0_data_bits_45 = 8'h0; // @[SimTarget.scala 43:26:@49490.4]
  assign accel_io_memStreams_gathers_0_data_bits_46 = 8'h0; // @[SimTarget.scala 43:26:@49491.4]
  assign accel_io_memStreams_gathers_0_data_bits_47 = 8'h0; // @[SimTarget.scala 43:26:@49492.4]
  assign accel_io_memStreams_gathers_0_data_bits_48 = 8'h0; // @[SimTarget.scala 43:26:@49493.4]
  assign accel_io_memStreams_gathers_0_data_bits_49 = 8'h0; // @[SimTarget.scala 43:26:@49494.4]
  assign accel_io_memStreams_gathers_0_data_bits_50 = 8'h0; // @[SimTarget.scala 43:26:@49495.4]
  assign accel_io_memStreams_gathers_0_data_bits_51 = 8'h0; // @[SimTarget.scala 43:26:@49496.4]
  assign accel_io_memStreams_gathers_0_data_bits_52 = 8'h0; // @[SimTarget.scala 43:26:@49497.4]
  assign accel_io_memStreams_gathers_0_data_bits_53 = 8'h0; // @[SimTarget.scala 43:26:@49498.4]
  assign accel_io_memStreams_gathers_0_data_bits_54 = 8'h0; // @[SimTarget.scala 43:26:@49499.4]
  assign accel_io_memStreams_gathers_0_data_bits_55 = 8'h0; // @[SimTarget.scala 43:26:@49500.4]
  assign accel_io_memStreams_gathers_0_data_bits_56 = 8'h0; // @[SimTarget.scala 43:26:@49501.4]
  assign accel_io_memStreams_gathers_0_data_bits_57 = 8'h0; // @[SimTarget.scala 43:26:@49502.4]
  assign accel_io_memStreams_gathers_0_data_bits_58 = 8'h0; // @[SimTarget.scala 43:26:@49503.4]
  assign accel_io_memStreams_gathers_0_data_bits_59 = 8'h0; // @[SimTarget.scala 43:26:@49504.4]
  assign accel_io_memStreams_gathers_0_data_bits_60 = 8'h0; // @[SimTarget.scala 43:26:@49505.4]
  assign accel_io_memStreams_gathers_0_data_bits_61 = 8'h0; // @[SimTarget.scala 43:26:@49506.4]
  assign accel_io_memStreams_gathers_0_data_bits_62 = 8'h0; // @[SimTarget.scala 43:26:@49507.4]
  assign accel_io_memStreams_gathers_0_data_bits_63 = 8'h0; // @[SimTarget.scala 43:26:@49508.4]
  assign accel_io_memStreams_scatters_0_cmd_ready = 1'h0; // @[SimTarget.scala 43:26:@49444.4]
  assign accel_io_memStreams_scatters_0_wresp_valid = 1'h0; // @[SimTarget.scala 43:26:@49313.4]
  assign accel_io_memStreams_scatters_0_wresp_bits = 1'h0; // @[SimTarget.scala 43:26:@49312.4]
  assign accel_io_axiStreamsIn_0_TVALID = 1'h0;
  assign accel_io_axiStreamsIn_0_TDATA = 256'h0;
  assign accel_io_axiStreamsIn_0_TSTRB = 32'h0;
  assign accel_io_axiStreamsIn_0_TKEEP = 32'h0;
  assign accel_io_axiStreamsIn_0_TLAST = 1'h0;
  assign accel_io_axiStreamsIn_0_TID = 8'h0;
  assign accel_io_axiStreamsIn_0_TDEST = 8'h0;
  assign accel_io_axiStreamsIn_0_TUSER = 32'h0;
  assign accel_io_axiStreamsOut_0_TREADY = 1'h0;
  assign accel_io_heap_0_resp_valid = Fringe_io_heap_0_resp_valid; // @[SimTarget.scala 44:20:@49723.4]
  assign accel_io_heap_0_resp_bits_allocDealloc = Fringe_io_heap_0_resp_bits_allocDealloc; // @[SimTarget.scala 44:20:@49722.4]
  assign accel_io_heap_0_resp_bits_sizeAddr = Fringe_io_heap_0_resp_bits_sizeAddr; // @[SimTarget.scala 44:20:@49721.4]
  assign accel_io_argIns_0 = Fringe_io_argIns_0; // @[SimTarget.scala 30:23:@49307.4]
  assign accel_io_argOuts_0_port_ready = 1'h1; // @[SimTarget.scala 37:32:@49310.4]
  assign accel_io_argOuts_0_echo = Fringe_io_argEchos_0; // @[SimTarget.scala 40:26:@49311.4]
  assign Fringe_clock = clock; // @[:@48291.4]
  assign Fringe_reset = reset; // @[:@48292.4]
  assign Fringe_io_raddr = io_raddr; // @[SimTarget.scala 20:21:@49094.4]
  assign Fringe_io_wen = io_wen; // @[SimTarget.scala 21:21:@49095.4]
  assign Fringe_io_waddr = io_waddr; // @[SimTarget.scala 22:21:@49096.4]
  assign Fringe_io_wdata = io_wdata; // @[SimTarget.scala 23:21:@49097.4]
  assign Fringe_io_done = accel_io_done; // @[SimTarget.scala 46:20:@49728.4]
  assign Fringe_io_argOuts_0_valid = accel_io_argOuts_0_port_valid; // @[SimTarget.scala 36:28:@49309.4]
  assign Fringe_io_argOuts_0_bits = accel_io_argOuts_0_port_bits; // @[SimTarget.scala 35:27:@49308.4]
  assign Fringe_io_heap_0_req_valid = accel_io_heap_0_req_valid; // @[SimTarget.scala 44:20:@49726.4]
  assign Fringe_io_heap_0_req_bits_allocDealloc = accel_io_heap_0_req_bits_allocDealloc; // @[SimTarget.scala 44:20:@49725.4]
  assign Fringe_io_heap_0_req_bits_sizeAddr = accel_io_heap_0_req_bits_sizeAddr; // @[SimTarget.scala 44:20:@49724.4]
endmodule
