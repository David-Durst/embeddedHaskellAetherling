// Latency = 4
module Top(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  input  [7:0] I_2,
  input  [7:0] I_3,
  output [7:0] O_0_0_0,
  output [7:0] O_1_0_0,
  output [7:0] O_2_0_0,
  output [7:0] O_3_0_0
);
  wire dontcare;
  wire [31:0] io_output_counts_1;
  wire [31:0] io_output_counts_0;

  x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1 sampler_box ( // @[m_x55_ctr_0.scala 26:17:@1721.4]
    .clock(clock), // @[:@1296.4]
    .reset('b0), // @[:@1297.4]
    .io_in_x316_TREADY(dontcare), // @[:@1298.4]
    .io_in_x316_TDATA({I_0,I_1,I_2,I_3}), // @[:@1298.4]
    .io_in_x316_TID(8'h0),
    .io_in_x316_TDEST(8'h0),
    .io_in_x317_TVALID(valid_down), // @[:@1298.4]
    .io_in_x317_TDATA({O_0_0_0,O_1_0_0,O_2_0_0,O_3_0_0}), // @[:@1298.4]
    .io_in_x317_TREADY(1'b1), // @[:@1298.4]
    .io_sigsIn_datapathEn(valid_up), // @[:@1298.4]
    .io_sigsIn_backpressure(1'b1), // @[:@20563.4]
    .io_sigsIn_break(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_1(io_output_counts_1), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_0(io_output_counts_0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_0(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_1(1'b0), // @[:@20563.4]
    .io_rr('b1) // @[:@1298.4]
  );

  wire dontcare2;

  wire io_output_oobs_0;
  wire io_output_oobs_1;
  x324_ctrchain cchain ( // @[:@2879.2]
    .clock(clock), // @[:@2880.4]
    .reset(1'b0), // @[:@2881.4]
    .io_input_reset(1'b0), // @[:@2882.4]
    .io_input_enable(valid_up), // @[:@2882.4]
    .io_output_counts_1(io_output_counts_1), // @[:@2882.4]
    .io_output_counts_0(io_output_counts_0), // @[:@2882.4]
    .io_output_oobs_0(io_output_oobs_0), // @[:@2882.4]
    .io_output_oobs_1(io_output_oobs_1), // @[:@2882.4]
    .io_output_done(dontcare2) // @[:@2882.4]
  );

endmodule

module SRAMVerilogSim
#(
    parameter WORDS = 1024,
    parameter AWIDTH = 10,
    parameter DWIDTH = 32)
(
    input clk,
    input [AWIDTH-1:0] raddr,
    input [AWIDTH-1:0] waddr,
    input raddrEn,
    input waddrEn,
    input wen,
    input [DWIDTH-1:0] wdata,
    input backpressure,
    output reg [DWIDTH-1:0] rdata
);

    reg [DWIDTH-1:0] mem [0:WORDS-1];

    always @(posedge clk) begin
      if (wen) mem[waddr] <= wdata;
      if (backpressure) rdata <= mem[raddr];
    end

endmodule
module RetimeShiftRegister
#(
    parameter WIDTH = 1,
    parameter STAGES = 1)
(
    input clock,
    input reset,
    input flow,
    input [WIDTH-1:0] init,
    input [WIDTH-1:0] in,
    output reg [WIDTH-1:0] out
);
  integer i;
  reg [WIDTH-1:0] sr[STAGES:0]; // Create 'STAGES' number of register, each 'WIDTH' bits wide

   /* synopsys dc_tcl_script_begin
    set_ungroup [current_design] true
    set_flatten true -effort high -phase true -design [current_design]
    set_dont_retime [current_design] false
    set_optimize_registers true -design [current_design]
    */
  always @(posedge clock) begin
    if (reset) begin
      for(i=0; i<STAGES; i=i+1) begin
        sr[i] <= init;
      end
    end else begin
      if (flow) begin 
        sr[0] <= in;
        for(i=1; i<STAGES; i=i+1) begin
          sr[i] <= sr[i-1];
        end
      end
    end
  end

  always @(*) begin
    out = sr[STAGES-1];
  end
endmodule
module FF( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  output [31:0] io_rPort_0_output_0, // @[:@6.4]
  input  [31:0] io_wPort_0_data_0, // @[:@6.4]
  input         io_wPort_0_reset, // @[:@6.4]
  input         io_wPort_0_en_0 // @[:@6.4]
);
  reg [31:0] ff; // @[MemPrimitives.scala 173:19:@21.4]
  reg [31:0] _RAND_0;
  wire [31:0] _T_68; // @[MemPrimitives.scala 177:32:@23.4]
  wire [31:0] _T_69; // @[MemPrimitives.scala 177:12:@24.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 177:32:@23.4]
  assign _T_69 = io_wPort_0_reset ? 32'h0 : _T_68; // @[MemPrimitives.scala 177:12:@24.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 178:34:@26.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 32'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 32'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SRFF( // @[:@28.2]
  input   clock, // @[:@29.4]
  input   reset, // @[:@30.4]
  input   io_input_set, // @[:@31.4]
  input   io_input_reset, // @[:@31.4]
  input   io_input_asyn_reset, // @[:@31.4]
  output  io_output // @[:@31.4]
);
  reg  _T_15; // @[SRFF.scala 20:21:@33.4]
  reg [31:0] _RAND_0;
  wire  _T_19; // @[SRFF.scala 21:74:@34.4]
  wire  _T_20; // @[SRFF.scala 21:48:@35.4]
  wire  _T_21; // @[SRFF.scala 21:14:@36.4]
  assign _T_19 = io_input_reset ? 1'h0 : _T_15; // @[SRFF.scala 21:74:@34.4]
  assign _T_20 = io_input_set ? 1'h1 : _T_19; // @[SRFF.scala 21:48:@35.4]
  assign _T_21 = io_input_asyn_reset ? 1'h0 : _T_20; // @[SRFF.scala 21:14:@36.4]
  assign io_output = io_input_asyn_reset ? 1'h0 : _T_15; // @[SRFF.scala 22:15:@39.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_15 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_15 <= 1'h0;
    end else begin
      if (io_input_asyn_reset) begin
        _T_15 <= 1'h0;
      end else begin
        if (io_input_set) begin
          _T_15 <= 1'h1;
        end else begin
          if (io_input_reset) begin
            _T_15 <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module SingleCounter( // @[:@41.2]
  input   clock, // @[:@42.4]
  input   reset, // @[:@43.4]
  input   io_input_reset, // @[:@44.4]
  output  io_output_done // @[:@44.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@57.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@57.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@57.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@57.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@57.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@57.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@73.4]
  wire [12:0] _T_48; // @[Counter.scala 287:52:@101.4]
  wire [13:0] _T_50; // @[Counter.scala 291:33:@102.4]
  wire [12:0] _T_51; // @[Counter.scala 291:33:@103.4]
  wire [12:0] _T_52; // @[Counter.scala 291:33:@104.4]
  wire  _T_57; // @[Counter.scala 293:18:@106.4]
  wire [12:0] _T_68; // @[Counter.scala 299:115:@114.4]
  wire [12:0] _T_71; // @[Counter.scala 299:152:@117.4]
  wire [12:0] _T_72; // @[Counter.scala 299:74:@118.4]
  FF bases_0 ( // @[Counter.scala 261:53:@57.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@73.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@101.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@102.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@103.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@104.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh3f); // @[Counter.scala 293:18:@106.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@114.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@117.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 299:74:@118.4]
  assign io_output_done = $signed(_T_52) >= $signed(32'sh3f); // @[Counter.scala 333:20:@127.4]
  assign bases_0_clock = clock; // @[:@58.4]
  assign bases_0_reset = reset; // @[:@59.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 299:31:@120.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@99.4]
  assign bases_0_io_wPort_0_en_0 = 1'h1; // @[Counter.scala 284:29:@100.4]
  assign SRFF_clock = clock; // @[:@74.4]
  assign SRFF_reset = reset; // @[:@75.4]
  assign SRFF_io_input_set = io_input_reset == 1'h0; // @[Counter.scala 264:23:@78.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@80.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@81.4]
endmodule
module RetimeWrapper( // @[:@144.2]
  input   clock, // @[:@145.4]
  input   reset, // @[:@146.4]
  input   io_flow, // @[:@147.4]
  input   io_in, // @[:@147.4]
  output  io_out // @[:@147.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@149.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@149.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@162.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@161.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@160.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@159.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@158.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@156.4]
endmodule
module RootController_sm( // @[:@312.2]
  input   clock, // @[:@313.4]
  input   reset, // @[:@314.4]
  input   io_enable, // @[:@315.4]
  output  io_done, // @[:@315.4]
  input   io_rst, // @[:@315.4]
  input   io_ctrDone, // @[:@315.4]
  output  io_ctrInc, // @[:@315.4]
  input   io_doneIn_0, // @[:@315.4]
  output  io_enableOut_0, // @[:@315.4]
  output  io_childAck_0 // @[:@315.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@318.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@321.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@338.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@433.4]
  wire  finished; // @[Controllers.scala 81:26:@324.4]
  wire  synchronize; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  wire  _T_122; // @[Controllers.scala 128:33:@371.4]
  wire  _T_124; // @[Controllers.scala 128:54:@372.4]
  wire  _T_125; // @[Controllers.scala 128:52:@373.4]
  wire  _T_126; // @[Controllers.scala 128:66:@374.4]
  wire  _T_128; // @[Controllers.scala 128:98:@376.4]
  wire  _T_129; // @[Controllers.scala 128:96:@377.4]
  wire  _T_131; // @[Controllers.scala 128:123:@378.4]
  wire  _T_133; // @[Controllers.scala 129:48:@381.4]
  wire  _T_138; // @[Controllers.scala 130:52:@386.4]
  wire  _T_139; // @[Controllers.scala 130:50:@387.4]
  wire  _T_147; // @[Controllers.scala 130:129:@393.4]
  wire  _T_150; // @[Controllers.scala 131:45:@396.4]
  wire  _T_154; // @[Controllers.scala 213:68:@402.4]
  wire  _T_156; // @[Controllers.scala 213:90:@404.4]
  wire  _T_158; // @[Controllers.scala 213:132:@406.4]
  wire  _T_159; // @[Controllers.scala 213:130:@407.4]
  wire  _T_160; // @[Controllers.scala 213:156:@408.4]
  reg  _T_166; // @[package.scala 48:56:@412.4]
  reg [31:0] _RAND_0;
  reg  _T_180; // @[package.scala 48:56:@430.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@318.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@321.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@338.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@357.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@416.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@433.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  assign finished = done_0_io_output | io_done; // @[Controllers.scala 81:26:@324.4]
  assign synchronize = RetimeWrapper_io_out; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  assign _T_122 = done_0_io_output == 1'h0; // @[Controllers.scala 128:33:@371.4]
  assign _T_124 = io_ctrDone == 1'h0; // @[Controllers.scala 128:54:@372.4]
  assign _T_125 = _T_122 & _T_124; // @[Controllers.scala 128:52:@373.4]
  assign _T_126 = _T_125 & io_enable; // @[Controllers.scala 128:66:@374.4]
  assign _T_128 = ~ iterDone_0_io_output; // @[Controllers.scala 128:98:@376.4]
  assign _T_129 = _T_126 & _T_128; // @[Controllers.scala 128:96:@377.4]
  assign _T_131 = io_doneIn_0 == 1'h0; // @[Controllers.scala 128:123:@378.4]
  assign _T_133 = io_doneIn_0 | io_rst; // @[Controllers.scala 129:48:@381.4]
  assign _T_138 = synchronize == 1'h0; // @[Controllers.scala 130:52:@386.4]
  assign _T_139 = io_doneIn_0 & _T_138; // @[Controllers.scala 130:50:@387.4]
  assign _T_147 = finished == 1'h0; // @[Controllers.scala 130:129:@393.4]
  assign _T_150 = io_rst == 1'h0; // @[Controllers.scala 131:45:@396.4]
  assign _T_154 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@402.4]
  assign _T_156 = _T_154 & _T_128; // @[Controllers.scala 213:90:@404.4]
  assign _T_158 = ~ done_0_io_output; // @[Controllers.scala 213:132:@406.4]
  assign _T_159 = _T_156 & _T_158; // @[Controllers.scala 213:130:@407.4]
  assign _T_160 = ~ io_ctrDone; // @[Controllers.scala 213:156:@408.4]
  assign io_done = RetimeWrapper_2_io_out; // @[Controllers.scala 245:13:@440.4]
  assign io_ctrInc = io_doneIn_0; // @[Controllers.scala 122:17:@356.4]
  assign io_enableOut_0 = _T_159 & _T_160; // @[Controllers.scala 213:55:@410.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@401.4]
  assign active_0_clock = clock; // @[:@319.4]
  assign active_0_reset = reset; // @[:@320.4]
  assign active_0_io_input_set = _T_129 & _T_131; // @[Controllers.scala 128:30:@380.4]
  assign active_0_io_input_reset = _T_133 | done_0_io_output; // @[Controllers.scala 129:32:@385.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@326.4]
  assign done_0_clock = clock; // @[:@322.4]
  assign done_0_reset = reset; // @[:@323.4]
  assign done_0_io_input_set = io_ctrDone & _T_150; // @[Controllers.scala 131:28:@399.4]
  assign done_0_io_input_reset = io_rst | done_0_io_output; // @[Controllers.scala 86:33:@336.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@327.4]
  assign iterDone_0_clock = clock; // @[:@339.4]
  assign iterDone_0_reset = reset; // @[:@340.4]
  assign iterDone_0_io_input_set = _T_139 & _T_147; // @[Controllers.scala 130:32:@395.4]
  assign iterDone_0_io_input_reset = synchronize | io_rst; // @[Controllers.scala 92:37:@350.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@341.4]
  assign RetimeWrapper_clock = clock; // @[:@358.4]
  assign RetimeWrapper_reset = reset; // @[:@359.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@361.4]
  assign RetimeWrapper_io_in = io_doneIn_0; // @[package.scala 94:16:@360.4]
  assign RetimeWrapper_1_clock = clock; // @[:@417.4]
  assign RetimeWrapper_1_reset = reset; // @[:@418.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@420.4]
  assign RetimeWrapper_1_io_in = done_0_io_output & _T_166; // @[package.scala 94:16:@419.4]
  assign RetimeWrapper_2_clock = clock; // @[:@434.4]
  assign RetimeWrapper_2_reset = reset; // @[:@435.4]
  assign RetimeWrapper_2_io_flow = io_enable; // @[package.scala 95:18:@437.4]
  assign RetimeWrapper_2_io_in = done_0_io_output & _T_180; // @[package.scala 94:16:@436.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_166 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_180 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_166 <= 1'h0;
    end else begin
      _T_166 <= _T_122;
    end
    if (reset) begin
      _T_180 <= 1'h0;
    end else begin
      _T_180 <= _T_122;
    end
  end
endmodule
module x543_outr_UnitPipe_sm( // @[:@2390.2]
  input   clock, // @[:@2391.4]
  input   reset, // @[:@2392.4]
  input   io_enable, // @[:@2393.4]
  output  io_done, // @[:@2393.4]
  input   io_parentAck, // @[:@2393.4]
  input   io_doneIn_0, // @[:@2393.4]
  output  io_enableOut_0, // @[:@2393.4]
  output  io_childAck_0, // @[:@2393.4]
  input   io_ctrCopyDone_0 // @[:@2393.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@2396.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@2396.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@2396.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@2396.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@2396.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@2396.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@2399.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@2399.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@2399.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@2399.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@2399.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@2399.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@2416.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@2416.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@2416.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@2416.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@2416.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@2416.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@2447.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@2447.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@2447.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@2447.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@2447.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@2461.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@2461.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@2461.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@2461.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@2461.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@2479.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@2479.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@2479.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@2479.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@2479.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@2516.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@2516.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@2516.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@2516.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@2516.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@2533.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@2533.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@2533.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@2533.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@2533.4]
  wire  _T_105; // @[Controllers.scala 165:35:@2431.4]
  wire  _T_107; // @[Controllers.scala 165:60:@2432.4]
  wire  _T_108; // @[Controllers.scala 165:58:@2433.4]
  wire  _T_110; // @[Controllers.scala 165:76:@2434.4]
  wire  _T_111; // @[Controllers.scala 165:74:@2435.4]
  wire  _T_115; // @[Controllers.scala 165:109:@2438.4]
  wire  _T_118; // @[Controllers.scala 165:141:@2440.4]
  wire  _T_126; // @[package.scala 96:25:@2452.4 package.scala 96:25:@2453.4]
  wire  _T_130; // @[Controllers.scala 167:54:@2455.4]
  wire  _T_131; // @[Controllers.scala 167:52:@2456.4]
  wire  _T_138; // @[package.scala 96:25:@2466.4 package.scala 96:25:@2467.4]
  wire  _T_156; // @[package.scala 96:25:@2484.4 package.scala 96:25:@2485.4]
  wire  _T_160; // @[Controllers.scala 169:67:@2487.4]
  wire  _T_161; // @[Controllers.scala 169:86:@2488.4]
  wire  _T_174; // @[Controllers.scala 213:68:@2502.4]
  wire  _T_176; // @[Controllers.scala 213:90:@2504.4]
  wire  _T_178; // @[Controllers.scala 213:132:@2506.4]
  reg  _T_186; // @[package.scala 48:56:@2512.4]
  reg [31:0] _RAND_0;
  wire  _T_187; // @[package.scala 100:41:@2514.4]
  reg  _T_200; // @[package.scala 48:56:@2530.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@2396.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@2399.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@2416.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@2447.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@2461.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@2479.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@2516.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@2533.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_105 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@2431.4]
  assign _T_107 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@2432.4]
  assign _T_108 = _T_105 & _T_107; // @[Controllers.scala 165:58:@2433.4]
  assign _T_110 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@2434.4]
  assign _T_111 = _T_108 & _T_110; // @[Controllers.scala 165:74:@2435.4]
  assign _T_115 = _T_111 & io_enable; // @[Controllers.scala 165:109:@2438.4]
  assign _T_118 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@2440.4]
  assign _T_126 = RetimeWrapper_io_out; // @[package.scala 96:25:@2452.4 package.scala 96:25:@2453.4]
  assign _T_130 = _T_126 == 1'h0; // @[Controllers.scala 167:54:@2455.4]
  assign _T_131 = io_doneIn_0 | _T_130; // @[Controllers.scala 167:52:@2456.4]
  assign _T_138 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@2466.4 package.scala 96:25:@2467.4]
  assign _T_156 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@2484.4 package.scala 96:25:@2485.4]
  assign _T_160 = _T_156 == 1'h0; // @[Controllers.scala 169:67:@2487.4]
  assign _T_161 = _T_160 & io_enable; // @[Controllers.scala 169:86:@2488.4]
  assign _T_174 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@2502.4]
  assign _T_176 = _T_174 & _T_105; // @[Controllers.scala 213:90:@2504.4]
  assign _T_178 = ~ done_0_io_output; // @[Controllers.scala 213:132:@2506.4]
  assign _T_187 = done_0_io_output & _T_186; // @[package.scala 100:41:@2514.4]
  assign io_done = RetimeWrapper_4_io_out; // @[Controllers.scala 245:13:@2540.4]
  assign io_enableOut_0 = _T_176 & _T_178; // @[Controllers.scala 213:55:@2510.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@2501.4]
  assign active_0_clock = clock; // @[:@2397.4]
  assign active_0_reset = reset; // @[:@2398.4]
  assign active_0_io_input_set = _T_115 & _T_118; // @[Controllers.scala 165:32:@2442.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@2446.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@2404.4]
  assign done_0_clock = clock; // @[:@2400.4]
  assign done_0_reset = reset; // @[:@2401.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_161; // @[Controllers.scala 169:30:@2492.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@2414.4 Controllers.scala 170:32:@2499.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@2405.4]
  assign iterDone_0_clock = clock; // @[:@2417.4]
  assign iterDone_0_reset = reset; // @[:@2418.4]
  assign iterDone_0_io_input_set = _T_131 & io_enable; // @[Controllers.scala 167:34:@2460.4]
  assign iterDone_0_io_input_reset = _T_138 | io_parentAck; // @[Controllers.scala 92:37:@2428.4 Controllers.scala 168:36:@2476.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@2419.4]
  assign RetimeWrapper_clock = clock; // @[:@2448.4]
  assign RetimeWrapper_reset = reset; // @[:@2449.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@2451.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@2450.4]
  assign RetimeWrapper_1_clock = clock; // @[:@2462.4]
  assign RetimeWrapper_1_reset = reset; // @[:@2463.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@2465.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@2464.4]
  assign RetimeWrapper_2_clock = clock; // @[:@2480.4]
  assign RetimeWrapper_2_reset = reset; // @[:@2481.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@2483.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@2482.4]
  assign RetimeWrapper_3_clock = clock; // @[:@2517.4]
  assign RetimeWrapper_3_reset = reset; // @[:@2518.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@2520.4]
  assign RetimeWrapper_3_io_in = _T_187 | io_parentAck; // @[package.scala 94:16:@2519.4]
  assign RetimeWrapper_4_clock = clock; // @[:@2534.4]
  assign RetimeWrapper_4_reset = reset; // @[:@2535.4]
  assign RetimeWrapper_4_io_flow = io_enable; // @[package.scala 95:18:@2537.4]
  assign RetimeWrapper_4_io_in = done_0_io_output & _T_200; // @[package.scala 94:16:@2536.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_186 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_200 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_186 <= 1'h0;
    end else begin
      _T_186 <= _T_110;
    end
    if (reset) begin
      _T_200 <= 1'h0;
    end else begin
      _T_200 <= _T_110;
    end
  end
endmodule
module SingleCounter_1( // @[:@2661.2]
  input         clock, // @[:@2662.4]
  input         reset, // @[:@2663.4]
  input         io_input_reset, // @[:@2664.4]
  input         io_input_enable, // @[:@2664.4]
  output [31:0] io_output_count_0, // @[:@2664.4]
  output        io_output_oobs_0, // @[:@2664.4]
  output        io_output_done, // @[:@2664.4]
  output        io_output_saturated // @[:@2664.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@2677.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@2677.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@2677.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@2677.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@2677.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@2677.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@2693.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@2693.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@2693.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@2693.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@2693.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@2693.4]
  wire  _T_36; // @[Counter.scala 264:45:@2696.4]
  wire [12:0] _T_48; // @[Counter.scala 287:52:@2721.4]
  wire [13:0] _T_50; // @[Counter.scala 291:33:@2722.4]
  wire [12:0] _T_51; // @[Counter.scala 291:33:@2723.4]
  wire [12:0] _T_52; // @[Counter.scala 291:33:@2724.4]
  wire  _T_57; // @[Counter.scala 293:18:@2726.4]
  wire [12:0] _T_68; // @[Counter.scala 299:115:@2734.4]
  wire [12:0] _T_71; // @[Counter.scala 299:152:@2737.4]
  wire [12:0] _T_72; // @[Counter.scala 299:74:@2738.4]
  wire  _T_75; // @[Counter.scala 322:102:@2742.4]
  wire  _T_77; // @[Counter.scala 322:130:@2743.4]
  FF bases_0 ( // @[Counter.scala 261:53:@2677.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@2693.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@2696.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@2721.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@2722.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@2723.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@2724.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh780); // @[Counter.scala 293:18:@2726.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@2734.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@2737.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 299:74:@2738.4]
  assign _T_75 = $signed(_T_48) < $signed(32'sh0); // @[Counter.scala 322:102:@2742.4]
  assign _T_77 = $signed(_T_48) >= $signed(32'sh780); // @[Counter.scala 322:130:@2743.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@2741.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@2745.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@2747.4]
  assign io_output_saturated = $signed(_T_52) >= $signed(32'sh780); // @[Counter.scala 340:25:@2750.4]
  assign bases_0_clock = clock; // @[:@2678.4]
  assign bases_0_reset = reset; // @[:@2679.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 299:31:@2740.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@2719.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@2720.4]
  assign SRFF_clock = clock; // @[:@2694.4]
  assign SRFF_reset = reset; // @[:@2695.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@2698.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@2700.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@2701.4]
endmodule
module SingleCounter_2( // @[:@2790.2]
  input         clock, // @[:@2791.4]
  input         reset, // @[:@2792.4]
  input         io_setup_saturate, // @[:@2793.4]
  input         io_input_reset, // @[:@2793.4]
  input         io_input_enable, // @[:@2793.4]
  output [31:0] io_output_count_0, // @[:@2793.4]
  output        io_output_oobs_0, // @[:@2793.4]
  output        io_output_done // @[:@2793.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@2806.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@2806.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@2806.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@2806.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@2806.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@2806.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@2822.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@2822.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@2822.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@2822.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@2822.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@2822.4]
  wire  _T_36; // @[Counter.scala 264:45:@2825.4]
  wire [12:0] _T_48; // @[Counter.scala 287:52:@2850.4]
  wire [13:0] _T_50; // @[Counter.scala 291:33:@2851.4]
  wire [12:0] _T_51; // @[Counter.scala 291:33:@2852.4]
  wire [12:0] _T_52; // @[Counter.scala 291:33:@2853.4]
  wire  _T_57; // @[Counter.scala 293:18:@2855.4]
  wire [12:0] _T_68; // @[Counter.scala 299:115:@2863.4]
  wire [12:0] _T_70; // @[Counter.scala 299:85:@2865.4]
  wire [12:0] _T_71; // @[Counter.scala 299:152:@2866.4]
  wire [12:0] _T_72; // @[Counter.scala 299:74:@2867.4]
  wire  _T_75; // @[Counter.scala 322:102:@2871.4]
  wire  _T_77; // @[Counter.scala 322:130:@2872.4]
  FF bases_0 ( // @[Counter.scala 261:53:@2806.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@2822.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@2825.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@2850.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh4); // @[Counter.scala 291:33:@2851.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh4); // @[Counter.scala 291:33:@2852.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@2853.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh400); // @[Counter.scala 293:18:@2855.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@2863.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 32'h0; // @[Counter.scala 299:85:@2865.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@2866.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 299:74:@2867.4]
  assign _T_75 = $signed(_T_48) < $signed(32'sh0); // @[Counter.scala 322:102:@2871.4]
  assign _T_77 = $signed(_T_48) >= $signed(32'sh400); // @[Counter.scala 322:130:@2872.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@2870.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@2874.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@2876.4]
  assign bases_0_clock = clock; // @[:@2807.4]
  assign bases_0_reset = reset; // @[:@2808.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 299:31:@2869.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@2848.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@2849.4]
  assign SRFF_clock = clock; // @[:@2823.4]
  assign SRFF_reset = reset; // @[:@2824.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@2827.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@2829.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@2830.4]
endmodule
module x324_ctrchain( // @[:@2881.2]
  input         clock, // @[:@2882.4]
  input         reset, // @[:@2883.4]
  input         io_input_reset, // @[:@2884.4]
  input         io_input_enable, // @[:@2884.4]
  output [31:0] io_output_counts_1, // @[:@2884.4]
  output [31:0] io_output_counts_0, // @[:@2884.4]
  output        io_output_oobs_0, // @[:@2884.4]
  output        io_output_oobs_1, // @[:@2884.4]
  output        io_output_done // @[:@2884.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 513:46:@2886.4]
  wire  ctrs_0_reset; // @[Counter.scala 513:46:@2886.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 513:46:@2886.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 513:46:@2886.4]
  wire [31:0] ctrs_0_io_output_count_0; // @[Counter.scala 513:46:@2886.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 513:46:@2886.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 513:46:@2886.4]
  wire  ctrs_0_io_output_saturated; // @[Counter.scala 513:46:@2886.4]
  wire  ctrs_1_clock; // @[Counter.scala 513:46:@2889.4]
  wire  ctrs_1_reset; // @[Counter.scala 513:46:@2889.4]
  wire  ctrs_1_io_setup_saturate; // @[Counter.scala 513:46:@2889.4]
  wire  ctrs_1_io_input_reset; // @[Counter.scala 513:46:@2889.4]
  wire  ctrs_1_io_input_enable; // @[Counter.scala 513:46:@2889.4]
  wire [31:0] ctrs_1_io_output_count_0; // @[Counter.scala 513:46:@2889.4]
  wire  ctrs_1_io_output_oobs_0; // @[Counter.scala 513:46:@2889.4]
  wire  ctrs_1_io_output_done; // @[Counter.scala 513:46:@2889.4]
  wire  isDone; // @[Counter.scala 541:51:@2906.4]
  reg  wasDone; // @[Counter.scala 542:24:@2907.4]
  reg [31:0] _RAND_0;
  wire  _T_64; // @[Counter.scala 546:69:@2915.4]
  wire  _T_66; // @[Counter.scala 546:80:@2916.4]
  reg  doneLatch; // @[Counter.scala 550:26:@2921.4]
  reg [31:0] _RAND_1;
  wire  _T_73; // @[Counter.scala 551:48:@2922.4]
  wire  _T_74; // @[Counter.scala 551:19:@2923.4]
  SingleCounter_1 ctrs_0 ( // @[Counter.scala 513:46:@2886.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done),
    .io_output_saturated(ctrs_0_io_output_saturated)
  );
  SingleCounter_2 ctrs_1 ( // @[Counter.scala 513:46:@2889.4]
    .clock(ctrs_1_clock),
    .reset(ctrs_1_reset),
    .io_setup_saturate(ctrs_1_io_setup_saturate),
    .io_input_reset(ctrs_1_io_input_reset),
    .io_input_enable(ctrs_1_io_input_enable),
    .io_output_count_0(ctrs_1_io_output_count_0),
    .io_output_oobs_0(ctrs_1_io_output_oobs_0),
    .io_output_done(ctrs_1_io_output_done)
  );
  assign isDone = ctrs_0_io_output_done & ctrs_1_io_output_done; // @[Counter.scala 541:51:@2906.4]
  assign _T_64 = io_input_enable & isDone; // @[Counter.scala 546:69:@2915.4]
  assign _T_66 = wasDone == 1'h0; // @[Counter.scala 546:80:@2916.4]
  assign _T_73 = isDone ? 1'h1 : doneLatch; // @[Counter.scala 551:48:@2922.4]
  assign _T_74 = io_input_reset ? 1'h0 : _T_73; // @[Counter.scala 551:19:@2923.4]
  assign io_output_counts_1 = ctrs_1_io_output_count_0; // @[Counter.scala 557:32:@2928.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 557:32:@2925.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@2927.4]
  assign io_output_oobs_1 = ctrs_1_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@2930.4]
  assign io_output_done = _T_64 & _T_66; // @[Counter.scala 546:18:@2918.4]
  assign ctrs_0_clock = clock; // @[:@2887.4]
  assign ctrs_0_reset = reset; // @[:@2888.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@2895.4]
  assign ctrs_0_io_input_enable = ctrs_1_io_output_done & io_input_enable; // @[Counter.scala 526:29:@2902.4]
  assign ctrs_1_clock = clock; // @[:@2890.4]
  assign ctrs_1_reset = reset; // @[:@2891.4]
  assign ctrs_1_io_setup_saturate = ctrs_0_io_output_saturated; // @[Counter.scala 532:31:@2905.4]
  assign ctrs_1_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@2899.4]
  assign ctrs_1_io_input_enable = io_input_enable; // @[Counter.scala 524:33:@2900.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= isDone;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (isDone) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module RetimeWrapper_12( // @[:@2970.2]
  input   clock, // @[:@2971.4]
  input   reset, // @[:@2972.4]
  input   io_flow, // @[:@2973.4]
  input   io_in, // @[:@2973.4]
  output  io_out // @[:@2973.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@2975.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@2975.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@2975.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@2975.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@2975.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@2975.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(63)) sr ( // @[RetimeShiftRegister.scala 15:20:@2975.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@2988.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@2987.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@2986.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@2985.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@2984.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@2982.4]
endmodule
module RetimeWrapper_16( // @[:@3098.2]
  input   clock, // @[:@3099.4]
  input   reset, // @[:@3100.4]
  input   io_flow, // @[:@3101.4]
  input   io_in, // @[:@3101.4]
  output  io_out // @[:@3101.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3103.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3103.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3103.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3103.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3103.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3103.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(62)) sr ( // @[RetimeShiftRegister.scala 15:20:@3103.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3116.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3115.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3114.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3113.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3112.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3110.4]
endmodule
module x542_inr_Foreach_SAMPLER_BOX_sm( // @[:@3118.2]
  input   clock, // @[:@3119.4]
  input   reset, // @[:@3120.4]
  input   io_enable, // @[:@3121.4]
  output  io_done, // @[:@3121.4]
  output  io_doneLatch, // @[:@3121.4]
  input   io_ctrDone, // @[:@3121.4]
  output  io_datapathEn, // @[:@3121.4]
  output  io_ctrInc, // @[:@3121.4]
  output  io_ctrRst, // @[:@3121.4]
  input   io_parentAck, // @[:@3121.4]
  input   io_backpressure, // @[:@3121.4]
  input   io_break // @[:@3121.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@3123.4]
  wire  active_reset; // @[Controllers.scala 261:22:@3123.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@3123.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@3123.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@3123.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@3123.4]
  wire  done_clock; // @[Controllers.scala 262:20:@3126.4]
  wire  done_reset; // @[Controllers.scala 262:20:@3126.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@3126.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@3126.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@3126.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@3126.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3160.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3160.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3160.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@3160.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@3160.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@3182.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@3182.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@3182.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@3182.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@3182.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@3194.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@3194.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@3194.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@3194.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@3194.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@3202.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@3202.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@3202.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@3202.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@3202.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@3218.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@3218.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@3218.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@3218.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@3218.4]
  wire  _T_80; // @[Controllers.scala 264:48:@3131.4]
  wire  _T_81; // @[Controllers.scala 264:46:@3132.4]
  wire  _T_82; // @[Controllers.scala 264:62:@3133.4]
  wire  _T_83; // @[Controllers.scala 264:60:@3134.4]
  wire  _T_100; // @[package.scala 100:49:@3151.4]
  reg  _T_103; // @[package.scala 48:56:@3152.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@3165.4 package.scala 96:25:@3166.4]
  wire  _T_110; // @[package.scala 100:49:@3167.4]
  reg  _T_113; // @[package.scala 48:56:@3168.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@3170.4]
  wire  _T_118; // @[Controllers.scala 283:41:@3175.4]
  wire  _T_119; // @[Controllers.scala 283:59:@3176.4]
  wire  _T_121; // @[Controllers.scala 284:37:@3179.4]
  wire  _T_124; // @[package.scala 96:25:@3187.4 package.scala 96:25:@3188.4]
  wire  _T_126; // @[package.scala 100:49:@3189.4]
  reg  _T_129; // @[package.scala 48:56:@3190.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@3212.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@3214.4]
  reg  _T_153; // @[package.scala 48:56:@3215.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@3223.4 package.scala 96:25:@3224.4]
  wire  _T_158; // @[Controllers.scala 292:61:@3225.4]
  wire  _T_159; // @[Controllers.scala 292:24:@3226.4]
  SRFF active ( // @[Controllers.scala 261:22:@3123.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@3126.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_12 RetimeWrapper ( // @[package.scala 93:22:@3160.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_12 RetimeWrapper_1 ( // @[package.scala 93:22:@3182.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@3194.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@3202.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_16 RetimeWrapper_4 ( // @[package.scala 93:22:@3218.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@3131.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@3132.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@3133.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@3134.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@3151.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@3165.4 package.scala 96:25:@3166.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@3167.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@3170.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@3175.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@3176.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@3179.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@3187.4 package.scala 96:25:@3188.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@3189.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@3214.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@3223.4 package.scala 96:25:@3224.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@3225.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@3226.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@3193.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@3228.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@3178.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@3181.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@3173.4]
  assign active_clock = clock; // @[:@3124.4]
  assign active_reset = reset; // @[:@3125.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@3136.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@3140.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@3141.4]
  assign done_clock = clock; // @[:@3127.4]
  assign done_reset = reset; // @[:@3128.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@3156.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@3149.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@3150.4]
  assign RetimeWrapper_clock = clock; // @[:@3161.4]
  assign RetimeWrapper_reset = reset; // @[:@3162.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@3164.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@3163.4]
  assign RetimeWrapper_1_clock = clock; // @[:@3183.4]
  assign RetimeWrapper_1_reset = reset; // @[:@3184.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@3186.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@3185.4]
  assign RetimeWrapper_2_clock = clock; // @[:@3195.4]
  assign RetimeWrapper_2_reset = reset; // @[:@3196.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@3198.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@3197.4]
  assign RetimeWrapper_3_clock = clock; // @[:@3203.4]
  assign RetimeWrapper_3_reset = reset; // @[:@3204.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@3206.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@3205.4]
  assign RetimeWrapper_4_clock = clock; // @[:@3219.4]
  assign RetimeWrapper_4_reset = reset; // @[:@3220.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@3222.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@3221.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module SimBlackBoxesfix2fixBox( // @[:@3335.2]
  input  [31:0] io_a, // @[:@3338.4]
  output [31:0] io_b // @[:@3338.4]
);
  assign io_b = io_a; // @[SimBlackBoxes.scala 99:40:@3351.4]
endmodule
module _( // @[:@3353.2]
  input  [31:0] io_b, // @[:@3356.4]
  output [31:0] io_result // @[:@3356.4]
);
  wire [31:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@3361.4]
  wire [31:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@3361.4]
  SimBlackBoxesfix2fixBox SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@3361.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@3374.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@3369.4]
endmodule
module SRAM( // @[:@3433.2]
  input        clock, // @[:@3434.4]
  input  [7:0] io_raddr, // @[:@3436.4]
  input        io_wen, // @[:@3436.4]
  input  [7:0] io_waddr, // @[:@3436.4]
  input  [7:0] io_wdata, // @[:@3436.4]
  output [7:0] io_rdata, // @[:@3436.4]
  input        io_backpressure // @[:@3436.4]
);
  wire [7:0] SRAMVerilogSim_rdata; // @[SRAM.scala 143:23:@3438.4]
  wire [7:0] SRAMVerilogSim_wdata; // @[SRAM.scala 143:23:@3438.4]
  wire  SRAMVerilogSim_backpressure; // @[SRAM.scala 143:23:@3438.4]
  wire  SRAMVerilogSim_wen; // @[SRAM.scala 143:23:@3438.4]
  wire  SRAMVerilogSim_waddrEn; // @[SRAM.scala 143:23:@3438.4]
  wire  SRAMVerilogSim_raddrEn; // @[SRAM.scala 143:23:@3438.4]
  wire [7:0] SRAMVerilogSim_waddr; // @[SRAM.scala 143:23:@3438.4]
  wire [7:0] SRAMVerilogSim_raddr; // @[SRAM.scala 143:23:@3438.4]
  wire  SRAMVerilogSim_clk; // @[SRAM.scala 143:23:@3438.4]
  SRAMVerilogSim #(.DWIDTH(8), .WORDS(171), .AWIDTH(8)) SRAMVerilogSim ( // @[SRAM.scala 143:23:@3438.4]
    .rdata(SRAMVerilogSim_rdata),
    .wdata(SRAMVerilogSim_wdata),
    .backpressure(SRAMVerilogSim_backpressure),
    .wen(SRAMVerilogSim_wen),
    .waddrEn(SRAMVerilogSim_waddrEn),
    .raddrEn(SRAMVerilogSim_raddrEn),
    .waddr(SRAMVerilogSim_waddr),
    .raddr(SRAMVerilogSim_raddr),
    .clk(SRAMVerilogSim_clk)
  );
  assign io_rdata = SRAMVerilogSim_rdata; // @[SRAM.scala 153:16:@3458.4]
  assign SRAMVerilogSim_wdata = io_wdata; // @[SRAM.scala 148:20:@3452.4]
  assign SRAMVerilogSim_backpressure = io_backpressure; // @[SRAM.scala 149:27:@3453.4]
  assign SRAMVerilogSim_wen = io_wen; // @[SRAM.scala 146:18:@3450.4]
  assign SRAMVerilogSim_waddrEn = 1'h1; // @[SRAM.scala 151:22:@3455.4]
  assign SRAMVerilogSim_raddrEn = 1'h1; // @[SRAM.scala 150:22:@3454.4]
  assign SRAMVerilogSim_waddr = io_waddr; // @[SRAM.scala 147:20:@3451.4]
  assign SRAMVerilogSim_raddr = io_raddr; // @[SRAM.scala 145:20:@3449.4]
  assign SRAMVerilogSim_clk = clock; // @[SRAM.scala 144:18:@3448.4]
endmodule
module RetimeWrapper_20( // @[:@3472.2]
  input        clock, // @[:@3473.4]
  input        reset, // @[:@3474.4]
  input        io_flow, // @[:@3475.4]
  input  [7:0] io_in, // @[:@3475.4]
  output [7:0] io_out // @[:@3475.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@3477.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@3477.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@3477.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3477.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3477.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3477.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@3477.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3490.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3489.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@3488.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3487.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3486.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3484.4]
endmodule
module Mem1D_4( // @[:@3492.2]
  input        clock, // @[:@3493.4]
  input        reset, // @[:@3494.4]
  input  [7:0] io_r_ofs_0, // @[:@3495.4]
  input        io_r_backpressure, // @[:@3495.4]
  input  [7:0] io_w_ofs_0, // @[:@3495.4]
  input  [7:0] io_w_data_0, // @[:@3495.4]
  input        io_w_en_0, // @[:@3495.4]
  output [7:0] io_output // @[:@3495.4]
);
  wire  SRAM_clock; // @[MemPrimitives.scala 567:21:@3499.4]
  wire [7:0] SRAM_io_raddr; // @[MemPrimitives.scala 567:21:@3499.4]
  wire  SRAM_io_wen; // @[MemPrimitives.scala 567:21:@3499.4]
  wire [7:0] SRAM_io_waddr; // @[MemPrimitives.scala 567:21:@3499.4]
  wire [7:0] SRAM_io_wdata; // @[MemPrimitives.scala 567:21:@3499.4]
  wire [7:0] SRAM_io_rdata; // @[MemPrimitives.scala 567:21:@3499.4]
  wire  SRAM_io_backpressure; // @[MemPrimitives.scala 567:21:@3499.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3502.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3502.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3502.4]
  wire [7:0] RetimeWrapper_io_in; // @[package.scala 93:22:@3502.4]
  wire [7:0] RetimeWrapper_io_out; // @[package.scala 93:22:@3502.4]
  wire  wInBound; // @[MemPrimitives.scala 554:32:@3497.4]
  SRAM SRAM ( // @[MemPrimitives.scala 567:21:@3499.4]
    .clock(SRAM_clock),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata(SRAM_io_wdata),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  RetimeWrapper_20 RetimeWrapper ( // @[package.scala 93:22:@3502.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign wInBound = io_w_ofs_0 <= 8'hab; // @[MemPrimitives.scala 554:32:@3497.4]
  assign io_output = SRAM_io_rdata; // @[MemPrimitives.scala 574:17:@3515.4]
  assign SRAM_clock = clock; // @[:@3500.4]
  assign SRAM_io_raddr = RetimeWrapper_io_out; // @[MemPrimitives.scala 568:37:@3509.4]
  assign SRAM_io_wen = io_w_en_0 & wInBound; // @[MemPrimitives.scala 571:22:@3512.4]
  assign SRAM_io_waddr = io_w_ofs_0; // @[MemPrimitives.scala 570:22:@3510.4]
  assign SRAM_io_wdata = io_w_data_0; // @[MemPrimitives.scala 572:22:@3513.4]
  assign SRAM_io_backpressure = io_r_backpressure; // @[MemPrimitives.scala 573:30:@3514.4]
  assign RetimeWrapper_clock = clock; // @[:@3503.4]
  assign RetimeWrapper_reset = reset; // @[:@3504.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@3506.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@3505.4]
endmodule
module StickySelects( // @[:@5817.2]
  input   clock, // @[:@5818.4]
  input   reset, // @[:@5819.4]
  input   io_ins_0, // @[:@5820.4]
  input   io_ins_1, // @[:@5820.4]
  input   io_ins_2, // @[:@5820.4]
  input   io_ins_3, // @[:@5820.4]
  input   io_ins_4, // @[:@5820.4]
  input   io_ins_5, // @[:@5820.4]
  input   io_ins_6, // @[:@5820.4]
  input   io_ins_7, // @[:@5820.4]
  input   io_ins_8, // @[:@5820.4]
  output  io_outs_0, // @[:@5820.4]
  output  io_outs_1, // @[:@5820.4]
  output  io_outs_2, // @[:@5820.4]
  output  io_outs_3, // @[:@5820.4]
  output  io_outs_4, // @[:@5820.4]
  output  io_outs_5, // @[:@5820.4]
  output  io_outs_6, // @[:@5820.4]
  output  io_outs_7, // @[:@5820.4]
  output  io_outs_8 // @[:@5820.4]
);
  reg  _T_19; // @[StickySelects.scala 21:22:@5822.4]
  reg [31:0] _RAND_0;
  wire  _T_20; // @[StickySelects.scala 22:54:@5823.4]
  wire  _T_21; // @[StickySelects.scala 22:54:@5824.4]
  wire  _T_22; // @[StickySelects.scala 22:54:@5825.4]
  wire  _T_23; // @[StickySelects.scala 22:54:@5826.4]
  wire  _T_24; // @[StickySelects.scala 22:54:@5827.4]
  wire  _T_25; // @[StickySelects.scala 22:54:@5828.4]
  wire  _T_26; // @[StickySelects.scala 22:54:@5829.4]
  wire  _T_28; // @[StickySelects.scala 24:52:@5830.4]
  wire  _T_29; // @[StickySelects.scala 24:21:@5831.4]
  reg  _T_32; // @[StickySelects.scala 21:22:@5833.4]
  reg [31:0] _RAND_1;
  wire  _T_33; // @[StickySelects.scala 22:54:@5834.4]
  wire  _T_34; // @[StickySelects.scala 22:54:@5835.4]
  wire  _T_35; // @[StickySelects.scala 22:54:@5836.4]
  wire  _T_36; // @[StickySelects.scala 22:54:@5837.4]
  wire  _T_37; // @[StickySelects.scala 22:54:@5838.4]
  wire  _T_38; // @[StickySelects.scala 22:54:@5839.4]
  wire  _T_39; // @[StickySelects.scala 22:54:@5840.4]
  wire  _T_41; // @[StickySelects.scala 24:52:@5841.4]
  wire  _T_42; // @[StickySelects.scala 24:21:@5842.4]
  reg  _T_45; // @[StickySelects.scala 21:22:@5844.4]
  reg [31:0] _RAND_2;
  wire  _T_46; // @[StickySelects.scala 22:54:@5845.4]
  wire  _T_47; // @[StickySelects.scala 22:54:@5846.4]
  wire  _T_48; // @[StickySelects.scala 22:54:@5847.4]
  wire  _T_49; // @[StickySelects.scala 22:54:@5848.4]
  wire  _T_50; // @[StickySelects.scala 22:54:@5849.4]
  wire  _T_51; // @[StickySelects.scala 22:54:@5850.4]
  wire  _T_52; // @[StickySelects.scala 22:54:@5851.4]
  wire  _T_54; // @[StickySelects.scala 24:52:@5852.4]
  wire  _T_55; // @[StickySelects.scala 24:21:@5853.4]
  reg  _T_58; // @[StickySelects.scala 21:22:@5855.4]
  reg [31:0] _RAND_3;
  wire  _T_60; // @[StickySelects.scala 22:54:@5857.4]
  wire  _T_61; // @[StickySelects.scala 22:54:@5858.4]
  wire  _T_62; // @[StickySelects.scala 22:54:@5859.4]
  wire  _T_63; // @[StickySelects.scala 22:54:@5860.4]
  wire  _T_64; // @[StickySelects.scala 22:54:@5861.4]
  wire  _T_65; // @[StickySelects.scala 22:54:@5862.4]
  wire  _T_67; // @[StickySelects.scala 24:52:@5863.4]
  wire  _T_68; // @[StickySelects.scala 24:21:@5864.4]
  reg  _T_71; // @[StickySelects.scala 21:22:@5866.4]
  reg [31:0] _RAND_4;
  wire  _T_74; // @[StickySelects.scala 22:54:@5869.4]
  wire  _T_75; // @[StickySelects.scala 22:54:@5870.4]
  wire  _T_76; // @[StickySelects.scala 22:54:@5871.4]
  wire  _T_77; // @[StickySelects.scala 22:54:@5872.4]
  wire  _T_78; // @[StickySelects.scala 22:54:@5873.4]
  wire  _T_80; // @[StickySelects.scala 24:52:@5874.4]
  wire  _T_81; // @[StickySelects.scala 24:21:@5875.4]
  reg  _T_84; // @[StickySelects.scala 21:22:@5877.4]
  reg [31:0] _RAND_5;
  wire  _T_88; // @[StickySelects.scala 22:54:@5881.4]
  wire  _T_89; // @[StickySelects.scala 22:54:@5882.4]
  wire  _T_90; // @[StickySelects.scala 22:54:@5883.4]
  wire  _T_91; // @[StickySelects.scala 22:54:@5884.4]
  wire  _T_93; // @[StickySelects.scala 24:52:@5885.4]
  wire  _T_94; // @[StickySelects.scala 24:21:@5886.4]
  reg  _T_97; // @[StickySelects.scala 21:22:@5888.4]
  reg [31:0] _RAND_6;
  wire  _T_102; // @[StickySelects.scala 22:54:@5893.4]
  wire  _T_103; // @[StickySelects.scala 22:54:@5894.4]
  wire  _T_104; // @[StickySelects.scala 22:54:@5895.4]
  wire  _T_106; // @[StickySelects.scala 24:52:@5896.4]
  wire  _T_107; // @[StickySelects.scala 24:21:@5897.4]
  reg  _T_110; // @[StickySelects.scala 21:22:@5899.4]
  reg [31:0] _RAND_7;
  wire  _T_116; // @[StickySelects.scala 22:54:@5905.4]
  wire  _T_117; // @[StickySelects.scala 22:54:@5906.4]
  wire  _T_119; // @[StickySelects.scala 24:52:@5907.4]
  wire  _T_120; // @[StickySelects.scala 24:21:@5908.4]
  reg  _T_123; // @[StickySelects.scala 21:22:@5910.4]
  reg [31:0] _RAND_8;
  wire  _T_130; // @[StickySelects.scala 22:54:@5917.4]
  wire  _T_132; // @[StickySelects.scala 24:52:@5918.4]
  wire  _T_133; // @[StickySelects.scala 24:21:@5919.4]
  assign _T_20 = io_ins_1 | io_ins_2; // @[StickySelects.scala 22:54:@5823.4]
  assign _T_21 = _T_20 | io_ins_3; // @[StickySelects.scala 22:54:@5824.4]
  assign _T_22 = _T_21 | io_ins_4; // @[StickySelects.scala 22:54:@5825.4]
  assign _T_23 = _T_22 | io_ins_5; // @[StickySelects.scala 22:54:@5826.4]
  assign _T_24 = _T_23 | io_ins_6; // @[StickySelects.scala 22:54:@5827.4]
  assign _T_25 = _T_24 | io_ins_7; // @[StickySelects.scala 22:54:@5828.4]
  assign _T_26 = _T_25 | io_ins_8; // @[StickySelects.scala 22:54:@5829.4]
  assign _T_28 = io_ins_0 | _T_19; // @[StickySelects.scala 24:52:@5830.4]
  assign _T_29 = _T_26 ? 1'h0 : _T_28; // @[StickySelects.scala 24:21:@5831.4]
  assign _T_33 = io_ins_0 | io_ins_2; // @[StickySelects.scala 22:54:@5834.4]
  assign _T_34 = _T_33 | io_ins_3; // @[StickySelects.scala 22:54:@5835.4]
  assign _T_35 = _T_34 | io_ins_4; // @[StickySelects.scala 22:54:@5836.4]
  assign _T_36 = _T_35 | io_ins_5; // @[StickySelects.scala 22:54:@5837.4]
  assign _T_37 = _T_36 | io_ins_6; // @[StickySelects.scala 22:54:@5838.4]
  assign _T_38 = _T_37 | io_ins_7; // @[StickySelects.scala 22:54:@5839.4]
  assign _T_39 = _T_38 | io_ins_8; // @[StickySelects.scala 22:54:@5840.4]
  assign _T_41 = io_ins_1 | _T_32; // @[StickySelects.scala 24:52:@5841.4]
  assign _T_42 = _T_39 ? 1'h0 : _T_41; // @[StickySelects.scala 24:21:@5842.4]
  assign _T_46 = io_ins_0 | io_ins_1; // @[StickySelects.scala 22:54:@5845.4]
  assign _T_47 = _T_46 | io_ins_3; // @[StickySelects.scala 22:54:@5846.4]
  assign _T_48 = _T_47 | io_ins_4; // @[StickySelects.scala 22:54:@5847.4]
  assign _T_49 = _T_48 | io_ins_5; // @[StickySelects.scala 22:54:@5848.4]
  assign _T_50 = _T_49 | io_ins_6; // @[StickySelects.scala 22:54:@5849.4]
  assign _T_51 = _T_50 | io_ins_7; // @[StickySelects.scala 22:54:@5850.4]
  assign _T_52 = _T_51 | io_ins_8; // @[StickySelects.scala 22:54:@5851.4]
  assign _T_54 = io_ins_2 | _T_45; // @[StickySelects.scala 24:52:@5852.4]
  assign _T_55 = _T_52 ? 1'h0 : _T_54; // @[StickySelects.scala 24:21:@5853.4]
  assign _T_60 = _T_46 | io_ins_2; // @[StickySelects.scala 22:54:@5857.4]
  assign _T_61 = _T_60 | io_ins_4; // @[StickySelects.scala 22:54:@5858.4]
  assign _T_62 = _T_61 | io_ins_5; // @[StickySelects.scala 22:54:@5859.4]
  assign _T_63 = _T_62 | io_ins_6; // @[StickySelects.scala 22:54:@5860.4]
  assign _T_64 = _T_63 | io_ins_7; // @[StickySelects.scala 22:54:@5861.4]
  assign _T_65 = _T_64 | io_ins_8; // @[StickySelects.scala 22:54:@5862.4]
  assign _T_67 = io_ins_3 | _T_58; // @[StickySelects.scala 24:52:@5863.4]
  assign _T_68 = _T_65 ? 1'h0 : _T_67; // @[StickySelects.scala 24:21:@5864.4]
  assign _T_74 = _T_60 | io_ins_3; // @[StickySelects.scala 22:54:@5869.4]
  assign _T_75 = _T_74 | io_ins_5; // @[StickySelects.scala 22:54:@5870.4]
  assign _T_76 = _T_75 | io_ins_6; // @[StickySelects.scala 22:54:@5871.4]
  assign _T_77 = _T_76 | io_ins_7; // @[StickySelects.scala 22:54:@5872.4]
  assign _T_78 = _T_77 | io_ins_8; // @[StickySelects.scala 22:54:@5873.4]
  assign _T_80 = io_ins_4 | _T_71; // @[StickySelects.scala 24:52:@5874.4]
  assign _T_81 = _T_78 ? 1'h0 : _T_80; // @[StickySelects.scala 24:21:@5875.4]
  assign _T_88 = _T_74 | io_ins_4; // @[StickySelects.scala 22:54:@5881.4]
  assign _T_89 = _T_88 | io_ins_6; // @[StickySelects.scala 22:54:@5882.4]
  assign _T_90 = _T_89 | io_ins_7; // @[StickySelects.scala 22:54:@5883.4]
  assign _T_91 = _T_90 | io_ins_8; // @[StickySelects.scala 22:54:@5884.4]
  assign _T_93 = io_ins_5 | _T_84; // @[StickySelects.scala 24:52:@5885.4]
  assign _T_94 = _T_91 ? 1'h0 : _T_93; // @[StickySelects.scala 24:21:@5886.4]
  assign _T_102 = _T_88 | io_ins_5; // @[StickySelects.scala 22:54:@5893.4]
  assign _T_103 = _T_102 | io_ins_7; // @[StickySelects.scala 22:54:@5894.4]
  assign _T_104 = _T_103 | io_ins_8; // @[StickySelects.scala 22:54:@5895.4]
  assign _T_106 = io_ins_6 | _T_97; // @[StickySelects.scala 24:52:@5896.4]
  assign _T_107 = _T_104 ? 1'h0 : _T_106; // @[StickySelects.scala 24:21:@5897.4]
  assign _T_116 = _T_102 | io_ins_6; // @[StickySelects.scala 22:54:@5905.4]
  assign _T_117 = _T_116 | io_ins_8; // @[StickySelects.scala 22:54:@5906.4]
  assign _T_119 = io_ins_7 | _T_110; // @[StickySelects.scala 24:52:@5907.4]
  assign _T_120 = _T_117 ? 1'h0 : _T_119; // @[StickySelects.scala 24:21:@5908.4]
  assign _T_130 = _T_116 | io_ins_7; // @[StickySelects.scala 22:54:@5917.4]
  assign _T_132 = io_ins_8 | _T_123; // @[StickySelects.scala 24:52:@5918.4]
  assign _T_133 = _T_130 ? 1'h0 : _T_132; // @[StickySelects.scala 24:21:@5919.4]
  assign io_outs_0 = _T_26 ? 1'h0 : _T_28; // @[StickySelects.scala 28:52:@5921.4]
  assign io_outs_1 = _T_39 ? 1'h0 : _T_41; // @[StickySelects.scala 28:52:@5922.4]
  assign io_outs_2 = _T_52 ? 1'h0 : _T_54; // @[StickySelects.scala 28:52:@5923.4]
  assign io_outs_3 = _T_65 ? 1'h0 : _T_67; // @[StickySelects.scala 28:52:@5924.4]
  assign io_outs_4 = _T_78 ? 1'h0 : _T_80; // @[StickySelects.scala 28:52:@5925.4]
  assign io_outs_5 = _T_91 ? 1'h0 : _T_93; // @[StickySelects.scala 28:52:@5926.4]
  assign io_outs_6 = _T_104 ? 1'h0 : _T_106; // @[StickySelects.scala 28:52:@5927.4]
  assign io_outs_7 = _T_117 ? 1'h0 : _T_119; // @[StickySelects.scala 28:52:@5928.4]
  assign io_outs_8 = _T_130 ? 1'h0 : _T_132; // @[StickySelects.scala 28:52:@5929.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_32 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_45 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_58 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_71 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_84 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_97 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_110 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_123 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (_T_26) begin
        _T_19 <= 1'h0;
      end else begin
        _T_19 <= _T_28;
      end
    end
    if (reset) begin
      _T_32 <= 1'h0;
    end else begin
      if (_T_39) begin
        _T_32 <= 1'h0;
      end else begin
        _T_32 <= _T_41;
      end
    end
    if (reset) begin
      _T_45 <= 1'h0;
    end else begin
      if (_T_52) begin
        _T_45 <= 1'h0;
      end else begin
        _T_45 <= _T_54;
      end
    end
    if (reset) begin
      _T_58 <= 1'h0;
    end else begin
      if (_T_65) begin
        _T_58 <= 1'h0;
      end else begin
        _T_58 <= _T_67;
      end
    end
    if (reset) begin
      _T_71 <= 1'h0;
    end else begin
      if (_T_78) begin
        _T_71 <= 1'h0;
      end else begin
        _T_71 <= _T_80;
      end
    end
    if (reset) begin
      _T_84 <= 1'h0;
    end else begin
      if (_T_91) begin
        _T_84 <= 1'h0;
      end else begin
        _T_84 <= _T_93;
      end
    end
    if (reset) begin
      _T_97 <= 1'h0;
    end else begin
      if (_T_104) begin
        _T_97 <= 1'h0;
      end else begin
        _T_97 <= _T_106;
      end
    end
    if (reset) begin
      _T_110 <= 1'h0;
    end else begin
      if (_T_117) begin
        _T_110 <= 1'h0;
      end else begin
        _T_110 <= _T_119;
      end
    end
    if (reset) begin
      _T_123 <= 1'h0;
    end else begin
      if (_T_130) begin
        _T_123 <= 1'h0;
      end else begin
        _T_123 <= _T_132;
      end
    end
  end
endmodule
module RetimeWrapper_44( // @[:@8565.2]
  input   clock, // @[:@8566.4]
  input   reset, // @[:@8567.4]
  input   io_flow, // @[:@8568.4]
  input   io_in, // @[:@8568.4]
  output  io_out // @[:@8568.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@8570.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@8570.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@8570.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@8570.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@8570.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@8570.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@8570.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@8583.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@8582.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@8581.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@8580.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@8579.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@8577.4]
endmodule
module x329_lb_0( // @[:@15465.2]
  input        clock, // @[:@15466.4]
  input        reset, // @[:@15467.4]
  input  [2:0] io_rPort_17_banks_1, // @[:@15468.4]
  input  [2:0] io_rPort_17_banks_0, // @[:@15468.4]
  input  [7:0] io_rPort_17_ofs_0, // @[:@15468.4]
  input        io_rPort_17_en_0, // @[:@15468.4]
  input        io_rPort_17_backpressure, // @[:@15468.4]
  output [7:0] io_rPort_17_output_0, // @[:@15468.4]
  input  [2:0] io_rPort_16_banks_1, // @[:@15468.4]
  input  [2:0] io_rPort_16_banks_0, // @[:@15468.4]
  input  [7:0] io_rPort_16_ofs_0, // @[:@15468.4]
  input        io_rPort_16_en_0, // @[:@15468.4]
  input        io_rPort_16_backpressure, // @[:@15468.4]
  output [7:0] io_rPort_16_output_0, // @[:@15468.4]
  input  [2:0] io_rPort_15_banks_1, // @[:@15468.4]
  input  [2:0] io_rPort_15_banks_0, // @[:@15468.4]
  input  [7:0] io_rPort_15_ofs_0, // @[:@15468.4]
  input        io_rPort_15_en_0, // @[:@15468.4]
  input        io_rPort_15_backpressure, // @[:@15468.4]
  output [7:0] io_rPort_15_output_0, // @[:@15468.4]
  input  [2:0] io_rPort_14_banks_1, // @[:@15468.4]
  input  [2:0] io_rPort_14_banks_0, // @[:@15468.4]
  input  [7:0] io_rPort_14_ofs_0, // @[:@15468.4]
  input        io_rPort_14_en_0, // @[:@15468.4]
  input        io_rPort_14_backpressure, // @[:@15468.4]
  output [7:0] io_rPort_14_output_0, // @[:@15468.4]
  input  [2:0] io_rPort_13_banks_1, // @[:@15468.4]
  input  [2:0] io_rPort_13_banks_0, // @[:@15468.4]
  input  [7:0] io_rPort_13_ofs_0, // @[:@15468.4]
  input        io_rPort_13_en_0, // @[:@15468.4]
  input        io_rPort_13_backpressure, // @[:@15468.4]
  output [7:0] io_rPort_13_output_0, // @[:@15468.4]
  input  [2:0] io_rPort_12_banks_1, // @[:@15468.4]
  input  [2:0] io_rPort_12_banks_0, // @[:@15468.4]
  input  [7:0] io_rPort_12_ofs_0, // @[:@15468.4]
  input        io_rPort_12_en_0, // @[:@15468.4]
  input        io_rPort_12_backpressure, // @[:@15468.4]
  output [7:0] io_rPort_12_output_0, // @[:@15468.4]
  input  [2:0] io_rPort_11_banks_1, // @[:@15468.4]
  input  [2:0] io_rPort_11_banks_0, // @[:@15468.4]
  input  [7:0] io_rPort_11_ofs_0, // @[:@15468.4]
  input        io_rPort_11_en_0, // @[:@15468.4]
  input        io_rPort_11_backpressure, // @[:@15468.4]
  output [7:0] io_rPort_11_output_0, // @[:@15468.4]
  input  [2:0] io_rPort_10_banks_1, // @[:@15468.4]
  input  [2:0] io_rPort_10_banks_0, // @[:@15468.4]
  input  [7:0] io_rPort_10_ofs_0, // @[:@15468.4]
  input        io_rPort_10_en_0, // @[:@15468.4]
  input        io_rPort_10_backpressure, // @[:@15468.4]
  output [7:0] io_rPort_10_output_0, // @[:@15468.4]
  input  [2:0] io_rPort_9_banks_1, // @[:@15468.4]
  input  [2:0] io_rPort_9_banks_0, // @[:@15468.4]
  input  [7:0] io_rPort_9_ofs_0, // @[:@15468.4]
  input        io_rPort_9_en_0, // @[:@15468.4]
  input        io_rPort_9_backpressure, // @[:@15468.4]
  output [7:0] io_rPort_9_output_0, // @[:@15468.4]
  input  [2:0] io_rPort_8_banks_1, // @[:@15468.4]
  input  [2:0] io_rPort_8_banks_0, // @[:@15468.4]
  input  [7:0] io_rPort_8_ofs_0, // @[:@15468.4]
  input        io_rPort_8_en_0, // @[:@15468.4]
  input        io_rPort_8_backpressure, // @[:@15468.4]
  output [7:0] io_rPort_8_output_0, // @[:@15468.4]
  input  [2:0] io_rPort_7_banks_1, // @[:@15468.4]
  input  [2:0] io_rPort_7_banks_0, // @[:@15468.4]
  input  [7:0] io_rPort_7_ofs_0, // @[:@15468.4]
  input        io_rPort_7_en_0, // @[:@15468.4]
  input        io_rPort_7_backpressure, // @[:@15468.4]
  output [7:0] io_rPort_7_output_0, // @[:@15468.4]
  input  [2:0] io_rPort_6_banks_1, // @[:@15468.4]
  input  [2:0] io_rPort_6_banks_0, // @[:@15468.4]
  input  [7:0] io_rPort_6_ofs_0, // @[:@15468.4]
  input        io_rPort_6_en_0, // @[:@15468.4]
  input        io_rPort_6_backpressure, // @[:@15468.4]
  output [7:0] io_rPort_6_output_0, // @[:@15468.4]
  input  [2:0] io_rPort_5_banks_1, // @[:@15468.4]
  input  [2:0] io_rPort_5_banks_0, // @[:@15468.4]
  input  [7:0] io_rPort_5_ofs_0, // @[:@15468.4]
  input        io_rPort_5_en_0, // @[:@15468.4]
  input        io_rPort_5_backpressure, // @[:@15468.4]
  output [7:0] io_rPort_5_output_0, // @[:@15468.4]
  input  [2:0] io_rPort_4_banks_1, // @[:@15468.4]
  input  [2:0] io_rPort_4_banks_0, // @[:@15468.4]
  input  [7:0] io_rPort_4_ofs_0, // @[:@15468.4]
  input        io_rPort_4_en_0, // @[:@15468.4]
  input        io_rPort_4_backpressure, // @[:@15468.4]
  output [7:0] io_rPort_4_output_0, // @[:@15468.4]
  input  [2:0] io_rPort_3_banks_1, // @[:@15468.4]
  input  [2:0] io_rPort_3_banks_0, // @[:@15468.4]
  input  [7:0] io_rPort_3_ofs_0, // @[:@15468.4]
  input        io_rPort_3_en_0, // @[:@15468.4]
  input        io_rPort_3_backpressure, // @[:@15468.4]
  output [7:0] io_rPort_3_output_0, // @[:@15468.4]
  input  [2:0] io_rPort_2_banks_1, // @[:@15468.4]
  input  [2:0] io_rPort_2_banks_0, // @[:@15468.4]
  input  [7:0] io_rPort_2_ofs_0, // @[:@15468.4]
  input        io_rPort_2_en_0, // @[:@15468.4]
  input        io_rPort_2_backpressure, // @[:@15468.4]
  output [7:0] io_rPort_2_output_0, // @[:@15468.4]
  input  [2:0] io_rPort_1_banks_1, // @[:@15468.4]
  input  [2:0] io_rPort_1_banks_0, // @[:@15468.4]
  input  [7:0] io_rPort_1_ofs_0, // @[:@15468.4]
  input        io_rPort_1_en_0, // @[:@15468.4]
  input        io_rPort_1_backpressure, // @[:@15468.4]
  output [7:0] io_rPort_1_output_0, // @[:@15468.4]
  input  [2:0] io_rPort_0_banks_1, // @[:@15468.4]
  input  [2:0] io_rPort_0_banks_0, // @[:@15468.4]
  input  [7:0] io_rPort_0_ofs_0, // @[:@15468.4]
  input        io_rPort_0_en_0, // @[:@15468.4]
  input        io_rPort_0_backpressure, // @[:@15468.4]
  output [7:0] io_rPort_0_output_0, // @[:@15468.4]
  input  [2:0] io_wPort_3_banks_1, // @[:@15468.4]
  input  [2:0] io_wPort_3_banks_0, // @[:@15468.4]
  input  [7:0] io_wPort_3_ofs_0, // @[:@15468.4]
  input  [7:0] io_wPort_3_data_0, // @[:@15468.4]
  input        io_wPort_3_en_0, // @[:@15468.4]
  input  [2:0] io_wPort_2_banks_1, // @[:@15468.4]
  input  [2:0] io_wPort_2_banks_0, // @[:@15468.4]
  input  [7:0] io_wPort_2_ofs_0, // @[:@15468.4]
  input  [7:0] io_wPort_2_data_0, // @[:@15468.4]
  input        io_wPort_2_en_0, // @[:@15468.4]
  input  [2:0] io_wPort_1_banks_1, // @[:@15468.4]
  input  [2:0] io_wPort_1_banks_0, // @[:@15468.4]
  input  [7:0] io_wPort_1_ofs_0, // @[:@15468.4]
  input  [7:0] io_wPort_1_data_0, // @[:@15468.4]
  input        io_wPort_1_en_0, // @[:@15468.4]
  input  [2:0] io_wPort_0_banks_1, // @[:@15468.4]
  input  [2:0] io_wPort_0_banks_0, // @[:@15468.4]
  input  [7:0] io_wPort_0_ofs_0, // @[:@15468.4]
  input  [7:0] io_wPort_0_data_0, // @[:@15468.4]
  input        io_wPort_0_en_0 // @[:@15468.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@15611.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@15611.4]
  wire [7:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15611.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15611.4]
  wire [7:0] Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15611.4]
  wire [7:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@15611.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@15611.4]
  wire [7:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@15611.4]
  wire  Mem1D_1_clock; // @[MemPrimitives.scala 64:21:@15627.4]
  wire  Mem1D_1_reset; // @[MemPrimitives.scala 64:21:@15627.4]
  wire [7:0] Mem1D_1_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15627.4]
  wire  Mem1D_1_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15627.4]
  wire [7:0] Mem1D_1_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15627.4]
  wire [7:0] Mem1D_1_io_w_data_0; // @[MemPrimitives.scala 64:21:@15627.4]
  wire  Mem1D_1_io_w_en_0; // @[MemPrimitives.scala 64:21:@15627.4]
  wire [7:0] Mem1D_1_io_output; // @[MemPrimitives.scala 64:21:@15627.4]
  wire  Mem1D_2_clock; // @[MemPrimitives.scala 64:21:@15643.4]
  wire  Mem1D_2_reset; // @[MemPrimitives.scala 64:21:@15643.4]
  wire [7:0] Mem1D_2_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15643.4]
  wire  Mem1D_2_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15643.4]
  wire [7:0] Mem1D_2_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15643.4]
  wire [7:0] Mem1D_2_io_w_data_0; // @[MemPrimitives.scala 64:21:@15643.4]
  wire  Mem1D_2_io_w_en_0; // @[MemPrimitives.scala 64:21:@15643.4]
  wire [7:0] Mem1D_2_io_output; // @[MemPrimitives.scala 64:21:@15643.4]
  wire  Mem1D_3_clock; // @[MemPrimitives.scala 64:21:@15659.4]
  wire  Mem1D_3_reset; // @[MemPrimitives.scala 64:21:@15659.4]
  wire [7:0] Mem1D_3_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15659.4]
  wire  Mem1D_3_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15659.4]
  wire [7:0] Mem1D_3_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15659.4]
  wire [7:0] Mem1D_3_io_w_data_0; // @[MemPrimitives.scala 64:21:@15659.4]
  wire  Mem1D_3_io_w_en_0; // @[MemPrimitives.scala 64:21:@15659.4]
  wire [7:0] Mem1D_3_io_output; // @[MemPrimitives.scala 64:21:@15659.4]
  wire  Mem1D_4_clock; // @[MemPrimitives.scala 64:21:@15675.4]
  wire  Mem1D_4_reset; // @[MemPrimitives.scala 64:21:@15675.4]
  wire [7:0] Mem1D_4_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15675.4]
  wire  Mem1D_4_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15675.4]
  wire [7:0] Mem1D_4_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15675.4]
  wire [7:0] Mem1D_4_io_w_data_0; // @[MemPrimitives.scala 64:21:@15675.4]
  wire  Mem1D_4_io_w_en_0; // @[MemPrimitives.scala 64:21:@15675.4]
  wire [7:0] Mem1D_4_io_output; // @[MemPrimitives.scala 64:21:@15675.4]
  wire  Mem1D_5_clock; // @[MemPrimitives.scala 64:21:@15691.4]
  wire  Mem1D_5_reset; // @[MemPrimitives.scala 64:21:@15691.4]
  wire [7:0] Mem1D_5_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15691.4]
  wire  Mem1D_5_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15691.4]
  wire [7:0] Mem1D_5_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15691.4]
  wire [7:0] Mem1D_5_io_w_data_0; // @[MemPrimitives.scala 64:21:@15691.4]
  wire  Mem1D_5_io_w_en_0; // @[MemPrimitives.scala 64:21:@15691.4]
  wire [7:0] Mem1D_5_io_output; // @[MemPrimitives.scala 64:21:@15691.4]
  wire  Mem1D_6_clock; // @[MemPrimitives.scala 64:21:@15707.4]
  wire  Mem1D_6_reset; // @[MemPrimitives.scala 64:21:@15707.4]
  wire [7:0] Mem1D_6_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15707.4]
  wire  Mem1D_6_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15707.4]
  wire [7:0] Mem1D_6_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15707.4]
  wire [7:0] Mem1D_6_io_w_data_0; // @[MemPrimitives.scala 64:21:@15707.4]
  wire  Mem1D_6_io_w_en_0; // @[MemPrimitives.scala 64:21:@15707.4]
  wire [7:0] Mem1D_6_io_output; // @[MemPrimitives.scala 64:21:@15707.4]
  wire  Mem1D_7_clock; // @[MemPrimitives.scala 64:21:@15723.4]
  wire  Mem1D_7_reset; // @[MemPrimitives.scala 64:21:@15723.4]
  wire [7:0] Mem1D_7_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15723.4]
  wire  Mem1D_7_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15723.4]
  wire [7:0] Mem1D_7_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15723.4]
  wire [7:0] Mem1D_7_io_w_data_0; // @[MemPrimitives.scala 64:21:@15723.4]
  wire  Mem1D_7_io_w_en_0; // @[MemPrimitives.scala 64:21:@15723.4]
  wire [7:0] Mem1D_7_io_output; // @[MemPrimitives.scala 64:21:@15723.4]
  wire  Mem1D_8_clock; // @[MemPrimitives.scala 64:21:@15739.4]
  wire  Mem1D_8_reset; // @[MemPrimitives.scala 64:21:@15739.4]
  wire [7:0] Mem1D_8_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15739.4]
  wire  Mem1D_8_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15739.4]
  wire [7:0] Mem1D_8_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15739.4]
  wire [7:0] Mem1D_8_io_w_data_0; // @[MemPrimitives.scala 64:21:@15739.4]
  wire  Mem1D_8_io_w_en_0; // @[MemPrimitives.scala 64:21:@15739.4]
  wire [7:0] Mem1D_8_io_output; // @[MemPrimitives.scala 64:21:@15739.4]
  wire  Mem1D_9_clock; // @[MemPrimitives.scala 64:21:@15755.4]
  wire  Mem1D_9_reset; // @[MemPrimitives.scala 64:21:@15755.4]
  wire [7:0] Mem1D_9_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15755.4]
  wire  Mem1D_9_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15755.4]
  wire [7:0] Mem1D_9_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15755.4]
  wire [7:0] Mem1D_9_io_w_data_0; // @[MemPrimitives.scala 64:21:@15755.4]
  wire  Mem1D_9_io_w_en_0; // @[MemPrimitives.scala 64:21:@15755.4]
  wire [7:0] Mem1D_9_io_output; // @[MemPrimitives.scala 64:21:@15755.4]
  wire  Mem1D_10_clock; // @[MemPrimitives.scala 64:21:@15771.4]
  wire  Mem1D_10_reset; // @[MemPrimitives.scala 64:21:@15771.4]
  wire [7:0] Mem1D_10_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15771.4]
  wire  Mem1D_10_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15771.4]
  wire [7:0] Mem1D_10_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15771.4]
  wire [7:0] Mem1D_10_io_w_data_0; // @[MemPrimitives.scala 64:21:@15771.4]
  wire  Mem1D_10_io_w_en_0; // @[MemPrimitives.scala 64:21:@15771.4]
  wire [7:0] Mem1D_10_io_output; // @[MemPrimitives.scala 64:21:@15771.4]
  wire  Mem1D_11_clock; // @[MemPrimitives.scala 64:21:@15787.4]
  wire  Mem1D_11_reset; // @[MemPrimitives.scala 64:21:@15787.4]
  wire [7:0] Mem1D_11_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15787.4]
  wire  Mem1D_11_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15787.4]
  wire [7:0] Mem1D_11_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15787.4]
  wire [7:0] Mem1D_11_io_w_data_0; // @[MemPrimitives.scala 64:21:@15787.4]
  wire  Mem1D_11_io_w_en_0; // @[MemPrimitives.scala 64:21:@15787.4]
  wire [7:0] Mem1D_11_io_output; // @[MemPrimitives.scala 64:21:@15787.4]
  wire  Mem1D_12_clock; // @[MemPrimitives.scala 64:21:@15803.4]
  wire  Mem1D_12_reset; // @[MemPrimitives.scala 64:21:@15803.4]
  wire [7:0] Mem1D_12_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15803.4]
  wire  Mem1D_12_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15803.4]
  wire [7:0] Mem1D_12_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15803.4]
  wire [7:0] Mem1D_12_io_w_data_0; // @[MemPrimitives.scala 64:21:@15803.4]
  wire  Mem1D_12_io_w_en_0; // @[MemPrimitives.scala 64:21:@15803.4]
  wire [7:0] Mem1D_12_io_output; // @[MemPrimitives.scala 64:21:@15803.4]
  wire  Mem1D_13_clock; // @[MemPrimitives.scala 64:21:@15819.4]
  wire  Mem1D_13_reset; // @[MemPrimitives.scala 64:21:@15819.4]
  wire [7:0] Mem1D_13_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15819.4]
  wire  Mem1D_13_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15819.4]
  wire [7:0] Mem1D_13_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15819.4]
  wire [7:0] Mem1D_13_io_w_data_0; // @[MemPrimitives.scala 64:21:@15819.4]
  wire  Mem1D_13_io_w_en_0; // @[MemPrimitives.scala 64:21:@15819.4]
  wire [7:0] Mem1D_13_io_output; // @[MemPrimitives.scala 64:21:@15819.4]
  wire  Mem1D_14_clock; // @[MemPrimitives.scala 64:21:@15835.4]
  wire  Mem1D_14_reset; // @[MemPrimitives.scala 64:21:@15835.4]
  wire [7:0] Mem1D_14_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15835.4]
  wire  Mem1D_14_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15835.4]
  wire [7:0] Mem1D_14_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15835.4]
  wire [7:0] Mem1D_14_io_w_data_0; // @[MemPrimitives.scala 64:21:@15835.4]
  wire  Mem1D_14_io_w_en_0; // @[MemPrimitives.scala 64:21:@15835.4]
  wire [7:0] Mem1D_14_io_output; // @[MemPrimitives.scala 64:21:@15835.4]
  wire  Mem1D_15_clock; // @[MemPrimitives.scala 64:21:@15851.4]
  wire  Mem1D_15_reset; // @[MemPrimitives.scala 64:21:@15851.4]
  wire [7:0] Mem1D_15_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15851.4]
  wire  Mem1D_15_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15851.4]
  wire [7:0] Mem1D_15_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15851.4]
  wire [7:0] Mem1D_15_io_w_data_0; // @[MemPrimitives.scala 64:21:@15851.4]
  wire  Mem1D_15_io_w_en_0; // @[MemPrimitives.scala 64:21:@15851.4]
  wire [7:0] Mem1D_15_io_output; // @[MemPrimitives.scala 64:21:@15851.4]
  wire  Mem1D_16_clock; // @[MemPrimitives.scala 64:21:@15867.4]
  wire  Mem1D_16_reset; // @[MemPrimitives.scala 64:21:@15867.4]
  wire [7:0] Mem1D_16_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15867.4]
  wire  Mem1D_16_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15867.4]
  wire [7:0] Mem1D_16_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15867.4]
  wire [7:0] Mem1D_16_io_w_data_0; // @[MemPrimitives.scala 64:21:@15867.4]
  wire  Mem1D_16_io_w_en_0; // @[MemPrimitives.scala 64:21:@15867.4]
  wire [7:0] Mem1D_16_io_output; // @[MemPrimitives.scala 64:21:@15867.4]
  wire  Mem1D_17_clock; // @[MemPrimitives.scala 64:21:@15883.4]
  wire  Mem1D_17_reset; // @[MemPrimitives.scala 64:21:@15883.4]
  wire [7:0] Mem1D_17_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15883.4]
  wire  Mem1D_17_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15883.4]
  wire [7:0] Mem1D_17_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15883.4]
  wire [7:0] Mem1D_17_io_w_data_0; // @[MemPrimitives.scala 64:21:@15883.4]
  wire  Mem1D_17_io_w_en_0; // @[MemPrimitives.scala 64:21:@15883.4]
  wire [7:0] Mem1D_17_io_output; // @[MemPrimitives.scala 64:21:@15883.4]
  wire  Mem1D_18_clock; // @[MemPrimitives.scala 64:21:@15899.4]
  wire  Mem1D_18_reset; // @[MemPrimitives.scala 64:21:@15899.4]
  wire [7:0] Mem1D_18_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15899.4]
  wire  Mem1D_18_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15899.4]
  wire [7:0] Mem1D_18_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15899.4]
  wire [7:0] Mem1D_18_io_w_data_0; // @[MemPrimitives.scala 64:21:@15899.4]
  wire  Mem1D_18_io_w_en_0; // @[MemPrimitives.scala 64:21:@15899.4]
  wire [7:0] Mem1D_18_io_output; // @[MemPrimitives.scala 64:21:@15899.4]
  wire  Mem1D_19_clock; // @[MemPrimitives.scala 64:21:@15915.4]
  wire  Mem1D_19_reset; // @[MemPrimitives.scala 64:21:@15915.4]
  wire [7:0] Mem1D_19_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15915.4]
  wire  Mem1D_19_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15915.4]
  wire [7:0] Mem1D_19_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15915.4]
  wire [7:0] Mem1D_19_io_w_data_0; // @[MemPrimitives.scala 64:21:@15915.4]
  wire  Mem1D_19_io_w_en_0; // @[MemPrimitives.scala 64:21:@15915.4]
  wire [7:0] Mem1D_19_io_output; // @[MemPrimitives.scala 64:21:@15915.4]
  wire  Mem1D_20_clock; // @[MemPrimitives.scala 64:21:@15931.4]
  wire  Mem1D_20_reset; // @[MemPrimitives.scala 64:21:@15931.4]
  wire [7:0] Mem1D_20_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15931.4]
  wire  Mem1D_20_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15931.4]
  wire [7:0] Mem1D_20_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15931.4]
  wire [7:0] Mem1D_20_io_w_data_0; // @[MemPrimitives.scala 64:21:@15931.4]
  wire  Mem1D_20_io_w_en_0; // @[MemPrimitives.scala 64:21:@15931.4]
  wire [7:0] Mem1D_20_io_output; // @[MemPrimitives.scala 64:21:@15931.4]
  wire  Mem1D_21_clock; // @[MemPrimitives.scala 64:21:@15947.4]
  wire  Mem1D_21_reset; // @[MemPrimitives.scala 64:21:@15947.4]
  wire [7:0] Mem1D_21_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15947.4]
  wire  Mem1D_21_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15947.4]
  wire [7:0] Mem1D_21_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15947.4]
  wire [7:0] Mem1D_21_io_w_data_0; // @[MemPrimitives.scala 64:21:@15947.4]
  wire  Mem1D_21_io_w_en_0; // @[MemPrimitives.scala 64:21:@15947.4]
  wire [7:0] Mem1D_21_io_output; // @[MemPrimitives.scala 64:21:@15947.4]
  wire  Mem1D_22_clock; // @[MemPrimitives.scala 64:21:@15963.4]
  wire  Mem1D_22_reset; // @[MemPrimitives.scala 64:21:@15963.4]
  wire [7:0] Mem1D_22_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15963.4]
  wire  Mem1D_22_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15963.4]
  wire [7:0] Mem1D_22_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15963.4]
  wire [7:0] Mem1D_22_io_w_data_0; // @[MemPrimitives.scala 64:21:@15963.4]
  wire  Mem1D_22_io_w_en_0; // @[MemPrimitives.scala 64:21:@15963.4]
  wire [7:0] Mem1D_22_io_output; // @[MemPrimitives.scala 64:21:@15963.4]
  wire  Mem1D_23_clock; // @[MemPrimitives.scala 64:21:@15979.4]
  wire  Mem1D_23_reset; // @[MemPrimitives.scala 64:21:@15979.4]
  wire [7:0] Mem1D_23_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15979.4]
  wire  Mem1D_23_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15979.4]
  wire [7:0] Mem1D_23_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15979.4]
  wire [7:0] Mem1D_23_io_w_data_0; // @[MemPrimitives.scala 64:21:@15979.4]
  wire  Mem1D_23_io_w_en_0; // @[MemPrimitives.scala 64:21:@15979.4]
  wire [7:0] Mem1D_23_io_output; // @[MemPrimitives.scala 64:21:@15979.4]
  wire  StickySelects_clock; // @[MemPrimitives.scala 121:29:@16487.4]
  wire  StickySelects_reset; // @[MemPrimitives.scala 121:29:@16487.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 121:29:@16487.4]
  wire  StickySelects_io_ins_1; // @[MemPrimitives.scala 121:29:@16487.4]
  wire  StickySelects_io_ins_2; // @[MemPrimitives.scala 121:29:@16487.4]
  wire  StickySelects_io_ins_3; // @[MemPrimitives.scala 121:29:@16487.4]
  wire  StickySelects_io_ins_4; // @[MemPrimitives.scala 121:29:@16487.4]
  wire  StickySelects_io_ins_5; // @[MemPrimitives.scala 121:29:@16487.4]
  wire  StickySelects_io_ins_6; // @[MemPrimitives.scala 121:29:@16487.4]
  wire  StickySelects_io_ins_7; // @[MemPrimitives.scala 121:29:@16487.4]
  wire  StickySelects_io_ins_8; // @[MemPrimitives.scala 121:29:@16487.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 121:29:@16487.4]
  wire  StickySelects_io_outs_1; // @[MemPrimitives.scala 121:29:@16487.4]
  wire  StickySelects_io_outs_2; // @[MemPrimitives.scala 121:29:@16487.4]
  wire  StickySelects_io_outs_3; // @[MemPrimitives.scala 121:29:@16487.4]
  wire  StickySelects_io_outs_4; // @[MemPrimitives.scala 121:29:@16487.4]
  wire  StickySelects_io_outs_5; // @[MemPrimitives.scala 121:29:@16487.4]
  wire  StickySelects_io_outs_6; // @[MemPrimitives.scala 121:29:@16487.4]
  wire  StickySelects_io_outs_7; // @[MemPrimitives.scala 121:29:@16487.4]
  wire  StickySelects_io_outs_8; // @[MemPrimitives.scala 121:29:@16487.4]
  wire  StickySelects_1_clock; // @[MemPrimitives.scala 121:29:@16576.4]
  wire  StickySelects_1_reset; // @[MemPrimitives.scala 121:29:@16576.4]
  wire  StickySelects_1_io_ins_0; // @[MemPrimitives.scala 121:29:@16576.4]
  wire  StickySelects_1_io_ins_1; // @[MemPrimitives.scala 121:29:@16576.4]
  wire  StickySelects_1_io_ins_2; // @[MemPrimitives.scala 121:29:@16576.4]
  wire  StickySelects_1_io_ins_3; // @[MemPrimitives.scala 121:29:@16576.4]
  wire  StickySelects_1_io_ins_4; // @[MemPrimitives.scala 121:29:@16576.4]
  wire  StickySelects_1_io_ins_5; // @[MemPrimitives.scala 121:29:@16576.4]
  wire  StickySelects_1_io_ins_6; // @[MemPrimitives.scala 121:29:@16576.4]
  wire  StickySelects_1_io_ins_7; // @[MemPrimitives.scala 121:29:@16576.4]
  wire  StickySelects_1_io_ins_8; // @[MemPrimitives.scala 121:29:@16576.4]
  wire  StickySelects_1_io_outs_0; // @[MemPrimitives.scala 121:29:@16576.4]
  wire  StickySelects_1_io_outs_1; // @[MemPrimitives.scala 121:29:@16576.4]
  wire  StickySelects_1_io_outs_2; // @[MemPrimitives.scala 121:29:@16576.4]
  wire  StickySelects_1_io_outs_3; // @[MemPrimitives.scala 121:29:@16576.4]
  wire  StickySelects_1_io_outs_4; // @[MemPrimitives.scala 121:29:@16576.4]
  wire  StickySelects_1_io_outs_5; // @[MemPrimitives.scala 121:29:@16576.4]
  wire  StickySelects_1_io_outs_6; // @[MemPrimitives.scala 121:29:@16576.4]
  wire  StickySelects_1_io_outs_7; // @[MemPrimitives.scala 121:29:@16576.4]
  wire  StickySelects_1_io_outs_8; // @[MemPrimitives.scala 121:29:@16576.4]
  wire  StickySelects_2_clock; // @[MemPrimitives.scala 121:29:@16665.4]
  wire  StickySelects_2_reset; // @[MemPrimitives.scala 121:29:@16665.4]
  wire  StickySelects_2_io_ins_0; // @[MemPrimitives.scala 121:29:@16665.4]
  wire  StickySelects_2_io_ins_1; // @[MemPrimitives.scala 121:29:@16665.4]
  wire  StickySelects_2_io_ins_2; // @[MemPrimitives.scala 121:29:@16665.4]
  wire  StickySelects_2_io_ins_3; // @[MemPrimitives.scala 121:29:@16665.4]
  wire  StickySelects_2_io_ins_4; // @[MemPrimitives.scala 121:29:@16665.4]
  wire  StickySelects_2_io_ins_5; // @[MemPrimitives.scala 121:29:@16665.4]
  wire  StickySelects_2_io_ins_6; // @[MemPrimitives.scala 121:29:@16665.4]
  wire  StickySelects_2_io_ins_7; // @[MemPrimitives.scala 121:29:@16665.4]
  wire  StickySelects_2_io_ins_8; // @[MemPrimitives.scala 121:29:@16665.4]
  wire  StickySelects_2_io_outs_0; // @[MemPrimitives.scala 121:29:@16665.4]
  wire  StickySelects_2_io_outs_1; // @[MemPrimitives.scala 121:29:@16665.4]
  wire  StickySelects_2_io_outs_2; // @[MemPrimitives.scala 121:29:@16665.4]
  wire  StickySelects_2_io_outs_3; // @[MemPrimitives.scala 121:29:@16665.4]
  wire  StickySelects_2_io_outs_4; // @[MemPrimitives.scala 121:29:@16665.4]
  wire  StickySelects_2_io_outs_5; // @[MemPrimitives.scala 121:29:@16665.4]
  wire  StickySelects_2_io_outs_6; // @[MemPrimitives.scala 121:29:@16665.4]
  wire  StickySelects_2_io_outs_7; // @[MemPrimitives.scala 121:29:@16665.4]
  wire  StickySelects_2_io_outs_8; // @[MemPrimitives.scala 121:29:@16665.4]
  wire  StickySelects_3_clock; // @[MemPrimitives.scala 121:29:@16754.4]
  wire  StickySelects_3_reset; // @[MemPrimitives.scala 121:29:@16754.4]
  wire  StickySelects_3_io_ins_0; // @[MemPrimitives.scala 121:29:@16754.4]
  wire  StickySelects_3_io_ins_1; // @[MemPrimitives.scala 121:29:@16754.4]
  wire  StickySelects_3_io_ins_2; // @[MemPrimitives.scala 121:29:@16754.4]
  wire  StickySelects_3_io_ins_3; // @[MemPrimitives.scala 121:29:@16754.4]
  wire  StickySelects_3_io_ins_4; // @[MemPrimitives.scala 121:29:@16754.4]
  wire  StickySelects_3_io_ins_5; // @[MemPrimitives.scala 121:29:@16754.4]
  wire  StickySelects_3_io_ins_6; // @[MemPrimitives.scala 121:29:@16754.4]
  wire  StickySelects_3_io_ins_7; // @[MemPrimitives.scala 121:29:@16754.4]
  wire  StickySelects_3_io_ins_8; // @[MemPrimitives.scala 121:29:@16754.4]
  wire  StickySelects_3_io_outs_0; // @[MemPrimitives.scala 121:29:@16754.4]
  wire  StickySelects_3_io_outs_1; // @[MemPrimitives.scala 121:29:@16754.4]
  wire  StickySelects_3_io_outs_2; // @[MemPrimitives.scala 121:29:@16754.4]
  wire  StickySelects_3_io_outs_3; // @[MemPrimitives.scala 121:29:@16754.4]
  wire  StickySelects_3_io_outs_4; // @[MemPrimitives.scala 121:29:@16754.4]
  wire  StickySelects_3_io_outs_5; // @[MemPrimitives.scala 121:29:@16754.4]
  wire  StickySelects_3_io_outs_6; // @[MemPrimitives.scala 121:29:@16754.4]
  wire  StickySelects_3_io_outs_7; // @[MemPrimitives.scala 121:29:@16754.4]
  wire  StickySelects_3_io_outs_8; // @[MemPrimitives.scala 121:29:@16754.4]
  wire  StickySelects_4_clock; // @[MemPrimitives.scala 121:29:@16843.4]
  wire  StickySelects_4_reset; // @[MemPrimitives.scala 121:29:@16843.4]
  wire  StickySelects_4_io_ins_0; // @[MemPrimitives.scala 121:29:@16843.4]
  wire  StickySelects_4_io_ins_1; // @[MemPrimitives.scala 121:29:@16843.4]
  wire  StickySelects_4_io_ins_2; // @[MemPrimitives.scala 121:29:@16843.4]
  wire  StickySelects_4_io_ins_3; // @[MemPrimitives.scala 121:29:@16843.4]
  wire  StickySelects_4_io_ins_4; // @[MemPrimitives.scala 121:29:@16843.4]
  wire  StickySelects_4_io_ins_5; // @[MemPrimitives.scala 121:29:@16843.4]
  wire  StickySelects_4_io_ins_6; // @[MemPrimitives.scala 121:29:@16843.4]
  wire  StickySelects_4_io_ins_7; // @[MemPrimitives.scala 121:29:@16843.4]
  wire  StickySelects_4_io_ins_8; // @[MemPrimitives.scala 121:29:@16843.4]
  wire  StickySelects_4_io_outs_0; // @[MemPrimitives.scala 121:29:@16843.4]
  wire  StickySelects_4_io_outs_1; // @[MemPrimitives.scala 121:29:@16843.4]
  wire  StickySelects_4_io_outs_2; // @[MemPrimitives.scala 121:29:@16843.4]
  wire  StickySelects_4_io_outs_3; // @[MemPrimitives.scala 121:29:@16843.4]
  wire  StickySelects_4_io_outs_4; // @[MemPrimitives.scala 121:29:@16843.4]
  wire  StickySelects_4_io_outs_5; // @[MemPrimitives.scala 121:29:@16843.4]
  wire  StickySelects_4_io_outs_6; // @[MemPrimitives.scala 121:29:@16843.4]
  wire  StickySelects_4_io_outs_7; // @[MemPrimitives.scala 121:29:@16843.4]
  wire  StickySelects_4_io_outs_8; // @[MemPrimitives.scala 121:29:@16843.4]
  wire  StickySelects_5_clock; // @[MemPrimitives.scala 121:29:@16932.4]
  wire  StickySelects_5_reset; // @[MemPrimitives.scala 121:29:@16932.4]
  wire  StickySelects_5_io_ins_0; // @[MemPrimitives.scala 121:29:@16932.4]
  wire  StickySelects_5_io_ins_1; // @[MemPrimitives.scala 121:29:@16932.4]
  wire  StickySelects_5_io_ins_2; // @[MemPrimitives.scala 121:29:@16932.4]
  wire  StickySelects_5_io_ins_3; // @[MemPrimitives.scala 121:29:@16932.4]
  wire  StickySelects_5_io_ins_4; // @[MemPrimitives.scala 121:29:@16932.4]
  wire  StickySelects_5_io_ins_5; // @[MemPrimitives.scala 121:29:@16932.4]
  wire  StickySelects_5_io_ins_6; // @[MemPrimitives.scala 121:29:@16932.4]
  wire  StickySelects_5_io_ins_7; // @[MemPrimitives.scala 121:29:@16932.4]
  wire  StickySelects_5_io_ins_8; // @[MemPrimitives.scala 121:29:@16932.4]
  wire  StickySelects_5_io_outs_0; // @[MemPrimitives.scala 121:29:@16932.4]
  wire  StickySelects_5_io_outs_1; // @[MemPrimitives.scala 121:29:@16932.4]
  wire  StickySelects_5_io_outs_2; // @[MemPrimitives.scala 121:29:@16932.4]
  wire  StickySelects_5_io_outs_3; // @[MemPrimitives.scala 121:29:@16932.4]
  wire  StickySelects_5_io_outs_4; // @[MemPrimitives.scala 121:29:@16932.4]
  wire  StickySelects_5_io_outs_5; // @[MemPrimitives.scala 121:29:@16932.4]
  wire  StickySelects_5_io_outs_6; // @[MemPrimitives.scala 121:29:@16932.4]
  wire  StickySelects_5_io_outs_7; // @[MemPrimitives.scala 121:29:@16932.4]
  wire  StickySelects_5_io_outs_8; // @[MemPrimitives.scala 121:29:@16932.4]
  wire  StickySelects_6_clock; // @[MemPrimitives.scala 121:29:@17021.4]
  wire  StickySelects_6_reset; // @[MemPrimitives.scala 121:29:@17021.4]
  wire  StickySelects_6_io_ins_0; // @[MemPrimitives.scala 121:29:@17021.4]
  wire  StickySelects_6_io_ins_1; // @[MemPrimitives.scala 121:29:@17021.4]
  wire  StickySelects_6_io_ins_2; // @[MemPrimitives.scala 121:29:@17021.4]
  wire  StickySelects_6_io_ins_3; // @[MemPrimitives.scala 121:29:@17021.4]
  wire  StickySelects_6_io_ins_4; // @[MemPrimitives.scala 121:29:@17021.4]
  wire  StickySelects_6_io_ins_5; // @[MemPrimitives.scala 121:29:@17021.4]
  wire  StickySelects_6_io_ins_6; // @[MemPrimitives.scala 121:29:@17021.4]
  wire  StickySelects_6_io_ins_7; // @[MemPrimitives.scala 121:29:@17021.4]
  wire  StickySelects_6_io_ins_8; // @[MemPrimitives.scala 121:29:@17021.4]
  wire  StickySelects_6_io_outs_0; // @[MemPrimitives.scala 121:29:@17021.4]
  wire  StickySelects_6_io_outs_1; // @[MemPrimitives.scala 121:29:@17021.4]
  wire  StickySelects_6_io_outs_2; // @[MemPrimitives.scala 121:29:@17021.4]
  wire  StickySelects_6_io_outs_3; // @[MemPrimitives.scala 121:29:@17021.4]
  wire  StickySelects_6_io_outs_4; // @[MemPrimitives.scala 121:29:@17021.4]
  wire  StickySelects_6_io_outs_5; // @[MemPrimitives.scala 121:29:@17021.4]
  wire  StickySelects_6_io_outs_6; // @[MemPrimitives.scala 121:29:@17021.4]
  wire  StickySelects_6_io_outs_7; // @[MemPrimitives.scala 121:29:@17021.4]
  wire  StickySelects_6_io_outs_8; // @[MemPrimitives.scala 121:29:@17021.4]
  wire  StickySelects_7_clock; // @[MemPrimitives.scala 121:29:@17110.4]
  wire  StickySelects_7_reset; // @[MemPrimitives.scala 121:29:@17110.4]
  wire  StickySelects_7_io_ins_0; // @[MemPrimitives.scala 121:29:@17110.4]
  wire  StickySelects_7_io_ins_1; // @[MemPrimitives.scala 121:29:@17110.4]
  wire  StickySelects_7_io_ins_2; // @[MemPrimitives.scala 121:29:@17110.4]
  wire  StickySelects_7_io_ins_3; // @[MemPrimitives.scala 121:29:@17110.4]
  wire  StickySelects_7_io_ins_4; // @[MemPrimitives.scala 121:29:@17110.4]
  wire  StickySelects_7_io_ins_5; // @[MemPrimitives.scala 121:29:@17110.4]
  wire  StickySelects_7_io_ins_6; // @[MemPrimitives.scala 121:29:@17110.4]
  wire  StickySelects_7_io_ins_7; // @[MemPrimitives.scala 121:29:@17110.4]
  wire  StickySelects_7_io_ins_8; // @[MemPrimitives.scala 121:29:@17110.4]
  wire  StickySelects_7_io_outs_0; // @[MemPrimitives.scala 121:29:@17110.4]
  wire  StickySelects_7_io_outs_1; // @[MemPrimitives.scala 121:29:@17110.4]
  wire  StickySelects_7_io_outs_2; // @[MemPrimitives.scala 121:29:@17110.4]
  wire  StickySelects_7_io_outs_3; // @[MemPrimitives.scala 121:29:@17110.4]
  wire  StickySelects_7_io_outs_4; // @[MemPrimitives.scala 121:29:@17110.4]
  wire  StickySelects_7_io_outs_5; // @[MemPrimitives.scala 121:29:@17110.4]
  wire  StickySelects_7_io_outs_6; // @[MemPrimitives.scala 121:29:@17110.4]
  wire  StickySelects_7_io_outs_7; // @[MemPrimitives.scala 121:29:@17110.4]
  wire  StickySelects_7_io_outs_8; // @[MemPrimitives.scala 121:29:@17110.4]
  wire  StickySelects_8_clock; // @[MemPrimitives.scala 121:29:@17199.4]
  wire  StickySelects_8_reset; // @[MemPrimitives.scala 121:29:@17199.4]
  wire  StickySelects_8_io_ins_0; // @[MemPrimitives.scala 121:29:@17199.4]
  wire  StickySelects_8_io_ins_1; // @[MemPrimitives.scala 121:29:@17199.4]
  wire  StickySelects_8_io_ins_2; // @[MemPrimitives.scala 121:29:@17199.4]
  wire  StickySelects_8_io_ins_3; // @[MemPrimitives.scala 121:29:@17199.4]
  wire  StickySelects_8_io_ins_4; // @[MemPrimitives.scala 121:29:@17199.4]
  wire  StickySelects_8_io_ins_5; // @[MemPrimitives.scala 121:29:@17199.4]
  wire  StickySelects_8_io_ins_6; // @[MemPrimitives.scala 121:29:@17199.4]
  wire  StickySelects_8_io_ins_7; // @[MemPrimitives.scala 121:29:@17199.4]
  wire  StickySelects_8_io_ins_8; // @[MemPrimitives.scala 121:29:@17199.4]
  wire  StickySelects_8_io_outs_0; // @[MemPrimitives.scala 121:29:@17199.4]
  wire  StickySelects_8_io_outs_1; // @[MemPrimitives.scala 121:29:@17199.4]
  wire  StickySelects_8_io_outs_2; // @[MemPrimitives.scala 121:29:@17199.4]
  wire  StickySelects_8_io_outs_3; // @[MemPrimitives.scala 121:29:@17199.4]
  wire  StickySelects_8_io_outs_4; // @[MemPrimitives.scala 121:29:@17199.4]
  wire  StickySelects_8_io_outs_5; // @[MemPrimitives.scala 121:29:@17199.4]
  wire  StickySelects_8_io_outs_6; // @[MemPrimitives.scala 121:29:@17199.4]
  wire  StickySelects_8_io_outs_7; // @[MemPrimitives.scala 121:29:@17199.4]
  wire  StickySelects_8_io_outs_8; // @[MemPrimitives.scala 121:29:@17199.4]
  wire  StickySelects_9_clock; // @[MemPrimitives.scala 121:29:@17288.4]
  wire  StickySelects_9_reset; // @[MemPrimitives.scala 121:29:@17288.4]
  wire  StickySelects_9_io_ins_0; // @[MemPrimitives.scala 121:29:@17288.4]
  wire  StickySelects_9_io_ins_1; // @[MemPrimitives.scala 121:29:@17288.4]
  wire  StickySelects_9_io_ins_2; // @[MemPrimitives.scala 121:29:@17288.4]
  wire  StickySelects_9_io_ins_3; // @[MemPrimitives.scala 121:29:@17288.4]
  wire  StickySelects_9_io_ins_4; // @[MemPrimitives.scala 121:29:@17288.4]
  wire  StickySelects_9_io_ins_5; // @[MemPrimitives.scala 121:29:@17288.4]
  wire  StickySelects_9_io_ins_6; // @[MemPrimitives.scala 121:29:@17288.4]
  wire  StickySelects_9_io_ins_7; // @[MemPrimitives.scala 121:29:@17288.4]
  wire  StickySelects_9_io_ins_8; // @[MemPrimitives.scala 121:29:@17288.4]
  wire  StickySelects_9_io_outs_0; // @[MemPrimitives.scala 121:29:@17288.4]
  wire  StickySelects_9_io_outs_1; // @[MemPrimitives.scala 121:29:@17288.4]
  wire  StickySelects_9_io_outs_2; // @[MemPrimitives.scala 121:29:@17288.4]
  wire  StickySelects_9_io_outs_3; // @[MemPrimitives.scala 121:29:@17288.4]
  wire  StickySelects_9_io_outs_4; // @[MemPrimitives.scala 121:29:@17288.4]
  wire  StickySelects_9_io_outs_5; // @[MemPrimitives.scala 121:29:@17288.4]
  wire  StickySelects_9_io_outs_6; // @[MemPrimitives.scala 121:29:@17288.4]
  wire  StickySelects_9_io_outs_7; // @[MemPrimitives.scala 121:29:@17288.4]
  wire  StickySelects_9_io_outs_8; // @[MemPrimitives.scala 121:29:@17288.4]
  wire  StickySelects_10_clock; // @[MemPrimitives.scala 121:29:@17377.4]
  wire  StickySelects_10_reset; // @[MemPrimitives.scala 121:29:@17377.4]
  wire  StickySelects_10_io_ins_0; // @[MemPrimitives.scala 121:29:@17377.4]
  wire  StickySelects_10_io_ins_1; // @[MemPrimitives.scala 121:29:@17377.4]
  wire  StickySelects_10_io_ins_2; // @[MemPrimitives.scala 121:29:@17377.4]
  wire  StickySelects_10_io_ins_3; // @[MemPrimitives.scala 121:29:@17377.4]
  wire  StickySelects_10_io_ins_4; // @[MemPrimitives.scala 121:29:@17377.4]
  wire  StickySelects_10_io_ins_5; // @[MemPrimitives.scala 121:29:@17377.4]
  wire  StickySelects_10_io_ins_6; // @[MemPrimitives.scala 121:29:@17377.4]
  wire  StickySelects_10_io_ins_7; // @[MemPrimitives.scala 121:29:@17377.4]
  wire  StickySelects_10_io_ins_8; // @[MemPrimitives.scala 121:29:@17377.4]
  wire  StickySelects_10_io_outs_0; // @[MemPrimitives.scala 121:29:@17377.4]
  wire  StickySelects_10_io_outs_1; // @[MemPrimitives.scala 121:29:@17377.4]
  wire  StickySelects_10_io_outs_2; // @[MemPrimitives.scala 121:29:@17377.4]
  wire  StickySelects_10_io_outs_3; // @[MemPrimitives.scala 121:29:@17377.4]
  wire  StickySelects_10_io_outs_4; // @[MemPrimitives.scala 121:29:@17377.4]
  wire  StickySelects_10_io_outs_5; // @[MemPrimitives.scala 121:29:@17377.4]
  wire  StickySelects_10_io_outs_6; // @[MemPrimitives.scala 121:29:@17377.4]
  wire  StickySelects_10_io_outs_7; // @[MemPrimitives.scala 121:29:@17377.4]
  wire  StickySelects_10_io_outs_8; // @[MemPrimitives.scala 121:29:@17377.4]
  wire  StickySelects_11_clock; // @[MemPrimitives.scala 121:29:@17466.4]
  wire  StickySelects_11_reset; // @[MemPrimitives.scala 121:29:@17466.4]
  wire  StickySelects_11_io_ins_0; // @[MemPrimitives.scala 121:29:@17466.4]
  wire  StickySelects_11_io_ins_1; // @[MemPrimitives.scala 121:29:@17466.4]
  wire  StickySelects_11_io_ins_2; // @[MemPrimitives.scala 121:29:@17466.4]
  wire  StickySelects_11_io_ins_3; // @[MemPrimitives.scala 121:29:@17466.4]
  wire  StickySelects_11_io_ins_4; // @[MemPrimitives.scala 121:29:@17466.4]
  wire  StickySelects_11_io_ins_5; // @[MemPrimitives.scala 121:29:@17466.4]
  wire  StickySelects_11_io_ins_6; // @[MemPrimitives.scala 121:29:@17466.4]
  wire  StickySelects_11_io_ins_7; // @[MemPrimitives.scala 121:29:@17466.4]
  wire  StickySelects_11_io_ins_8; // @[MemPrimitives.scala 121:29:@17466.4]
  wire  StickySelects_11_io_outs_0; // @[MemPrimitives.scala 121:29:@17466.4]
  wire  StickySelects_11_io_outs_1; // @[MemPrimitives.scala 121:29:@17466.4]
  wire  StickySelects_11_io_outs_2; // @[MemPrimitives.scala 121:29:@17466.4]
  wire  StickySelects_11_io_outs_3; // @[MemPrimitives.scala 121:29:@17466.4]
  wire  StickySelects_11_io_outs_4; // @[MemPrimitives.scala 121:29:@17466.4]
  wire  StickySelects_11_io_outs_5; // @[MemPrimitives.scala 121:29:@17466.4]
  wire  StickySelects_11_io_outs_6; // @[MemPrimitives.scala 121:29:@17466.4]
  wire  StickySelects_11_io_outs_7; // @[MemPrimitives.scala 121:29:@17466.4]
  wire  StickySelects_11_io_outs_8; // @[MemPrimitives.scala 121:29:@17466.4]
  wire  StickySelects_12_clock; // @[MemPrimitives.scala 121:29:@17555.4]
  wire  StickySelects_12_reset; // @[MemPrimitives.scala 121:29:@17555.4]
  wire  StickySelects_12_io_ins_0; // @[MemPrimitives.scala 121:29:@17555.4]
  wire  StickySelects_12_io_ins_1; // @[MemPrimitives.scala 121:29:@17555.4]
  wire  StickySelects_12_io_ins_2; // @[MemPrimitives.scala 121:29:@17555.4]
  wire  StickySelects_12_io_ins_3; // @[MemPrimitives.scala 121:29:@17555.4]
  wire  StickySelects_12_io_ins_4; // @[MemPrimitives.scala 121:29:@17555.4]
  wire  StickySelects_12_io_ins_5; // @[MemPrimitives.scala 121:29:@17555.4]
  wire  StickySelects_12_io_ins_6; // @[MemPrimitives.scala 121:29:@17555.4]
  wire  StickySelects_12_io_ins_7; // @[MemPrimitives.scala 121:29:@17555.4]
  wire  StickySelects_12_io_ins_8; // @[MemPrimitives.scala 121:29:@17555.4]
  wire  StickySelects_12_io_outs_0; // @[MemPrimitives.scala 121:29:@17555.4]
  wire  StickySelects_12_io_outs_1; // @[MemPrimitives.scala 121:29:@17555.4]
  wire  StickySelects_12_io_outs_2; // @[MemPrimitives.scala 121:29:@17555.4]
  wire  StickySelects_12_io_outs_3; // @[MemPrimitives.scala 121:29:@17555.4]
  wire  StickySelects_12_io_outs_4; // @[MemPrimitives.scala 121:29:@17555.4]
  wire  StickySelects_12_io_outs_5; // @[MemPrimitives.scala 121:29:@17555.4]
  wire  StickySelects_12_io_outs_6; // @[MemPrimitives.scala 121:29:@17555.4]
  wire  StickySelects_12_io_outs_7; // @[MemPrimitives.scala 121:29:@17555.4]
  wire  StickySelects_12_io_outs_8; // @[MemPrimitives.scala 121:29:@17555.4]
  wire  StickySelects_13_clock; // @[MemPrimitives.scala 121:29:@17644.4]
  wire  StickySelects_13_reset; // @[MemPrimitives.scala 121:29:@17644.4]
  wire  StickySelects_13_io_ins_0; // @[MemPrimitives.scala 121:29:@17644.4]
  wire  StickySelects_13_io_ins_1; // @[MemPrimitives.scala 121:29:@17644.4]
  wire  StickySelects_13_io_ins_2; // @[MemPrimitives.scala 121:29:@17644.4]
  wire  StickySelects_13_io_ins_3; // @[MemPrimitives.scala 121:29:@17644.4]
  wire  StickySelects_13_io_ins_4; // @[MemPrimitives.scala 121:29:@17644.4]
  wire  StickySelects_13_io_ins_5; // @[MemPrimitives.scala 121:29:@17644.4]
  wire  StickySelects_13_io_ins_6; // @[MemPrimitives.scala 121:29:@17644.4]
  wire  StickySelects_13_io_ins_7; // @[MemPrimitives.scala 121:29:@17644.4]
  wire  StickySelects_13_io_ins_8; // @[MemPrimitives.scala 121:29:@17644.4]
  wire  StickySelects_13_io_outs_0; // @[MemPrimitives.scala 121:29:@17644.4]
  wire  StickySelects_13_io_outs_1; // @[MemPrimitives.scala 121:29:@17644.4]
  wire  StickySelects_13_io_outs_2; // @[MemPrimitives.scala 121:29:@17644.4]
  wire  StickySelects_13_io_outs_3; // @[MemPrimitives.scala 121:29:@17644.4]
  wire  StickySelects_13_io_outs_4; // @[MemPrimitives.scala 121:29:@17644.4]
  wire  StickySelects_13_io_outs_5; // @[MemPrimitives.scala 121:29:@17644.4]
  wire  StickySelects_13_io_outs_6; // @[MemPrimitives.scala 121:29:@17644.4]
  wire  StickySelects_13_io_outs_7; // @[MemPrimitives.scala 121:29:@17644.4]
  wire  StickySelects_13_io_outs_8; // @[MemPrimitives.scala 121:29:@17644.4]
  wire  StickySelects_14_clock; // @[MemPrimitives.scala 121:29:@17733.4]
  wire  StickySelects_14_reset; // @[MemPrimitives.scala 121:29:@17733.4]
  wire  StickySelects_14_io_ins_0; // @[MemPrimitives.scala 121:29:@17733.4]
  wire  StickySelects_14_io_ins_1; // @[MemPrimitives.scala 121:29:@17733.4]
  wire  StickySelects_14_io_ins_2; // @[MemPrimitives.scala 121:29:@17733.4]
  wire  StickySelects_14_io_ins_3; // @[MemPrimitives.scala 121:29:@17733.4]
  wire  StickySelects_14_io_ins_4; // @[MemPrimitives.scala 121:29:@17733.4]
  wire  StickySelects_14_io_ins_5; // @[MemPrimitives.scala 121:29:@17733.4]
  wire  StickySelects_14_io_ins_6; // @[MemPrimitives.scala 121:29:@17733.4]
  wire  StickySelects_14_io_ins_7; // @[MemPrimitives.scala 121:29:@17733.4]
  wire  StickySelects_14_io_ins_8; // @[MemPrimitives.scala 121:29:@17733.4]
  wire  StickySelects_14_io_outs_0; // @[MemPrimitives.scala 121:29:@17733.4]
  wire  StickySelects_14_io_outs_1; // @[MemPrimitives.scala 121:29:@17733.4]
  wire  StickySelects_14_io_outs_2; // @[MemPrimitives.scala 121:29:@17733.4]
  wire  StickySelects_14_io_outs_3; // @[MemPrimitives.scala 121:29:@17733.4]
  wire  StickySelects_14_io_outs_4; // @[MemPrimitives.scala 121:29:@17733.4]
  wire  StickySelects_14_io_outs_5; // @[MemPrimitives.scala 121:29:@17733.4]
  wire  StickySelects_14_io_outs_6; // @[MemPrimitives.scala 121:29:@17733.4]
  wire  StickySelects_14_io_outs_7; // @[MemPrimitives.scala 121:29:@17733.4]
  wire  StickySelects_14_io_outs_8; // @[MemPrimitives.scala 121:29:@17733.4]
  wire  StickySelects_15_clock; // @[MemPrimitives.scala 121:29:@17822.4]
  wire  StickySelects_15_reset; // @[MemPrimitives.scala 121:29:@17822.4]
  wire  StickySelects_15_io_ins_0; // @[MemPrimitives.scala 121:29:@17822.4]
  wire  StickySelects_15_io_ins_1; // @[MemPrimitives.scala 121:29:@17822.4]
  wire  StickySelects_15_io_ins_2; // @[MemPrimitives.scala 121:29:@17822.4]
  wire  StickySelects_15_io_ins_3; // @[MemPrimitives.scala 121:29:@17822.4]
  wire  StickySelects_15_io_ins_4; // @[MemPrimitives.scala 121:29:@17822.4]
  wire  StickySelects_15_io_ins_5; // @[MemPrimitives.scala 121:29:@17822.4]
  wire  StickySelects_15_io_ins_6; // @[MemPrimitives.scala 121:29:@17822.4]
  wire  StickySelects_15_io_ins_7; // @[MemPrimitives.scala 121:29:@17822.4]
  wire  StickySelects_15_io_ins_8; // @[MemPrimitives.scala 121:29:@17822.4]
  wire  StickySelects_15_io_outs_0; // @[MemPrimitives.scala 121:29:@17822.4]
  wire  StickySelects_15_io_outs_1; // @[MemPrimitives.scala 121:29:@17822.4]
  wire  StickySelects_15_io_outs_2; // @[MemPrimitives.scala 121:29:@17822.4]
  wire  StickySelects_15_io_outs_3; // @[MemPrimitives.scala 121:29:@17822.4]
  wire  StickySelects_15_io_outs_4; // @[MemPrimitives.scala 121:29:@17822.4]
  wire  StickySelects_15_io_outs_5; // @[MemPrimitives.scala 121:29:@17822.4]
  wire  StickySelects_15_io_outs_6; // @[MemPrimitives.scala 121:29:@17822.4]
  wire  StickySelects_15_io_outs_7; // @[MemPrimitives.scala 121:29:@17822.4]
  wire  StickySelects_15_io_outs_8; // @[MemPrimitives.scala 121:29:@17822.4]
  wire  StickySelects_16_clock; // @[MemPrimitives.scala 121:29:@17911.4]
  wire  StickySelects_16_reset; // @[MemPrimitives.scala 121:29:@17911.4]
  wire  StickySelects_16_io_ins_0; // @[MemPrimitives.scala 121:29:@17911.4]
  wire  StickySelects_16_io_ins_1; // @[MemPrimitives.scala 121:29:@17911.4]
  wire  StickySelects_16_io_ins_2; // @[MemPrimitives.scala 121:29:@17911.4]
  wire  StickySelects_16_io_ins_3; // @[MemPrimitives.scala 121:29:@17911.4]
  wire  StickySelects_16_io_ins_4; // @[MemPrimitives.scala 121:29:@17911.4]
  wire  StickySelects_16_io_ins_5; // @[MemPrimitives.scala 121:29:@17911.4]
  wire  StickySelects_16_io_ins_6; // @[MemPrimitives.scala 121:29:@17911.4]
  wire  StickySelects_16_io_ins_7; // @[MemPrimitives.scala 121:29:@17911.4]
  wire  StickySelects_16_io_ins_8; // @[MemPrimitives.scala 121:29:@17911.4]
  wire  StickySelects_16_io_outs_0; // @[MemPrimitives.scala 121:29:@17911.4]
  wire  StickySelects_16_io_outs_1; // @[MemPrimitives.scala 121:29:@17911.4]
  wire  StickySelects_16_io_outs_2; // @[MemPrimitives.scala 121:29:@17911.4]
  wire  StickySelects_16_io_outs_3; // @[MemPrimitives.scala 121:29:@17911.4]
  wire  StickySelects_16_io_outs_4; // @[MemPrimitives.scala 121:29:@17911.4]
  wire  StickySelects_16_io_outs_5; // @[MemPrimitives.scala 121:29:@17911.4]
  wire  StickySelects_16_io_outs_6; // @[MemPrimitives.scala 121:29:@17911.4]
  wire  StickySelects_16_io_outs_7; // @[MemPrimitives.scala 121:29:@17911.4]
  wire  StickySelects_16_io_outs_8; // @[MemPrimitives.scala 121:29:@17911.4]
  wire  StickySelects_17_clock; // @[MemPrimitives.scala 121:29:@18000.4]
  wire  StickySelects_17_reset; // @[MemPrimitives.scala 121:29:@18000.4]
  wire  StickySelects_17_io_ins_0; // @[MemPrimitives.scala 121:29:@18000.4]
  wire  StickySelects_17_io_ins_1; // @[MemPrimitives.scala 121:29:@18000.4]
  wire  StickySelects_17_io_ins_2; // @[MemPrimitives.scala 121:29:@18000.4]
  wire  StickySelects_17_io_ins_3; // @[MemPrimitives.scala 121:29:@18000.4]
  wire  StickySelects_17_io_ins_4; // @[MemPrimitives.scala 121:29:@18000.4]
  wire  StickySelects_17_io_ins_5; // @[MemPrimitives.scala 121:29:@18000.4]
  wire  StickySelects_17_io_ins_6; // @[MemPrimitives.scala 121:29:@18000.4]
  wire  StickySelects_17_io_ins_7; // @[MemPrimitives.scala 121:29:@18000.4]
  wire  StickySelects_17_io_ins_8; // @[MemPrimitives.scala 121:29:@18000.4]
  wire  StickySelects_17_io_outs_0; // @[MemPrimitives.scala 121:29:@18000.4]
  wire  StickySelects_17_io_outs_1; // @[MemPrimitives.scala 121:29:@18000.4]
  wire  StickySelects_17_io_outs_2; // @[MemPrimitives.scala 121:29:@18000.4]
  wire  StickySelects_17_io_outs_3; // @[MemPrimitives.scala 121:29:@18000.4]
  wire  StickySelects_17_io_outs_4; // @[MemPrimitives.scala 121:29:@18000.4]
  wire  StickySelects_17_io_outs_5; // @[MemPrimitives.scala 121:29:@18000.4]
  wire  StickySelects_17_io_outs_6; // @[MemPrimitives.scala 121:29:@18000.4]
  wire  StickySelects_17_io_outs_7; // @[MemPrimitives.scala 121:29:@18000.4]
  wire  StickySelects_17_io_outs_8; // @[MemPrimitives.scala 121:29:@18000.4]
  wire  StickySelects_18_clock; // @[MemPrimitives.scala 121:29:@18089.4]
  wire  StickySelects_18_reset; // @[MemPrimitives.scala 121:29:@18089.4]
  wire  StickySelects_18_io_ins_0; // @[MemPrimitives.scala 121:29:@18089.4]
  wire  StickySelects_18_io_ins_1; // @[MemPrimitives.scala 121:29:@18089.4]
  wire  StickySelects_18_io_ins_2; // @[MemPrimitives.scala 121:29:@18089.4]
  wire  StickySelects_18_io_ins_3; // @[MemPrimitives.scala 121:29:@18089.4]
  wire  StickySelects_18_io_ins_4; // @[MemPrimitives.scala 121:29:@18089.4]
  wire  StickySelects_18_io_ins_5; // @[MemPrimitives.scala 121:29:@18089.4]
  wire  StickySelects_18_io_ins_6; // @[MemPrimitives.scala 121:29:@18089.4]
  wire  StickySelects_18_io_ins_7; // @[MemPrimitives.scala 121:29:@18089.4]
  wire  StickySelects_18_io_ins_8; // @[MemPrimitives.scala 121:29:@18089.4]
  wire  StickySelects_18_io_outs_0; // @[MemPrimitives.scala 121:29:@18089.4]
  wire  StickySelects_18_io_outs_1; // @[MemPrimitives.scala 121:29:@18089.4]
  wire  StickySelects_18_io_outs_2; // @[MemPrimitives.scala 121:29:@18089.4]
  wire  StickySelects_18_io_outs_3; // @[MemPrimitives.scala 121:29:@18089.4]
  wire  StickySelects_18_io_outs_4; // @[MemPrimitives.scala 121:29:@18089.4]
  wire  StickySelects_18_io_outs_5; // @[MemPrimitives.scala 121:29:@18089.4]
  wire  StickySelects_18_io_outs_6; // @[MemPrimitives.scala 121:29:@18089.4]
  wire  StickySelects_18_io_outs_7; // @[MemPrimitives.scala 121:29:@18089.4]
  wire  StickySelects_18_io_outs_8; // @[MemPrimitives.scala 121:29:@18089.4]
  wire  StickySelects_19_clock; // @[MemPrimitives.scala 121:29:@18178.4]
  wire  StickySelects_19_reset; // @[MemPrimitives.scala 121:29:@18178.4]
  wire  StickySelects_19_io_ins_0; // @[MemPrimitives.scala 121:29:@18178.4]
  wire  StickySelects_19_io_ins_1; // @[MemPrimitives.scala 121:29:@18178.4]
  wire  StickySelects_19_io_ins_2; // @[MemPrimitives.scala 121:29:@18178.4]
  wire  StickySelects_19_io_ins_3; // @[MemPrimitives.scala 121:29:@18178.4]
  wire  StickySelects_19_io_ins_4; // @[MemPrimitives.scala 121:29:@18178.4]
  wire  StickySelects_19_io_ins_5; // @[MemPrimitives.scala 121:29:@18178.4]
  wire  StickySelects_19_io_ins_6; // @[MemPrimitives.scala 121:29:@18178.4]
  wire  StickySelects_19_io_ins_7; // @[MemPrimitives.scala 121:29:@18178.4]
  wire  StickySelects_19_io_ins_8; // @[MemPrimitives.scala 121:29:@18178.4]
  wire  StickySelects_19_io_outs_0; // @[MemPrimitives.scala 121:29:@18178.4]
  wire  StickySelects_19_io_outs_1; // @[MemPrimitives.scala 121:29:@18178.4]
  wire  StickySelects_19_io_outs_2; // @[MemPrimitives.scala 121:29:@18178.4]
  wire  StickySelects_19_io_outs_3; // @[MemPrimitives.scala 121:29:@18178.4]
  wire  StickySelects_19_io_outs_4; // @[MemPrimitives.scala 121:29:@18178.4]
  wire  StickySelects_19_io_outs_5; // @[MemPrimitives.scala 121:29:@18178.4]
  wire  StickySelects_19_io_outs_6; // @[MemPrimitives.scala 121:29:@18178.4]
  wire  StickySelects_19_io_outs_7; // @[MemPrimitives.scala 121:29:@18178.4]
  wire  StickySelects_19_io_outs_8; // @[MemPrimitives.scala 121:29:@18178.4]
  wire  StickySelects_20_clock; // @[MemPrimitives.scala 121:29:@18267.4]
  wire  StickySelects_20_reset; // @[MemPrimitives.scala 121:29:@18267.4]
  wire  StickySelects_20_io_ins_0; // @[MemPrimitives.scala 121:29:@18267.4]
  wire  StickySelects_20_io_ins_1; // @[MemPrimitives.scala 121:29:@18267.4]
  wire  StickySelects_20_io_ins_2; // @[MemPrimitives.scala 121:29:@18267.4]
  wire  StickySelects_20_io_ins_3; // @[MemPrimitives.scala 121:29:@18267.4]
  wire  StickySelects_20_io_ins_4; // @[MemPrimitives.scala 121:29:@18267.4]
  wire  StickySelects_20_io_ins_5; // @[MemPrimitives.scala 121:29:@18267.4]
  wire  StickySelects_20_io_ins_6; // @[MemPrimitives.scala 121:29:@18267.4]
  wire  StickySelects_20_io_ins_7; // @[MemPrimitives.scala 121:29:@18267.4]
  wire  StickySelects_20_io_ins_8; // @[MemPrimitives.scala 121:29:@18267.4]
  wire  StickySelects_20_io_outs_0; // @[MemPrimitives.scala 121:29:@18267.4]
  wire  StickySelects_20_io_outs_1; // @[MemPrimitives.scala 121:29:@18267.4]
  wire  StickySelects_20_io_outs_2; // @[MemPrimitives.scala 121:29:@18267.4]
  wire  StickySelects_20_io_outs_3; // @[MemPrimitives.scala 121:29:@18267.4]
  wire  StickySelects_20_io_outs_4; // @[MemPrimitives.scala 121:29:@18267.4]
  wire  StickySelects_20_io_outs_5; // @[MemPrimitives.scala 121:29:@18267.4]
  wire  StickySelects_20_io_outs_6; // @[MemPrimitives.scala 121:29:@18267.4]
  wire  StickySelects_20_io_outs_7; // @[MemPrimitives.scala 121:29:@18267.4]
  wire  StickySelects_20_io_outs_8; // @[MemPrimitives.scala 121:29:@18267.4]
  wire  StickySelects_21_clock; // @[MemPrimitives.scala 121:29:@18356.4]
  wire  StickySelects_21_reset; // @[MemPrimitives.scala 121:29:@18356.4]
  wire  StickySelects_21_io_ins_0; // @[MemPrimitives.scala 121:29:@18356.4]
  wire  StickySelects_21_io_ins_1; // @[MemPrimitives.scala 121:29:@18356.4]
  wire  StickySelects_21_io_ins_2; // @[MemPrimitives.scala 121:29:@18356.4]
  wire  StickySelects_21_io_ins_3; // @[MemPrimitives.scala 121:29:@18356.4]
  wire  StickySelects_21_io_ins_4; // @[MemPrimitives.scala 121:29:@18356.4]
  wire  StickySelects_21_io_ins_5; // @[MemPrimitives.scala 121:29:@18356.4]
  wire  StickySelects_21_io_ins_6; // @[MemPrimitives.scala 121:29:@18356.4]
  wire  StickySelects_21_io_ins_7; // @[MemPrimitives.scala 121:29:@18356.4]
  wire  StickySelects_21_io_ins_8; // @[MemPrimitives.scala 121:29:@18356.4]
  wire  StickySelects_21_io_outs_0; // @[MemPrimitives.scala 121:29:@18356.4]
  wire  StickySelects_21_io_outs_1; // @[MemPrimitives.scala 121:29:@18356.4]
  wire  StickySelects_21_io_outs_2; // @[MemPrimitives.scala 121:29:@18356.4]
  wire  StickySelects_21_io_outs_3; // @[MemPrimitives.scala 121:29:@18356.4]
  wire  StickySelects_21_io_outs_4; // @[MemPrimitives.scala 121:29:@18356.4]
  wire  StickySelects_21_io_outs_5; // @[MemPrimitives.scala 121:29:@18356.4]
  wire  StickySelects_21_io_outs_6; // @[MemPrimitives.scala 121:29:@18356.4]
  wire  StickySelects_21_io_outs_7; // @[MemPrimitives.scala 121:29:@18356.4]
  wire  StickySelects_21_io_outs_8; // @[MemPrimitives.scala 121:29:@18356.4]
  wire  StickySelects_22_clock; // @[MemPrimitives.scala 121:29:@18445.4]
  wire  StickySelects_22_reset; // @[MemPrimitives.scala 121:29:@18445.4]
  wire  StickySelects_22_io_ins_0; // @[MemPrimitives.scala 121:29:@18445.4]
  wire  StickySelects_22_io_ins_1; // @[MemPrimitives.scala 121:29:@18445.4]
  wire  StickySelects_22_io_ins_2; // @[MemPrimitives.scala 121:29:@18445.4]
  wire  StickySelects_22_io_ins_3; // @[MemPrimitives.scala 121:29:@18445.4]
  wire  StickySelects_22_io_ins_4; // @[MemPrimitives.scala 121:29:@18445.4]
  wire  StickySelects_22_io_ins_5; // @[MemPrimitives.scala 121:29:@18445.4]
  wire  StickySelects_22_io_ins_6; // @[MemPrimitives.scala 121:29:@18445.4]
  wire  StickySelects_22_io_ins_7; // @[MemPrimitives.scala 121:29:@18445.4]
  wire  StickySelects_22_io_ins_8; // @[MemPrimitives.scala 121:29:@18445.4]
  wire  StickySelects_22_io_outs_0; // @[MemPrimitives.scala 121:29:@18445.4]
  wire  StickySelects_22_io_outs_1; // @[MemPrimitives.scala 121:29:@18445.4]
  wire  StickySelects_22_io_outs_2; // @[MemPrimitives.scala 121:29:@18445.4]
  wire  StickySelects_22_io_outs_3; // @[MemPrimitives.scala 121:29:@18445.4]
  wire  StickySelects_22_io_outs_4; // @[MemPrimitives.scala 121:29:@18445.4]
  wire  StickySelects_22_io_outs_5; // @[MemPrimitives.scala 121:29:@18445.4]
  wire  StickySelects_22_io_outs_6; // @[MemPrimitives.scala 121:29:@18445.4]
  wire  StickySelects_22_io_outs_7; // @[MemPrimitives.scala 121:29:@18445.4]
  wire  StickySelects_22_io_outs_8; // @[MemPrimitives.scala 121:29:@18445.4]
  wire  StickySelects_23_clock; // @[MemPrimitives.scala 121:29:@18534.4]
  wire  StickySelects_23_reset; // @[MemPrimitives.scala 121:29:@18534.4]
  wire  StickySelects_23_io_ins_0; // @[MemPrimitives.scala 121:29:@18534.4]
  wire  StickySelects_23_io_ins_1; // @[MemPrimitives.scala 121:29:@18534.4]
  wire  StickySelects_23_io_ins_2; // @[MemPrimitives.scala 121:29:@18534.4]
  wire  StickySelects_23_io_ins_3; // @[MemPrimitives.scala 121:29:@18534.4]
  wire  StickySelects_23_io_ins_4; // @[MemPrimitives.scala 121:29:@18534.4]
  wire  StickySelects_23_io_ins_5; // @[MemPrimitives.scala 121:29:@18534.4]
  wire  StickySelects_23_io_ins_6; // @[MemPrimitives.scala 121:29:@18534.4]
  wire  StickySelects_23_io_ins_7; // @[MemPrimitives.scala 121:29:@18534.4]
  wire  StickySelects_23_io_ins_8; // @[MemPrimitives.scala 121:29:@18534.4]
  wire  StickySelects_23_io_outs_0; // @[MemPrimitives.scala 121:29:@18534.4]
  wire  StickySelects_23_io_outs_1; // @[MemPrimitives.scala 121:29:@18534.4]
  wire  StickySelects_23_io_outs_2; // @[MemPrimitives.scala 121:29:@18534.4]
  wire  StickySelects_23_io_outs_3; // @[MemPrimitives.scala 121:29:@18534.4]
  wire  StickySelects_23_io_outs_4; // @[MemPrimitives.scala 121:29:@18534.4]
  wire  StickySelects_23_io_outs_5; // @[MemPrimitives.scala 121:29:@18534.4]
  wire  StickySelects_23_io_outs_6; // @[MemPrimitives.scala 121:29:@18534.4]
  wire  StickySelects_23_io_outs_7; // @[MemPrimitives.scala 121:29:@18534.4]
  wire  StickySelects_23_io_outs_8; // @[MemPrimitives.scala 121:29:@18534.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@18624.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@18624.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@18624.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@18624.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@18624.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@18632.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@18632.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@18632.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@18632.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@18632.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@18640.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@18640.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@18640.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@18640.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@18640.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@18648.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@18648.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@18648.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@18648.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@18648.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@18656.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@18656.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@18656.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@18656.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@18656.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@18664.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@18664.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@18664.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@18664.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@18664.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@18672.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@18672.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@18672.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@18672.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@18672.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@18680.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@18680.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@18680.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@18680.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@18680.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@18688.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@18688.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@18688.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@18688.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@18688.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@18696.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@18696.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@18696.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@18696.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@18696.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@18704.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@18704.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@18704.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@18704.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@18704.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@18712.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@18712.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@18712.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@18712.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@18712.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@18768.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@18768.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@18768.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@18768.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@18768.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@18776.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@18776.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@18776.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@18776.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@18776.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@18784.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@18784.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@18784.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@18784.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@18784.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@18792.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@18792.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@18792.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@18792.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@18792.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@18800.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@18800.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@18800.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@18800.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@18800.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@18808.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@18808.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@18808.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@18808.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@18808.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@18816.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@18816.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@18816.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@18816.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@18816.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@18824.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@18824.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@18824.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@18824.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@18824.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@18832.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@18832.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@18832.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@18832.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@18832.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@18840.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@18840.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@18840.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@18840.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@18840.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@18848.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@18848.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@18848.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@18848.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@18848.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@18856.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@18856.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@18856.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@18856.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@18856.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@18912.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@18912.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@18912.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@18912.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@18912.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@18920.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@18920.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@18920.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@18920.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@18920.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@18928.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@18928.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@18928.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@18928.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@18928.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@18936.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@18936.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@18936.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@18936.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@18936.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@18944.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@18944.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@18944.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@18944.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@18944.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@18952.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@18952.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@18952.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@18952.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@18952.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@18960.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@18960.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@18960.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@18960.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@18960.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@18968.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@18968.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@18968.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@18968.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@18968.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@18976.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@18976.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@18976.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@18976.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@18976.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@18984.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@18984.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@18984.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@18984.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@18984.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@18992.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@18992.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@18992.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@18992.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@18992.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@19000.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@19000.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@19000.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@19000.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@19000.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@19056.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@19056.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@19056.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@19056.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@19056.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@19064.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@19064.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@19064.4]
  wire  RetimeWrapper_37_io_in; // @[package.scala 93:22:@19064.4]
  wire  RetimeWrapper_37_io_out; // @[package.scala 93:22:@19064.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@19072.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@19072.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@19072.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@19072.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@19072.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@19080.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@19080.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@19080.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@19080.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@19080.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@19088.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@19088.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@19088.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@19088.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@19088.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@19096.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@19096.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@19096.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@19096.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@19096.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@19104.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@19104.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@19104.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@19104.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@19104.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@19112.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@19112.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@19112.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@19112.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@19112.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@19120.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@19120.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@19120.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@19120.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@19120.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@19128.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@19128.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@19128.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@19128.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@19128.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@19136.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@19136.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@19136.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@19136.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@19136.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@19144.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@19144.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@19144.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@19144.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@19144.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@19200.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@19200.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@19200.4]
  wire  RetimeWrapper_48_io_in; // @[package.scala 93:22:@19200.4]
  wire  RetimeWrapper_48_io_out; // @[package.scala 93:22:@19200.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@19208.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@19208.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@19208.4]
  wire  RetimeWrapper_49_io_in; // @[package.scala 93:22:@19208.4]
  wire  RetimeWrapper_49_io_out; // @[package.scala 93:22:@19208.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@19216.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@19216.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@19216.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@19216.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@19216.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@19224.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@19224.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@19224.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@19224.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@19224.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@19232.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@19232.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@19232.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@19232.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@19232.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@19240.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@19240.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@19240.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@19240.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@19240.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@19248.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@19248.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@19248.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@19248.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@19248.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@19256.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@19256.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@19256.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@19256.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@19256.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@19264.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@19264.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@19264.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@19264.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@19264.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@19272.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@19272.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@19272.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@19272.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@19272.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@19280.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@19280.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@19280.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@19280.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@19280.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@19288.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@19288.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@19288.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@19288.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@19288.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@19344.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@19344.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@19344.4]
  wire  RetimeWrapper_60_io_in; // @[package.scala 93:22:@19344.4]
  wire  RetimeWrapper_60_io_out; // @[package.scala 93:22:@19344.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@19352.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@19352.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@19352.4]
  wire  RetimeWrapper_61_io_in; // @[package.scala 93:22:@19352.4]
  wire  RetimeWrapper_61_io_out; // @[package.scala 93:22:@19352.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@19360.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@19360.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@19360.4]
  wire  RetimeWrapper_62_io_in; // @[package.scala 93:22:@19360.4]
  wire  RetimeWrapper_62_io_out; // @[package.scala 93:22:@19360.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@19368.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@19368.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@19368.4]
  wire  RetimeWrapper_63_io_in; // @[package.scala 93:22:@19368.4]
  wire  RetimeWrapper_63_io_out; // @[package.scala 93:22:@19368.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@19376.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@19376.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@19376.4]
  wire  RetimeWrapper_64_io_in; // @[package.scala 93:22:@19376.4]
  wire  RetimeWrapper_64_io_out; // @[package.scala 93:22:@19376.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@19384.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@19384.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@19384.4]
  wire  RetimeWrapper_65_io_in; // @[package.scala 93:22:@19384.4]
  wire  RetimeWrapper_65_io_out; // @[package.scala 93:22:@19384.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@19392.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@19392.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@19392.4]
  wire  RetimeWrapper_66_io_in; // @[package.scala 93:22:@19392.4]
  wire  RetimeWrapper_66_io_out; // @[package.scala 93:22:@19392.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@19400.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@19400.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@19400.4]
  wire  RetimeWrapper_67_io_in; // @[package.scala 93:22:@19400.4]
  wire  RetimeWrapper_67_io_out; // @[package.scala 93:22:@19400.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@19408.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@19408.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@19408.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@19408.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@19408.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@19416.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@19416.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@19416.4]
  wire  RetimeWrapper_69_io_in; // @[package.scala 93:22:@19416.4]
  wire  RetimeWrapper_69_io_out; // @[package.scala 93:22:@19416.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@19424.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@19424.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@19424.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@19424.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@19424.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@19432.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@19432.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@19432.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@19432.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@19432.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@19488.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@19488.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@19488.4]
  wire  RetimeWrapper_72_io_in; // @[package.scala 93:22:@19488.4]
  wire  RetimeWrapper_72_io_out; // @[package.scala 93:22:@19488.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@19496.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@19496.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@19496.4]
  wire  RetimeWrapper_73_io_in; // @[package.scala 93:22:@19496.4]
  wire  RetimeWrapper_73_io_out; // @[package.scala 93:22:@19496.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@19504.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@19504.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@19504.4]
  wire  RetimeWrapper_74_io_in; // @[package.scala 93:22:@19504.4]
  wire  RetimeWrapper_74_io_out; // @[package.scala 93:22:@19504.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@19512.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@19512.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@19512.4]
  wire  RetimeWrapper_75_io_in; // @[package.scala 93:22:@19512.4]
  wire  RetimeWrapper_75_io_out; // @[package.scala 93:22:@19512.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@19520.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@19520.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@19520.4]
  wire  RetimeWrapper_76_io_in; // @[package.scala 93:22:@19520.4]
  wire  RetimeWrapper_76_io_out; // @[package.scala 93:22:@19520.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@19528.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@19528.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@19528.4]
  wire  RetimeWrapper_77_io_in; // @[package.scala 93:22:@19528.4]
  wire  RetimeWrapper_77_io_out; // @[package.scala 93:22:@19528.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@19536.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@19536.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@19536.4]
  wire  RetimeWrapper_78_io_in; // @[package.scala 93:22:@19536.4]
  wire  RetimeWrapper_78_io_out; // @[package.scala 93:22:@19536.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@19544.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@19544.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@19544.4]
  wire  RetimeWrapper_79_io_in; // @[package.scala 93:22:@19544.4]
  wire  RetimeWrapper_79_io_out; // @[package.scala 93:22:@19544.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@19552.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@19552.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@19552.4]
  wire  RetimeWrapper_80_io_in; // @[package.scala 93:22:@19552.4]
  wire  RetimeWrapper_80_io_out; // @[package.scala 93:22:@19552.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@19560.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@19560.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@19560.4]
  wire  RetimeWrapper_81_io_in; // @[package.scala 93:22:@19560.4]
  wire  RetimeWrapper_81_io_out; // @[package.scala 93:22:@19560.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@19568.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@19568.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@19568.4]
  wire  RetimeWrapper_82_io_in; // @[package.scala 93:22:@19568.4]
  wire  RetimeWrapper_82_io_out; // @[package.scala 93:22:@19568.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@19576.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@19576.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@19576.4]
  wire  RetimeWrapper_83_io_in; // @[package.scala 93:22:@19576.4]
  wire  RetimeWrapper_83_io_out; // @[package.scala 93:22:@19576.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@19632.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@19632.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@19632.4]
  wire  RetimeWrapper_84_io_in; // @[package.scala 93:22:@19632.4]
  wire  RetimeWrapper_84_io_out; // @[package.scala 93:22:@19632.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@19640.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@19640.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@19640.4]
  wire  RetimeWrapper_85_io_in; // @[package.scala 93:22:@19640.4]
  wire  RetimeWrapper_85_io_out; // @[package.scala 93:22:@19640.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@19648.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@19648.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@19648.4]
  wire  RetimeWrapper_86_io_in; // @[package.scala 93:22:@19648.4]
  wire  RetimeWrapper_86_io_out; // @[package.scala 93:22:@19648.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@19656.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@19656.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@19656.4]
  wire  RetimeWrapper_87_io_in; // @[package.scala 93:22:@19656.4]
  wire  RetimeWrapper_87_io_out; // @[package.scala 93:22:@19656.4]
  wire  RetimeWrapper_88_clock; // @[package.scala 93:22:@19664.4]
  wire  RetimeWrapper_88_reset; // @[package.scala 93:22:@19664.4]
  wire  RetimeWrapper_88_io_flow; // @[package.scala 93:22:@19664.4]
  wire  RetimeWrapper_88_io_in; // @[package.scala 93:22:@19664.4]
  wire  RetimeWrapper_88_io_out; // @[package.scala 93:22:@19664.4]
  wire  RetimeWrapper_89_clock; // @[package.scala 93:22:@19672.4]
  wire  RetimeWrapper_89_reset; // @[package.scala 93:22:@19672.4]
  wire  RetimeWrapper_89_io_flow; // @[package.scala 93:22:@19672.4]
  wire  RetimeWrapper_89_io_in; // @[package.scala 93:22:@19672.4]
  wire  RetimeWrapper_89_io_out; // @[package.scala 93:22:@19672.4]
  wire  RetimeWrapper_90_clock; // @[package.scala 93:22:@19680.4]
  wire  RetimeWrapper_90_reset; // @[package.scala 93:22:@19680.4]
  wire  RetimeWrapper_90_io_flow; // @[package.scala 93:22:@19680.4]
  wire  RetimeWrapper_90_io_in; // @[package.scala 93:22:@19680.4]
  wire  RetimeWrapper_90_io_out; // @[package.scala 93:22:@19680.4]
  wire  RetimeWrapper_91_clock; // @[package.scala 93:22:@19688.4]
  wire  RetimeWrapper_91_reset; // @[package.scala 93:22:@19688.4]
  wire  RetimeWrapper_91_io_flow; // @[package.scala 93:22:@19688.4]
  wire  RetimeWrapper_91_io_in; // @[package.scala 93:22:@19688.4]
  wire  RetimeWrapper_91_io_out; // @[package.scala 93:22:@19688.4]
  wire  RetimeWrapper_92_clock; // @[package.scala 93:22:@19696.4]
  wire  RetimeWrapper_92_reset; // @[package.scala 93:22:@19696.4]
  wire  RetimeWrapper_92_io_flow; // @[package.scala 93:22:@19696.4]
  wire  RetimeWrapper_92_io_in; // @[package.scala 93:22:@19696.4]
  wire  RetimeWrapper_92_io_out; // @[package.scala 93:22:@19696.4]
  wire  RetimeWrapper_93_clock; // @[package.scala 93:22:@19704.4]
  wire  RetimeWrapper_93_reset; // @[package.scala 93:22:@19704.4]
  wire  RetimeWrapper_93_io_flow; // @[package.scala 93:22:@19704.4]
  wire  RetimeWrapper_93_io_in; // @[package.scala 93:22:@19704.4]
  wire  RetimeWrapper_93_io_out; // @[package.scala 93:22:@19704.4]
  wire  RetimeWrapper_94_clock; // @[package.scala 93:22:@19712.4]
  wire  RetimeWrapper_94_reset; // @[package.scala 93:22:@19712.4]
  wire  RetimeWrapper_94_io_flow; // @[package.scala 93:22:@19712.4]
  wire  RetimeWrapper_94_io_in; // @[package.scala 93:22:@19712.4]
  wire  RetimeWrapper_94_io_out; // @[package.scala 93:22:@19712.4]
  wire  RetimeWrapper_95_clock; // @[package.scala 93:22:@19720.4]
  wire  RetimeWrapper_95_reset; // @[package.scala 93:22:@19720.4]
  wire  RetimeWrapper_95_io_flow; // @[package.scala 93:22:@19720.4]
  wire  RetimeWrapper_95_io_in; // @[package.scala 93:22:@19720.4]
  wire  RetimeWrapper_95_io_out; // @[package.scala 93:22:@19720.4]
  wire  RetimeWrapper_96_clock; // @[package.scala 93:22:@19776.4]
  wire  RetimeWrapper_96_reset; // @[package.scala 93:22:@19776.4]
  wire  RetimeWrapper_96_io_flow; // @[package.scala 93:22:@19776.4]
  wire  RetimeWrapper_96_io_in; // @[package.scala 93:22:@19776.4]
  wire  RetimeWrapper_96_io_out; // @[package.scala 93:22:@19776.4]
  wire  RetimeWrapper_97_clock; // @[package.scala 93:22:@19784.4]
  wire  RetimeWrapper_97_reset; // @[package.scala 93:22:@19784.4]
  wire  RetimeWrapper_97_io_flow; // @[package.scala 93:22:@19784.4]
  wire  RetimeWrapper_97_io_in; // @[package.scala 93:22:@19784.4]
  wire  RetimeWrapper_97_io_out; // @[package.scala 93:22:@19784.4]
  wire  RetimeWrapper_98_clock; // @[package.scala 93:22:@19792.4]
  wire  RetimeWrapper_98_reset; // @[package.scala 93:22:@19792.4]
  wire  RetimeWrapper_98_io_flow; // @[package.scala 93:22:@19792.4]
  wire  RetimeWrapper_98_io_in; // @[package.scala 93:22:@19792.4]
  wire  RetimeWrapper_98_io_out; // @[package.scala 93:22:@19792.4]
  wire  RetimeWrapper_99_clock; // @[package.scala 93:22:@19800.4]
  wire  RetimeWrapper_99_reset; // @[package.scala 93:22:@19800.4]
  wire  RetimeWrapper_99_io_flow; // @[package.scala 93:22:@19800.4]
  wire  RetimeWrapper_99_io_in; // @[package.scala 93:22:@19800.4]
  wire  RetimeWrapper_99_io_out; // @[package.scala 93:22:@19800.4]
  wire  RetimeWrapper_100_clock; // @[package.scala 93:22:@19808.4]
  wire  RetimeWrapper_100_reset; // @[package.scala 93:22:@19808.4]
  wire  RetimeWrapper_100_io_flow; // @[package.scala 93:22:@19808.4]
  wire  RetimeWrapper_100_io_in; // @[package.scala 93:22:@19808.4]
  wire  RetimeWrapper_100_io_out; // @[package.scala 93:22:@19808.4]
  wire  RetimeWrapper_101_clock; // @[package.scala 93:22:@19816.4]
  wire  RetimeWrapper_101_reset; // @[package.scala 93:22:@19816.4]
  wire  RetimeWrapper_101_io_flow; // @[package.scala 93:22:@19816.4]
  wire  RetimeWrapper_101_io_in; // @[package.scala 93:22:@19816.4]
  wire  RetimeWrapper_101_io_out; // @[package.scala 93:22:@19816.4]
  wire  RetimeWrapper_102_clock; // @[package.scala 93:22:@19824.4]
  wire  RetimeWrapper_102_reset; // @[package.scala 93:22:@19824.4]
  wire  RetimeWrapper_102_io_flow; // @[package.scala 93:22:@19824.4]
  wire  RetimeWrapper_102_io_in; // @[package.scala 93:22:@19824.4]
  wire  RetimeWrapper_102_io_out; // @[package.scala 93:22:@19824.4]
  wire  RetimeWrapper_103_clock; // @[package.scala 93:22:@19832.4]
  wire  RetimeWrapper_103_reset; // @[package.scala 93:22:@19832.4]
  wire  RetimeWrapper_103_io_flow; // @[package.scala 93:22:@19832.4]
  wire  RetimeWrapper_103_io_in; // @[package.scala 93:22:@19832.4]
  wire  RetimeWrapper_103_io_out; // @[package.scala 93:22:@19832.4]
  wire  RetimeWrapper_104_clock; // @[package.scala 93:22:@19840.4]
  wire  RetimeWrapper_104_reset; // @[package.scala 93:22:@19840.4]
  wire  RetimeWrapper_104_io_flow; // @[package.scala 93:22:@19840.4]
  wire  RetimeWrapper_104_io_in; // @[package.scala 93:22:@19840.4]
  wire  RetimeWrapper_104_io_out; // @[package.scala 93:22:@19840.4]
  wire  RetimeWrapper_105_clock; // @[package.scala 93:22:@19848.4]
  wire  RetimeWrapper_105_reset; // @[package.scala 93:22:@19848.4]
  wire  RetimeWrapper_105_io_flow; // @[package.scala 93:22:@19848.4]
  wire  RetimeWrapper_105_io_in; // @[package.scala 93:22:@19848.4]
  wire  RetimeWrapper_105_io_out; // @[package.scala 93:22:@19848.4]
  wire  RetimeWrapper_106_clock; // @[package.scala 93:22:@19856.4]
  wire  RetimeWrapper_106_reset; // @[package.scala 93:22:@19856.4]
  wire  RetimeWrapper_106_io_flow; // @[package.scala 93:22:@19856.4]
  wire  RetimeWrapper_106_io_in; // @[package.scala 93:22:@19856.4]
  wire  RetimeWrapper_106_io_out; // @[package.scala 93:22:@19856.4]
  wire  RetimeWrapper_107_clock; // @[package.scala 93:22:@19864.4]
  wire  RetimeWrapper_107_reset; // @[package.scala 93:22:@19864.4]
  wire  RetimeWrapper_107_io_flow; // @[package.scala 93:22:@19864.4]
  wire  RetimeWrapper_107_io_in; // @[package.scala 93:22:@19864.4]
  wire  RetimeWrapper_107_io_out; // @[package.scala 93:22:@19864.4]
  wire  RetimeWrapper_108_clock; // @[package.scala 93:22:@19920.4]
  wire  RetimeWrapper_108_reset; // @[package.scala 93:22:@19920.4]
  wire  RetimeWrapper_108_io_flow; // @[package.scala 93:22:@19920.4]
  wire  RetimeWrapper_108_io_in; // @[package.scala 93:22:@19920.4]
  wire  RetimeWrapper_108_io_out; // @[package.scala 93:22:@19920.4]
  wire  RetimeWrapper_109_clock; // @[package.scala 93:22:@19928.4]
  wire  RetimeWrapper_109_reset; // @[package.scala 93:22:@19928.4]
  wire  RetimeWrapper_109_io_flow; // @[package.scala 93:22:@19928.4]
  wire  RetimeWrapper_109_io_in; // @[package.scala 93:22:@19928.4]
  wire  RetimeWrapper_109_io_out; // @[package.scala 93:22:@19928.4]
  wire  RetimeWrapper_110_clock; // @[package.scala 93:22:@19936.4]
  wire  RetimeWrapper_110_reset; // @[package.scala 93:22:@19936.4]
  wire  RetimeWrapper_110_io_flow; // @[package.scala 93:22:@19936.4]
  wire  RetimeWrapper_110_io_in; // @[package.scala 93:22:@19936.4]
  wire  RetimeWrapper_110_io_out; // @[package.scala 93:22:@19936.4]
  wire  RetimeWrapper_111_clock; // @[package.scala 93:22:@19944.4]
  wire  RetimeWrapper_111_reset; // @[package.scala 93:22:@19944.4]
  wire  RetimeWrapper_111_io_flow; // @[package.scala 93:22:@19944.4]
  wire  RetimeWrapper_111_io_in; // @[package.scala 93:22:@19944.4]
  wire  RetimeWrapper_111_io_out; // @[package.scala 93:22:@19944.4]
  wire  RetimeWrapper_112_clock; // @[package.scala 93:22:@19952.4]
  wire  RetimeWrapper_112_reset; // @[package.scala 93:22:@19952.4]
  wire  RetimeWrapper_112_io_flow; // @[package.scala 93:22:@19952.4]
  wire  RetimeWrapper_112_io_in; // @[package.scala 93:22:@19952.4]
  wire  RetimeWrapper_112_io_out; // @[package.scala 93:22:@19952.4]
  wire  RetimeWrapper_113_clock; // @[package.scala 93:22:@19960.4]
  wire  RetimeWrapper_113_reset; // @[package.scala 93:22:@19960.4]
  wire  RetimeWrapper_113_io_flow; // @[package.scala 93:22:@19960.4]
  wire  RetimeWrapper_113_io_in; // @[package.scala 93:22:@19960.4]
  wire  RetimeWrapper_113_io_out; // @[package.scala 93:22:@19960.4]
  wire  RetimeWrapper_114_clock; // @[package.scala 93:22:@19968.4]
  wire  RetimeWrapper_114_reset; // @[package.scala 93:22:@19968.4]
  wire  RetimeWrapper_114_io_flow; // @[package.scala 93:22:@19968.4]
  wire  RetimeWrapper_114_io_in; // @[package.scala 93:22:@19968.4]
  wire  RetimeWrapper_114_io_out; // @[package.scala 93:22:@19968.4]
  wire  RetimeWrapper_115_clock; // @[package.scala 93:22:@19976.4]
  wire  RetimeWrapper_115_reset; // @[package.scala 93:22:@19976.4]
  wire  RetimeWrapper_115_io_flow; // @[package.scala 93:22:@19976.4]
  wire  RetimeWrapper_115_io_in; // @[package.scala 93:22:@19976.4]
  wire  RetimeWrapper_115_io_out; // @[package.scala 93:22:@19976.4]
  wire  RetimeWrapper_116_clock; // @[package.scala 93:22:@19984.4]
  wire  RetimeWrapper_116_reset; // @[package.scala 93:22:@19984.4]
  wire  RetimeWrapper_116_io_flow; // @[package.scala 93:22:@19984.4]
  wire  RetimeWrapper_116_io_in; // @[package.scala 93:22:@19984.4]
  wire  RetimeWrapper_116_io_out; // @[package.scala 93:22:@19984.4]
  wire  RetimeWrapper_117_clock; // @[package.scala 93:22:@19992.4]
  wire  RetimeWrapper_117_reset; // @[package.scala 93:22:@19992.4]
  wire  RetimeWrapper_117_io_flow; // @[package.scala 93:22:@19992.4]
  wire  RetimeWrapper_117_io_in; // @[package.scala 93:22:@19992.4]
  wire  RetimeWrapper_117_io_out; // @[package.scala 93:22:@19992.4]
  wire  RetimeWrapper_118_clock; // @[package.scala 93:22:@20000.4]
  wire  RetimeWrapper_118_reset; // @[package.scala 93:22:@20000.4]
  wire  RetimeWrapper_118_io_flow; // @[package.scala 93:22:@20000.4]
  wire  RetimeWrapper_118_io_in; // @[package.scala 93:22:@20000.4]
  wire  RetimeWrapper_118_io_out; // @[package.scala 93:22:@20000.4]
  wire  RetimeWrapper_119_clock; // @[package.scala 93:22:@20008.4]
  wire  RetimeWrapper_119_reset; // @[package.scala 93:22:@20008.4]
  wire  RetimeWrapper_119_io_flow; // @[package.scala 93:22:@20008.4]
  wire  RetimeWrapper_119_io_in; // @[package.scala 93:22:@20008.4]
  wire  RetimeWrapper_119_io_out; // @[package.scala 93:22:@20008.4]
  wire  RetimeWrapper_120_clock; // @[package.scala 93:22:@20064.4]
  wire  RetimeWrapper_120_reset; // @[package.scala 93:22:@20064.4]
  wire  RetimeWrapper_120_io_flow; // @[package.scala 93:22:@20064.4]
  wire  RetimeWrapper_120_io_in; // @[package.scala 93:22:@20064.4]
  wire  RetimeWrapper_120_io_out; // @[package.scala 93:22:@20064.4]
  wire  RetimeWrapper_121_clock; // @[package.scala 93:22:@20072.4]
  wire  RetimeWrapper_121_reset; // @[package.scala 93:22:@20072.4]
  wire  RetimeWrapper_121_io_flow; // @[package.scala 93:22:@20072.4]
  wire  RetimeWrapper_121_io_in; // @[package.scala 93:22:@20072.4]
  wire  RetimeWrapper_121_io_out; // @[package.scala 93:22:@20072.4]
  wire  RetimeWrapper_122_clock; // @[package.scala 93:22:@20080.4]
  wire  RetimeWrapper_122_reset; // @[package.scala 93:22:@20080.4]
  wire  RetimeWrapper_122_io_flow; // @[package.scala 93:22:@20080.4]
  wire  RetimeWrapper_122_io_in; // @[package.scala 93:22:@20080.4]
  wire  RetimeWrapper_122_io_out; // @[package.scala 93:22:@20080.4]
  wire  RetimeWrapper_123_clock; // @[package.scala 93:22:@20088.4]
  wire  RetimeWrapper_123_reset; // @[package.scala 93:22:@20088.4]
  wire  RetimeWrapper_123_io_flow; // @[package.scala 93:22:@20088.4]
  wire  RetimeWrapper_123_io_in; // @[package.scala 93:22:@20088.4]
  wire  RetimeWrapper_123_io_out; // @[package.scala 93:22:@20088.4]
  wire  RetimeWrapper_124_clock; // @[package.scala 93:22:@20096.4]
  wire  RetimeWrapper_124_reset; // @[package.scala 93:22:@20096.4]
  wire  RetimeWrapper_124_io_flow; // @[package.scala 93:22:@20096.4]
  wire  RetimeWrapper_124_io_in; // @[package.scala 93:22:@20096.4]
  wire  RetimeWrapper_124_io_out; // @[package.scala 93:22:@20096.4]
  wire  RetimeWrapper_125_clock; // @[package.scala 93:22:@20104.4]
  wire  RetimeWrapper_125_reset; // @[package.scala 93:22:@20104.4]
  wire  RetimeWrapper_125_io_flow; // @[package.scala 93:22:@20104.4]
  wire  RetimeWrapper_125_io_in; // @[package.scala 93:22:@20104.4]
  wire  RetimeWrapper_125_io_out; // @[package.scala 93:22:@20104.4]
  wire  RetimeWrapper_126_clock; // @[package.scala 93:22:@20112.4]
  wire  RetimeWrapper_126_reset; // @[package.scala 93:22:@20112.4]
  wire  RetimeWrapper_126_io_flow; // @[package.scala 93:22:@20112.4]
  wire  RetimeWrapper_126_io_in; // @[package.scala 93:22:@20112.4]
  wire  RetimeWrapper_126_io_out; // @[package.scala 93:22:@20112.4]
  wire  RetimeWrapper_127_clock; // @[package.scala 93:22:@20120.4]
  wire  RetimeWrapper_127_reset; // @[package.scala 93:22:@20120.4]
  wire  RetimeWrapper_127_io_flow; // @[package.scala 93:22:@20120.4]
  wire  RetimeWrapper_127_io_in; // @[package.scala 93:22:@20120.4]
  wire  RetimeWrapper_127_io_out; // @[package.scala 93:22:@20120.4]
  wire  RetimeWrapper_128_clock; // @[package.scala 93:22:@20128.4]
  wire  RetimeWrapper_128_reset; // @[package.scala 93:22:@20128.4]
  wire  RetimeWrapper_128_io_flow; // @[package.scala 93:22:@20128.4]
  wire  RetimeWrapper_128_io_in; // @[package.scala 93:22:@20128.4]
  wire  RetimeWrapper_128_io_out; // @[package.scala 93:22:@20128.4]
  wire  RetimeWrapper_129_clock; // @[package.scala 93:22:@20136.4]
  wire  RetimeWrapper_129_reset; // @[package.scala 93:22:@20136.4]
  wire  RetimeWrapper_129_io_flow; // @[package.scala 93:22:@20136.4]
  wire  RetimeWrapper_129_io_in; // @[package.scala 93:22:@20136.4]
  wire  RetimeWrapper_129_io_out; // @[package.scala 93:22:@20136.4]
  wire  RetimeWrapper_130_clock; // @[package.scala 93:22:@20144.4]
  wire  RetimeWrapper_130_reset; // @[package.scala 93:22:@20144.4]
  wire  RetimeWrapper_130_io_flow; // @[package.scala 93:22:@20144.4]
  wire  RetimeWrapper_130_io_in; // @[package.scala 93:22:@20144.4]
  wire  RetimeWrapper_130_io_out; // @[package.scala 93:22:@20144.4]
  wire  RetimeWrapper_131_clock; // @[package.scala 93:22:@20152.4]
  wire  RetimeWrapper_131_reset; // @[package.scala 93:22:@20152.4]
  wire  RetimeWrapper_131_io_flow; // @[package.scala 93:22:@20152.4]
  wire  RetimeWrapper_131_io_in; // @[package.scala 93:22:@20152.4]
  wire  RetimeWrapper_131_io_out; // @[package.scala 93:22:@20152.4]
  wire  RetimeWrapper_132_clock; // @[package.scala 93:22:@20208.4]
  wire  RetimeWrapper_132_reset; // @[package.scala 93:22:@20208.4]
  wire  RetimeWrapper_132_io_flow; // @[package.scala 93:22:@20208.4]
  wire  RetimeWrapper_132_io_in; // @[package.scala 93:22:@20208.4]
  wire  RetimeWrapper_132_io_out; // @[package.scala 93:22:@20208.4]
  wire  RetimeWrapper_133_clock; // @[package.scala 93:22:@20216.4]
  wire  RetimeWrapper_133_reset; // @[package.scala 93:22:@20216.4]
  wire  RetimeWrapper_133_io_flow; // @[package.scala 93:22:@20216.4]
  wire  RetimeWrapper_133_io_in; // @[package.scala 93:22:@20216.4]
  wire  RetimeWrapper_133_io_out; // @[package.scala 93:22:@20216.4]
  wire  RetimeWrapper_134_clock; // @[package.scala 93:22:@20224.4]
  wire  RetimeWrapper_134_reset; // @[package.scala 93:22:@20224.4]
  wire  RetimeWrapper_134_io_flow; // @[package.scala 93:22:@20224.4]
  wire  RetimeWrapper_134_io_in; // @[package.scala 93:22:@20224.4]
  wire  RetimeWrapper_134_io_out; // @[package.scala 93:22:@20224.4]
  wire  RetimeWrapper_135_clock; // @[package.scala 93:22:@20232.4]
  wire  RetimeWrapper_135_reset; // @[package.scala 93:22:@20232.4]
  wire  RetimeWrapper_135_io_flow; // @[package.scala 93:22:@20232.4]
  wire  RetimeWrapper_135_io_in; // @[package.scala 93:22:@20232.4]
  wire  RetimeWrapper_135_io_out; // @[package.scala 93:22:@20232.4]
  wire  RetimeWrapper_136_clock; // @[package.scala 93:22:@20240.4]
  wire  RetimeWrapper_136_reset; // @[package.scala 93:22:@20240.4]
  wire  RetimeWrapper_136_io_flow; // @[package.scala 93:22:@20240.4]
  wire  RetimeWrapper_136_io_in; // @[package.scala 93:22:@20240.4]
  wire  RetimeWrapper_136_io_out; // @[package.scala 93:22:@20240.4]
  wire  RetimeWrapper_137_clock; // @[package.scala 93:22:@20248.4]
  wire  RetimeWrapper_137_reset; // @[package.scala 93:22:@20248.4]
  wire  RetimeWrapper_137_io_flow; // @[package.scala 93:22:@20248.4]
  wire  RetimeWrapper_137_io_in; // @[package.scala 93:22:@20248.4]
  wire  RetimeWrapper_137_io_out; // @[package.scala 93:22:@20248.4]
  wire  RetimeWrapper_138_clock; // @[package.scala 93:22:@20256.4]
  wire  RetimeWrapper_138_reset; // @[package.scala 93:22:@20256.4]
  wire  RetimeWrapper_138_io_flow; // @[package.scala 93:22:@20256.4]
  wire  RetimeWrapper_138_io_in; // @[package.scala 93:22:@20256.4]
  wire  RetimeWrapper_138_io_out; // @[package.scala 93:22:@20256.4]
  wire  RetimeWrapper_139_clock; // @[package.scala 93:22:@20264.4]
  wire  RetimeWrapper_139_reset; // @[package.scala 93:22:@20264.4]
  wire  RetimeWrapper_139_io_flow; // @[package.scala 93:22:@20264.4]
  wire  RetimeWrapper_139_io_in; // @[package.scala 93:22:@20264.4]
  wire  RetimeWrapper_139_io_out; // @[package.scala 93:22:@20264.4]
  wire  RetimeWrapper_140_clock; // @[package.scala 93:22:@20272.4]
  wire  RetimeWrapper_140_reset; // @[package.scala 93:22:@20272.4]
  wire  RetimeWrapper_140_io_flow; // @[package.scala 93:22:@20272.4]
  wire  RetimeWrapper_140_io_in; // @[package.scala 93:22:@20272.4]
  wire  RetimeWrapper_140_io_out; // @[package.scala 93:22:@20272.4]
  wire  RetimeWrapper_141_clock; // @[package.scala 93:22:@20280.4]
  wire  RetimeWrapper_141_reset; // @[package.scala 93:22:@20280.4]
  wire  RetimeWrapper_141_io_flow; // @[package.scala 93:22:@20280.4]
  wire  RetimeWrapper_141_io_in; // @[package.scala 93:22:@20280.4]
  wire  RetimeWrapper_141_io_out; // @[package.scala 93:22:@20280.4]
  wire  RetimeWrapper_142_clock; // @[package.scala 93:22:@20288.4]
  wire  RetimeWrapper_142_reset; // @[package.scala 93:22:@20288.4]
  wire  RetimeWrapper_142_io_flow; // @[package.scala 93:22:@20288.4]
  wire  RetimeWrapper_142_io_in; // @[package.scala 93:22:@20288.4]
  wire  RetimeWrapper_142_io_out; // @[package.scala 93:22:@20288.4]
  wire  RetimeWrapper_143_clock; // @[package.scala 93:22:@20296.4]
  wire  RetimeWrapper_143_reset; // @[package.scala 93:22:@20296.4]
  wire  RetimeWrapper_143_io_flow; // @[package.scala 93:22:@20296.4]
  wire  RetimeWrapper_143_io_in; // @[package.scala 93:22:@20296.4]
  wire  RetimeWrapper_143_io_out; // @[package.scala 93:22:@20296.4]
  wire  RetimeWrapper_144_clock; // @[package.scala 93:22:@20352.4]
  wire  RetimeWrapper_144_reset; // @[package.scala 93:22:@20352.4]
  wire  RetimeWrapper_144_io_flow; // @[package.scala 93:22:@20352.4]
  wire  RetimeWrapper_144_io_in; // @[package.scala 93:22:@20352.4]
  wire  RetimeWrapper_144_io_out; // @[package.scala 93:22:@20352.4]
  wire  RetimeWrapper_145_clock; // @[package.scala 93:22:@20360.4]
  wire  RetimeWrapper_145_reset; // @[package.scala 93:22:@20360.4]
  wire  RetimeWrapper_145_io_flow; // @[package.scala 93:22:@20360.4]
  wire  RetimeWrapper_145_io_in; // @[package.scala 93:22:@20360.4]
  wire  RetimeWrapper_145_io_out; // @[package.scala 93:22:@20360.4]
  wire  RetimeWrapper_146_clock; // @[package.scala 93:22:@20368.4]
  wire  RetimeWrapper_146_reset; // @[package.scala 93:22:@20368.4]
  wire  RetimeWrapper_146_io_flow; // @[package.scala 93:22:@20368.4]
  wire  RetimeWrapper_146_io_in; // @[package.scala 93:22:@20368.4]
  wire  RetimeWrapper_146_io_out; // @[package.scala 93:22:@20368.4]
  wire  RetimeWrapper_147_clock; // @[package.scala 93:22:@20376.4]
  wire  RetimeWrapper_147_reset; // @[package.scala 93:22:@20376.4]
  wire  RetimeWrapper_147_io_flow; // @[package.scala 93:22:@20376.4]
  wire  RetimeWrapper_147_io_in; // @[package.scala 93:22:@20376.4]
  wire  RetimeWrapper_147_io_out; // @[package.scala 93:22:@20376.4]
  wire  RetimeWrapper_148_clock; // @[package.scala 93:22:@20384.4]
  wire  RetimeWrapper_148_reset; // @[package.scala 93:22:@20384.4]
  wire  RetimeWrapper_148_io_flow; // @[package.scala 93:22:@20384.4]
  wire  RetimeWrapper_148_io_in; // @[package.scala 93:22:@20384.4]
  wire  RetimeWrapper_148_io_out; // @[package.scala 93:22:@20384.4]
  wire  RetimeWrapper_149_clock; // @[package.scala 93:22:@20392.4]
  wire  RetimeWrapper_149_reset; // @[package.scala 93:22:@20392.4]
  wire  RetimeWrapper_149_io_flow; // @[package.scala 93:22:@20392.4]
  wire  RetimeWrapper_149_io_in; // @[package.scala 93:22:@20392.4]
  wire  RetimeWrapper_149_io_out; // @[package.scala 93:22:@20392.4]
  wire  RetimeWrapper_150_clock; // @[package.scala 93:22:@20400.4]
  wire  RetimeWrapper_150_reset; // @[package.scala 93:22:@20400.4]
  wire  RetimeWrapper_150_io_flow; // @[package.scala 93:22:@20400.4]
  wire  RetimeWrapper_150_io_in; // @[package.scala 93:22:@20400.4]
  wire  RetimeWrapper_150_io_out; // @[package.scala 93:22:@20400.4]
  wire  RetimeWrapper_151_clock; // @[package.scala 93:22:@20408.4]
  wire  RetimeWrapper_151_reset; // @[package.scala 93:22:@20408.4]
  wire  RetimeWrapper_151_io_flow; // @[package.scala 93:22:@20408.4]
  wire  RetimeWrapper_151_io_in; // @[package.scala 93:22:@20408.4]
  wire  RetimeWrapper_151_io_out; // @[package.scala 93:22:@20408.4]
  wire  RetimeWrapper_152_clock; // @[package.scala 93:22:@20416.4]
  wire  RetimeWrapper_152_reset; // @[package.scala 93:22:@20416.4]
  wire  RetimeWrapper_152_io_flow; // @[package.scala 93:22:@20416.4]
  wire  RetimeWrapper_152_io_in; // @[package.scala 93:22:@20416.4]
  wire  RetimeWrapper_152_io_out; // @[package.scala 93:22:@20416.4]
  wire  RetimeWrapper_153_clock; // @[package.scala 93:22:@20424.4]
  wire  RetimeWrapper_153_reset; // @[package.scala 93:22:@20424.4]
  wire  RetimeWrapper_153_io_flow; // @[package.scala 93:22:@20424.4]
  wire  RetimeWrapper_153_io_in; // @[package.scala 93:22:@20424.4]
  wire  RetimeWrapper_153_io_out; // @[package.scala 93:22:@20424.4]
  wire  RetimeWrapper_154_clock; // @[package.scala 93:22:@20432.4]
  wire  RetimeWrapper_154_reset; // @[package.scala 93:22:@20432.4]
  wire  RetimeWrapper_154_io_flow; // @[package.scala 93:22:@20432.4]
  wire  RetimeWrapper_154_io_in; // @[package.scala 93:22:@20432.4]
  wire  RetimeWrapper_154_io_out; // @[package.scala 93:22:@20432.4]
  wire  RetimeWrapper_155_clock; // @[package.scala 93:22:@20440.4]
  wire  RetimeWrapper_155_reset; // @[package.scala 93:22:@20440.4]
  wire  RetimeWrapper_155_io_flow; // @[package.scala 93:22:@20440.4]
  wire  RetimeWrapper_155_io_in; // @[package.scala 93:22:@20440.4]
  wire  RetimeWrapper_155_io_out; // @[package.scala 93:22:@20440.4]
  wire  RetimeWrapper_156_clock; // @[package.scala 93:22:@20496.4]
  wire  RetimeWrapper_156_reset; // @[package.scala 93:22:@20496.4]
  wire  RetimeWrapper_156_io_flow; // @[package.scala 93:22:@20496.4]
  wire  RetimeWrapper_156_io_in; // @[package.scala 93:22:@20496.4]
  wire  RetimeWrapper_156_io_out; // @[package.scala 93:22:@20496.4]
  wire  RetimeWrapper_157_clock; // @[package.scala 93:22:@20504.4]
  wire  RetimeWrapper_157_reset; // @[package.scala 93:22:@20504.4]
  wire  RetimeWrapper_157_io_flow; // @[package.scala 93:22:@20504.4]
  wire  RetimeWrapper_157_io_in; // @[package.scala 93:22:@20504.4]
  wire  RetimeWrapper_157_io_out; // @[package.scala 93:22:@20504.4]
  wire  RetimeWrapper_158_clock; // @[package.scala 93:22:@20512.4]
  wire  RetimeWrapper_158_reset; // @[package.scala 93:22:@20512.4]
  wire  RetimeWrapper_158_io_flow; // @[package.scala 93:22:@20512.4]
  wire  RetimeWrapper_158_io_in; // @[package.scala 93:22:@20512.4]
  wire  RetimeWrapper_158_io_out; // @[package.scala 93:22:@20512.4]
  wire  RetimeWrapper_159_clock; // @[package.scala 93:22:@20520.4]
  wire  RetimeWrapper_159_reset; // @[package.scala 93:22:@20520.4]
  wire  RetimeWrapper_159_io_flow; // @[package.scala 93:22:@20520.4]
  wire  RetimeWrapper_159_io_in; // @[package.scala 93:22:@20520.4]
  wire  RetimeWrapper_159_io_out; // @[package.scala 93:22:@20520.4]
  wire  RetimeWrapper_160_clock; // @[package.scala 93:22:@20528.4]
  wire  RetimeWrapper_160_reset; // @[package.scala 93:22:@20528.4]
  wire  RetimeWrapper_160_io_flow; // @[package.scala 93:22:@20528.4]
  wire  RetimeWrapper_160_io_in; // @[package.scala 93:22:@20528.4]
  wire  RetimeWrapper_160_io_out; // @[package.scala 93:22:@20528.4]
  wire  RetimeWrapper_161_clock; // @[package.scala 93:22:@20536.4]
  wire  RetimeWrapper_161_reset; // @[package.scala 93:22:@20536.4]
  wire  RetimeWrapper_161_io_flow; // @[package.scala 93:22:@20536.4]
  wire  RetimeWrapper_161_io_in; // @[package.scala 93:22:@20536.4]
  wire  RetimeWrapper_161_io_out; // @[package.scala 93:22:@20536.4]
  wire  RetimeWrapper_162_clock; // @[package.scala 93:22:@20544.4]
  wire  RetimeWrapper_162_reset; // @[package.scala 93:22:@20544.4]
  wire  RetimeWrapper_162_io_flow; // @[package.scala 93:22:@20544.4]
  wire  RetimeWrapper_162_io_in; // @[package.scala 93:22:@20544.4]
  wire  RetimeWrapper_162_io_out; // @[package.scala 93:22:@20544.4]
  wire  RetimeWrapper_163_clock; // @[package.scala 93:22:@20552.4]
  wire  RetimeWrapper_163_reset; // @[package.scala 93:22:@20552.4]
  wire  RetimeWrapper_163_io_flow; // @[package.scala 93:22:@20552.4]
  wire  RetimeWrapper_163_io_in; // @[package.scala 93:22:@20552.4]
  wire  RetimeWrapper_163_io_out; // @[package.scala 93:22:@20552.4]
  wire  RetimeWrapper_164_clock; // @[package.scala 93:22:@20560.4]
  wire  RetimeWrapper_164_reset; // @[package.scala 93:22:@20560.4]
  wire  RetimeWrapper_164_io_flow; // @[package.scala 93:22:@20560.4]
  wire  RetimeWrapper_164_io_in; // @[package.scala 93:22:@20560.4]
  wire  RetimeWrapper_164_io_out; // @[package.scala 93:22:@20560.4]
  wire  RetimeWrapper_165_clock; // @[package.scala 93:22:@20568.4]
  wire  RetimeWrapper_165_reset; // @[package.scala 93:22:@20568.4]
  wire  RetimeWrapper_165_io_flow; // @[package.scala 93:22:@20568.4]
  wire  RetimeWrapper_165_io_in; // @[package.scala 93:22:@20568.4]
  wire  RetimeWrapper_165_io_out; // @[package.scala 93:22:@20568.4]
  wire  RetimeWrapper_166_clock; // @[package.scala 93:22:@20576.4]
  wire  RetimeWrapper_166_reset; // @[package.scala 93:22:@20576.4]
  wire  RetimeWrapper_166_io_flow; // @[package.scala 93:22:@20576.4]
  wire  RetimeWrapper_166_io_in; // @[package.scala 93:22:@20576.4]
  wire  RetimeWrapper_166_io_out; // @[package.scala 93:22:@20576.4]
  wire  RetimeWrapper_167_clock; // @[package.scala 93:22:@20584.4]
  wire  RetimeWrapper_167_reset; // @[package.scala 93:22:@20584.4]
  wire  RetimeWrapper_167_io_flow; // @[package.scala 93:22:@20584.4]
  wire  RetimeWrapper_167_io_in; // @[package.scala 93:22:@20584.4]
  wire  RetimeWrapper_167_io_out; // @[package.scala 93:22:@20584.4]
  wire  RetimeWrapper_168_clock; // @[package.scala 93:22:@20640.4]
  wire  RetimeWrapper_168_reset; // @[package.scala 93:22:@20640.4]
  wire  RetimeWrapper_168_io_flow; // @[package.scala 93:22:@20640.4]
  wire  RetimeWrapper_168_io_in; // @[package.scala 93:22:@20640.4]
  wire  RetimeWrapper_168_io_out; // @[package.scala 93:22:@20640.4]
  wire  RetimeWrapper_169_clock; // @[package.scala 93:22:@20648.4]
  wire  RetimeWrapper_169_reset; // @[package.scala 93:22:@20648.4]
  wire  RetimeWrapper_169_io_flow; // @[package.scala 93:22:@20648.4]
  wire  RetimeWrapper_169_io_in; // @[package.scala 93:22:@20648.4]
  wire  RetimeWrapper_169_io_out; // @[package.scala 93:22:@20648.4]
  wire  RetimeWrapper_170_clock; // @[package.scala 93:22:@20656.4]
  wire  RetimeWrapper_170_reset; // @[package.scala 93:22:@20656.4]
  wire  RetimeWrapper_170_io_flow; // @[package.scala 93:22:@20656.4]
  wire  RetimeWrapper_170_io_in; // @[package.scala 93:22:@20656.4]
  wire  RetimeWrapper_170_io_out; // @[package.scala 93:22:@20656.4]
  wire  RetimeWrapper_171_clock; // @[package.scala 93:22:@20664.4]
  wire  RetimeWrapper_171_reset; // @[package.scala 93:22:@20664.4]
  wire  RetimeWrapper_171_io_flow; // @[package.scala 93:22:@20664.4]
  wire  RetimeWrapper_171_io_in; // @[package.scala 93:22:@20664.4]
  wire  RetimeWrapper_171_io_out; // @[package.scala 93:22:@20664.4]
  wire  RetimeWrapper_172_clock; // @[package.scala 93:22:@20672.4]
  wire  RetimeWrapper_172_reset; // @[package.scala 93:22:@20672.4]
  wire  RetimeWrapper_172_io_flow; // @[package.scala 93:22:@20672.4]
  wire  RetimeWrapper_172_io_in; // @[package.scala 93:22:@20672.4]
  wire  RetimeWrapper_172_io_out; // @[package.scala 93:22:@20672.4]
  wire  RetimeWrapper_173_clock; // @[package.scala 93:22:@20680.4]
  wire  RetimeWrapper_173_reset; // @[package.scala 93:22:@20680.4]
  wire  RetimeWrapper_173_io_flow; // @[package.scala 93:22:@20680.4]
  wire  RetimeWrapper_173_io_in; // @[package.scala 93:22:@20680.4]
  wire  RetimeWrapper_173_io_out; // @[package.scala 93:22:@20680.4]
  wire  RetimeWrapper_174_clock; // @[package.scala 93:22:@20688.4]
  wire  RetimeWrapper_174_reset; // @[package.scala 93:22:@20688.4]
  wire  RetimeWrapper_174_io_flow; // @[package.scala 93:22:@20688.4]
  wire  RetimeWrapper_174_io_in; // @[package.scala 93:22:@20688.4]
  wire  RetimeWrapper_174_io_out; // @[package.scala 93:22:@20688.4]
  wire  RetimeWrapper_175_clock; // @[package.scala 93:22:@20696.4]
  wire  RetimeWrapper_175_reset; // @[package.scala 93:22:@20696.4]
  wire  RetimeWrapper_175_io_flow; // @[package.scala 93:22:@20696.4]
  wire  RetimeWrapper_175_io_in; // @[package.scala 93:22:@20696.4]
  wire  RetimeWrapper_175_io_out; // @[package.scala 93:22:@20696.4]
  wire  RetimeWrapper_176_clock; // @[package.scala 93:22:@20704.4]
  wire  RetimeWrapper_176_reset; // @[package.scala 93:22:@20704.4]
  wire  RetimeWrapper_176_io_flow; // @[package.scala 93:22:@20704.4]
  wire  RetimeWrapper_176_io_in; // @[package.scala 93:22:@20704.4]
  wire  RetimeWrapper_176_io_out; // @[package.scala 93:22:@20704.4]
  wire  RetimeWrapper_177_clock; // @[package.scala 93:22:@20712.4]
  wire  RetimeWrapper_177_reset; // @[package.scala 93:22:@20712.4]
  wire  RetimeWrapper_177_io_flow; // @[package.scala 93:22:@20712.4]
  wire  RetimeWrapper_177_io_in; // @[package.scala 93:22:@20712.4]
  wire  RetimeWrapper_177_io_out; // @[package.scala 93:22:@20712.4]
  wire  RetimeWrapper_178_clock; // @[package.scala 93:22:@20720.4]
  wire  RetimeWrapper_178_reset; // @[package.scala 93:22:@20720.4]
  wire  RetimeWrapper_178_io_flow; // @[package.scala 93:22:@20720.4]
  wire  RetimeWrapper_178_io_in; // @[package.scala 93:22:@20720.4]
  wire  RetimeWrapper_178_io_out; // @[package.scala 93:22:@20720.4]
  wire  RetimeWrapper_179_clock; // @[package.scala 93:22:@20728.4]
  wire  RetimeWrapper_179_reset; // @[package.scala 93:22:@20728.4]
  wire  RetimeWrapper_179_io_flow; // @[package.scala 93:22:@20728.4]
  wire  RetimeWrapper_179_io_in; // @[package.scala 93:22:@20728.4]
  wire  RetimeWrapper_179_io_out; // @[package.scala 93:22:@20728.4]
  wire  RetimeWrapper_180_clock; // @[package.scala 93:22:@20784.4]
  wire  RetimeWrapper_180_reset; // @[package.scala 93:22:@20784.4]
  wire  RetimeWrapper_180_io_flow; // @[package.scala 93:22:@20784.4]
  wire  RetimeWrapper_180_io_in; // @[package.scala 93:22:@20784.4]
  wire  RetimeWrapper_180_io_out; // @[package.scala 93:22:@20784.4]
  wire  RetimeWrapper_181_clock; // @[package.scala 93:22:@20792.4]
  wire  RetimeWrapper_181_reset; // @[package.scala 93:22:@20792.4]
  wire  RetimeWrapper_181_io_flow; // @[package.scala 93:22:@20792.4]
  wire  RetimeWrapper_181_io_in; // @[package.scala 93:22:@20792.4]
  wire  RetimeWrapper_181_io_out; // @[package.scala 93:22:@20792.4]
  wire  RetimeWrapper_182_clock; // @[package.scala 93:22:@20800.4]
  wire  RetimeWrapper_182_reset; // @[package.scala 93:22:@20800.4]
  wire  RetimeWrapper_182_io_flow; // @[package.scala 93:22:@20800.4]
  wire  RetimeWrapper_182_io_in; // @[package.scala 93:22:@20800.4]
  wire  RetimeWrapper_182_io_out; // @[package.scala 93:22:@20800.4]
  wire  RetimeWrapper_183_clock; // @[package.scala 93:22:@20808.4]
  wire  RetimeWrapper_183_reset; // @[package.scala 93:22:@20808.4]
  wire  RetimeWrapper_183_io_flow; // @[package.scala 93:22:@20808.4]
  wire  RetimeWrapper_183_io_in; // @[package.scala 93:22:@20808.4]
  wire  RetimeWrapper_183_io_out; // @[package.scala 93:22:@20808.4]
  wire  RetimeWrapper_184_clock; // @[package.scala 93:22:@20816.4]
  wire  RetimeWrapper_184_reset; // @[package.scala 93:22:@20816.4]
  wire  RetimeWrapper_184_io_flow; // @[package.scala 93:22:@20816.4]
  wire  RetimeWrapper_184_io_in; // @[package.scala 93:22:@20816.4]
  wire  RetimeWrapper_184_io_out; // @[package.scala 93:22:@20816.4]
  wire  RetimeWrapper_185_clock; // @[package.scala 93:22:@20824.4]
  wire  RetimeWrapper_185_reset; // @[package.scala 93:22:@20824.4]
  wire  RetimeWrapper_185_io_flow; // @[package.scala 93:22:@20824.4]
  wire  RetimeWrapper_185_io_in; // @[package.scala 93:22:@20824.4]
  wire  RetimeWrapper_185_io_out; // @[package.scala 93:22:@20824.4]
  wire  RetimeWrapper_186_clock; // @[package.scala 93:22:@20832.4]
  wire  RetimeWrapper_186_reset; // @[package.scala 93:22:@20832.4]
  wire  RetimeWrapper_186_io_flow; // @[package.scala 93:22:@20832.4]
  wire  RetimeWrapper_186_io_in; // @[package.scala 93:22:@20832.4]
  wire  RetimeWrapper_186_io_out; // @[package.scala 93:22:@20832.4]
  wire  RetimeWrapper_187_clock; // @[package.scala 93:22:@20840.4]
  wire  RetimeWrapper_187_reset; // @[package.scala 93:22:@20840.4]
  wire  RetimeWrapper_187_io_flow; // @[package.scala 93:22:@20840.4]
  wire  RetimeWrapper_187_io_in; // @[package.scala 93:22:@20840.4]
  wire  RetimeWrapper_187_io_out; // @[package.scala 93:22:@20840.4]
  wire  RetimeWrapper_188_clock; // @[package.scala 93:22:@20848.4]
  wire  RetimeWrapper_188_reset; // @[package.scala 93:22:@20848.4]
  wire  RetimeWrapper_188_io_flow; // @[package.scala 93:22:@20848.4]
  wire  RetimeWrapper_188_io_in; // @[package.scala 93:22:@20848.4]
  wire  RetimeWrapper_188_io_out; // @[package.scala 93:22:@20848.4]
  wire  RetimeWrapper_189_clock; // @[package.scala 93:22:@20856.4]
  wire  RetimeWrapper_189_reset; // @[package.scala 93:22:@20856.4]
  wire  RetimeWrapper_189_io_flow; // @[package.scala 93:22:@20856.4]
  wire  RetimeWrapper_189_io_in; // @[package.scala 93:22:@20856.4]
  wire  RetimeWrapper_189_io_out; // @[package.scala 93:22:@20856.4]
  wire  RetimeWrapper_190_clock; // @[package.scala 93:22:@20864.4]
  wire  RetimeWrapper_190_reset; // @[package.scala 93:22:@20864.4]
  wire  RetimeWrapper_190_io_flow; // @[package.scala 93:22:@20864.4]
  wire  RetimeWrapper_190_io_in; // @[package.scala 93:22:@20864.4]
  wire  RetimeWrapper_190_io_out; // @[package.scala 93:22:@20864.4]
  wire  RetimeWrapper_191_clock; // @[package.scala 93:22:@20872.4]
  wire  RetimeWrapper_191_reset; // @[package.scala 93:22:@20872.4]
  wire  RetimeWrapper_191_io_flow; // @[package.scala 93:22:@20872.4]
  wire  RetimeWrapper_191_io_in; // @[package.scala 93:22:@20872.4]
  wire  RetimeWrapper_191_io_out; // @[package.scala 93:22:@20872.4]
  wire  RetimeWrapper_192_clock; // @[package.scala 93:22:@20928.4]
  wire  RetimeWrapper_192_reset; // @[package.scala 93:22:@20928.4]
  wire  RetimeWrapper_192_io_flow; // @[package.scala 93:22:@20928.4]
  wire  RetimeWrapper_192_io_in; // @[package.scala 93:22:@20928.4]
  wire  RetimeWrapper_192_io_out; // @[package.scala 93:22:@20928.4]
  wire  RetimeWrapper_193_clock; // @[package.scala 93:22:@20936.4]
  wire  RetimeWrapper_193_reset; // @[package.scala 93:22:@20936.4]
  wire  RetimeWrapper_193_io_flow; // @[package.scala 93:22:@20936.4]
  wire  RetimeWrapper_193_io_in; // @[package.scala 93:22:@20936.4]
  wire  RetimeWrapper_193_io_out; // @[package.scala 93:22:@20936.4]
  wire  RetimeWrapper_194_clock; // @[package.scala 93:22:@20944.4]
  wire  RetimeWrapper_194_reset; // @[package.scala 93:22:@20944.4]
  wire  RetimeWrapper_194_io_flow; // @[package.scala 93:22:@20944.4]
  wire  RetimeWrapper_194_io_in; // @[package.scala 93:22:@20944.4]
  wire  RetimeWrapper_194_io_out; // @[package.scala 93:22:@20944.4]
  wire  RetimeWrapper_195_clock; // @[package.scala 93:22:@20952.4]
  wire  RetimeWrapper_195_reset; // @[package.scala 93:22:@20952.4]
  wire  RetimeWrapper_195_io_flow; // @[package.scala 93:22:@20952.4]
  wire  RetimeWrapper_195_io_in; // @[package.scala 93:22:@20952.4]
  wire  RetimeWrapper_195_io_out; // @[package.scala 93:22:@20952.4]
  wire  RetimeWrapper_196_clock; // @[package.scala 93:22:@20960.4]
  wire  RetimeWrapper_196_reset; // @[package.scala 93:22:@20960.4]
  wire  RetimeWrapper_196_io_flow; // @[package.scala 93:22:@20960.4]
  wire  RetimeWrapper_196_io_in; // @[package.scala 93:22:@20960.4]
  wire  RetimeWrapper_196_io_out; // @[package.scala 93:22:@20960.4]
  wire  RetimeWrapper_197_clock; // @[package.scala 93:22:@20968.4]
  wire  RetimeWrapper_197_reset; // @[package.scala 93:22:@20968.4]
  wire  RetimeWrapper_197_io_flow; // @[package.scala 93:22:@20968.4]
  wire  RetimeWrapper_197_io_in; // @[package.scala 93:22:@20968.4]
  wire  RetimeWrapper_197_io_out; // @[package.scala 93:22:@20968.4]
  wire  RetimeWrapper_198_clock; // @[package.scala 93:22:@20976.4]
  wire  RetimeWrapper_198_reset; // @[package.scala 93:22:@20976.4]
  wire  RetimeWrapper_198_io_flow; // @[package.scala 93:22:@20976.4]
  wire  RetimeWrapper_198_io_in; // @[package.scala 93:22:@20976.4]
  wire  RetimeWrapper_198_io_out; // @[package.scala 93:22:@20976.4]
  wire  RetimeWrapper_199_clock; // @[package.scala 93:22:@20984.4]
  wire  RetimeWrapper_199_reset; // @[package.scala 93:22:@20984.4]
  wire  RetimeWrapper_199_io_flow; // @[package.scala 93:22:@20984.4]
  wire  RetimeWrapper_199_io_in; // @[package.scala 93:22:@20984.4]
  wire  RetimeWrapper_199_io_out; // @[package.scala 93:22:@20984.4]
  wire  RetimeWrapper_200_clock; // @[package.scala 93:22:@20992.4]
  wire  RetimeWrapper_200_reset; // @[package.scala 93:22:@20992.4]
  wire  RetimeWrapper_200_io_flow; // @[package.scala 93:22:@20992.4]
  wire  RetimeWrapper_200_io_in; // @[package.scala 93:22:@20992.4]
  wire  RetimeWrapper_200_io_out; // @[package.scala 93:22:@20992.4]
  wire  RetimeWrapper_201_clock; // @[package.scala 93:22:@21000.4]
  wire  RetimeWrapper_201_reset; // @[package.scala 93:22:@21000.4]
  wire  RetimeWrapper_201_io_flow; // @[package.scala 93:22:@21000.4]
  wire  RetimeWrapper_201_io_in; // @[package.scala 93:22:@21000.4]
  wire  RetimeWrapper_201_io_out; // @[package.scala 93:22:@21000.4]
  wire  RetimeWrapper_202_clock; // @[package.scala 93:22:@21008.4]
  wire  RetimeWrapper_202_reset; // @[package.scala 93:22:@21008.4]
  wire  RetimeWrapper_202_io_flow; // @[package.scala 93:22:@21008.4]
  wire  RetimeWrapper_202_io_in; // @[package.scala 93:22:@21008.4]
  wire  RetimeWrapper_202_io_out; // @[package.scala 93:22:@21008.4]
  wire  RetimeWrapper_203_clock; // @[package.scala 93:22:@21016.4]
  wire  RetimeWrapper_203_reset; // @[package.scala 93:22:@21016.4]
  wire  RetimeWrapper_203_io_flow; // @[package.scala 93:22:@21016.4]
  wire  RetimeWrapper_203_io_in; // @[package.scala 93:22:@21016.4]
  wire  RetimeWrapper_203_io_out; // @[package.scala 93:22:@21016.4]
  wire  RetimeWrapper_204_clock; // @[package.scala 93:22:@21072.4]
  wire  RetimeWrapper_204_reset; // @[package.scala 93:22:@21072.4]
  wire  RetimeWrapper_204_io_flow; // @[package.scala 93:22:@21072.4]
  wire  RetimeWrapper_204_io_in; // @[package.scala 93:22:@21072.4]
  wire  RetimeWrapper_204_io_out; // @[package.scala 93:22:@21072.4]
  wire  RetimeWrapper_205_clock; // @[package.scala 93:22:@21080.4]
  wire  RetimeWrapper_205_reset; // @[package.scala 93:22:@21080.4]
  wire  RetimeWrapper_205_io_flow; // @[package.scala 93:22:@21080.4]
  wire  RetimeWrapper_205_io_in; // @[package.scala 93:22:@21080.4]
  wire  RetimeWrapper_205_io_out; // @[package.scala 93:22:@21080.4]
  wire  RetimeWrapper_206_clock; // @[package.scala 93:22:@21088.4]
  wire  RetimeWrapper_206_reset; // @[package.scala 93:22:@21088.4]
  wire  RetimeWrapper_206_io_flow; // @[package.scala 93:22:@21088.4]
  wire  RetimeWrapper_206_io_in; // @[package.scala 93:22:@21088.4]
  wire  RetimeWrapper_206_io_out; // @[package.scala 93:22:@21088.4]
  wire  RetimeWrapper_207_clock; // @[package.scala 93:22:@21096.4]
  wire  RetimeWrapper_207_reset; // @[package.scala 93:22:@21096.4]
  wire  RetimeWrapper_207_io_flow; // @[package.scala 93:22:@21096.4]
  wire  RetimeWrapper_207_io_in; // @[package.scala 93:22:@21096.4]
  wire  RetimeWrapper_207_io_out; // @[package.scala 93:22:@21096.4]
  wire  RetimeWrapper_208_clock; // @[package.scala 93:22:@21104.4]
  wire  RetimeWrapper_208_reset; // @[package.scala 93:22:@21104.4]
  wire  RetimeWrapper_208_io_flow; // @[package.scala 93:22:@21104.4]
  wire  RetimeWrapper_208_io_in; // @[package.scala 93:22:@21104.4]
  wire  RetimeWrapper_208_io_out; // @[package.scala 93:22:@21104.4]
  wire  RetimeWrapper_209_clock; // @[package.scala 93:22:@21112.4]
  wire  RetimeWrapper_209_reset; // @[package.scala 93:22:@21112.4]
  wire  RetimeWrapper_209_io_flow; // @[package.scala 93:22:@21112.4]
  wire  RetimeWrapper_209_io_in; // @[package.scala 93:22:@21112.4]
  wire  RetimeWrapper_209_io_out; // @[package.scala 93:22:@21112.4]
  wire  RetimeWrapper_210_clock; // @[package.scala 93:22:@21120.4]
  wire  RetimeWrapper_210_reset; // @[package.scala 93:22:@21120.4]
  wire  RetimeWrapper_210_io_flow; // @[package.scala 93:22:@21120.4]
  wire  RetimeWrapper_210_io_in; // @[package.scala 93:22:@21120.4]
  wire  RetimeWrapper_210_io_out; // @[package.scala 93:22:@21120.4]
  wire  RetimeWrapper_211_clock; // @[package.scala 93:22:@21128.4]
  wire  RetimeWrapper_211_reset; // @[package.scala 93:22:@21128.4]
  wire  RetimeWrapper_211_io_flow; // @[package.scala 93:22:@21128.4]
  wire  RetimeWrapper_211_io_in; // @[package.scala 93:22:@21128.4]
  wire  RetimeWrapper_211_io_out; // @[package.scala 93:22:@21128.4]
  wire  RetimeWrapper_212_clock; // @[package.scala 93:22:@21136.4]
  wire  RetimeWrapper_212_reset; // @[package.scala 93:22:@21136.4]
  wire  RetimeWrapper_212_io_flow; // @[package.scala 93:22:@21136.4]
  wire  RetimeWrapper_212_io_in; // @[package.scala 93:22:@21136.4]
  wire  RetimeWrapper_212_io_out; // @[package.scala 93:22:@21136.4]
  wire  RetimeWrapper_213_clock; // @[package.scala 93:22:@21144.4]
  wire  RetimeWrapper_213_reset; // @[package.scala 93:22:@21144.4]
  wire  RetimeWrapper_213_io_flow; // @[package.scala 93:22:@21144.4]
  wire  RetimeWrapper_213_io_in; // @[package.scala 93:22:@21144.4]
  wire  RetimeWrapper_213_io_out; // @[package.scala 93:22:@21144.4]
  wire  RetimeWrapper_214_clock; // @[package.scala 93:22:@21152.4]
  wire  RetimeWrapper_214_reset; // @[package.scala 93:22:@21152.4]
  wire  RetimeWrapper_214_io_flow; // @[package.scala 93:22:@21152.4]
  wire  RetimeWrapper_214_io_in; // @[package.scala 93:22:@21152.4]
  wire  RetimeWrapper_214_io_out; // @[package.scala 93:22:@21152.4]
  wire  RetimeWrapper_215_clock; // @[package.scala 93:22:@21160.4]
  wire  RetimeWrapper_215_reset; // @[package.scala 93:22:@21160.4]
  wire  RetimeWrapper_215_io_flow; // @[package.scala 93:22:@21160.4]
  wire  RetimeWrapper_215_io_in; // @[package.scala 93:22:@21160.4]
  wire  RetimeWrapper_215_io_out; // @[package.scala 93:22:@21160.4]
  wire  _T_700; // @[MemPrimitives.scala 82:210:@15995.4]
  wire  _T_702; // @[MemPrimitives.scala 82:210:@15996.4]
  wire  _T_703; // @[MemPrimitives.scala 82:228:@15997.4]
  wire  _T_704; // @[MemPrimitives.scala 83:102:@15998.4]
  wire  _T_706; // @[MemPrimitives.scala 82:210:@15999.4]
  wire  _T_708; // @[MemPrimitives.scala 82:210:@16000.4]
  wire  _T_709; // @[MemPrimitives.scala 82:228:@16001.4]
  wire  _T_710; // @[MemPrimitives.scala 83:102:@16002.4]
  wire [16:0] _T_712; // @[Cat.scala 30:58:@16004.4]
  wire [16:0] _T_714; // @[Cat.scala 30:58:@16006.4]
  wire [16:0] _T_715; // @[Mux.scala 31:69:@16007.4]
  wire  _T_720; // @[MemPrimitives.scala 82:210:@16014.4]
  wire  _T_722; // @[MemPrimitives.scala 82:210:@16015.4]
  wire  _T_723; // @[MemPrimitives.scala 82:228:@16016.4]
  wire  _T_724; // @[MemPrimitives.scala 83:102:@16017.4]
  wire  _T_726; // @[MemPrimitives.scala 82:210:@16018.4]
  wire  _T_728; // @[MemPrimitives.scala 82:210:@16019.4]
  wire  _T_729; // @[MemPrimitives.scala 82:228:@16020.4]
  wire  _T_730; // @[MemPrimitives.scala 83:102:@16021.4]
  wire [16:0] _T_732; // @[Cat.scala 30:58:@16023.4]
  wire [16:0] _T_734; // @[Cat.scala 30:58:@16025.4]
  wire [16:0] _T_735; // @[Mux.scala 31:69:@16026.4]
  wire  _T_742; // @[MemPrimitives.scala 82:210:@16034.4]
  wire  _T_743; // @[MemPrimitives.scala 82:228:@16035.4]
  wire  _T_744; // @[MemPrimitives.scala 83:102:@16036.4]
  wire  _T_748; // @[MemPrimitives.scala 82:210:@16038.4]
  wire  _T_749; // @[MemPrimitives.scala 82:228:@16039.4]
  wire  _T_750; // @[MemPrimitives.scala 83:102:@16040.4]
  wire [16:0] _T_752; // @[Cat.scala 30:58:@16042.4]
  wire [16:0] _T_754; // @[Cat.scala 30:58:@16044.4]
  wire [16:0] _T_755; // @[Mux.scala 31:69:@16045.4]
  wire  _T_762; // @[MemPrimitives.scala 82:210:@16053.4]
  wire  _T_763; // @[MemPrimitives.scala 82:228:@16054.4]
  wire  _T_764; // @[MemPrimitives.scala 83:102:@16055.4]
  wire  _T_768; // @[MemPrimitives.scala 82:210:@16057.4]
  wire  _T_769; // @[MemPrimitives.scala 82:228:@16058.4]
  wire  _T_770; // @[MemPrimitives.scala 83:102:@16059.4]
  wire [16:0] _T_772; // @[Cat.scala 30:58:@16061.4]
  wire [16:0] _T_774; // @[Cat.scala 30:58:@16063.4]
  wire [16:0] _T_775; // @[Mux.scala 31:69:@16064.4]
  wire  _T_782; // @[MemPrimitives.scala 82:210:@16072.4]
  wire  _T_783; // @[MemPrimitives.scala 82:228:@16073.4]
  wire  _T_784; // @[MemPrimitives.scala 83:102:@16074.4]
  wire  _T_788; // @[MemPrimitives.scala 82:210:@16076.4]
  wire  _T_789; // @[MemPrimitives.scala 82:228:@16077.4]
  wire  _T_790; // @[MemPrimitives.scala 83:102:@16078.4]
  wire [16:0] _T_792; // @[Cat.scala 30:58:@16080.4]
  wire [16:0] _T_794; // @[Cat.scala 30:58:@16082.4]
  wire [16:0] _T_795; // @[Mux.scala 31:69:@16083.4]
  wire  _T_802; // @[MemPrimitives.scala 82:210:@16091.4]
  wire  _T_803; // @[MemPrimitives.scala 82:228:@16092.4]
  wire  _T_804; // @[MemPrimitives.scala 83:102:@16093.4]
  wire  _T_808; // @[MemPrimitives.scala 82:210:@16095.4]
  wire  _T_809; // @[MemPrimitives.scala 82:228:@16096.4]
  wire  _T_810; // @[MemPrimitives.scala 83:102:@16097.4]
  wire [16:0] _T_812; // @[Cat.scala 30:58:@16099.4]
  wire [16:0] _T_814; // @[Cat.scala 30:58:@16101.4]
  wire [16:0] _T_815; // @[Mux.scala 31:69:@16102.4]
  wire  _T_820; // @[MemPrimitives.scala 82:210:@16109.4]
  wire  _T_823; // @[MemPrimitives.scala 82:228:@16111.4]
  wire  _T_824; // @[MemPrimitives.scala 83:102:@16112.4]
  wire  _T_826; // @[MemPrimitives.scala 82:210:@16113.4]
  wire  _T_829; // @[MemPrimitives.scala 82:228:@16115.4]
  wire  _T_830; // @[MemPrimitives.scala 83:102:@16116.4]
  wire [16:0] _T_832; // @[Cat.scala 30:58:@16118.4]
  wire [16:0] _T_834; // @[Cat.scala 30:58:@16120.4]
  wire [16:0] _T_835; // @[Mux.scala 31:69:@16121.4]
  wire  _T_840; // @[MemPrimitives.scala 82:210:@16128.4]
  wire  _T_843; // @[MemPrimitives.scala 82:228:@16130.4]
  wire  _T_844; // @[MemPrimitives.scala 83:102:@16131.4]
  wire  _T_846; // @[MemPrimitives.scala 82:210:@16132.4]
  wire  _T_849; // @[MemPrimitives.scala 82:228:@16134.4]
  wire  _T_850; // @[MemPrimitives.scala 83:102:@16135.4]
  wire [16:0] _T_852; // @[Cat.scala 30:58:@16137.4]
  wire [16:0] _T_854; // @[Cat.scala 30:58:@16139.4]
  wire [16:0] _T_855; // @[Mux.scala 31:69:@16140.4]
  wire  _T_863; // @[MemPrimitives.scala 82:228:@16149.4]
  wire  _T_864; // @[MemPrimitives.scala 83:102:@16150.4]
  wire  _T_869; // @[MemPrimitives.scala 82:228:@16153.4]
  wire  _T_870; // @[MemPrimitives.scala 83:102:@16154.4]
  wire [16:0] _T_872; // @[Cat.scala 30:58:@16156.4]
  wire [16:0] _T_874; // @[Cat.scala 30:58:@16158.4]
  wire [16:0] _T_875; // @[Mux.scala 31:69:@16159.4]
  wire  _T_883; // @[MemPrimitives.scala 82:228:@16168.4]
  wire  _T_884; // @[MemPrimitives.scala 83:102:@16169.4]
  wire  _T_889; // @[MemPrimitives.scala 82:228:@16172.4]
  wire  _T_890; // @[MemPrimitives.scala 83:102:@16173.4]
  wire [16:0] _T_892; // @[Cat.scala 30:58:@16175.4]
  wire [16:0] _T_894; // @[Cat.scala 30:58:@16177.4]
  wire [16:0] _T_895; // @[Mux.scala 31:69:@16178.4]
  wire  _T_903; // @[MemPrimitives.scala 82:228:@16187.4]
  wire  _T_904; // @[MemPrimitives.scala 83:102:@16188.4]
  wire  _T_909; // @[MemPrimitives.scala 82:228:@16191.4]
  wire  _T_910; // @[MemPrimitives.scala 83:102:@16192.4]
  wire [16:0] _T_912; // @[Cat.scala 30:58:@16194.4]
  wire [16:0] _T_914; // @[Cat.scala 30:58:@16196.4]
  wire [16:0] _T_915; // @[Mux.scala 31:69:@16197.4]
  wire  _T_923; // @[MemPrimitives.scala 82:228:@16206.4]
  wire  _T_924; // @[MemPrimitives.scala 83:102:@16207.4]
  wire  _T_929; // @[MemPrimitives.scala 82:228:@16210.4]
  wire  _T_930; // @[MemPrimitives.scala 83:102:@16211.4]
  wire [16:0] _T_932; // @[Cat.scala 30:58:@16213.4]
  wire [16:0] _T_934; // @[Cat.scala 30:58:@16215.4]
  wire [16:0] _T_935; // @[Mux.scala 31:69:@16216.4]
  wire  _T_940; // @[MemPrimitives.scala 82:210:@16223.4]
  wire  _T_943; // @[MemPrimitives.scala 82:228:@16225.4]
  wire  _T_944; // @[MemPrimitives.scala 83:102:@16226.4]
  wire  _T_946; // @[MemPrimitives.scala 82:210:@16227.4]
  wire  _T_949; // @[MemPrimitives.scala 82:228:@16229.4]
  wire  _T_950; // @[MemPrimitives.scala 83:102:@16230.4]
  wire [16:0] _T_952; // @[Cat.scala 30:58:@16232.4]
  wire [16:0] _T_954; // @[Cat.scala 30:58:@16234.4]
  wire [16:0] _T_955; // @[Mux.scala 31:69:@16235.4]
  wire  _T_960; // @[MemPrimitives.scala 82:210:@16242.4]
  wire  _T_963; // @[MemPrimitives.scala 82:228:@16244.4]
  wire  _T_964; // @[MemPrimitives.scala 83:102:@16245.4]
  wire  _T_966; // @[MemPrimitives.scala 82:210:@16246.4]
  wire  _T_969; // @[MemPrimitives.scala 82:228:@16248.4]
  wire  _T_970; // @[MemPrimitives.scala 83:102:@16249.4]
  wire [16:0] _T_972; // @[Cat.scala 30:58:@16251.4]
  wire [16:0] _T_974; // @[Cat.scala 30:58:@16253.4]
  wire [16:0] _T_975; // @[Mux.scala 31:69:@16254.4]
  wire  _T_983; // @[MemPrimitives.scala 82:228:@16263.4]
  wire  _T_984; // @[MemPrimitives.scala 83:102:@16264.4]
  wire  _T_989; // @[MemPrimitives.scala 82:228:@16267.4]
  wire  _T_990; // @[MemPrimitives.scala 83:102:@16268.4]
  wire [16:0] _T_992; // @[Cat.scala 30:58:@16270.4]
  wire [16:0] _T_994; // @[Cat.scala 30:58:@16272.4]
  wire [16:0] _T_995; // @[Mux.scala 31:69:@16273.4]
  wire  _T_1003; // @[MemPrimitives.scala 82:228:@16282.4]
  wire  _T_1004; // @[MemPrimitives.scala 83:102:@16283.4]
  wire  _T_1009; // @[MemPrimitives.scala 82:228:@16286.4]
  wire  _T_1010; // @[MemPrimitives.scala 83:102:@16287.4]
  wire [16:0] _T_1012; // @[Cat.scala 30:58:@16289.4]
  wire [16:0] _T_1014; // @[Cat.scala 30:58:@16291.4]
  wire [16:0] _T_1015; // @[Mux.scala 31:69:@16292.4]
  wire  _T_1023; // @[MemPrimitives.scala 82:228:@16301.4]
  wire  _T_1024; // @[MemPrimitives.scala 83:102:@16302.4]
  wire  _T_1029; // @[MemPrimitives.scala 82:228:@16305.4]
  wire  _T_1030; // @[MemPrimitives.scala 83:102:@16306.4]
  wire [16:0] _T_1032; // @[Cat.scala 30:58:@16308.4]
  wire [16:0] _T_1034; // @[Cat.scala 30:58:@16310.4]
  wire [16:0] _T_1035; // @[Mux.scala 31:69:@16311.4]
  wire  _T_1043; // @[MemPrimitives.scala 82:228:@16320.4]
  wire  _T_1044; // @[MemPrimitives.scala 83:102:@16321.4]
  wire  _T_1049; // @[MemPrimitives.scala 82:228:@16324.4]
  wire  _T_1050; // @[MemPrimitives.scala 83:102:@16325.4]
  wire [16:0] _T_1052; // @[Cat.scala 30:58:@16327.4]
  wire [16:0] _T_1054; // @[Cat.scala 30:58:@16329.4]
  wire [16:0] _T_1055; // @[Mux.scala 31:69:@16330.4]
  wire  _T_1060; // @[MemPrimitives.scala 82:210:@16337.4]
  wire  _T_1063; // @[MemPrimitives.scala 82:228:@16339.4]
  wire  _T_1064; // @[MemPrimitives.scala 83:102:@16340.4]
  wire  _T_1066; // @[MemPrimitives.scala 82:210:@16341.4]
  wire  _T_1069; // @[MemPrimitives.scala 82:228:@16343.4]
  wire  _T_1070; // @[MemPrimitives.scala 83:102:@16344.4]
  wire [16:0] _T_1072; // @[Cat.scala 30:58:@16346.4]
  wire [16:0] _T_1074; // @[Cat.scala 30:58:@16348.4]
  wire [16:0] _T_1075; // @[Mux.scala 31:69:@16349.4]
  wire  _T_1080; // @[MemPrimitives.scala 82:210:@16356.4]
  wire  _T_1083; // @[MemPrimitives.scala 82:228:@16358.4]
  wire  _T_1084; // @[MemPrimitives.scala 83:102:@16359.4]
  wire  _T_1086; // @[MemPrimitives.scala 82:210:@16360.4]
  wire  _T_1089; // @[MemPrimitives.scala 82:228:@16362.4]
  wire  _T_1090; // @[MemPrimitives.scala 83:102:@16363.4]
  wire [16:0] _T_1092; // @[Cat.scala 30:58:@16365.4]
  wire [16:0] _T_1094; // @[Cat.scala 30:58:@16367.4]
  wire [16:0] _T_1095; // @[Mux.scala 31:69:@16368.4]
  wire  _T_1103; // @[MemPrimitives.scala 82:228:@16377.4]
  wire  _T_1104; // @[MemPrimitives.scala 83:102:@16378.4]
  wire  _T_1109; // @[MemPrimitives.scala 82:228:@16381.4]
  wire  _T_1110; // @[MemPrimitives.scala 83:102:@16382.4]
  wire [16:0] _T_1112; // @[Cat.scala 30:58:@16384.4]
  wire [16:0] _T_1114; // @[Cat.scala 30:58:@16386.4]
  wire [16:0] _T_1115; // @[Mux.scala 31:69:@16387.4]
  wire  _T_1123; // @[MemPrimitives.scala 82:228:@16396.4]
  wire  _T_1124; // @[MemPrimitives.scala 83:102:@16397.4]
  wire  _T_1129; // @[MemPrimitives.scala 82:228:@16400.4]
  wire  _T_1130; // @[MemPrimitives.scala 83:102:@16401.4]
  wire [16:0] _T_1132; // @[Cat.scala 30:58:@16403.4]
  wire [16:0] _T_1134; // @[Cat.scala 30:58:@16405.4]
  wire [16:0] _T_1135; // @[Mux.scala 31:69:@16406.4]
  wire  _T_1143; // @[MemPrimitives.scala 82:228:@16415.4]
  wire  _T_1144; // @[MemPrimitives.scala 83:102:@16416.4]
  wire  _T_1149; // @[MemPrimitives.scala 82:228:@16419.4]
  wire  _T_1150; // @[MemPrimitives.scala 83:102:@16420.4]
  wire [16:0] _T_1152; // @[Cat.scala 30:58:@16422.4]
  wire [16:0] _T_1154; // @[Cat.scala 30:58:@16424.4]
  wire [16:0] _T_1155; // @[Mux.scala 31:69:@16425.4]
  wire  _T_1163; // @[MemPrimitives.scala 82:228:@16434.4]
  wire  _T_1164; // @[MemPrimitives.scala 83:102:@16435.4]
  wire  _T_1169; // @[MemPrimitives.scala 82:228:@16438.4]
  wire  _T_1170; // @[MemPrimitives.scala 83:102:@16439.4]
  wire [16:0] _T_1172; // @[Cat.scala 30:58:@16441.4]
  wire [16:0] _T_1174; // @[Cat.scala 30:58:@16443.4]
  wire [16:0] _T_1175; // @[Mux.scala 31:69:@16444.4]
  wire  _T_1180; // @[MemPrimitives.scala 110:210:@16451.4]
  wire  _T_1182; // @[MemPrimitives.scala 110:210:@16452.4]
  wire  _T_1183; // @[MemPrimitives.scala 110:228:@16453.4]
  wire  _T_1186; // @[MemPrimitives.scala 110:210:@16455.4]
  wire  _T_1188; // @[MemPrimitives.scala 110:210:@16456.4]
  wire  _T_1189; // @[MemPrimitives.scala 110:228:@16457.4]
  wire  _T_1192; // @[MemPrimitives.scala 110:210:@16459.4]
  wire  _T_1194; // @[MemPrimitives.scala 110:210:@16460.4]
  wire  _T_1195; // @[MemPrimitives.scala 110:228:@16461.4]
  wire  _T_1198; // @[MemPrimitives.scala 110:210:@16463.4]
  wire  _T_1200; // @[MemPrimitives.scala 110:210:@16464.4]
  wire  _T_1201; // @[MemPrimitives.scala 110:228:@16465.4]
  wire  _T_1204; // @[MemPrimitives.scala 110:210:@16467.4]
  wire  _T_1206; // @[MemPrimitives.scala 110:210:@16468.4]
  wire  _T_1207; // @[MemPrimitives.scala 110:228:@16469.4]
  wire  _T_1210; // @[MemPrimitives.scala 110:210:@16471.4]
  wire  _T_1212; // @[MemPrimitives.scala 110:210:@16472.4]
  wire  _T_1213; // @[MemPrimitives.scala 110:228:@16473.4]
  wire  _T_1216; // @[MemPrimitives.scala 110:210:@16475.4]
  wire  _T_1218; // @[MemPrimitives.scala 110:210:@16476.4]
  wire  _T_1219; // @[MemPrimitives.scala 110:228:@16477.4]
  wire  _T_1222; // @[MemPrimitives.scala 110:210:@16479.4]
  wire  _T_1224; // @[MemPrimitives.scala 110:210:@16480.4]
  wire  _T_1225; // @[MemPrimitives.scala 110:228:@16481.4]
  wire  _T_1228; // @[MemPrimitives.scala 110:210:@16483.4]
  wire  _T_1230; // @[MemPrimitives.scala 110:210:@16484.4]
  wire  _T_1231; // @[MemPrimitives.scala 110:228:@16485.4]
  wire  _T_1233; // @[MemPrimitives.scala 123:41:@16499.4]
  wire  _T_1234; // @[MemPrimitives.scala 123:41:@16500.4]
  wire  _T_1235; // @[MemPrimitives.scala 123:41:@16501.4]
  wire  _T_1236; // @[MemPrimitives.scala 123:41:@16502.4]
  wire  _T_1237; // @[MemPrimitives.scala 123:41:@16503.4]
  wire  _T_1238; // @[MemPrimitives.scala 123:41:@16504.4]
  wire  _T_1239; // @[MemPrimitives.scala 123:41:@16505.4]
  wire  _T_1240; // @[MemPrimitives.scala 123:41:@16506.4]
  wire  _T_1241; // @[MemPrimitives.scala 123:41:@16507.4]
  wire [9:0] _T_1243; // @[Cat.scala 30:58:@16509.4]
  wire [9:0] _T_1245; // @[Cat.scala 30:58:@16511.4]
  wire [9:0] _T_1247; // @[Cat.scala 30:58:@16513.4]
  wire [9:0] _T_1249; // @[Cat.scala 30:58:@16515.4]
  wire [9:0] _T_1251; // @[Cat.scala 30:58:@16517.4]
  wire [9:0] _T_1253; // @[Cat.scala 30:58:@16519.4]
  wire [9:0] _T_1255; // @[Cat.scala 30:58:@16521.4]
  wire [9:0] _T_1257; // @[Cat.scala 30:58:@16523.4]
  wire [9:0] _T_1259; // @[Cat.scala 30:58:@16525.4]
  wire [9:0] _T_1260; // @[Mux.scala 31:69:@16526.4]
  wire [9:0] _T_1261; // @[Mux.scala 31:69:@16527.4]
  wire [9:0] _T_1262; // @[Mux.scala 31:69:@16528.4]
  wire [9:0] _T_1263; // @[Mux.scala 31:69:@16529.4]
  wire [9:0] _T_1264; // @[Mux.scala 31:69:@16530.4]
  wire [9:0] _T_1265; // @[Mux.scala 31:69:@16531.4]
  wire [9:0] _T_1266; // @[Mux.scala 31:69:@16532.4]
  wire [9:0] _T_1267; // @[Mux.scala 31:69:@16533.4]
  wire  _T_1272; // @[MemPrimitives.scala 110:210:@16540.4]
  wire  _T_1274; // @[MemPrimitives.scala 110:210:@16541.4]
  wire  _T_1275; // @[MemPrimitives.scala 110:228:@16542.4]
  wire  _T_1278; // @[MemPrimitives.scala 110:210:@16544.4]
  wire  _T_1280; // @[MemPrimitives.scala 110:210:@16545.4]
  wire  _T_1281; // @[MemPrimitives.scala 110:228:@16546.4]
  wire  _T_1284; // @[MemPrimitives.scala 110:210:@16548.4]
  wire  _T_1286; // @[MemPrimitives.scala 110:210:@16549.4]
  wire  _T_1287; // @[MemPrimitives.scala 110:228:@16550.4]
  wire  _T_1290; // @[MemPrimitives.scala 110:210:@16552.4]
  wire  _T_1292; // @[MemPrimitives.scala 110:210:@16553.4]
  wire  _T_1293; // @[MemPrimitives.scala 110:228:@16554.4]
  wire  _T_1296; // @[MemPrimitives.scala 110:210:@16556.4]
  wire  _T_1298; // @[MemPrimitives.scala 110:210:@16557.4]
  wire  _T_1299; // @[MemPrimitives.scala 110:228:@16558.4]
  wire  _T_1302; // @[MemPrimitives.scala 110:210:@16560.4]
  wire  _T_1304; // @[MemPrimitives.scala 110:210:@16561.4]
  wire  _T_1305; // @[MemPrimitives.scala 110:228:@16562.4]
  wire  _T_1308; // @[MemPrimitives.scala 110:210:@16564.4]
  wire  _T_1310; // @[MemPrimitives.scala 110:210:@16565.4]
  wire  _T_1311; // @[MemPrimitives.scala 110:228:@16566.4]
  wire  _T_1314; // @[MemPrimitives.scala 110:210:@16568.4]
  wire  _T_1316; // @[MemPrimitives.scala 110:210:@16569.4]
  wire  _T_1317; // @[MemPrimitives.scala 110:228:@16570.4]
  wire  _T_1320; // @[MemPrimitives.scala 110:210:@16572.4]
  wire  _T_1322; // @[MemPrimitives.scala 110:210:@16573.4]
  wire  _T_1323; // @[MemPrimitives.scala 110:228:@16574.4]
  wire  _T_1325; // @[MemPrimitives.scala 123:41:@16588.4]
  wire  _T_1326; // @[MemPrimitives.scala 123:41:@16589.4]
  wire  _T_1327; // @[MemPrimitives.scala 123:41:@16590.4]
  wire  _T_1328; // @[MemPrimitives.scala 123:41:@16591.4]
  wire  _T_1329; // @[MemPrimitives.scala 123:41:@16592.4]
  wire  _T_1330; // @[MemPrimitives.scala 123:41:@16593.4]
  wire  _T_1331; // @[MemPrimitives.scala 123:41:@16594.4]
  wire  _T_1332; // @[MemPrimitives.scala 123:41:@16595.4]
  wire  _T_1333; // @[MemPrimitives.scala 123:41:@16596.4]
  wire [9:0] _T_1335; // @[Cat.scala 30:58:@16598.4]
  wire [9:0] _T_1337; // @[Cat.scala 30:58:@16600.4]
  wire [9:0] _T_1339; // @[Cat.scala 30:58:@16602.4]
  wire [9:0] _T_1341; // @[Cat.scala 30:58:@16604.4]
  wire [9:0] _T_1343; // @[Cat.scala 30:58:@16606.4]
  wire [9:0] _T_1345; // @[Cat.scala 30:58:@16608.4]
  wire [9:0] _T_1347; // @[Cat.scala 30:58:@16610.4]
  wire [9:0] _T_1349; // @[Cat.scala 30:58:@16612.4]
  wire [9:0] _T_1351; // @[Cat.scala 30:58:@16614.4]
  wire [9:0] _T_1352; // @[Mux.scala 31:69:@16615.4]
  wire [9:0] _T_1353; // @[Mux.scala 31:69:@16616.4]
  wire [9:0] _T_1354; // @[Mux.scala 31:69:@16617.4]
  wire [9:0] _T_1355; // @[Mux.scala 31:69:@16618.4]
  wire [9:0] _T_1356; // @[Mux.scala 31:69:@16619.4]
  wire [9:0] _T_1357; // @[Mux.scala 31:69:@16620.4]
  wire [9:0] _T_1358; // @[Mux.scala 31:69:@16621.4]
  wire [9:0] _T_1359; // @[Mux.scala 31:69:@16622.4]
  wire  _T_1366; // @[MemPrimitives.scala 110:210:@16630.4]
  wire  _T_1367; // @[MemPrimitives.scala 110:228:@16631.4]
  wire  _T_1372; // @[MemPrimitives.scala 110:210:@16634.4]
  wire  _T_1373; // @[MemPrimitives.scala 110:228:@16635.4]
  wire  _T_1378; // @[MemPrimitives.scala 110:210:@16638.4]
  wire  _T_1379; // @[MemPrimitives.scala 110:228:@16639.4]
  wire  _T_1384; // @[MemPrimitives.scala 110:210:@16642.4]
  wire  _T_1385; // @[MemPrimitives.scala 110:228:@16643.4]
  wire  _T_1390; // @[MemPrimitives.scala 110:210:@16646.4]
  wire  _T_1391; // @[MemPrimitives.scala 110:228:@16647.4]
  wire  _T_1396; // @[MemPrimitives.scala 110:210:@16650.4]
  wire  _T_1397; // @[MemPrimitives.scala 110:228:@16651.4]
  wire  _T_1402; // @[MemPrimitives.scala 110:210:@16654.4]
  wire  _T_1403; // @[MemPrimitives.scala 110:228:@16655.4]
  wire  _T_1408; // @[MemPrimitives.scala 110:210:@16658.4]
  wire  _T_1409; // @[MemPrimitives.scala 110:228:@16659.4]
  wire  _T_1414; // @[MemPrimitives.scala 110:210:@16662.4]
  wire  _T_1415; // @[MemPrimitives.scala 110:228:@16663.4]
  wire  _T_1417; // @[MemPrimitives.scala 123:41:@16677.4]
  wire  _T_1418; // @[MemPrimitives.scala 123:41:@16678.4]
  wire  _T_1419; // @[MemPrimitives.scala 123:41:@16679.4]
  wire  _T_1420; // @[MemPrimitives.scala 123:41:@16680.4]
  wire  _T_1421; // @[MemPrimitives.scala 123:41:@16681.4]
  wire  _T_1422; // @[MemPrimitives.scala 123:41:@16682.4]
  wire  _T_1423; // @[MemPrimitives.scala 123:41:@16683.4]
  wire  _T_1424; // @[MemPrimitives.scala 123:41:@16684.4]
  wire  _T_1425; // @[MemPrimitives.scala 123:41:@16685.4]
  wire [9:0] _T_1427; // @[Cat.scala 30:58:@16687.4]
  wire [9:0] _T_1429; // @[Cat.scala 30:58:@16689.4]
  wire [9:0] _T_1431; // @[Cat.scala 30:58:@16691.4]
  wire [9:0] _T_1433; // @[Cat.scala 30:58:@16693.4]
  wire [9:0] _T_1435; // @[Cat.scala 30:58:@16695.4]
  wire [9:0] _T_1437; // @[Cat.scala 30:58:@16697.4]
  wire [9:0] _T_1439; // @[Cat.scala 30:58:@16699.4]
  wire [9:0] _T_1441; // @[Cat.scala 30:58:@16701.4]
  wire [9:0] _T_1443; // @[Cat.scala 30:58:@16703.4]
  wire [9:0] _T_1444; // @[Mux.scala 31:69:@16704.4]
  wire [9:0] _T_1445; // @[Mux.scala 31:69:@16705.4]
  wire [9:0] _T_1446; // @[Mux.scala 31:69:@16706.4]
  wire [9:0] _T_1447; // @[Mux.scala 31:69:@16707.4]
  wire [9:0] _T_1448; // @[Mux.scala 31:69:@16708.4]
  wire [9:0] _T_1449; // @[Mux.scala 31:69:@16709.4]
  wire [9:0] _T_1450; // @[Mux.scala 31:69:@16710.4]
  wire [9:0] _T_1451; // @[Mux.scala 31:69:@16711.4]
  wire  _T_1458; // @[MemPrimitives.scala 110:210:@16719.4]
  wire  _T_1459; // @[MemPrimitives.scala 110:228:@16720.4]
  wire  _T_1464; // @[MemPrimitives.scala 110:210:@16723.4]
  wire  _T_1465; // @[MemPrimitives.scala 110:228:@16724.4]
  wire  _T_1470; // @[MemPrimitives.scala 110:210:@16727.4]
  wire  _T_1471; // @[MemPrimitives.scala 110:228:@16728.4]
  wire  _T_1476; // @[MemPrimitives.scala 110:210:@16731.4]
  wire  _T_1477; // @[MemPrimitives.scala 110:228:@16732.4]
  wire  _T_1482; // @[MemPrimitives.scala 110:210:@16735.4]
  wire  _T_1483; // @[MemPrimitives.scala 110:228:@16736.4]
  wire  _T_1488; // @[MemPrimitives.scala 110:210:@16739.4]
  wire  _T_1489; // @[MemPrimitives.scala 110:228:@16740.4]
  wire  _T_1494; // @[MemPrimitives.scala 110:210:@16743.4]
  wire  _T_1495; // @[MemPrimitives.scala 110:228:@16744.4]
  wire  _T_1500; // @[MemPrimitives.scala 110:210:@16747.4]
  wire  _T_1501; // @[MemPrimitives.scala 110:228:@16748.4]
  wire  _T_1506; // @[MemPrimitives.scala 110:210:@16751.4]
  wire  _T_1507; // @[MemPrimitives.scala 110:228:@16752.4]
  wire  _T_1509; // @[MemPrimitives.scala 123:41:@16766.4]
  wire  _T_1510; // @[MemPrimitives.scala 123:41:@16767.4]
  wire  _T_1511; // @[MemPrimitives.scala 123:41:@16768.4]
  wire  _T_1512; // @[MemPrimitives.scala 123:41:@16769.4]
  wire  _T_1513; // @[MemPrimitives.scala 123:41:@16770.4]
  wire  _T_1514; // @[MemPrimitives.scala 123:41:@16771.4]
  wire  _T_1515; // @[MemPrimitives.scala 123:41:@16772.4]
  wire  _T_1516; // @[MemPrimitives.scala 123:41:@16773.4]
  wire  _T_1517; // @[MemPrimitives.scala 123:41:@16774.4]
  wire [9:0] _T_1519; // @[Cat.scala 30:58:@16776.4]
  wire [9:0] _T_1521; // @[Cat.scala 30:58:@16778.4]
  wire [9:0] _T_1523; // @[Cat.scala 30:58:@16780.4]
  wire [9:0] _T_1525; // @[Cat.scala 30:58:@16782.4]
  wire [9:0] _T_1527; // @[Cat.scala 30:58:@16784.4]
  wire [9:0] _T_1529; // @[Cat.scala 30:58:@16786.4]
  wire [9:0] _T_1531; // @[Cat.scala 30:58:@16788.4]
  wire [9:0] _T_1533; // @[Cat.scala 30:58:@16790.4]
  wire [9:0] _T_1535; // @[Cat.scala 30:58:@16792.4]
  wire [9:0] _T_1536; // @[Mux.scala 31:69:@16793.4]
  wire [9:0] _T_1537; // @[Mux.scala 31:69:@16794.4]
  wire [9:0] _T_1538; // @[Mux.scala 31:69:@16795.4]
  wire [9:0] _T_1539; // @[Mux.scala 31:69:@16796.4]
  wire [9:0] _T_1540; // @[Mux.scala 31:69:@16797.4]
  wire [9:0] _T_1541; // @[Mux.scala 31:69:@16798.4]
  wire [9:0] _T_1542; // @[Mux.scala 31:69:@16799.4]
  wire [9:0] _T_1543; // @[Mux.scala 31:69:@16800.4]
  wire  _T_1550; // @[MemPrimitives.scala 110:210:@16808.4]
  wire  _T_1551; // @[MemPrimitives.scala 110:228:@16809.4]
  wire  _T_1556; // @[MemPrimitives.scala 110:210:@16812.4]
  wire  _T_1557; // @[MemPrimitives.scala 110:228:@16813.4]
  wire  _T_1562; // @[MemPrimitives.scala 110:210:@16816.4]
  wire  _T_1563; // @[MemPrimitives.scala 110:228:@16817.4]
  wire  _T_1568; // @[MemPrimitives.scala 110:210:@16820.4]
  wire  _T_1569; // @[MemPrimitives.scala 110:228:@16821.4]
  wire  _T_1574; // @[MemPrimitives.scala 110:210:@16824.4]
  wire  _T_1575; // @[MemPrimitives.scala 110:228:@16825.4]
  wire  _T_1580; // @[MemPrimitives.scala 110:210:@16828.4]
  wire  _T_1581; // @[MemPrimitives.scala 110:228:@16829.4]
  wire  _T_1586; // @[MemPrimitives.scala 110:210:@16832.4]
  wire  _T_1587; // @[MemPrimitives.scala 110:228:@16833.4]
  wire  _T_1592; // @[MemPrimitives.scala 110:210:@16836.4]
  wire  _T_1593; // @[MemPrimitives.scala 110:228:@16837.4]
  wire  _T_1598; // @[MemPrimitives.scala 110:210:@16840.4]
  wire  _T_1599; // @[MemPrimitives.scala 110:228:@16841.4]
  wire  _T_1601; // @[MemPrimitives.scala 123:41:@16855.4]
  wire  _T_1602; // @[MemPrimitives.scala 123:41:@16856.4]
  wire  _T_1603; // @[MemPrimitives.scala 123:41:@16857.4]
  wire  _T_1604; // @[MemPrimitives.scala 123:41:@16858.4]
  wire  _T_1605; // @[MemPrimitives.scala 123:41:@16859.4]
  wire  _T_1606; // @[MemPrimitives.scala 123:41:@16860.4]
  wire  _T_1607; // @[MemPrimitives.scala 123:41:@16861.4]
  wire  _T_1608; // @[MemPrimitives.scala 123:41:@16862.4]
  wire  _T_1609; // @[MemPrimitives.scala 123:41:@16863.4]
  wire [9:0] _T_1611; // @[Cat.scala 30:58:@16865.4]
  wire [9:0] _T_1613; // @[Cat.scala 30:58:@16867.4]
  wire [9:0] _T_1615; // @[Cat.scala 30:58:@16869.4]
  wire [9:0] _T_1617; // @[Cat.scala 30:58:@16871.4]
  wire [9:0] _T_1619; // @[Cat.scala 30:58:@16873.4]
  wire [9:0] _T_1621; // @[Cat.scala 30:58:@16875.4]
  wire [9:0] _T_1623; // @[Cat.scala 30:58:@16877.4]
  wire [9:0] _T_1625; // @[Cat.scala 30:58:@16879.4]
  wire [9:0] _T_1627; // @[Cat.scala 30:58:@16881.4]
  wire [9:0] _T_1628; // @[Mux.scala 31:69:@16882.4]
  wire [9:0] _T_1629; // @[Mux.scala 31:69:@16883.4]
  wire [9:0] _T_1630; // @[Mux.scala 31:69:@16884.4]
  wire [9:0] _T_1631; // @[Mux.scala 31:69:@16885.4]
  wire [9:0] _T_1632; // @[Mux.scala 31:69:@16886.4]
  wire [9:0] _T_1633; // @[Mux.scala 31:69:@16887.4]
  wire [9:0] _T_1634; // @[Mux.scala 31:69:@16888.4]
  wire [9:0] _T_1635; // @[Mux.scala 31:69:@16889.4]
  wire  _T_1642; // @[MemPrimitives.scala 110:210:@16897.4]
  wire  _T_1643; // @[MemPrimitives.scala 110:228:@16898.4]
  wire  _T_1648; // @[MemPrimitives.scala 110:210:@16901.4]
  wire  _T_1649; // @[MemPrimitives.scala 110:228:@16902.4]
  wire  _T_1654; // @[MemPrimitives.scala 110:210:@16905.4]
  wire  _T_1655; // @[MemPrimitives.scala 110:228:@16906.4]
  wire  _T_1660; // @[MemPrimitives.scala 110:210:@16909.4]
  wire  _T_1661; // @[MemPrimitives.scala 110:228:@16910.4]
  wire  _T_1666; // @[MemPrimitives.scala 110:210:@16913.4]
  wire  _T_1667; // @[MemPrimitives.scala 110:228:@16914.4]
  wire  _T_1672; // @[MemPrimitives.scala 110:210:@16917.4]
  wire  _T_1673; // @[MemPrimitives.scala 110:228:@16918.4]
  wire  _T_1678; // @[MemPrimitives.scala 110:210:@16921.4]
  wire  _T_1679; // @[MemPrimitives.scala 110:228:@16922.4]
  wire  _T_1684; // @[MemPrimitives.scala 110:210:@16925.4]
  wire  _T_1685; // @[MemPrimitives.scala 110:228:@16926.4]
  wire  _T_1690; // @[MemPrimitives.scala 110:210:@16929.4]
  wire  _T_1691; // @[MemPrimitives.scala 110:228:@16930.4]
  wire  _T_1693; // @[MemPrimitives.scala 123:41:@16944.4]
  wire  _T_1694; // @[MemPrimitives.scala 123:41:@16945.4]
  wire  _T_1695; // @[MemPrimitives.scala 123:41:@16946.4]
  wire  _T_1696; // @[MemPrimitives.scala 123:41:@16947.4]
  wire  _T_1697; // @[MemPrimitives.scala 123:41:@16948.4]
  wire  _T_1698; // @[MemPrimitives.scala 123:41:@16949.4]
  wire  _T_1699; // @[MemPrimitives.scala 123:41:@16950.4]
  wire  _T_1700; // @[MemPrimitives.scala 123:41:@16951.4]
  wire  _T_1701; // @[MemPrimitives.scala 123:41:@16952.4]
  wire [9:0] _T_1703; // @[Cat.scala 30:58:@16954.4]
  wire [9:0] _T_1705; // @[Cat.scala 30:58:@16956.4]
  wire [9:0] _T_1707; // @[Cat.scala 30:58:@16958.4]
  wire [9:0] _T_1709; // @[Cat.scala 30:58:@16960.4]
  wire [9:0] _T_1711; // @[Cat.scala 30:58:@16962.4]
  wire [9:0] _T_1713; // @[Cat.scala 30:58:@16964.4]
  wire [9:0] _T_1715; // @[Cat.scala 30:58:@16966.4]
  wire [9:0] _T_1717; // @[Cat.scala 30:58:@16968.4]
  wire [9:0] _T_1719; // @[Cat.scala 30:58:@16970.4]
  wire [9:0] _T_1720; // @[Mux.scala 31:69:@16971.4]
  wire [9:0] _T_1721; // @[Mux.scala 31:69:@16972.4]
  wire [9:0] _T_1722; // @[Mux.scala 31:69:@16973.4]
  wire [9:0] _T_1723; // @[Mux.scala 31:69:@16974.4]
  wire [9:0] _T_1724; // @[Mux.scala 31:69:@16975.4]
  wire [9:0] _T_1725; // @[Mux.scala 31:69:@16976.4]
  wire [9:0] _T_1726; // @[Mux.scala 31:69:@16977.4]
  wire [9:0] _T_1727; // @[Mux.scala 31:69:@16978.4]
  wire  _T_1732; // @[MemPrimitives.scala 110:210:@16985.4]
  wire  _T_1735; // @[MemPrimitives.scala 110:228:@16987.4]
  wire  _T_1738; // @[MemPrimitives.scala 110:210:@16989.4]
  wire  _T_1741; // @[MemPrimitives.scala 110:228:@16991.4]
  wire  _T_1744; // @[MemPrimitives.scala 110:210:@16993.4]
  wire  _T_1747; // @[MemPrimitives.scala 110:228:@16995.4]
  wire  _T_1750; // @[MemPrimitives.scala 110:210:@16997.4]
  wire  _T_1753; // @[MemPrimitives.scala 110:228:@16999.4]
  wire  _T_1756; // @[MemPrimitives.scala 110:210:@17001.4]
  wire  _T_1759; // @[MemPrimitives.scala 110:228:@17003.4]
  wire  _T_1762; // @[MemPrimitives.scala 110:210:@17005.4]
  wire  _T_1765; // @[MemPrimitives.scala 110:228:@17007.4]
  wire  _T_1768; // @[MemPrimitives.scala 110:210:@17009.4]
  wire  _T_1771; // @[MemPrimitives.scala 110:228:@17011.4]
  wire  _T_1774; // @[MemPrimitives.scala 110:210:@17013.4]
  wire  _T_1777; // @[MemPrimitives.scala 110:228:@17015.4]
  wire  _T_1780; // @[MemPrimitives.scala 110:210:@17017.4]
  wire  _T_1783; // @[MemPrimitives.scala 110:228:@17019.4]
  wire  _T_1785; // @[MemPrimitives.scala 123:41:@17033.4]
  wire  _T_1786; // @[MemPrimitives.scala 123:41:@17034.4]
  wire  _T_1787; // @[MemPrimitives.scala 123:41:@17035.4]
  wire  _T_1788; // @[MemPrimitives.scala 123:41:@17036.4]
  wire  _T_1789; // @[MemPrimitives.scala 123:41:@17037.4]
  wire  _T_1790; // @[MemPrimitives.scala 123:41:@17038.4]
  wire  _T_1791; // @[MemPrimitives.scala 123:41:@17039.4]
  wire  _T_1792; // @[MemPrimitives.scala 123:41:@17040.4]
  wire  _T_1793; // @[MemPrimitives.scala 123:41:@17041.4]
  wire [9:0] _T_1795; // @[Cat.scala 30:58:@17043.4]
  wire [9:0] _T_1797; // @[Cat.scala 30:58:@17045.4]
  wire [9:0] _T_1799; // @[Cat.scala 30:58:@17047.4]
  wire [9:0] _T_1801; // @[Cat.scala 30:58:@17049.4]
  wire [9:0] _T_1803; // @[Cat.scala 30:58:@17051.4]
  wire [9:0] _T_1805; // @[Cat.scala 30:58:@17053.4]
  wire [9:0] _T_1807; // @[Cat.scala 30:58:@17055.4]
  wire [9:0] _T_1809; // @[Cat.scala 30:58:@17057.4]
  wire [9:0] _T_1811; // @[Cat.scala 30:58:@17059.4]
  wire [9:0] _T_1812; // @[Mux.scala 31:69:@17060.4]
  wire [9:0] _T_1813; // @[Mux.scala 31:69:@17061.4]
  wire [9:0] _T_1814; // @[Mux.scala 31:69:@17062.4]
  wire [9:0] _T_1815; // @[Mux.scala 31:69:@17063.4]
  wire [9:0] _T_1816; // @[Mux.scala 31:69:@17064.4]
  wire [9:0] _T_1817; // @[Mux.scala 31:69:@17065.4]
  wire [9:0] _T_1818; // @[Mux.scala 31:69:@17066.4]
  wire [9:0] _T_1819; // @[Mux.scala 31:69:@17067.4]
  wire  _T_1824; // @[MemPrimitives.scala 110:210:@17074.4]
  wire  _T_1827; // @[MemPrimitives.scala 110:228:@17076.4]
  wire  _T_1830; // @[MemPrimitives.scala 110:210:@17078.4]
  wire  _T_1833; // @[MemPrimitives.scala 110:228:@17080.4]
  wire  _T_1836; // @[MemPrimitives.scala 110:210:@17082.4]
  wire  _T_1839; // @[MemPrimitives.scala 110:228:@17084.4]
  wire  _T_1842; // @[MemPrimitives.scala 110:210:@17086.4]
  wire  _T_1845; // @[MemPrimitives.scala 110:228:@17088.4]
  wire  _T_1848; // @[MemPrimitives.scala 110:210:@17090.4]
  wire  _T_1851; // @[MemPrimitives.scala 110:228:@17092.4]
  wire  _T_1854; // @[MemPrimitives.scala 110:210:@17094.4]
  wire  _T_1857; // @[MemPrimitives.scala 110:228:@17096.4]
  wire  _T_1860; // @[MemPrimitives.scala 110:210:@17098.4]
  wire  _T_1863; // @[MemPrimitives.scala 110:228:@17100.4]
  wire  _T_1866; // @[MemPrimitives.scala 110:210:@17102.4]
  wire  _T_1869; // @[MemPrimitives.scala 110:228:@17104.4]
  wire  _T_1872; // @[MemPrimitives.scala 110:210:@17106.4]
  wire  _T_1875; // @[MemPrimitives.scala 110:228:@17108.4]
  wire  _T_1877; // @[MemPrimitives.scala 123:41:@17122.4]
  wire  _T_1878; // @[MemPrimitives.scala 123:41:@17123.4]
  wire  _T_1879; // @[MemPrimitives.scala 123:41:@17124.4]
  wire  _T_1880; // @[MemPrimitives.scala 123:41:@17125.4]
  wire  _T_1881; // @[MemPrimitives.scala 123:41:@17126.4]
  wire  _T_1882; // @[MemPrimitives.scala 123:41:@17127.4]
  wire  _T_1883; // @[MemPrimitives.scala 123:41:@17128.4]
  wire  _T_1884; // @[MemPrimitives.scala 123:41:@17129.4]
  wire  _T_1885; // @[MemPrimitives.scala 123:41:@17130.4]
  wire [9:0] _T_1887; // @[Cat.scala 30:58:@17132.4]
  wire [9:0] _T_1889; // @[Cat.scala 30:58:@17134.4]
  wire [9:0] _T_1891; // @[Cat.scala 30:58:@17136.4]
  wire [9:0] _T_1893; // @[Cat.scala 30:58:@17138.4]
  wire [9:0] _T_1895; // @[Cat.scala 30:58:@17140.4]
  wire [9:0] _T_1897; // @[Cat.scala 30:58:@17142.4]
  wire [9:0] _T_1899; // @[Cat.scala 30:58:@17144.4]
  wire [9:0] _T_1901; // @[Cat.scala 30:58:@17146.4]
  wire [9:0] _T_1903; // @[Cat.scala 30:58:@17148.4]
  wire [9:0] _T_1904; // @[Mux.scala 31:69:@17149.4]
  wire [9:0] _T_1905; // @[Mux.scala 31:69:@17150.4]
  wire [9:0] _T_1906; // @[Mux.scala 31:69:@17151.4]
  wire [9:0] _T_1907; // @[Mux.scala 31:69:@17152.4]
  wire [9:0] _T_1908; // @[Mux.scala 31:69:@17153.4]
  wire [9:0] _T_1909; // @[Mux.scala 31:69:@17154.4]
  wire [9:0] _T_1910; // @[Mux.scala 31:69:@17155.4]
  wire [9:0] _T_1911; // @[Mux.scala 31:69:@17156.4]
  wire  _T_1919; // @[MemPrimitives.scala 110:228:@17165.4]
  wire  _T_1925; // @[MemPrimitives.scala 110:228:@17169.4]
  wire  _T_1931; // @[MemPrimitives.scala 110:228:@17173.4]
  wire  _T_1937; // @[MemPrimitives.scala 110:228:@17177.4]
  wire  _T_1943; // @[MemPrimitives.scala 110:228:@17181.4]
  wire  _T_1949; // @[MemPrimitives.scala 110:228:@17185.4]
  wire  _T_1955; // @[MemPrimitives.scala 110:228:@17189.4]
  wire  _T_1961; // @[MemPrimitives.scala 110:228:@17193.4]
  wire  _T_1967; // @[MemPrimitives.scala 110:228:@17197.4]
  wire  _T_1969; // @[MemPrimitives.scala 123:41:@17211.4]
  wire  _T_1970; // @[MemPrimitives.scala 123:41:@17212.4]
  wire  _T_1971; // @[MemPrimitives.scala 123:41:@17213.4]
  wire  _T_1972; // @[MemPrimitives.scala 123:41:@17214.4]
  wire  _T_1973; // @[MemPrimitives.scala 123:41:@17215.4]
  wire  _T_1974; // @[MemPrimitives.scala 123:41:@17216.4]
  wire  _T_1975; // @[MemPrimitives.scala 123:41:@17217.4]
  wire  _T_1976; // @[MemPrimitives.scala 123:41:@17218.4]
  wire  _T_1977; // @[MemPrimitives.scala 123:41:@17219.4]
  wire [9:0] _T_1979; // @[Cat.scala 30:58:@17221.4]
  wire [9:0] _T_1981; // @[Cat.scala 30:58:@17223.4]
  wire [9:0] _T_1983; // @[Cat.scala 30:58:@17225.4]
  wire [9:0] _T_1985; // @[Cat.scala 30:58:@17227.4]
  wire [9:0] _T_1987; // @[Cat.scala 30:58:@17229.4]
  wire [9:0] _T_1989; // @[Cat.scala 30:58:@17231.4]
  wire [9:0] _T_1991; // @[Cat.scala 30:58:@17233.4]
  wire [9:0] _T_1993; // @[Cat.scala 30:58:@17235.4]
  wire [9:0] _T_1995; // @[Cat.scala 30:58:@17237.4]
  wire [9:0] _T_1996; // @[Mux.scala 31:69:@17238.4]
  wire [9:0] _T_1997; // @[Mux.scala 31:69:@17239.4]
  wire [9:0] _T_1998; // @[Mux.scala 31:69:@17240.4]
  wire [9:0] _T_1999; // @[Mux.scala 31:69:@17241.4]
  wire [9:0] _T_2000; // @[Mux.scala 31:69:@17242.4]
  wire [9:0] _T_2001; // @[Mux.scala 31:69:@17243.4]
  wire [9:0] _T_2002; // @[Mux.scala 31:69:@17244.4]
  wire [9:0] _T_2003; // @[Mux.scala 31:69:@17245.4]
  wire  _T_2011; // @[MemPrimitives.scala 110:228:@17254.4]
  wire  _T_2017; // @[MemPrimitives.scala 110:228:@17258.4]
  wire  _T_2023; // @[MemPrimitives.scala 110:228:@17262.4]
  wire  _T_2029; // @[MemPrimitives.scala 110:228:@17266.4]
  wire  _T_2035; // @[MemPrimitives.scala 110:228:@17270.4]
  wire  _T_2041; // @[MemPrimitives.scala 110:228:@17274.4]
  wire  _T_2047; // @[MemPrimitives.scala 110:228:@17278.4]
  wire  _T_2053; // @[MemPrimitives.scala 110:228:@17282.4]
  wire  _T_2059; // @[MemPrimitives.scala 110:228:@17286.4]
  wire  _T_2061; // @[MemPrimitives.scala 123:41:@17300.4]
  wire  _T_2062; // @[MemPrimitives.scala 123:41:@17301.4]
  wire  _T_2063; // @[MemPrimitives.scala 123:41:@17302.4]
  wire  _T_2064; // @[MemPrimitives.scala 123:41:@17303.4]
  wire  _T_2065; // @[MemPrimitives.scala 123:41:@17304.4]
  wire  _T_2066; // @[MemPrimitives.scala 123:41:@17305.4]
  wire  _T_2067; // @[MemPrimitives.scala 123:41:@17306.4]
  wire  _T_2068; // @[MemPrimitives.scala 123:41:@17307.4]
  wire  _T_2069; // @[MemPrimitives.scala 123:41:@17308.4]
  wire [9:0] _T_2071; // @[Cat.scala 30:58:@17310.4]
  wire [9:0] _T_2073; // @[Cat.scala 30:58:@17312.4]
  wire [9:0] _T_2075; // @[Cat.scala 30:58:@17314.4]
  wire [9:0] _T_2077; // @[Cat.scala 30:58:@17316.4]
  wire [9:0] _T_2079; // @[Cat.scala 30:58:@17318.4]
  wire [9:0] _T_2081; // @[Cat.scala 30:58:@17320.4]
  wire [9:0] _T_2083; // @[Cat.scala 30:58:@17322.4]
  wire [9:0] _T_2085; // @[Cat.scala 30:58:@17324.4]
  wire [9:0] _T_2087; // @[Cat.scala 30:58:@17326.4]
  wire [9:0] _T_2088; // @[Mux.scala 31:69:@17327.4]
  wire [9:0] _T_2089; // @[Mux.scala 31:69:@17328.4]
  wire [9:0] _T_2090; // @[Mux.scala 31:69:@17329.4]
  wire [9:0] _T_2091; // @[Mux.scala 31:69:@17330.4]
  wire [9:0] _T_2092; // @[Mux.scala 31:69:@17331.4]
  wire [9:0] _T_2093; // @[Mux.scala 31:69:@17332.4]
  wire [9:0] _T_2094; // @[Mux.scala 31:69:@17333.4]
  wire [9:0] _T_2095; // @[Mux.scala 31:69:@17334.4]
  wire  _T_2103; // @[MemPrimitives.scala 110:228:@17343.4]
  wire  _T_2109; // @[MemPrimitives.scala 110:228:@17347.4]
  wire  _T_2115; // @[MemPrimitives.scala 110:228:@17351.4]
  wire  _T_2121; // @[MemPrimitives.scala 110:228:@17355.4]
  wire  _T_2127; // @[MemPrimitives.scala 110:228:@17359.4]
  wire  _T_2133; // @[MemPrimitives.scala 110:228:@17363.4]
  wire  _T_2139; // @[MemPrimitives.scala 110:228:@17367.4]
  wire  _T_2145; // @[MemPrimitives.scala 110:228:@17371.4]
  wire  _T_2151; // @[MemPrimitives.scala 110:228:@17375.4]
  wire  _T_2153; // @[MemPrimitives.scala 123:41:@17389.4]
  wire  _T_2154; // @[MemPrimitives.scala 123:41:@17390.4]
  wire  _T_2155; // @[MemPrimitives.scala 123:41:@17391.4]
  wire  _T_2156; // @[MemPrimitives.scala 123:41:@17392.4]
  wire  _T_2157; // @[MemPrimitives.scala 123:41:@17393.4]
  wire  _T_2158; // @[MemPrimitives.scala 123:41:@17394.4]
  wire  _T_2159; // @[MemPrimitives.scala 123:41:@17395.4]
  wire  _T_2160; // @[MemPrimitives.scala 123:41:@17396.4]
  wire  _T_2161; // @[MemPrimitives.scala 123:41:@17397.4]
  wire [9:0] _T_2163; // @[Cat.scala 30:58:@17399.4]
  wire [9:0] _T_2165; // @[Cat.scala 30:58:@17401.4]
  wire [9:0] _T_2167; // @[Cat.scala 30:58:@17403.4]
  wire [9:0] _T_2169; // @[Cat.scala 30:58:@17405.4]
  wire [9:0] _T_2171; // @[Cat.scala 30:58:@17407.4]
  wire [9:0] _T_2173; // @[Cat.scala 30:58:@17409.4]
  wire [9:0] _T_2175; // @[Cat.scala 30:58:@17411.4]
  wire [9:0] _T_2177; // @[Cat.scala 30:58:@17413.4]
  wire [9:0] _T_2179; // @[Cat.scala 30:58:@17415.4]
  wire [9:0] _T_2180; // @[Mux.scala 31:69:@17416.4]
  wire [9:0] _T_2181; // @[Mux.scala 31:69:@17417.4]
  wire [9:0] _T_2182; // @[Mux.scala 31:69:@17418.4]
  wire [9:0] _T_2183; // @[Mux.scala 31:69:@17419.4]
  wire [9:0] _T_2184; // @[Mux.scala 31:69:@17420.4]
  wire [9:0] _T_2185; // @[Mux.scala 31:69:@17421.4]
  wire [9:0] _T_2186; // @[Mux.scala 31:69:@17422.4]
  wire [9:0] _T_2187; // @[Mux.scala 31:69:@17423.4]
  wire  _T_2195; // @[MemPrimitives.scala 110:228:@17432.4]
  wire  _T_2201; // @[MemPrimitives.scala 110:228:@17436.4]
  wire  _T_2207; // @[MemPrimitives.scala 110:228:@17440.4]
  wire  _T_2213; // @[MemPrimitives.scala 110:228:@17444.4]
  wire  _T_2219; // @[MemPrimitives.scala 110:228:@17448.4]
  wire  _T_2225; // @[MemPrimitives.scala 110:228:@17452.4]
  wire  _T_2231; // @[MemPrimitives.scala 110:228:@17456.4]
  wire  _T_2237; // @[MemPrimitives.scala 110:228:@17460.4]
  wire  _T_2243; // @[MemPrimitives.scala 110:228:@17464.4]
  wire  _T_2245; // @[MemPrimitives.scala 123:41:@17478.4]
  wire  _T_2246; // @[MemPrimitives.scala 123:41:@17479.4]
  wire  _T_2247; // @[MemPrimitives.scala 123:41:@17480.4]
  wire  _T_2248; // @[MemPrimitives.scala 123:41:@17481.4]
  wire  _T_2249; // @[MemPrimitives.scala 123:41:@17482.4]
  wire  _T_2250; // @[MemPrimitives.scala 123:41:@17483.4]
  wire  _T_2251; // @[MemPrimitives.scala 123:41:@17484.4]
  wire  _T_2252; // @[MemPrimitives.scala 123:41:@17485.4]
  wire  _T_2253; // @[MemPrimitives.scala 123:41:@17486.4]
  wire [9:0] _T_2255; // @[Cat.scala 30:58:@17488.4]
  wire [9:0] _T_2257; // @[Cat.scala 30:58:@17490.4]
  wire [9:0] _T_2259; // @[Cat.scala 30:58:@17492.4]
  wire [9:0] _T_2261; // @[Cat.scala 30:58:@17494.4]
  wire [9:0] _T_2263; // @[Cat.scala 30:58:@17496.4]
  wire [9:0] _T_2265; // @[Cat.scala 30:58:@17498.4]
  wire [9:0] _T_2267; // @[Cat.scala 30:58:@17500.4]
  wire [9:0] _T_2269; // @[Cat.scala 30:58:@17502.4]
  wire [9:0] _T_2271; // @[Cat.scala 30:58:@17504.4]
  wire [9:0] _T_2272; // @[Mux.scala 31:69:@17505.4]
  wire [9:0] _T_2273; // @[Mux.scala 31:69:@17506.4]
  wire [9:0] _T_2274; // @[Mux.scala 31:69:@17507.4]
  wire [9:0] _T_2275; // @[Mux.scala 31:69:@17508.4]
  wire [9:0] _T_2276; // @[Mux.scala 31:69:@17509.4]
  wire [9:0] _T_2277; // @[Mux.scala 31:69:@17510.4]
  wire [9:0] _T_2278; // @[Mux.scala 31:69:@17511.4]
  wire [9:0] _T_2279; // @[Mux.scala 31:69:@17512.4]
  wire  _T_2284; // @[MemPrimitives.scala 110:210:@17519.4]
  wire  _T_2287; // @[MemPrimitives.scala 110:228:@17521.4]
  wire  _T_2290; // @[MemPrimitives.scala 110:210:@17523.4]
  wire  _T_2293; // @[MemPrimitives.scala 110:228:@17525.4]
  wire  _T_2296; // @[MemPrimitives.scala 110:210:@17527.4]
  wire  _T_2299; // @[MemPrimitives.scala 110:228:@17529.4]
  wire  _T_2302; // @[MemPrimitives.scala 110:210:@17531.4]
  wire  _T_2305; // @[MemPrimitives.scala 110:228:@17533.4]
  wire  _T_2308; // @[MemPrimitives.scala 110:210:@17535.4]
  wire  _T_2311; // @[MemPrimitives.scala 110:228:@17537.4]
  wire  _T_2314; // @[MemPrimitives.scala 110:210:@17539.4]
  wire  _T_2317; // @[MemPrimitives.scala 110:228:@17541.4]
  wire  _T_2320; // @[MemPrimitives.scala 110:210:@17543.4]
  wire  _T_2323; // @[MemPrimitives.scala 110:228:@17545.4]
  wire  _T_2326; // @[MemPrimitives.scala 110:210:@17547.4]
  wire  _T_2329; // @[MemPrimitives.scala 110:228:@17549.4]
  wire  _T_2332; // @[MemPrimitives.scala 110:210:@17551.4]
  wire  _T_2335; // @[MemPrimitives.scala 110:228:@17553.4]
  wire  _T_2337; // @[MemPrimitives.scala 123:41:@17567.4]
  wire  _T_2338; // @[MemPrimitives.scala 123:41:@17568.4]
  wire  _T_2339; // @[MemPrimitives.scala 123:41:@17569.4]
  wire  _T_2340; // @[MemPrimitives.scala 123:41:@17570.4]
  wire  _T_2341; // @[MemPrimitives.scala 123:41:@17571.4]
  wire  _T_2342; // @[MemPrimitives.scala 123:41:@17572.4]
  wire  _T_2343; // @[MemPrimitives.scala 123:41:@17573.4]
  wire  _T_2344; // @[MemPrimitives.scala 123:41:@17574.4]
  wire  _T_2345; // @[MemPrimitives.scala 123:41:@17575.4]
  wire [9:0] _T_2347; // @[Cat.scala 30:58:@17577.4]
  wire [9:0] _T_2349; // @[Cat.scala 30:58:@17579.4]
  wire [9:0] _T_2351; // @[Cat.scala 30:58:@17581.4]
  wire [9:0] _T_2353; // @[Cat.scala 30:58:@17583.4]
  wire [9:0] _T_2355; // @[Cat.scala 30:58:@17585.4]
  wire [9:0] _T_2357; // @[Cat.scala 30:58:@17587.4]
  wire [9:0] _T_2359; // @[Cat.scala 30:58:@17589.4]
  wire [9:0] _T_2361; // @[Cat.scala 30:58:@17591.4]
  wire [9:0] _T_2363; // @[Cat.scala 30:58:@17593.4]
  wire [9:0] _T_2364; // @[Mux.scala 31:69:@17594.4]
  wire [9:0] _T_2365; // @[Mux.scala 31:69:@17595.4]
  wire [9:0] _T_2366; // @[Mux.scala 31:69:@17596.4]
  wire [9:0] _T_2367; // @[Mux.scala 31:69:@17597.4]
  wire [9:0] _T_2368; // @[Mux.scala 31:69:@17598.4]
  wire [9:0] _T_2369; // @[Mux.scala 31:69:@17599.4]
  wire [9:0] _T_2370; // @[Mux.scala 31:69:@17600.4]
  wire [9:0] _T_2371; // @[Mux.scala 31:69:@17601.4]
  wire  _T_2376; // @[MemPrimitives.scala 110:210:@17608.4]
  wire  _T_2379; // @[MemPrimitives.scala 110:228:@17610.4]
  wire  _T_2382; // @[MemPrimitives.scala 110:210:@17612.4]
  wire  _T_2385; // @[MemPrimitives.scala 110:228:@17614.4]
  wire  _T_2388; // @[MemPrimitives.scala 110:210:@17616.4]
  wire  _T_2391; // @[MemPrimitives.scala 110:228:@17618.4]
  wire  _T_2394; // @[MemPrimitives.scala 110:210:@17620.4]
  wire  _T_2397; // @[MemPrimitives.scala 110:228:@17622.4]
  wire  _T_2400; // @[MemPrimitives.scala 110:210:@17624.4]
  wire  _T_2403; // @[MemPrimitives.scala 110:228:@17626.4]
  wire  _T_2406; // @[MemPrimitives.scala 110:210:@17628.4]
  wire  _T_2409; // @[MemPrimitives.scala 110:228:@17630.4]
  wire  _T_2412; // @[MemPrimitives.scala 110:210:@17632.4]
  wire  _T_2415; // @[MemPrimitives.scala 110:228:@17634.4]
  wire  _T_2418; // @[MemPrimitives.scala 110:210:@17636.4]
  wire  _T_2421; // @[MemPrimitives.scala 110:228:@17638.4]
  wire  _T_2424; // @[MemPrimitives.scala 110:210:@17640.4]
  wire  _T_2427; // @[MemPrimitives.scala 110:228:@17642.4]
  wire  _T_2429; // @[MemPrimitives.scala 123:41:@17656.4]
  wire  _T_2430; // @[MemPrimitives.scala 123:41:@17657.4]
  wire  _T_2431; // @[MemPrimitives.scala 123:41:@17658.4]
  wire  _T_2432; // @[MemPrimitives.scala 123:41:@17659.4]
  wire  _T_2433; // @[MemPrimitives.scala 123:41:@17660.4]
  wire  _T_2434; // @[MemPrimitives.scala 123:41:@17661.4]
  wire  _T_2435; // @[MemPrimitives.scala 123:41:@17662.4]
  wire  _T_2436; // @[MemPrimitives.scala 123:41:@17663.4]
  wire  _T_2437; // @[MemPrimitives.scala 123:41:@17664.4]
  wire [9:0] _T_2439; // @[Cat.scala 30:58:@17666.4]
  wire [9:0] _T_2441; // @[Cat.scala 30:58:@17668.4]
  wire [9:0] _T_2443; // @[Cat.scala 30:58:@17670.4]
  wire [9:0] _T_2445; // @[Cat.scala 30:58:@17672.4]
  wire [9:0] _T_2447; // @[Cat.scala 30:58:@17674.4]
  wire [9:0] _T_2449; // @[Cat.scala 30:58:@17676.4]
  wire [9:0] _T_2451; // @[Cat.scala 30:58:@17678.4]
  wire [9:0] _T_2453; // @[Cat.scala 30:58:@17680.4]
  wire [9:0] _T_2455; // @[Cat.scala 30:58:@17682.4]
  wire [9:0] _T_2456; // @[Mux.scala 31:69:@17683.4]
  wire [9:0] _T_2457; // @[Mux.scala 31:69:@17684.4]
  wire [9:0] _T_2458; // @[Mux.scala 31:69:@17685.4]
  wire [9:0] _T_2459; // @[Mux.scala 31:69:@17686.4]
  wire [9:0] _T_2460; // @[Mux.scala 31:69:@17687.4]
  wire [9:0] _T_2461; // @[Mux.scala 31:69:@17688.4]
  wire [9:0] _T_2462; // @[Mux.scala 31:69:@17689.4]
  wire [9:0] _T_2463; // @[Mux.scala 31:69:@17690.4]
  wire  _T_2471; // @[MemPrimitives.scala 110:228:@17699.4]
  wire  _T_2477; // @[MemPrimitives.scala 110:228:@17703.4]
  wire  _T_2483; // @[MemPrimitives.scala 110:228:@17707.4]
  wire  _T_2489; // @[MemPrimitives.scala 110:228:@17711.4]
  wire  _T_2495; // @[MemPrimitives.scala 110:228:@17715.4]
  wire  _T_2501; // @[MemPrimitives.scala 110:228:@17719.4]
  wire  _T_2507; // @[MemPrimitives.scala 110:228:@17723.4]
  wire  _T_2513; // @[MemPrimitives.scala 110:228:@17727.4]
  wire  _T_2519; // @[MemPrimitives.scala 110:228:@17731.4]
  wire  _T_2521; // @[MemPrimitives.scala 123:41:@17745.4]
  wire  _T_2522; // @[MemPrimitives.scala 123:41:@17746.4]
  wire  _T_2523; // @[MemPrimitives.scala 123:41:@17747.4]
  wire  _T_2524; // @[MemPrimitives.scala 123:41:@17748.4]
  wire  _T_2525; // @[MemPrimitives.scala 123:41:@17749.4]
  wire  _T_2526; // @[MemPrimitives.scala 123:41:@17750.4]
  wire  _T_2527; // @[MemPrimitives.scala 123:41:@17751.4]
  wire  _T_2528; // @[MemPrimitives.scala 123:41:@17752.4]
  wire  _T_2529; // @[MemPrimitives.scala 123:41:@17753.4]
  wire [9:0] _T_2531; // @[Cat.scala 30:58:@17755.4]
  wire [9:0] _T_2533; // @[Cat.scala 30:58:@17757.4]
  wire [9:0] _T_2535; // @[Cat.scala 30:58:@17759.4]
  wire [9:0] _T_2537; // @[Cat.scala 30:58:@17761.4]
  wire [9:0] _T_2539; // @[Cat.scala 30:58:@17763.4]
  wire [9:0] _T_2541; // @[Cat.scala 30:58:@17765.4]
  wire [9:0] _T_2543; // @[Cat.scala 30:58:@17767.4]
  wire [9:0] _T_2545; // @[Cat.scala 30:58:@17769.4]
  wire [9:0] _T_2547; // @[Cat.scala 30:58:@17771.4]
  wire [9:0] _T_2548; // @[Mux.scala 31:69:@17772.4]
  wire [9:0] _T_2549; // @[Mux.scala 31:69:@17773.4]
  wire [9:0] _T_2550; // @[Mux.scala 31:69:@17774.4]
  wire [9:0] _T_2551; // @[Mux.scala 31:69:@17775.4]
  wire [9:0] _T_2552; // @[Mux.scala 31:69:@17776.4]
  wire [9:0] _T_2553; // @[Mux.scala 31:69:@17777.4]
  wire [9:0] _T_2554; // @[Mux.scala 31:69:@17778.4]
  wire [9:0] _T_2555; // @[Mux.scala 31:69:@17779.4]
  wire  _T_2563; // @[MemPrimitives.scala 110:228:@17788.4]
  wire  _T_2569; // @[MemPrimitives.scala 110:228:@17792.4]
  wire  _T_2575; // @[MemPrimitives.scala 110:228:@17796.4]
  wire  _T_2581; // @[MemPrimitives.scala 110:228:@17800.4]
  wire  _T_2587; // @[MemPrimitives.scala 110:228:@17804.4]
  wire  _T_2593; // @[MemPrimitives.scala 110:228:@17808.4]
  wire  _T_2599; // @[MemPrimitives.scala 110:228:@17812.4]
  wire  _T_2605; // @[MemPrimitives.scala 110:228:@17816.4]
  wire  _T_2611; // @[MemPrimitives.scala 110:228:@17820.4]
  wire  _T_2613; // @[MemPrimitives.scala 123:41:@17834.4]
  wire  _T_2614; // @[MemPrimitives.scala 123:41:@17835.4]
  wire  _T_2615; // @[MemPrimitives.scala 123:41:@17836.4]
  wire  _T_2616; // @[MemPrimitives.scala 123:41:@17837.4]
  wire  _T_2617; // @[MemPrimitives.scala 123:41:@17838.4]
  wire  _T_2618; // @[MemPrimitives.scala 123:41:@17839.4]
  wire  _T_2619; // @[MemPrimitives.scala 123:41:@17840.4]
  wire  _T_2620; // @[MemPrimitives.scala 123:41:@17841.4]
  wire  _T_2621; // @[MemPrimitives.scala 123:41:@17842.4]
  wire [9:0] _T_2623; // @[Cat.scala 30:58:@17844.4]
  wire [9:0] _T_2625; // @[Cat.scala 30:58:@17846.4]
  wire [9:0] _T_2627; // @[Cat.scala 30:58:@17848.4]
  wire [9:0] _T_2629; // @[Cat.scala 30:58:@17850.4]
  wire [9:0] _T_2631; // @[Cat.scala 30:58:@17852.4]
  wire [9:0] _T_2633; // @[Cat.scala 30:58:@17854.4]
  wire [9:0] _T_2635; // @[Cat.scala 30:58:@17856.4]
  wire [9:0] _T_2637; // @[Cat.scala 30:58:@17858.4]
  wire [9:0] _T_2639; // @[Cat.scala 30:58:@17860.4]
  wire [9:0] _T_2640; // @[Mux.scala 31:69:@17861.4]
  wire [9:0] _T_2641; // @[Mux.scala 31:69:@17862.4]
  wire [9:0] _T_2642; // @[Mux.scala 31:69:@17863.4]
  wire [9:0] _T_2643; // @[Mux.scala 31:69:@17864.4]
  wire [9:0] _T_2644; // @[Mux.scala 31:69:@17865.4]
  wire [9:0] _T_2645; // @[Mux.scala 31:69:@17866.4]
  wire [9:0] _T_2646; // @[Mux.scala 31:69:@17867.4]
  wire [9:0] _T_2647; // @[Mux.scala 31:69:@17868.4]
  wire  _T_2655; // @[MemPrimitives.scala 110:228:@17877.4]
  wire  _T_2661; // @[MemPrimitives.scala 110:228:@17881.4]
  wire  _T_2667; // @[MemPrimitives.scala 110:228:@17885.4]
  wire  _T_2673; // @[MemPrimitives.scala 110:228:@17889.4]
  wire  _T_2679; // @[MemPrimitives.scala 110:228:@17893.4]
  wire  _T_2685; // @[MemPrimitives.scala 110:228:@17897.4]
  wire  _T_2691; // @[MemPrimitives.scala 110:228:@17901.4]
  wire  _T_2697; // @[MemPrimitives.scala 110:228:@17905.4]
  wire  _T_2703; // @[MemPrimitives.scala 110:228:@17909.4]
  wire  _T_2705; // @[MemPrimitives.scala 123:41:@17923.4]
  wire  _T_2706; // @[MemPrimitives.scala 123:41:@17924.4]
  wire  _T_2707; // @[MemPrimitives.scala 123:41:@17925.4]
  wire  _T_2708; // @[MemPrimitives.scala 123:41:@17926.4]
  wire  _T_2709; // @[MemPrimitives.scala 123:41:@17927.4]
  wire  _T_2710; // @[MemPrimitives.scala 123:41:@17928.4]
  wire  _T_2711; // @[MemPrimitives.scala 123:41:@17929.4]
  wire  _T_2712; // @[MemPrimitives.scala 123:41:@17930.4]
  wire  _T_2713; // @[MemPrimitives.scala 123:41:@17931.4]
  wire [9:0] _T_2715; // @[Cat.scala 30:58:@17933.4]
  wire [9:0] _T_2717; // @[Cat.scala 30:58:@17935.4]
  wire [9:0] _T_2719; // @[Cat.scala 30:58:@17937.4]
  wire [9:0] _T_2721; // @[Cat.scala 30:58:@17939.4]
  wire [9:0] _T_2723; // @[Cat.scala 30:58:@17941.4]
  wire [9:0] _T_2725; // @[Cat.scala 30:58:@17943.4]
  wire [9:0] _T_2727; // @[Cat.scala 30:58:@17945.4]
  wire [9:0] _T_2729; // @[Cat.scala 30:58:@17947.4]
  wire [9:0] _T_2731; // @[Cat.scala 30:58:@17949.4]
  wire [9:0] _T_2732; // @[Mux.scala 31:69:@17950.4]
  wire [9:0] _T_2733; // @[Mux.scala 31:69:@17951.4]
  wire [9:0] _T_2734; // @[Mux.scala 31:69:@17952.4]
  wire [9:0] _T_2735; // @[Mux.scala 31:69:@17953.4]
  wire [9:0] _T_2736; // @[Mux.scala 31:69:@17954.4]
  wire [9:0] _T_2737; // @[Mux.scala 31:69:@17955.4]
  wire [9:0] _T_2738; // @[Mux.scala 31:69:@17956.4]
  wire [9:0] _T_2739; // @[Mux.scala 31:69:@17957.4]
  wire  _T_2747; // @[MemPrimitives.scala 110:228:@17966.4]
  wire  _T_2753; // @[MemPrimitives.scala 110:228:@17970.4]
  wire  _T_2759; // @[MemPrimitives.scala 110:228:@17974.4]
  wire  _T_2765; // @[MemPrimitives.scala 110:228:@17978.4]
  wire  _T_2771; // @[MemPrimitives.scala 110:228:@17982.4]
  wire  _T_2777; // @[MemPrimitives.scala 110:228:@17986.4]
  wire  _T_2783; // @[MemPrimitives.scala 110:228:@17990.4]
  wire  _T_2789; // @[MemPrimitives.scala 110:228:@17994.4]
  wire  _T_2795; // @[MemPrimitives.scala 110:228:@17998.4]
  wire  _T_2797; // @[MemPrimitives.scala 123:41:@18012.4]
  wire  _T_2798; // @[MemPrimitives.scala 123:41:@18013.4]
  wire  _T_2799; // @[MemPrimitives.scala 123:41:@18014.4]
  wire  _T_2800; // @[MemPrimitives.scala 123:41:@18015.4]
  wire  _T_2801; // @[MemPrimitives.scala 123:41:@18016.4]
  wire  _T_2802; // @[MemPrimitives.scala 123:41:@18017.4]
  wire  _T_2803; // @[MemPrimitives.scala 123:41:@18018.4]
  wire  _T_2804; // @[MemPrimitives.scala 123:41:@18019.4]
  wire  _T_2805; // @[MemPrimitives.scala 123:41:@18020.4]
  wire [9:0] _T_2807; // @[Cat.scala 30:58:@18022.4]
  wire [9:0] _T_2809; // @[Cat.scala 30:58:@18024.4]
  wire [9:0] _T_2811; // @[Cat.scala 30:58:@18026.4]
  wire [9:0] _T_2813; // @[Cat.scala 30:58:@18028.4]
  wire [9:0] _T_2815; // @[Cat.scala 30:58:@18030.4]
  wire [9:0] _T_2817; // @[Cat.scala 30:58:@18032.4]
  wire [9:0] _T_2819; // @[Cat.scala 30:58:@18034.4]
  wire [9:0] _T_2821; // @[Cat.scala 30:58:@18036.4]
  wire [9:0] _T_2823; // @[Cat.scala 30:58:@18038.4]
  wire [9:0] _T_2824; // @[Mux.scala 31:69:@18039.4]
  wire [9:0] _T_2825; // @[Mux.scala 31:69:@18040.4]
  wire [9:0] _T_2826; // @[Mux.scala 31:69:@18041.4]
  wire [9:0] _T_2827; // @[Mux.scala 31:69:@18042.4]
  wire [9:0] _T_2828; // @[Mux.scala 31:69:@18043.4]
  wire [9:0] _T_2829; // @[Mux.scala 31:69:@18044.4]
  wire [9:0] _T_2830; // @[Mux.scala 31:69:@18045.4]
  wire [9:0] _T_2831; // @[Mux.scala 31:69:@18046.4]
  wire  _T_2836; // @[MemPrimitives.scala 110:210:@18053.4]
  wire  _T_2839; // @[MemPrimitives.scala 110:228:@18055.4]
  wire  _T_2842; // @[MemPrimitives.scala 110:210:@18057.4]
  wire  _T_2845; // @[MemPrimitives.scala 110:228:@18059.4]
  wire  _T_2848; // @[MemPrimitives.scala 110:210:@18061.4]
  wire  _T_2851; // @[MemPrimitives.scala 110:228:@18063.4]
  wire  _T_2854; // @[MemPrimitives.scala 110:210:@18065.4]
  wire  _T_2857; // @[MemPrimitives.scala 110:228:@18067.4]
  wire  _T_2860; // @[MemPrimitives.scala 110:210:@18069.4]
  wire  _T_2863; // @[MemPrimitives.scala 110:228:@18071.4]
  wire  _T_2866; // @[MemPrimitives.scala 110:210:@18073.4]
  wire  _T_2869; // @[MemPrimitives.scala 110:228:@18075.4]
  wire  _T_2872; // @[MemPrimitives.scala 110:210:@18077.4]
  wire  _T_2875; // @[MemPrimitives.scala 110:228:@18079.4]
  wire  _T_2878; // @[MemPrimitives.scala 110:210:@18081.4]
  wire  _T_2881; // @[MemPrimitives.scala 110:228:@18083.4]
  wire  _T_2884; // @[MemPrimitives.scala 110:210:@18085.4]
  wire  _T_2887; // @[MemPrimitives.scala 110:228:@18087.4]
  wire  _T_2889; // @[MemPrimitives.scala 123:41:@18101.4]
  wire  _T_2890; // @[MemPrimitives.scala 123:41:@18102.4]
  wire  _T_2891; // @[MemPrimitives.scala 123:41:@18103.4]
  wire  _T_2892; // @[MemPrimitives.scala 123:41:@18104.4]
  wire  _T_2893; // @[MemPrimitives.scala 123:41:@18105.4]
  wire  _T_2894; // @[MemPrimitives.scala 123:41:@18106.4]
  wire  _T_2895; // @[MemPrimitives.scala 123:41:@18107.4]
  wire  _T_2896; // @[MemPrimitives.scala 123:41:@18108.4]
  wire  _T_2897; // @[MemPrimitives.scala 123:41:@18109.4]
  wire [9:0] _T_2899; // @[Cat.scala 30:58:@18111.4]
  wire [9:0] _T_2901; // @[Cat.scala 30:58:@18113.4]
  wire [9:0] _T_2903; // @[Cat.scala 30:58:@18115.4]
  wire [9:0] _T_2905; // @[Cat.scala 30:58:@18117.4]
  wire [9:0] _T_2907; // @[Cat.scala 30:58:@18119.4]
  wire [9:0] _T_2909; // @[Cat.scala 30:58:@18121.4]
  wire [9:0] _T_2911; // @[Cat.scala 30:58:@18123.4]
  wire [9:0] _T_2913; // @[Cat.scala 30:58:@18125.4]
  wire [9:0] _T_2915; // @[Cat.scala 30:58:@18127.4]
  wire [9:0] _T_2916; // @[Mux.scala 31:69:@18128.4]
  wire [9:0] _T_2917; // @[Mux.scala 31:69:@18129.4]
  wire [9:0] _T_2918; // @[Mux.scala 31:69:@18130.4]
  wire [9:0] _T_2919; // @[Mux.scala 31:69:@18131.4]
  wire [9:0] _T_2920; // @[Mux.scala 31:69:@18132.4]
  wire [9:0] _T_2921; // @[Mux.scala 31:69:@18133.4]
  wire [9:0] _T_2922; // @[Mux.scala 31:69:@18134.4]
  wire [9:0] _T_2923; // @[Mux.scala 31:69:@18135.4]
  wire  _T_2928; // @[MemPrimitives.scala 110:210:@18142.4]
  wire  _T_2931; // @[MemPrimitives.scala 110:228:@18144.4]
  wire  _T_2934; // @[MemPrimitives.scala 110:210:@18146.4]
  wire  _T_2937; // @[MemPrimitives.scala 110:228:@18148.4]
  wire  _T_2940; // @[MemPrimitives.scala 110:210:@18150.4]
  wire  _T_2943; // @[MemPrimitives.scala 110:228:@18152.4]
  wire  _T_2946; // @[MemPrimitives.scala 110:210:@18154.4]
  wire  _T_2949; // @[MemPrimitives.scala 110:228:@18156.4]
  wire  _T_2952; // @[MemPrimitives.scala 110:210:@18158.4]
  wire  _T_2955; // @[MemPrimitives.scala 110:228:@18160.4]
  wire  _T_2958; // @[MemPrimitives.scala 110:210:@18162.4]
  wire  _T_2961; // @[MemPrimitives.scala 110:228:@18164.4]
  wire  _T_2964; // @[MemPrimitives.scala 110:210:@18166.4]
  wire  _T_2967; // @[MemPrimitives.scala 110:228:@18168.4]
  wire  _T_2970; // @[MemPrimitives.scala 110:210:@18170.4]
  wire  _T_2973; // @[MemPrimitives.scala 110:228:@18172.4]
  wire  _T_2976; // @[MemPrimitives.scala 110:210:@18174.4]
  wire  _T_2979; // @[MemPrimitives.scala 110:228:@18176.4]
  wire  _T_2981; // @[MemPrimitives.scala 123:41:@18190.4]
  wire  _T_2982; // @[MemPrimitives.scala 123:41:@18191.4]
  wire  _T_2983; // @[MemPrimitives.scala 123:41:@18192.4]
  wire  _T_2984; // @[MemPrimitives.scala 123:41:@18193.4]
  wire  _T_2985; // @[MemPrimitives.scala 123:41:@18194.4]
  wire  _T_2986; // @[MemPrimitives.scala 123:41:@18195.4]
  wire  _T_2987; // @[MemPrimitives.scala 123:41:@18196.4]
  wire  _T_2988; // @[MemPrimitives.scala 123:41:@18197.4]
  wire  _T_2989; // @[MemPrimitives.scala 123:41:@18198.4]
  wire [9:0] _T_2991; // @[Cat.scala 30:58:@18200.4]
  wire [9:0] _T_2993; // @[Cat.scala 30:58:@18202.4]
  wire [9:0] _T_2995; // @[Cat.scala 30:58:@18204.4]
  wire [9:0] _T_2997; // @[Cat.scala 30:58:@18206.4]
  wire [9:0] _T_2999; // @[Cat.scala 30:58:@18208.4]
  wire [9:0] _T_3001; // @[Cat.scala 30:58:@18210.4]
  wire [9:0] _T_3003; // @[Cat.scala 30:58:@18212.4]
  wire [9:0] _T_3005; // @[Cat.scala 30:58:@18214.4]
  wire [9:0] _T_3007; // @[Cat.scala 30:58:@18216.4]
  wire [9:0] _T_3008; // @[Mux.scala 31:69:@18217.4]
  wire [9:0] _T_3009; // @[Mux.scala 31:69:@18218.4]
  wire [9:0] _T_3010; // @[Mux.scala 31:69:@18219.4]
  wire [9:0] _T_3011; // @[Mux.scala 31:69:@18220.4]
  wire [9:0] _T_3012; // @[Mux.scala 31:69:@18221.4]
  wire [9:0] _T_3013; // @[Mux.scala 31:69:@18222.4]
  wire [9:0] _T_3014; // @[Mux.scala 31:69:@18223.4]
  wire [9:0] _T_3015; // @[Mux.scala 31:69:@18224.4]
  wire  _T_3023; // @[MemPrimitives.scala 110:228:@18233.4]
  wire  _T_3029; // @[MemPrimitives.scala 110:228:@18237.4]
  wire  _T_3035; // @[MemPrimitives.scala 110:228:@18241.4]
  wire  _T_3041; // @[MemPrimitives.scala 110:228:@18245.4]
  wire  _T_3047; // @[MemPrimitives.scala 110:228:@18249.4]
  wire  _T_3053; // @[MemPrimitives.scala 110:228:@18253.4]
  wire  _T_3059; // @[MemPrimitives.scala 110:228:@18257.4]
  wire  _T_3065; // @[MemPrimitives.scala 110:228:@18261.4]
  wire  _T_3071; // @[MemPrimitives.scala 110:228:@18265.4]
  wire  _T_3073; // @[MemPrimitives.scala 123:41:@18279.4]
  wire  _T_3074; // @[MemPrimitives.scala 123:41:@18280.4]
  wire  _T_3075; // @[MemPrimitives.scala 123:41:@18281.4]
  wire  _T_3076; // @[MemPrimitives.scala 123:41:@18282.4]
  wire  _T_3077; // @[MemPrimitives.scala 123:41:@18283.4]
  wire  _T_3078; // @[MemPrimitives.scala 123:41:@18284.4]
  wire  _T_3079; // @[MemPrimitives.scala 123:41:@18285.4]
  wire  _T_3080; // @[MemPrimitives.scala 123:41:@18286.4]
  wire  _T_3081; // @[MemPrimitives.scala 123:41:@18287.4]
  wire [9:0] _T_3083; // @[Cat.scala 30:58:@18289.4]
  wire [9:0] _T_3085; // @[Cat.scala 30:58:@18291.4]
  wire [9:0] _T_3087; // @[Cat.scala 30:58:@18293.4]
  wire [9:0] _T_3089; // @[Cat.scala 30:58:@18295.4]
  wire [9:0] _T_3091; // @[Cat.scala 30:58:@18297.4]
  wire [9:0] _T_3093; // @[Cat.scala 30:58:@18299.4]
  wire [9:0] _T_3095; // @[Cat.scala 30:58:@18301.4]
  wire [9:0] _T_3097; // @[Cat.scala 30:58:@18303.4]
  wire [9:0] _T_3099; // @[Cat.scala 30:58:@18305.4]
  wire [9:0] _T_3100; // @[Mux.scala 31:69:@18306.4]
  wire [9:0] _T_3101; // @[Mux.scala 31:69:@18307.4]
  wire [9:0] _T_3102; // @[Mux.scala 31:69:@18308.4]
  wire [9:0] _T_3103; // @[Mux.scala 31:69:@18309.4]
  wire [9:0] _T_3104; // @[Mux.scala 31:69:@18310.4]
  wire [9:0] _T_3105; // @[Mux.scala 31:69:@18311.4]
  wire [9:0] _T_3106; // @[Mux.scala 31:69:@18312.4]
  wire [9:0] _T_3107; // @[Mux.scala 31:69:@18313.4]
  wire  _T_3115; // @[MemPrimitives.scala 110:228:@18322.4]
  wire  _T_3121; // @[MemPrimitives.scala 110:228:@18326.4]
  wire  _T_3127; // @[MemPrimitives.scala 110:228:@18330.4]
  wire  _T_3133; // @[MemPrimitives.scala 110:228:@18334.4]
  wire  _T_3139; // @[MemPrimitives.scala 110:228:@18338.4]
  wire  _T_3145; // @[MemPrimitives.scala 110:228:@18342.4]
  wire  _T_3151; // @[MemPrimitives.scala 110:228:@18346.4]
  wire  _T_3157; // @[MemPrimitives.scala 110:228:@18350.4]
  wire  _T_3163; // @[MemPrimitives.scala 110:228:@18354.4]
  wire  _T_3165; // @[MemPrimitives.scala 123:41:@18368.4]
  wire  _T_3166; // @[MemPrimitives.scala 123:41:@18369.4]
  wire  _T_3167; // @[MemPrimitives.scala 123:41:@18370.4]
  wire  _T_3168; // @[MemPrimitives.scala 123:41:@18371.4]
  wire  _T_3169; // @[MemPrimitives.scala 123:41:@18372.4]
  wire  _T_3170; // @[MemPrimitives.scala 123:41:@18373.4]
  wire  _T_3171; // @[MemPrimitives.scala 123:41:@18374.4]
  wire  _T_3172; // @[MemPrimitives.scala 123:41:@18375.4]
  wire  _T_3173; // @[MemPrimitives.scala 123:41:@18376.4]
  wire [9:0] _T_3175; // @[Cat.scala 30:58:@18378.4]
  wire [9:0] _T_3177; // @[Cat.scala 30:58:@18380.4]
  wire [9:0] _T_3179; // @[Cat.scala 30:58:@18382.4]
  wire [9:0] _T_3181; // @[Cat.scala 30:58:@18384.4]
  wire [9:0] _T_3183; // @[Cat.scala 30:58:@18386.4]
  wire [9:0] _T_3185; // @[Cat.scala 30:58:@18388.4]
  wire [9:0] _T_3187; // @[Cat.scala 30:58:@18390.4]
  wire [9:0] _T_3189; // @[Cat.scala 30:58:@18392.4]
  wire [9:0] _T_3191; // @[Cat.scala 30:58:@18394.4]
  wire [9:0] _T_3192; // @[Mux.scala 31:69:@18395.4]
  wire [9:0] _T_3193; // @[Mux.scala 31:69:@18396.4]
  wire [9:0] _T_3194; // @[Mux.scala 31:69:@18397.4]
  wire [9:0] _T_3195; // @[Mux.scala 31:69:@18398.4]
  wire [9:0] _T_3196; // @[Mux.scala 31:69:@18399.4]
  wire [9:0] _T_3197; // @[Mux.scala 31:69:@18400.4]
  wire [9:0] _T_3198; // @[Mux.scala 31:69:@18401.4]
  wire [9:0] _T_3199; // @[Mux.scala 31:69:@18402.4]
  wire  _T_3207; // @[MemPrimitives.scala 110:228:@18411.4]
  wire  _T_3213; // @[MemPrimitives.scala 110:228:@18415.4]
  wire  _T_3219; // @[MemPrimitives.scala 110:228:@18419.4]
  wire  _T_3225; // @[MemPrimitives.scala 110:228:@18423.4]
  wire  _T_3231; // @[MemPrimitives.scala 110:228:@18427.4]
  wire  _T_3237; // @[MemPrimitives.scala 110:228:@18431.4]
  wire  _T_3243; // @[MemPrimitives.scala 110:228:@18435.4]
  wire  _T_3249; // @[MemPrimitives.scala 110:228:@18439.4]
  wire  _T_3255; // @[MemPrimitives.scala 110:228:@18443.4]
  wire  _T_3257; // @[MemPrimitives.scala 123:41:@18457.4]
  wire  _T_3258; // @[MemPrimitives.scala 123:41:@18458.4]
  wire  _T_3259; // @[MemPrimitives.scala 123:41:@18459.4]
  wire  _T_3260; // @[MemPrimitives.scala 123:41:@18460.4]
  wire  _T_3261; // @[MemPrimitives.scala 123:41:@18461.4]
  wire  _T_3262; // @[MemPrimitives.scala 123:41:@18462.4]
  wire  _T_3263; // @[MemPrimitives.scala 123:41:@18463.4]
  wire  _T_3264; // @[MemPrimitives.scala 123:41:@18464.4]
  wire  _T_3265; // @[MemPrimitives.scala 123:41:@18465.4]
  wire [9:0] _T_3267; // @[Cat.scala 30:58:@18467.4]
  wire [9:0] _T_3269; // @[Cat.scala 30:58:@18469.4]
  wire [9:0] _T_3271; // @[Cat.scala 30:58:@18471.4]
  wire [9:0] _T_3273; // @[Cat.scala 30:58:@18473.4]
  wire [9:0] _T_3275; // @[Cat.scala 30:58:@18475.4]
  wire [9:0] _T_3277; // @[Cat.scala 30:58:@18477.4]
  wire [9:0] _T_3279; // @[Cat.scala 30:58:@18479.4]
  wire [9:0] _T_3281; // @[Cat.scala 30:58:@18481.4]
  wire [9:0] _T_3283; // @[Cat.scala 30:58:@18483.4]
  wire [9:0] _T_3284; // @[Mux.scala 31:69:@18484.4]
  wire [9:0] _T_3285; // @[Mux.scala 31:69:@18485.4]
  wire [9:0] _T_3286; // @[Mux.scala 31:69:@18486.4]
  wire [9:0] _T_3287; // @[Mux.scala 31:69:@18487.4]
  wire [9:0] _T_3288; // @[Mux.scala 31:69:@18488.4]
  wire [9:0] _T_3289; // @[Mux.scala 31:69:@18489.4]
  wire [9:0] _T_3290; // @[Mux.scala 31:69:@18490.4]
  wire [9:0] _T_3291; // @[Mux.scala 31:69:@18491.4]
  wire  _T_3299; // @[MemPrimitives.scala 110:228:@18500.4]
  wire  _T_3305; // @[MemPrimitives.scala 110:228:@18504.4]
  wire  _T_3311; // @[MemPrimitives.scala 110:228:@18508.4]
  wire  _T_3317; // @[MemPrimitives.scala 110:228:@18512.4]
  wire  _T_3323; // @[MemPrimitives.scala 110:228:@18516.4]
  wire  _T_3329; // @[MemPrimitives.scala 110:228:@18520.4]
  wire  _T_3335; // @[MemPrimitives.scala 110:228:@18524.4]
  wire  _T_3341; // @[MemPrimitives.scala 110:228:@18528.4]
  wire  _T_3347; // @[MemPrimitives.scala 110:228:@18532.4]
  wire  _T_3349; // @[MemPrimitives.scala 123:41:@18546.4]
  wire  _T_3350; // @[MemPrimitives.scala 123:41:@18547.4]
  wire  _T_3351; // @[MemPrimitives.scala 123:41:@18548.4]
  wire  _T_3352; // @[MemPrimitives.scala 123:41:@18549.4]
  wire  _T_3353; // @[MemPrimitives.scala 123:41:@18550.4]
  wire  _T_3354; // @[MemPrimitives.scala 123:41:@18551.4]
  wire  _T_3355; // @[MemPrimitives.scala 123:41:@18552.4]
  wire  _T_3356; // @[MemPrimitives.scala 123:41:@18553.4]
  wire  _T_3357; // @[MemPrimitives.scala 123:41:@18554.4]
  wire [9:0] _T_3359; // @[Cat.scala 30:58:@18556.4]
  wire [9:0] _T_3361; // @[Cat.scala 30:58:@18558.4]
  wire [9:0] _T_3363; // @[Cat.scala 30:58:@18560.4]
  wire [9:0] _T_3365; // @[Cat.scala 30:58:@18562.4]
  wire [9:0] _T_3367; // @[Cat.scala 30:58:@18564.4]
  wire [9:0] _T_3369; // @[Cat.scala 30:58:@18566.4]
  wire [9:0] _T_3371; // @[Cat.scala 30:58:@18568.4]
  wire [9:0] _T_3373; // @[Cat.scala 30:58:@18570.4]
  wire [9:0] _T_3375; // @[Cat.scala 30:58:@18572.4]
  wire [9:0] _T_3376; // @[Mux.scala 31:69:@18573.4]
  wire [9:0] _T_3377; // @[Mux.scala 31:69:@18574.4]
  wire [9:0] _T_3378; // @[Mux.scala 31:69:@18575.4]
  wire [9:0] _T_3379; // @[Mux.scala 31:69:@18576.4]
  wire [9:0] _T_3380; // @[Mux.scala 31:69:@18577.4]
  wire [9:0] _T_3381; // @[Mux.scala 31:69:@18578.4]
  wire [9:0] _T_3382; // @[Mux.scala 31:69:@18579.4]
  wire [9:0] _T_3383; // @[Mux.scala 31:69:@18580.4]
  wire  _T_3479; // @[package.scala 96:25:@18709.4 package.scala 96:25:@18710.4]
  wire [7:0] _T_3483; // @[Mux.scala 31:69:@18719.4]
  wire  _T_3476; // @[package.scala 96:25:@18701.4 package.scala 96:25:@18702.4]
  wire [7:0] _T_3484; // @[Mux.scala 31:69:@18720.4]
  wire  _T_3473; // @[package.scala 96:25:@18693.4 package.scala 96:25:@18694.4]
  wire [7:0] _T_3485; // @[Mux.scala 31:69:@18721.4]
  wire  _T_3470; // @[package.scala 96:25:@18685.4 package.scala 96:25:@18686.4]
  wire [7:0] _T_3486; // @[Mux.scala 31:69:@18722.4]
  wire  _T_3467; // @[package.scala 96:25:@18677.4 package.scala 96:25:@18678.4]
  wire [7:0] _T_3487; // @[Mux.scala 31:69:@18723.4]
  wire  _T_3464; // @[package.scala 96:25:@18669.4 package.scala 96:25:@18670.4]
  wire [7:0] _T_3488; // @[Mux.scala 31:69:@18724.4]
  wire  _T_3461; // @[package.scala 96:25:@18661.4 package.scala 96:25:@18662.4]
  wire [7:0] _T_3489; // @[Mux.scala 31:69:@18725.4]
  wire  _T_3458; // @[package.scala 96:25:@18653.4 package.scala 96:25:@18654.4]
  wire [7:0] _T_3490; // @[Mux.scala 31:69:@18726.4]
  wire  _T_3455; // @[package.scala 96:25:@18645.4 package.scala 96:25:@18646.4]
  wire [7:0] _T_3491; // @[Mux.scala 31:69:@18727.4]
  wire  _T_3452; // @[package.scala 96:25:@18637.4 package.scala 96:25:@18638.4]
  wire [7:0] _T_3492; // @[Mux.scala 31:69:@18728.4]
  wire  _T_3449; // @[package.scala 96:25:@18629.4 package.scala 96:25:@18630.4]
  wire  _T_3586; // @[package.scala 96:25:@18853.4 package.scala 96:25:@18854.4]
  wire [7:0] _T_3590; // @[Mux.scala 31:69:@18863.4]
  wire  _T_3583; // @[package.scala 96:25:@18845.4 package.scala 96:25:@18846.4]
  wire [7:0] _T_3591; // @[Mux.scala 31:69:@18864.4]
  wire  _T_3580; // @[package.scala 96:25:@18837.4 package.scala 96:25:@18838.4]
  wire [7:0] _T_3592; // @[Mux.scala 31:69:@18865.4]
  wire  _T_3577; // @[package.scala 96:25:@18829.4 package.scala 96:25:@18830.4]
  wire [7:0] _T_3593; // @[Mux.scala 31:69:@18866.4]
  wire  _T_3574; // @[package.scala 96:25:@18821.4 package.scala 96:25:@18822.4]
  wire [7:0] _T_3594; // @[Mux.scala 31:69:@18867.4]
  wire  _T_3571; // @[package.scala 96:25:@18813.4 package.scala 96:25:@18814.4]
  wire [7:0] _T_3595; // @[Mux.scala 31:69:@18868.4]
  wire  _T_3568; // @[package.scala 96:25:@18805.4 package.scala 96:25:@18806.4]
  wire [7:0] _T_3596; // @[Mux.scala 31:69:@18869.4]
  wire  _T_3565; // @[package.scala 96:25:@18797.4 package.scala 96:25:@18798.4]
  wire [7:0] _T_3597; // @[Mux.scala 31:69:@18870.4]
  wire  _T_3562; // @[package.scala 96:25:@18789.4 package.scala 96:25:@18790.4]
  wire [7:0] _T_3598; // @[Mux.scala 31:69:@18871.4]
  wire  _T_3559; // @[package.scala 96:25:@18781.4 package.scala 96:25:@18782.4]
  wire [7:0] _T_3599; // @[Mux.scala 31:69:@18872.4]
  wire  _T_3556; // @[package.scala 96:25:@18773.4 package.scala 96:25:@18774.4]
  wire  _T_3693; // @[package.scala 96:25:@18997.4 package.scala 96:25:@18998.4]
  wire [7:0] _T_3697; // @[Mux.scala 31:69:@19007.4]
  wire  _T_3690; // @[package.scala 96:25:@18989.4 package.scala 96:25:@18990.4]
  wire [7:0] _T_3698; // @[Mux.scala 31:69:@19008.4]
  wire  _T_3687; // @[package.scala 96:25:@18981.4 package.scala 96:25:@18982.4]
  wire [7:0] _T_3699; // @[Mux.scala 31:69:@19009.4]
  wire  _T_3684; // @[package.scala 96:25:@18973.4 package.scala 96:25:@18974.4]
  wire [7:0] _T_3700; // @[Mux.scala 31:69:@19010.4]
  wire  _T_3681; // @[package.scala 96:25:@18965.4 package.scala 96:25:@18966.4]
  wire [7:0] _T_3701; // @[Mux.scala 31:69:@19011.4]
  wire  _T_3678; // @[package.scala 96:25:@18957.4 package.scala 96:25:@18958.4]
  wire [7:0] _T_3702; // @[Mux.scala 31:69:@19012.4]
  wire  _T_3675; // @[package.scala 96:25:@18949.4 package.scala 96:25:@18950.4]
  wire [7:0] _T_3703; // @[Mux.scala 31:69:@19013.4]
  wire  _T_3672; // @[package.scala 96:25:@18941.4 package.scala 96:25:@18942.4]
  wire [7:0] _T_3704; // @[Mux.scala 31:69:@19014.4]
  wire  _T_3669; // @[package.scala 96:25:@18933.4 package.scala 96:25:@18934.4]
  wire [7:0] _T_3705; // @[Mux.scala 31:69:@19015.4]
  wire  _T_3666; // @[package.scala 96:25:@18925.4 package.scala 96:25:@18926.4]
  wire [7:0] _T_3706; // @[Mux.scala 31:69:@19016.4]
  wire  _T_3663; // @[package.scala 96:25:@18917.4 package.scala 96:25:@18918.4]
  wire  _T_3800; // @[package.scala 96:25:@19141.4 package.scala 96:25:@19142.4]
  wire [7:0] _T_3804; // @[Mux.scala 31:69:@19151.4]
  wire  _T_3797; // @[package.scala 96:25:@19133.4 package.scala 96:25:@19134.4]
  wire [7:0] _T_3805; // @[Mux.scala 31:69:@19152.4]
  wire  _T_3794; // @[package.scala 96:25:@19125.4 package.scala 96:25:@19126.4]
  wire [7:0] _T_3806; // @[Mux.scala 31:69:@19153.4]
  wire  _T_3791; // @[package.scala 96:25:@19117.4 package.scala 96:25:@19118.4]
  wire [7:0] _T_3807; // @[Mux.scala 31:69:@19154.4]
  wire  _T_3788; // @[package.scala 96:25:@19109.4 package.scala 96:25:@19110.4]
  wire [7:0] _T_3808; // @[Mux.scala 31:69:@19155.4]
  wire  _T_3785; // @[package.scala 96:25:@19101.4 package.scala 96:25:@19102.4]
  wire [7:0] _T_3809; // @[Mux.scala 31:69:@19156.4]
  wire  _T_3782; // @[package.scala 96:25:@19093.4 package.scala 96:25:@19094.4]
  wire [7:0] _T_3810; // @[Mux.scala 31:69:@19157.4]
  wire  _T_3779; // @[package.scala 96:25:@19085.4 package.scala 96:25:@19086.4]
  wire [7:0] _T_3811; // @[Mux.scala 31:69:@19158.4]
  wire  _T_3776; // @[package.scala 96:25:@19077.4 package.scala 96:25:@19078.4]
  wire [7:0] _T_3812; // @[Mux.scala 31:69:@19159.4]
  wire  _T_3773; // @[package.scala 96:25:@19069.4 package.scala 96:25:@19070.4]
  wire [7:0] _T_3813; // @[Mux.scala 31:69:@19160.4]
  wire  _T_3770; // @[package.scala 96:25:@19061.4 package.scala 96:25:@19062.4]
  wire  _T_3907; // @[package.scala 96:25:@19285.4 package.scala 96:25:@19286.4]
  wire [7:0] _T_3911; // @[Mux.scala 31:69:@19295.4]
  wire  _T_3904; // @[package.scala 96:25:@19277.4 package.scala 96:25:@19278.4]
  wire [7:0] _T_3912; // @[Mux.scala 31:69:@19296.4]
  wire  _T_3901; // @[package.scala 96:25:@19269.4 package.scala 96:25:@19270.4]
  wire [7:0] _T_3913; // @[Mux.scala 31:69:@19297.4]
  wire  _T_3898; // @[package.scala 96:25:@19261.4 package.scala 96:25:@19262.4]
  wire [7:0] _T_3914; // @[Mux.scala 31:69:@19298.4]
  wire  _T_3895; // @[package.scala 96:25:@19253.4 package.scala 96:25:@19254.4]
  wire [7:0] _T_3915; // @[Mux.scala 31:69:@19299.4]
  wire  _T_3892; // @[package.scala 96:25:@19245.4 package.scala 96:25:@19246.4]
  wire [7:0] _T_3916; // @[Mux.scala 31:69:@19300.4]
  wire  _T_3889; // @[package.scala 96:25:@19237.4 package.scala 96:25:@19238.4]
  wire [7:0] _T_3917; // @[Mux.scala 31:69:@19301.4]
  wire  _T_3886; // @[package.scala 96:25:@19229.4 package.scala 96:25:@19230.4]
  wire [7:0] _T_3918; // @[Mux.scala 31:69:@19302.4]
  wire  _T_3883; // @[package.scala 96:25:@19221.4 package.scala 96:25:@19222.4]
  wire [7:0] _T_3919; // @[Mux.scala 31:69:@19303.4]
  wire  _T_3880; // @[package.scala 96:25:@19213.4 package.scala 96:25:@19214.4]
  wire [7:0] _T_3920; // @[Mux.scala 31:69:@19304.4]
  wire  _T_3877; // @[package.scala 96:25:@19205.4 package.scala 96:25:@19206.4]
  wire  _T_4014; // @[package.scala 96:25:@19429.4 package.scala 96:25:@19430.4]
  wire [7:0] _T_4018; // @[Mux.scala 31:69:@19439.4]
  wire  _T_4011; // @[package.scala 96:25:@19421.4 package.scala 96:25:@19422.4]
  wire [7:0] _T_4019; // @[Mux.scala 31:69:@19440.4]
  wire  _T_4008; // @[package.scala 96:25:@19413.4 package.scala 96:25:@19414.4]
  wire [7:0] _T_4020; // @[Mux.scala 31:69:@19441.4]
  wire  _T_4005; // @[package.scala 96:25:@19405.4 package.scala 96:25:@19406.4]
  wire [7:0] _T_4021; // @[Mux.scala 31:69:@19442.4]
  wire  _T_4002; // @[package.scala 96:25:@19397.4 package.scala 96:25:@19398.4]
  wire [7:0] _T_4022; // @[Mux.scala 31:69:@19443.4]
  wire  _T_3999; // @[package.scala 96:25:@19389.4 package.scala 96:25:@19390.4]
  wire [7:0] _T_4023; // @[Mux.scala 31:69:@19444.4]
  wire  _T_3996; // @[package.scala 96:25:@19381.4 package.scala 96:25:@19382.4]
  wire [7:0] _T_4024; // @[Mux.scala 31:69:@19445.4]
  wire  _T_3993; // @[package.scala 96:25:@19373.4 package.scala 96:25:@19374.4]
  wire [7:0] _T_4025; // @[Mux.scala 31:69:@19446.4]
  wire  _T_3990; // @[package.scala 96:25:@19365.4 package.scala 96:25:@19366.4]
  wire [7:0] _T_4026; // @[Mux.scala 31:69:@19447.4]
  wire  _T_3987; // @[package.scala 96:25:@19357.4 package.scala 96:25:@19358.4]
  wire [7:0] _T_4027; // @[Mux.scala 31:69:@19448.4]
  wire  _T_3984; // @[package.scala 96:25:@19349.4 package.scala 96:25:@19350.4]
  wire  _T_4121; // @[package.scala 96:25:@19573.4 package.scala 96:25:@19574.4]
  wire [7:0] _T_4125; // @[Mux.scala 31:69:@19583.4]
  wire  _T_4118; // @[package.scala 96:25:@19565.4 package.scala 96:25:@19566.4]
  wire [7:0] _T_4126; // @[Mux.scala 31:69:@19584.4]
  wire  _T_4115; // @[package.scala 96:25:@19557.4 package.scala 96:25:@19558.4]
  wire [7:0] _T_4127; // @[Mux.scala 31:69:@19585.4]
  wire  _T_4112; // @[package.scala 96:25:@19549.4 package.scala 96:25:@19550.4]
  wire [7:0] _T_4128; // @[Mux.scala 31:69:@19586.4]
  wire  _T_4109; // @[package.scala 96:25:@19541.4 package.scala 96:25:@19542.4]
  wire [7:0] _T_4129; // @[Mux.scala 31:69:@19587.4]
  wire  _T_4106; // @[package.scala 96:25:@19533.4 package.scala 96:25:@19534.4]
  wire [7:0] _T_4130; // @[Mux.scala 31:69:@19588.4]
  wire  _T_4103; // @[package.scala 96:25:@19525.4 package.scala 96:25:@19526.4]
  wire [7:0] _T_4131; // @[Mux.scala 31:69:@19589.4]
  wire  _T_4100; // @[package.scala 96:25:@19517.4 package.scala 96:25:@19518.4]
  wire [7:0] _T_4132; // @[Mux.scala 31:69:@19590.4]
  wire  _T_4097; // @[package.scala 96:25:@19509.4 package.scala 96:25:@19510.4]
  wire [7:0] _T_4133; // @[Mux.scala 31:69:@19591.4]
  wire  _T_4094; // @[package.scala 96:25:@19501.4 package.scala 96:25:@19502.4]
  wire [7:0] _T_4134; // @[Mux.scala 31:69:@19592.4]
  wire  _T_4091; // @[package.scala 96:25:@19493.4 package.scala 96:25:@19494.4]
  wire  _T_4228; // @[package.scala 96:25:@19717.4 package.scala 96:25:@19718.4]
  wire [7:0] _T_4232; // @[Mux.scala 31:69:@19727.4]
  wire  _T_4225; // @[package.scala 96:25:@19709.4 package.scala 96:25:@19710.4]
  wire [7:0] _T_4233; // @[Mux.scala 31:69:@19728.4]
  wire  _T_4222; // @[package.scala 96:25:@19701.4 package.scala 96:25:@19702.4]
  wire [7:0] _T_4234; // @[Mux.scala 31:69:@19729.4]
  wire  _T_4219; // @[package.scala 96:25:@19693.4 package.scala 96:25:@19694.4]
  wire [7:0] _T_4235; // @[Mux.scala 31:69:@19730.4]
  wire  _T_4216; // @[package.scala 96:25:@19685.4 package.scala 96:25:@19686.4]
  wire [7:0] _T_4236; // @[Mux.scala 31:69:@19731.4]
  wire  _T_4213; // @[package.scala 96:25:@19677.4 package.scala 96:25:@19678.4]
  wire [7:0] _T_4237; // @[Mux.scala 31:69:@19732.4]
  wire  _T_4210; // @[package.scala 96:25:@19669.4 package.scala 96:25:@19670.4]
  wire [7:0] _T_4238; // @[Mux.scala 31:69:@19733.4]
  wire  _T_4207; // @[package.scala 96:25:@19661.4 package.scala 96:25:@19662.4]
  wire [7:0] _T_4239; // @[Mux.scala 31:69:@19734.4]
  wire  _T_4204; // @[package.scala 96:25:@19653.4 package.scala 96:25:@19654.4]
  wire [7:0] _T_4240; // @[Mux.scala 31:69:@19735.4]
  wire  _T_4201; // @[package.scala 96:25:@19645.4 package.scala 96:25:@19646.4]
  wire [7:0] _T_4241; // @[Mux.scala 31:69:@19736.4]
  wire  _T_4198; // @[package.scala 96:25:@19637.4 package.scala 96:25:@19638.4]
  wire  _T_4335; // @[package.scala 96:25:@19861.4 package.scala 96:25:@19862.4]
  wire [7:0] _T_4339; // @[Mux.scala 31:69:@19871.4]
  wire  _T_4332; // @[package.scala 96:25:@19853.4 package.scala 96:25:@19854.4]
  wire [7:0] _T_4340; // @[Mux.scala 31:69:@19872.4]
  wire  _T_4329; // @[package.scala 96:25:@19845.4 package.scala 96:25:@19846.4]
  wire [7:0] _T_4341; // @[Mux.scala 31:69:@19873.4]
  wire  _T_4326; // @[package.scala 96:25:@19837.4 package.scala 96:25:@19838.4]
  wire [7:0] _T_4342; // @[Mux.scala 31:69:@19874.4]
  wire  _T_4323; // @[package.scala 96:25:@19829.4 package.scala 96:25:@19830.4]
  wire [7:0] _T_4343; // @[Mux.scala 31:69:@19875.4]
  wire  _T_4320; // @[package.scala 96:25:@19821.4 package.scala 96:25:@19822.4]
  wire [7:0] _T_4344; // @[Mux.scala 31:69:@19876.4]
  wire  _T_4317; // @[package.scala 96:25:@19813.4 package.scala 96:25:@19814.4]
  wire [7:0] _T_4345; // @[Mux.scala 31:69:@19877.4]
  wire  _T_4314; // @[package.scala 96:25:@19805.4 package.scala 96:25:@19806.4]
  wire [7:0] _T_4346; // @[Mux.scala 31:69:@19878.4]
  wire  _T_4311; // @[package.scala 96:25:@19797.4 package.scala 96:25:@19798.4]
  wire [7:0] _T_4347; // @[Mux.scala 31:69:@19879.4]
  wire  _T_4308; // @[package.scala 96:25:@19789.4 package.scala 96:25:@19790.4]
  wire [7:0] _T_4348; // @[Mux.scala 31:69:@19880.4]
  wire  _T_4305; // @[package.scala 96:25:@19781.4 package.scala 96:25:@19782.4]
  wire  _T_4442; // @[package.scala 96:25:@20005.4 package.scala 96:25:@20006.4]
  wire [7:0] _T_4446; // @[Mux.scala 31:69:@20015.4]
  wire  _T_4439; // @[package.scala 96:25:@19997.4 package.scala 96:25:@19998.4]
  wire [7:0] _T_4447; // @[Mux.scala 31:69:@20016.4]
  wire  _T_4436; // @[package.scala 96:25:@19989.4 package.scala 96:25:@19990.4]
  wire [7:0] _T_4448; // @[Mux.scala 31:69:@20017.4]
  wire  _T_4433; // @[package.scala 96:25:@19981.4 package.scala 96:25:@19982.4]
  wire [7:0] _T_4449; // @[Mux.scala 31:69:@20018.4]
  wire  _T_4430; // @[package.scala 96:25:@19973.4 package.scala 96:25:@19974.4]
  wire [7:0] _T_4450; // @[Mux.scala 31:69:@20019.4]
  wire  _T_4427; // @[package.scala 96:25:@19965.4 package.scala 96:25:@19966.4]
  wire [7:0] _T_4451; // @[Mux.scala 31:69:@20020.4]
  wire  _T_4424; // @[package.scala 96:25:@19957.4 package.scala 96:25:@19958.4]
  wire [7:0] _T_4452; // @[Mux.scala 31:69:@20021.4]
  wire  _T_4421; // @[package.scala 96:25:@19949.4 package.scala 96:25:@19950.4]
  wire [7:0] _T_4453; // @[Mux.scala 31:69:@20022.4]
  wire  _T_4418; // @[package.scala 96:25:@19941.4 package.scala 96:25:@19942.4]
  wire [7:0] _T_4454; // @[Mux.scala 31:69:@20023.4]
  wire  _T_4415; // @[package.scala 96:25:@19933.4 package.scala 96:25:@19934.4]
  wire [7:0] _T_4455; // @[Mux.scala 31:69:@20024.4]
  wire  _T_4412; // @[package.scala 96:25:@19925.4 package.scala 96:25:@19926.4]
  wire  _T_4549; // @[package.scala 96:25:@20149.4 package.scala 96:25:@20150.4]
  wire [7:0] _T_4553; // @[Mux.scala 31:69:@20159.4]
  wire  _T_4546; // @[package.scala 96:25:@20141.4 package.scala 96:25:@20142.4]
  wire [7:0] _T_4554; // @[Mux.scala 31:69:@20160.4]
  wire  _T_4543; // @[package.scala 96:25:@20133.4 package.scala 96:25:@20134.4]
  wire [7:0] _T_4555; // @[Mux.scala 31:69:@20161.4]
  wire  _T_4540; // @[package.scala 96:25:@20125.4 package.scala 96:25:@20126.4]
  wire [7:0] _T_4556; // @[Mux.scala 31:69:@20162.4]
  wire  _T_4537; // @[package.scala 96:25:@20117.4 package.scala 96:25:@20118.4]
  wire [7:0] _T_4557; // @[Mux.scala 31:69:@20163.4]
  wire  _T_4534; // @[package.scala 96:25:@20109.4 package.scala 96:25:@20110.4]
  wire [7:0] _T_4558; // @[Mux.scala 31:69:@20164.4]
  wire  _T_4531; // @[package.scala 96:25:@20101.4 package.scala 96:25:@20102.4]
  wire [7:0] _T_4559; // @[Mux.scala 31:69:@20165.4]
  wire  _T_4528; // @[package.scala 96:25:@20093.4 package.scala 96:25:@20094.4]
  wire [7:0] _T_4560; // @[Mux.scala 31:69:@20166.4]
  wire  _T_4525; // @[package.scala 96:25:@20085.4 package.scala 96:25:@20086.4]
  wire [7:0] _T_4561; // @[Mux.scala 31:69:@20167.4]
  wire  _T_4522; // @[package.scala 96:25:@20077.4 package.scala 96:25:@20078.4]
  wire [7:0] _T_4562; // @[Mux.scala 31:69:@20168.4]
  wire  _T_4519; // @[package.scala 96:25:@20069.4 package.scala 96:25:@20070.4]
  wire  _T_4656; // @[package.scala 96:25:@20293.4 package.scala 96:25:@20294.4]
  wire [7:0] _T_4660; // @[Mux.scala 31:69:@20303.4]
  wire  _T_4653; // @[package.scala 96:25:@20285.4 package.scala 96:25:@20286.4]
  wire [7:0] _T_4661; // @[Mux.scala 31:69:@20304.4]
  wire  _T_4650; // @[package.scala 96:25:@20277.4 package.scala 96:25:@20278.4]
  wire [7:0] _T_4662; // @[Mux.scala 31:69:@20305.4]
  wire  _T_4647; // @[package.scala 96:25:@20269.4 package.scala 96:25:@20270.4]
  wire [7:0] _T_4663; // @[Mux.scala 31:69:@20306.4]
  wire  _T_4644; // @[package.scala 96:25:@20261.4 package.scala 96:25:@20262.4]
  wire [7:0] _T_4664; // @[Mux.scala 31:69:@20307.4]
  wire  _T_4641; // @[package.scala 96:25:@20253.4 package.scala 96:25:@20254.4]
  wire [7:0] _T_4665; // @[Mux.scala 31:69:@20308.4]
  wire  _T_4638; // @[package.scala 96:25:@20245.4 package.scala 96:25:@20246.4]
  wire [7:0] _T_4666; // @[Mux.scala 31:69:@20309.4]
  wire  _T_4635; // @[package.scala 96:25:@20237.4 package.scala 96:25:@20238.4]
  wire [7:0] _T_4667; // @[Mux.scala 31:69:@20310.4]
  wire  _T_4632; // @[package.scala 96:25:@20229.4 package.scala 96:25:@20230.4]
  wire [7:0] _T_4668; // @[Mux.scala 31:69:@20311.4]
  wire  _T_4629; // @[package.scala 96:25:@20221.4 package.scala 96:25:@20222.4]
  wire [7:0] _T_4669; // @[Mux.scala 31:69:@20312.4]
  wire  _T_4626; // @[package.scala 96:25:@20213.4 package.scala 96:25:@20214.4]
  wire  _T_4763; // @[package.scala 96:25:@20437.4 package.scala 96:25:@20438.4]
  wire [7:0] _T_4767; // @[Mux.scala 31:69:@20447.4]
  wire  _T_4760; // @[package.scala 96:25:@20429.4 package.scala 96:25:@20430.4]
  wire [7:0] _T_4768; // @[Mux.scala 31:69:@20448.4]
  wire  _T_4757; // @[package.scala 96:25:@20421.4 package.scala 96:25:@20422.4]
  wire [7:0] _T_4769; // @[Mux.scala 31:69:@20449.4]
  wire  _T_4754; // @[package.scala 96:25:@20413.4 package.scala 96:25:@20414.4]
  wire [7:0] _T_4770; // @[Mux.scala 31:69:@20450.4]
  wire  _T_4751; // @[package.scala 96:25:@20405.4 package.scala 96:25:@20406.4]
  wire [7:0] _T_4771; // @[Mux.scala 31:69:@20451.4]
  wire  _T_4748; // @[package.scala 96:25:@20397.4 package.scala 96:25:@20398.4]
  wire [7:0] _T_4772; // @[Mux.scala 31:69:@20452.4]
  wire  _T_4745; // @[package.scala 96:25:@20389.4 package.scala 96:25:@20390.4]
  wire [7:0] _T_4773; // @[Mux.scala 31:69:@20453.4]
  wire  _T_4742; // @[package.scala 96:25:@20381.4 package.scala 96:25:@20382.4]
  wire [7:0] _T_4774; // @[Mux.scala 31:69:@20454.4]
  wire  _T_4739; // @[package.scala 96:25:@20373.4 package.scala 96:25:@20374.4]
  wire [7:0] _T_4775; // @[Mux.scala 31:69:@20455.4]
  wire  _T_4736; // @[package.scala 96:25:@20365.4 package.scala 96:25:@20366.4]
  wire [7:0] _T_4776; // @[Mux.scala 31:69:@20456.4]
  wire  _T_4733; // @[package.scala 96:25:@20357.4 package.scala 96:25:@20358.4]
  wire  _T_4870; // @[package.scala 96:25:@20581.4 package.scala 96:25:@20582.4]
  wire [7:0] _T_4874; // @[Mux.scala 31:69:@20591.4]
  wire  _T_4867; // @[package.scala 96:25:@20573.4 package.scala 96:25:@20574.4]
  wire [7:0] _T_4875; // @[Mux.scala 31:69:@20592.4]
  wire  _T_4864; // @[package.scala 96:25:@20565.4 package.scala 96:25:@20566.4]
  wire [7:0] _T_4876; // @[Mux.scala 31:69:@20593.4]
  wire  _T_4861; // @[package.scala 96:25:@20557.4 package.scala 96:25:@20558.4]
  wire [7:0] _T_4877; // @[Mux.scala 31:69:@20594.4]
  wire  _T_4858; // @[package.scala 96:25:@20549.4 package.scala 96:25:@20550.4]
  wire [7:0] _T_4878; // @[Mux.scala 31:69:@20595.4]
  wire  _T_4855; // @[package.scala 96:25:@20541.4 package.scala 96:25:@20542.4]
  wire [7:0] _T_4879; // @[Mux.scala 31:69:@20596.4]
  wire  _T_4852; // @[package.scala 96:25:@20533.4 package.scala 96:25:@20534.4]
  wire [7:0] _T_4880; // @[Mux.scala 31:69:@20597.4]
  wire  _T_4849; // @[package.scala 96:25:@20525.4 package.scala 96:25:@20526.4]
  wire [7:0] _T_4881; // @[Mux.scala 31:69:@20598.4]
  wire  _T_4846; // @[package.scala 96:25:@20517.4 package.scala 96:25:@20518.4]
  wire [7:0] _T_4882; // @[Mux.scala 31:69:@20599.4]
  wire  _T_4843; // @[package.scala 96:25:@20509.4 package.scala 96:25:@20510.4]
  wire [7:0] _T_4883; // @[Mux.scala 31:69:@20600.4]
  wire  _T_4840; // @[package.scala 96:25:@20501.4 package.scala 96:25:@20502.4]
  wire  _T_4977; // @[package.scala 96:25:@20725.4 package.scala 96:25:@20726.4]
  wire [7:0] _T_4981; // @[Mux.scala 31:69:@20735.4]
  wire  _T_4974; // @[package.scala 96:25:@20717.4 package.scala 96:25:@20718.4]
  wire [7:0] _T_4982; // @[Mux.scala 31:69:@20736.4]
  wire  _T_4971; // @[package.scala 96:25:@20709.4 package.scala 96:25:@20710.4]
  wire [7:0] _T_4983; // @[Mux.scala 31:69:@20737.4]
  wire  _T_4968; // @[package.scala 96:25:@20701.4 package.scala 96:25:@20702.4]
  wire [7:0] _T_4984; // @[Mux.scala 31:69:@20738.4]
  wire  _T_4965; // @[package.scala 96:25:@20693.4 package.scala 96:25:@20694.4]
  wire [7:0] _T_4985; // @[Mux.scala 31:69:@20739.4]
  wire  _T_4962; // @[package.scala 96:25:@20685.4 package.scala 96:25:@20686.4]
  wire [7:0] _T_4986; // @[Mux.scala 31:69:@20740.4]
  wire  _T_4959; // @[package.scala 96:25:@20677.4 package.scala 96:25:@20678.4]
  wire [7:0] _T_4987; // @[Mux.scala 31:69:@20741.4]
  wire  _T_4956; // @[package.scala 96:25:@20669.4 package.scala 96:25:@20670.4]
  wire [7:0] _T_4988; // @[Mux.scala 31:69:@20742.4]
  wire  _T_4953; // @[package.scala 96:25:@20661.4 package.scala 96:25:@20662.4]
  wire [7:0] _T_4989; // @[Mux.scala 31:69:@20743.4]
  wire  _T_4950; // @[package.scala 96:25:@20653.4 package.scala 96:25:@20654.4]
  wire [7:0] _T_4990; // @[Mux.scala 31:69:@20744.4]
  wire  _T_4947; // @[package.scala 96:25:@20645.4 package.scala 96:25:@20646.4]
  wire  _T_5084; // @[package.scala 96:25:@20869.4 package.scala 96:25:@20870.4]
  wire [7:0] _T_5088; // @[Mux.scala 31:69:@20879.4]
  wire  _T_5081; // @[package.scala 96:25:@20861.4 package.scala 96:25:@20862.4]
  wire [7:0] _T_5089; // @[Mux.scala 31:69:@20880.4]
  wire  _T_5078; // @[package.scala 96:25:@20853.4 package.scala 96:25:@20854.4]
  wire [7:0] _T_5090; // @[Mux.scala 31:69:@20881.4]
  wire  _T_5075; // @[package.scala 96:25:@20845.4 package.scala 96:25:@20846.4]
  wire [7:0] _T_5091; // @[Mux.scala 31:69:@20882.4]
  wire  _T_5072; // @[package.scala 96:25:@20837.4 package.scala 96:25:@20838.4]
  wire [7:0] _T_5092; // @[Mux.scala 31:69:@20883.4]
  wire  _T_5069; // @[package.scala 96:25:@20829.4 package.scala 96:25:@20830.4]
  wire [7:0] _T_5093; // @[Mux.scala 31:69:@20884.4]
  wire  _T_5066; // @[package.scala 96:25:@20821.4 package.scala 96:25:@20822.4]
  wire [7:0] _T_5094; // @[Mux.scala 31:69:@20885.4]
  wire  _T_5063; // @[package.scala 96:25:@20813.4 package.scala 96:25:@20814.4]
  wire [7:0] _T_5095; // @[Mux.scala 31:69:@20886.4]
  wire  _T_5060; // @[package.scala 96:25:@20805.4 package.scala 96:25:@20806.4]
  wire [7:0] _T_5096; // @[Mux.scala 31:69:@20887.4]
  wire  _T_5057; // @[package.scala 96:25:@20797.4 package.scala 96:25:@20798.4]
  wire [7:0] _T_5097; // @[Mux.scala 31:69:@20888.4]
  wire  _T_5054; // @[package.scala 96:25:@20789.4 package.scala 96:25:@20790.4]
  wire  _T_5191; // @[package.scala 96:25:@21013.4 package.scala 96:25:@21014.4]
  wire [7:0] _T_5195; // @[Mux.scala 31:69:@21023.4]
  wire  _T_5188; // @[package.scala 96:25:@21005.4 package.scala 96:25:@21006.4]
  wire [7:0] _T_5196; // @[Mux.scala 31:69:@21024.4]
  wire  _T_5185; // @[package.scala 96:25:@20997.4 package.scala 96:25:@20998.4]
  wire [7:0] _T_5197; // @[Mux.scala 31:69:@21025.4]
  wire  _T_5182; // @[package.scala 96:25:@20989.4 package.scala 96:25:@20990.4]
  wire [7:0] _T_5198; // @[Mux.scala 31:69:@21026.4]
  wire  _T_5179; // @[package.scala 96:25:@20981.4 package.scala 96:25:@20982.4]
  wire [7:0] _T_5199; // @[Mux.scala 31:69:@21027.4]
  wire  _T_5176; // @[package.scala 96:25:@20973.4 package.scala 96:25:@20974.4]
  wire [7:0] _T_5200; // @[Mux.scala 31:69:@21028.4]
  wire  _T_5173; // @[package.scala 96:25:@20965.4 package.scala 96:25:@20966.4]
  wire [7:0] _T_5201; // @[Mux.scala 31:69:@21029.4]
  wire  _T_5170; // @[package.scala 96:25:@20957.4 package.scala 96:25:@20958.4]
  wire [7:0] _T_5202; // @[Mux.scala 31:69:@21030.4]
  wire  _T_5167; // @[package.scala 96:25:@20949.4 package.scala 96:25:@20950.4]
  wire [7:0] _T_5203; // @[Mux.scala 31:69:@21031.4]
  wire  _T_5164; // @[package.scala 96:25:@20941.4 package.scala 96:25:@20942.4]
  wire [7:0] _T_5204; // @[Mux.scala 31:69:@21032.4]
  wire  _T_5161; // @[package.scala 96:25:@20933.4 package.scala 96:25:@20934.4]
  wire  _T_5298; // @[package.scala 96:25:@21157.4 package.scala 96:25:@21158.4]
  wire [7:0] _T_5302; // @[Mux.scala 31:69:@21167.4]
  wire  _T_5295; // @[package.scala 96:25:@21149.4 package.scala 96:25:@21150.4]
  wire [7:0] _T_5303; // @[Mux.scala 31:69:@21168.4]
  wire  _T_5292; // @[package.scala 96:25:@21141.4 package.scala 96:25:@21142.4]
  wire [7:0] _T_5304; // @[Mux.scala 31:69:@21169.4]
  wire  _T_5289; // @[package.scala 96:25:@21133.4 package.scala 96:25:@21134.4]
  wire [7:0] _T_5305; // @[Mux.scala 31:69:@21170.4]
  wire  _T_5286; // @[package.scala 96:25:@21125.4 package.scala 96:25:@21126.4]
  wire [7:0] _T_5306; // @[Mux.scala 31:69:@21171.4]
  wire  _T_5283; // @[package.scala 96:25:@21117.4 package.scala 96:25:@21118.4]
  wire [7:0] _T_5307; // @[Mux.scala 31:69:@21172.4]
  wire  _T_5280; // @[package.scala 96:25:@21109.4 package.scala 96:25:@21110.4]
  wire [7:0] _T_5308; // @[Mux.scala 31:69:@21173.4]
  wire  _T_5277; // @[package.scala 96:25:@21101.4 package.scala 96:25:@21102.4]
  wire [7:0] _T_5309; // @[Mux.scala 31:69:@21174.4]
  wire  _T_5274; // @[package.scala 96:25:@21093.4 package.scala 96:25:@21094.4]
  wire [7:0] _T_5310; // @[Mux.scala 31:69:@21175.4]
  wire  _T_5271; // @[package.scala 96:25:@21085.4 package.scala 96:25:@21086.4]
  wire [7:0] _T_5311; // @[Mux.scala 31:69:@21176.4]
  wire  _T_5268; // @[package.scala 96:25:@21077.4 package.scala 96:25:@21078.4]
  Mem1D_4 Mem1D ( // @[MemPrimitives.scala 64:21:@15611.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  Mem1D_4 Mem1D_1 ( // @[MemPrimitives.scala 64:21:@15627.4]
    .clock(Mem1D_1_clock),
    .reset(Mem1D_1_reset),
    .io_r_ofs_0(Mem1D_1_io_r_ofs_0),
    .io_r_backpressure(Mem1D_1_io_r_backpressure),
    .io_w_ofs_0(Mem1D_1_io_w_ofs_0),
    .io_w_data_0(Mem1D_1_io_w_data_0),
    .io_w_en_0(Mem1D_1_io_w_en_0),
    .io_output(Mem1D_1_io_output)
  );
  Mem1D_4 Mem1D_2 ( // @[MemPrimitives.scala 64:21:@15643.4]
    .clock(Mem1D_2_clock),
    .reset(Mem1D_2_reset),
    .io_r_ofs_0(Mem1D_2_io_r_ofs_0),
    .io_r_backpressure(Mem1D_2_io_r_backpressure),
    .io_w_ofs_0(Mem1D_2_io_w_ofs_0),
    .io_w_data_0(Mem1D_2_io_w_data_0),
    .io_w_en_0(Mem1D_2_io_w_en_0),
    .io_output(Mem1D_2_io_output)
  );
  Mem1D_4 Mem1D_3 ( // @[MemPrimitives.scala 64:21:@15659.4]
    .clock(Mem1D_3_clock),
    .reset(Mem1D_3_reset),
    .io_r_ofs_0(Mem1D_3_io_r_ofs_0),
    .io_r_backpressure(Mem1D_3_io_r_backpressure),
    .io_w_ofs_0(Mem1D_3_io_w_ofs_0),
    .io_w_data_0(Mem1D_3_io_w_data_0),
    .io_w_en_0(Mem1D_3_io_w_en_0),
    .io_output(Mem1D_3_io_output)
  );
  Mem1D_4 Mem1D_4 ( // @[MemPrimitives.scala 64:21:@15675.4]
    .clock(Mem1D_4_clock),
    .reset(Mem1D_4_reset),
    .io_r_ofs_0(Mem1D_4_io_r_ofs_0),
    .io_r_backpressure(Mem1D_4_io_r_backpressure),
    .io_w_ofs_0(Mem1D_4_io_w_ofs_0),
    .io_w_data_0(Mem1D_4_io_w_data_0),
    .io_w_en_0(Mem1D_4_io_w_en_0),
    .io_output(Mem1D_4_io_output)
  );
  Mem1D_4 Mem1D_5 ( // @[MemPrimitives.scala 64:21:@15691.4]
    .clock(Mem1D_5_clock),
    .reset(Mem1D_5_reset),
    .io_r_ofs_0(Mem1D_5_io_r_ofs_0),
    .io_r_backpressure(Mem1D_5_io_r_backpressure),
    .io_w_ofs_0(Mem1D_5_io_w_ofs_0),
    .io_w_data_0(Mem1D_5_io_w_data_0),
    .io_w_en_0(Mem1D_5_io_w_en_0),
    .io_output(Mem1D_5_io_output)
  );
  Mem1D_4 Mem1D_6 ( // @[MemPrimitives.scala 64:21:@15707.4]
    .clock(Mem1D_6_clock),
    .reset(Mem1D_6_reset),
    .io_r_ofs_0(Mem1D_6_io_r_ofs_0),
    .io_r_backpressure(Mem1D_6_io_r_backpressure),
    .io_w_ofs_0(Mem1D_6_io_w_ofs_0),
    .io_w_data_0(Mem1D_6_io_w_data_0),
    .io_w_en_0(Mem1D_6_io_w_en_0),
    .io_output(Mem1D_6_io_output)
  );
  Mem1D_4 Mem1D_7 ( // @[MemPrimitives.scala 64:21:@15723.4]
    .clock(Mem1D_7_clock),
    .reset(Mem1D_7_reset),
    .io_r_ofs_0(Mem1D_7_io_r_ofs_0),
    .io_r_backpressure(Mem1D_7_io_r_backpressure),
    .io_w_ofs_0(Mem1D_7_io_w_ofs_0),
    .io_w_data_0(Mem1D_7_io_w_data_0),
    .io_w_en_0(Mem1D_7_io_w_en_0),
    .io_output(Mem1D_7_io_output)
  );
  Mem1D_4 Mem1D_8 ( // @[MemPrimitives.scala 64:21:@15739.4]
    .clock(Mem1D_8_clock),
    .reset(Mem1D_8_reset),
    .io_r_ofs_0(Mem1D_8_io_r_ofs_0),
    .io_r_backpressure(Mem1D_8_io_r_backpressure),
    .io_w_ofs_0(Mem1D_8_io_w_ofs_0),
    .io_w_data_0(Mem1D_8_io_w_data_0),
    .io_w_en_0(Mem1D_8_io_w_en_0),
    .io_output(Mem1D_8_io_output)
  );
  Mem1D_4 Mem1D_9 ( // @[MemPrimitives.scala 64:21:@15755.4]
    .clock(Mem1D_9_clock),
    .reset(Mem1D_9_reset),
    .io_r_ofs_0(Mem1D_9_io_r_ofs_0),
    .io_r_backpressure(Mem1D_9_io_r_backpressure),
    .io_w_ofs_0(Mem1D_9_io_w_ofs_0),
    .io_w_data_0(Mem1D_9_io_w_data_0),
    .io_w_en_0(Mem1D_9_io_w_en_0),
    .io_output(Mem1D_9_io_output)
  );
  Mem1D_4 Mem1D_10 ( // @[MemPrimitives.scala 64:21:@15771.4]
    .clock(Mem1D_10_clock),
    .reset(Mem1D_10_reset),
    .io_r_ofs_0(Mem1D_10_io_r_ofs_0),
    .io_r_backpressure(Mem1D_10_io_r_backpressure),
    .io_w_ofs_0(Mem1D_10_io_w_ofs_0),
    .io_w_data_0(Mem1D_10_io_w_data_0),
    .io_w_en_0(Mem1D_10_io_w_en_0),
    .io_output(Mem1D_10_io_output)
  );
  Mem1D_4 Mem1D_11 ( // @[MemPrimitives.scala 64:21:@15787.4]
    .clock(Mem1D_11_clock),
    .reset(Mem1D_11_reset),
    .io_r_ofs_0(Mem1D_11_io_r_ofs_0),
    .io_r_backpressure(Mem1D_11_io_r_backpressure),
    .io_w_ofs_0(Mem1D_11_io_w_ofs_0),
    .io_w_data_0(Mem1D_11_io_w_data_0),
    .io_w_en_0(Mem1D_11_io_w_en_0),
    .io_output(Mem1D_11_io_output)
  );
  Mem1D_4 Mem1D_12 ( // @[MemPrimitives.scala 64:21:@15803.4]
    .clock(Mem1D_12_clock),
    .reset(Mem1D_12_reset),
    .io_r_ofs_0(Mem1D_12_io_r_ofs_0),
    .io_r_backpressure(Mem1D_12_io_r_backpressure),
    .io_w_ofs_0(Mem1D_12_io_w_ofs_0),
    .io_w_data_0(Mem1D_12_io_w_data_0),
    .io_w_en_0(Mem1D_12_io_w_en_0),
    .io_output(Mem1D_12_io_output)
  );
  Mem1D_4 Mem1D_13 ( // @[MemPrimitives.scala 64:21:@15819.4]
    .clock(Mem1D_13_clock),
    .reset(Mem1D_13_reset),
    .io_r_ofs_0(Mem1D_13_io_r_ofs_0),
    .io_r_backpressure(Mem1D_13_io_r_backpressure),
    .io_w_ofs_0(Mem1D_13_io_w_ofs_0),
    .io_w_data_0(Mem1D_13_io_w_data_0),
    .io_w_en_0(Mem1D_13_io_w_en_0),
    .io_output(Mem1D_13_io_output)
  );
  Mem1D_4 Mem1D_14 ( // @[MemPrimitives.scala 64:21:@15835.4]
    .clock(Mem1D_14_clock),
    .reset(Mem1D_14_reset),
    .io_r_ofs_0(Mem1D_14_io_r_ofs_0),
    .io_r_backpressure(Mem1D_14_io_r_backpressure),
    .io_w_ofs_0(Mem1D_14_io_w_ofs_0),
    .io_w_data_0(Mem1D_14_io_w_data_0),
    .io_w_en_0(Mem1D_14_io_w_en_0),
    .io_output(Mem1D_14_io_output)
  );
  Mem1D_4 Mem1D_15 ( // @[MemPrimitives.scala 64:21:@15851.4]
    .clock(Mem1D_15_clock),
    .reset(Mem1D_15_reset),
    .io_r_ofs_0(Mem1D_15_io_r_ofs_0),
    .io_r_backpressure(Mem1D_15_io_r_backpressure),
    .io_w_ofs_0(Mem1D_15_io_w_ofs_0),
    .io_w_data_0(Mem1D_15_io_w_data_0),
    .io_w_en_0(Mem1D_15_io_w_en_0),
    .io_output(Mem1D_15_io_output)
  );
  Mem1D_4 Mem1D_16 ( // @[MemPrimitives.scala 64:21:@15867.4]
    .clock(Mem1D_16_clock),
    .reset(Mem1D_16_reset),
    .io_r_ofs_0(Mem1D_16_io_r_ofs_0),
    .io_r_backpressure(Mem1D_16_io_r_backpressure),
    .io_w_ofs_0(Mem1D_16_io_w_ofs_0),
    .io_w_data_0(Mem1D_16_io_w_data_0),
    .io_w_en_0(Mem1D_16_io_w_en_0),
    .io_output(Mem1D_16_io_output)
  );
  Mem1D_4 Mem1D_17 ( // @[MemPrimitives.scala 64:21:@15883.4]
    .clock(Mem1D_17_clock),
    .reset(Mem1D_17_reset),
    .io_r_ofs_0(Mem1D_17_io_r_ofs_0),
    .io_r_backpressure(Mem1D_17_io_r_backpressure),
    .io_w_ofs_0(Mem1D_17_io_w_ofs_0),
    .io_w_data_0(Mem1D_17_io_w_data_0),
    .io_w_en_0(Mem1D_17_io_w_en_0),
    .io_output(Mem1D_17_io_output)
  );
  Mem1D_4 Mem1D_18 ( // @[MemPrimitives.scala 64:21:@15899.4]
    .clock(Mem1D_18_clock),
    .reset(Mem1D_18_reset),
    .io_r_ofs_0(Mem1D_18_io_r_ofs_0),
    .io_r_backpressure(Mem1D_18_io_r_backpressure),
    .io_w_ofs_0(Mem1D_18_io_w_ofs_0),
    .io_w_data_0(Mem1D_18_io_w_data_0),
    .io_w_en_0(Mem1D_18_io_w_en_0),
    .io_output(Mem1D_18_io_output)
  );
  Mem1D_4 Mem1D_19 ( // @[MemPrimitives.scala 64:21:@15915.4]
    .clock(Mem1D_19_clock),
    .reset(Mem1D_19_reset),
    .io_r_ofs_0(Mem1D_19_io_r_ofs_0),
    .io_r_backpressure(Mem1D_19_io_r_backpressure),
    .io_w_ofs_0(Mem1D_19_io_w_ofs_0),
    .io_w_data_0(Mem1D_19_io_w_data_0),
    .io_w_en_0(Mem1D_19_io_w_en_0),
    .io_output(Mem1D_19_io_output)
  );
  Mem1D_4 Mem1D_20 ( // @[MemPrimitives.scala 64:21:@15931.4]
    .clock(Mem1D_20_clock),
    .reset(Mem1D_20_reset),
    .io_r_ofs_0(Mem1D_20_io_r_ofs_0),
    .io_r_backpressure(Mem1D_20_io_r_backpressure),
    .io_w_ofs_0(Mem1D_20_io_w_ofs_0),
    .io_w_data_0(Mem1D_20_io_w_data_0),
    .io_w_en_0(Mem1D_20_io_w_en_0),
    .io_output(Mem1D_20_io_output)
  );
  Mem1D_4 Mem1D_21 ( // @[MemPrimitives.scala 64:21:@15947.4]
    .clock(Mem1D_21_clock),
    .reset(Mem1D_21_reset),
    .io_r_ofs_0(Mem1D_21_io_r_ofs_0),
    .io_r_backpressure(Mem1D_21_io_r_backpressure),
    .io_w_ofs_0(Mem1D_21_io_w_ofs_0),
    .io_w_data_0(Mem1D_21_io_w_data_0),
    .io_w_en_0(Mem1D_21_io_w_en_0),
    .io_output(Mem1D_21_io_output)
  );
  Mem1D_4 Mem1D_22 ( // @[MemPrimitives.scala 64:21:@15963.4]
    .clock(Mem1D_22_clock),
    .reset(Mem1D_22_reset),
    .io_r_ofs_0(Mem1D_22_io_r_ofs_0),
    .io_r_backpressure(Mem1D_22_io_r_backpressure),
    .io_w_ofs_0(Mem1D_22_io_w_ofs_0),
    .io_w_data_0(Mem1D_22_io_w_data_0),
    .io_w_en_0(Mem1D_22_io_w_en_0),
    .io_output(Mem1D_22_io_output)
  );
  Mem1D_4 Mem1D_23 ( // @[MemPrimitives.scala 64:21:@15979.4]
    .clock(Mem1D_23_clock),
    .reset(Mem1D_23_reset),
    .io_r_ofs_0(Mem1D_23_io_r_ofs_0),
    .io_r_backpressure(Mem1D_23_io_r_backpressure),
    .io_w_ofs_0(Mem1D_23_io_w_ofs_0),
    .io_w_data_0(Mem1D_23_io_w_data_0),
    .io_w_en_0(Mem1D_23_io_w_en_0),
    .io_output(Mem1D_23_io_output)
  );
  StickySelects StickySelects ( // @[MemPrimitives.scala 121:29:@16487.4]
    .clock(StickySelects_clock),
    .reset(StickySelects_reset),
    .io_ins_0(StickySelects_io_ins_0),
    .io_ins_1(StickySelects_io_ins_1),
    .io_ins_2(StickySelects_io_ins_2),
    .io_ins_3(StickySelects_io_ins_3),
    .io_ins_4(StickySelects_io_ins_4),
    .io_ins_5(StickySelects_io_ins_5),
    .io_ins_6(StickySelects_io_ins_6),
    .io_ins_7(StickySelects_io_ins_7),
    .io_ins_8(StickySelects_io_ins_8),
    .io_outs_0(StickySelects_io_outs_0),
    .io_outs_1(StickySelects_io_outs_1),
    .io_outs_2(StickySelects_io_outs_2),
    .io_outs_3(StickySelects_io_outs_3),
    .io_outs_4(StickySelects_io_outs_4),
    .io_outs_5(StickySelects_io_outs_5),
    .io_outs_6(StickySelects_io_outs_6),
    .io_outs_7(StickySelects_io_outs_7),
    .io_outs_8(StickySelects_io_outs_8)
  );
  StickySelects StickySelects_1 ( // @[MemPrimitives.scala 121:29:@16576.4]
    .clock(StickySelects_1_clock),
    .reset(StickySelects_1_reset),
    .io_ins_0(StickySelects_1_io_ins_0),
    .io_ins_1(StickySelects_1_io_ins_1),
    .io_ins_2(StickySelects_1_io_ins_2),
    .io_ins_3(StickySelects_1_io_ins_3),
    .io_ins_4(StickySelects_1_io_ins_4),
    .io_ins_5(StickySelects_1_io_ins_5),
    .io_ins_6(StickySelects_1_io_ins_6),
    .io_ins_7(StickySelects_1_io_ins_7),
    .io_ins_8(StickySelects_1_io_ins_8),
    .io_outs_0(StickySelects_1_io_outs_0),
    .io_outs_1(StickySelects_1_io_outs_1),
    .io_outs_2(StickySelects_1_io_outs_2),
    .io_outs_3(StickySelects_1_io_outs_3),
    .io_outs_4(StickySelects_1_io_outs_4),
    .io_outs_5(StickySelects_1_io_outs_5),
    .io_outs_6(StickySelects_1_io_outs_6),
    .io_outs_7(StickySelects_1_io_outs_7),
    .io_outs_8(StickySelects_1_io_outs_8)
  );
  StickySelects StickySelects_2 ( // @[MemPrimitives.scala 121:29:@16665.4]
    .clock(StickySelects_2_clock),
    .reset(StickySelects_2_reset),
    .io_ins_0(StickySelects_2_io_ins_0),
    .io_ins_1(StickySelects_2_io_ins_1),
    .io_ins_2(StickySelects_2_io_ins_2),
    .io_ins_3(StickySelects_2_io_ins_3),
    .io_ins_4(StickySelects_2_io_ins_4),
    .io_ins_5(StickySelects_2_io_ins_5),
    .io_ins_6(StickySelects_2_io_ins_6),
    .io_ins_7(StickySelects_2_io_ins_7),
    .io_ins_8(StickySelects_2_io_ins_8),
    .io_outs_0(StickySelects_2_io_outs_0),
    .io_outs_1(StickySelects_2_io_outs_1),
    .io_outs_2(StickySelects_2_io_outs_2),
    .io_outs_3(StickySelects_2_io_outs_3),
    .io_outs_4(StickySelects_2_io_outs_4),
    .io_outs_5(StickySelects_2_io_outs_5),
    .io_outs_6(StickySelects_2_io_outs_6),
    .io_outs_7(StickySelects_2_io_outs_7),
    .io_outs_8(StickySelects_2_io_outs_8)
  );
  StickySelects StickySelects_3 ( // @[MemPrimitives.scala 121:29:@16754.4]
    .clock(StickySelects_3_clock),
    .reset(StickySelects_3_reset),
    .io_ins_0(StickySelects_3_io_ins_0),
    .io_ins_1(StickySelects_3_io_ins_1),
    .io_ins_2(StickySelects_3_io_ins_2),
    .io_ins_3(StickySelects_3_io_ins_3),
    .io_ins_4(StickySelects_3_io_ins_4),
    .io_ins_5(StickySelects_3_io_ins_5),
    .io_ins_6(StickySelects_3_io_ins_6),
    .io_ins_7(StickySelects_3_io_ins_7),
    .io_ins_8(StickySelects_3_io_ins_8),
    .io_outs_0(StickySelects_3_io_outs_0),
    .io_outs_1(StickySelects_3_io_outs_1),
    .io_outs_2(StickySelects_3_io_outs_2),
    .io_outs_3(StickySelects_3_io_outs_3),
    .io_outs_4(StickySelects_3_io_outs_4),
    .io_outs_5(StickySelects_3_io_outs_5),
    .io_outs_6(StickySelects_3_io_outs_6),
    .io_outs_7(StickySelects_3_io_outs_7),
    .io_outs_8(StickySelects_3_io_outs_8)
  );
  StickySelects StickySelects_4 ( // @[MemPrimitives.scala 121:29:@16843.4]
    .clock(StickySelects_4_clock),
    .reset(StickySelects_4_reset),
    .io_ins_0(StickySelects_4_io_ins_0),
    .io_ins_1(StickySelects_4_io_ins_1),
    .io_ins_2(StickySelects_4_io_ins_2),
    .io_ins_3(StickySelects_4_io_ins_3),
    .io_ins_4(StickySelects_4_io_ins_4),
    .io_ins_5(StickySelects_4_io_ins_5),
    .io_ins_6(StickySelects_4_io_ins_6),
    .io_ins_7(StickySelects_4_io_ins_7),
    .io_ins_8(StickySelects_4_io_ins_8),
    .io_outs_0(StickySelects_4_io_outs_0),
    .io_outs_1(StickySelects_4_io_outs_1),
    .io_outs_2(StickySelects_4_io_outs_2),
    .io_outs_3(StickySelects_4_io_outs_3),
    .io_outs_4(StickySelects_4_io_outs_4),
    .io_outs_5(StickySelects_4_io_outs_5),
    .io_outs_6(StickySelects_4_io_outs_6),
    .io_outs_7(StickySelects_4_io_outs_7),
    .io_outs_8(StickySelects_4_io_outs_8)
  );
  StickySelects StickySelects_5 ( // @[MemPrimitives.scala 121:29:@16932.4]
    .clock(StickySelects_5_clock),
    .reset(StickySelects_5_reset),
    .io_ins_0(StickySelects_5_io_ins_0),
    .io_ins_1(StickySelects_5_io_ins_1),
    .io_ins_2(StickySelects_5_io_ins_2),
    .io_ins_3(StickySelects_5_io_ins_3),
    .io_ins_4(StickySelects_5_io_ins_4),
    .io_ins_5(StickySelects_5_io_ins_5),
    .io_ins_6(StickySelects_5_io_ins_6),
    .io_ins_7(StickySelects_5_io_ins_7),
    .io_ins_8(StickySelects_5_io_ins_8),
    .io_outs_0(StickySelects_5_io_outs_0),
    .io_outs_1(StickySelects_5_io_outs_1),
    .io_outs_2(StickySelects_5_io_outs_2),
    .io_outs_3(StickySelects_5_io_outs_3),
    .io_outs_4(StickySelects_5_io_outs_4),
    .io_outs_5(StickySelects_5_io_outs_5),
    .io_outs_6(StickySelects_5_io_outs_6),
    .io_outs_7(StickySelects_5_io_outs_7),
    .io_outs_8(StickySelects_5_io_outs_8)
  );
  StickySelects StickySelects_6 ( // @[MemPrimitives.scala 121:29:@17021.4]
    .clock(StickySelects_6_clock),
    .reset(StickySelects_6_reset),
    .io_ins_0(StickySelects_6_io_ins_0),
    .io_ins_1(StickySelects_6_io_ins_1),
    .io_ins_2(StickySelects_6_io_ins_2),
    .io_ins_3(StickySelects_6_io_ins_3),
    .io_ins_4(StickySelects_6_io_ins_4),
    .io_ins_5(StickySelects_6_io_ins_5),
    .io_ins_6(StickySelects_6_io_ins_6),
    .io_ins_7(StickySelects_6_io_ins_7),
    .io_ins_8(StickySelects_6_io_ins_8),
    .io_outs_0(StickySelects_6_io_outs_0),
    .io_outs_1(StickySelects_6_io_outs_1),
    .io_outs_2(StickySelects_6_io_outs_2),
    .io_outs_3(StickySelects_6_io_outs_3),
    .io_outs_4(StickySelects_6_io_outs_4),
    .io_outs_5(StickySelects_6_io_outs_5),
    .io_outs_6(StickySelects_6_io_outs_6),
    .io_outs_7(StickySelects_6_io_outs_7),
    .io_outs_8(StickySelects_6_io_outs_8)
  );
  StickySelects StickySelects_7 ( // @[MemPrimitives.scala 121:29:@17110.4]
    .clock(StickySelects_7_clock),
    .reset(StickySelects_7_reset),
    .io_ins_0(StickySelects_7_io_ins_0),
    .io_ins_1(StickySelects_7_io_ins_1),
    .io_ins_2(StickySelects_7_io_ins_2),
    .io_ins_3(StickySelects_7_io_ins_3),
    .io_ins_4(StickySelects_7_io_ins_4),
    .io_ins_5(StickySelects_7_io_ins_5),
    .io_ins_6(StickySelects_7_io_ins_6),
    .io_ins_7(StickySelects_7_io_ins_7),
    .io_ins_8(StickySelects_7_io_ins_8),
    .io_outs_0(StickySelects_7_io_outs_0),
    .io_outs_1(StickySelects_7_io_outs_1),
    .io_outs_2(StickySelects_7_io_outs_2),
    .io_outs_3(StickySelects_7_io_outs_3),
    .io_outs_4(StickySelects_7_io_outs_4),
    .io_outs_5(StickySelects_7_io_outs_5),
    .io_outs_6(StickySelects_7_io_outs_6),
    .io_outs_7(StickySelects_7_io_outs_7),
    .io_outs_8(StickySelects_7_io_outs_8)
  );
  StickySelects StickySelects_8 ( // @[MemPrimitives.scala 121:29:@17199.4]
    .clock(StickySelects_8_clock),
    .reset(StickySelects_8_reset),
    .io_ins_0(StickySelects_8_io_ins_0),
    .io_ins_1(StickySelects_8_io_ins_1),
    .io_ins_2(StickySelects_8_io_ins_2),
    .io_ins_3(StickySelects_8_io_ins_3),
    .io_ins_4(StickySelects_8_io_ins_4),
    .io_ins_5(StickySelects_8_io_ins_5),
    .io_ins_6(StickySelects_8_io_ins_6),
    .io_ins_7(StickySelects_8_io_ins_7),
    .io_ins_8(StickySelects_8_io_ins_8),
    .io_outs_0(StickySelects_8_io_outs_0),
    .io_outs_1(StickySelects_8_io_outs_1),
    .io_outs_2(StickySelects_8_io_outs_2),
    .io_outs_3(StickySelects_8_io_outs_3),
    .io_outs_4(StickySelects_8_io_outs_4),
    .io_outs_5(StickySelects_8_io_outs_5),
    .io_outs_6(StickySelects_8_io_outs_6),
    .io_outs_7(StickySelects_8_io_outs_7),
    .io_outs_8(StickySelects_8_io_outs_8)
  );
  StickySelects StickySelects_9 ( // @[MemPrimitives.scala 121:29:@17288.4]
    .clock(StickySelects_9_clock),
    .reset(StickySelects_9_reset),
    .io_ins_0(StickySelects_9_io_ins_0),
    .io_ins_1(StickySelects_9_io_ins_1),
    .io_ins_2(StickySelects_9_io_ins_2),
    .io_ins_3(StickySelects_9_io_ins_3),
    .io_ins_4(StickySelects_9_io_ins_4),
    .io_ins_5(StickySelects_9_io_ins_5),
    .io_ins_6(StickySelects_9_io_ins_6),
    .io_ins_7(StickySelects_9_io_ins_7),
    .io_ins_8(StickySelects_9_io_ins_8),
    .io_outs_0(StickySelects_9_io_outs_0),
    .io_outs_1(StickySelects_9_io_outs_1),
    .io_outs_2(StickySelects_9_io_outs_2),
    .io_outs_3(StickySelects_9_io_outs_3),
    .io_outs_4(StickySelects_9_io_outs_4),
    .io_outs_5(StickySelects_9_io_outs_5),
    .io_outs_6(StickySelects_9_io_outs_6),
    .io_outs_7(StickySelects_9_io_outs_7),
    .io_outs_8(StickySelects_9_io_outs_8)
  );
  StickySelects StickySelects_10 ( // @[MemPrimitives.scala 121:29:@17377.4]
    .clock(StickySelects_10_clock),
    .reset(StickySelects_10_reset),
    .io_ins_0(StickySelects_10_io_ins_0),
    .io_ins_1(StickySelects_10_io_ins_1),
    .io_ins_2(StickySelects_10_io_ins_2),
    .io_ins_3(StickySelects_10_io_ins_3),
    .io_ins_4(StickySelects_10_io_ins_4),
    .io_ins_5(StickySelects_10_io_ins_5),
    .io_ins_6(StickySelects_10_io_ins_6),
    .io_ins_7(StickySelects_10_io_ins_7),
    .io_ins_8(StickySelects_10_io_ins_8),
    .io_outs_0(StickySelects_10_io_outs_0),
    .io_outs_1(StickySelects_10_io_outs_1),
    .io_outs_2(StickySelects_10_io_outs_2),
    .io_outs_3(StickySelects_10_io_outs_3),
    .io_outs_4(StickySelects_10_io_outs_4),
    .io_outs_5(StickySelects_10_io_outs_5),
    .io_outs_6(StickySelects_10_io_outs_6),
    .io_outs_7(StickySelects_10_io_outs_7),
    .io_outs_8(StickySelects_10_io_outs_8)
  );
  StickySelects StickySelects_11 ( // @[MemPrimitives.scala 121:29:@17466.4]
    .clock(StickySelects_11_clock),
    .reset(StickySelects_11_reset),
    .io_ins_0(StickySelects_11_io_ins_0),
    .io_ins_1(StickySelects_11_io_ins_1),
    .io_ins_2(StickySelects_11_io_ins_2),
    .io_ins_3(StickySelects_11_io_ins_3),
    .io_ins_4(StickySelects_11_io_ins_4),
    .io_ins_5(StickySelects_11_io_ins_5),
    .io_ins_6(StickySelects_11_io_ins_6),
    .io_ins_7(StickySelects_11_io_ins_7),
    .io_ins_8(StickySelects_11_io_ins_8),
    .io_outs_0(StickySelects_11_io_outs_0),
    .io_outs_1(StickySelects_11_io_outs_1),
    .io_outs_2(StickySelects_11_io_outs_2),
    .io_outs_3(StickySelects_11_io_outs_3),
    .io_outs_4(StickySelects_11_io_outs_4),
    .io_outs_5(StickySelects_11_io_outs_5),
    .io_outs_6(StickySelects_11_io_outs_6),
    .io_outs_7(StickySelects_11_io_outs_7),
    .io_outs_8(StickySelects_11_io_outs_8)
  );
  StickySelects StickySelects_12 ( // @[MemPrimitives.scala 121:29:@17555.4]
    .clock(StickySelects_12_clock),
    .reset(StickySelects_12_reset),
    .io_ins_0(StickySelects_12_io_ins_0),
    .io_ins_1(StickySelects_12_io_ins_1),
    .io_ins_2(StickySelects_12_io_ins_2),
    .io_ins_3(StickySelects_12_io_ins_3),
    .io_ins_4(StickySelects_12_io_ins_4),
    .io_ins_5(StickySelects_12_io_ins_5),
    .io_ins_6(StickySelects_12_io_ins_6),
    .io_ins_7(StickySelects_12_io_ins_7),
    .io_ins_8(StickySelects_12_io_ins_8),
    .io_outs_0(StickySelects_12_io_outs_0),
    .io_outs_1(StickySelects_12_io_outs_1),
    .io_outs_2(StickySelects_12_io_outs_2),
    .io_outs_3(StickySelects_12_io_outs_3),
    .io_outs_4(StickySelects_12_io_outs_4),
    .io_outs_5(StickySelects_12_io_outs_5),
    .io_outs_6(StickySelects_12_io_outs_6),
    .io_outs_7(StickySelects_12_io_outs_7),
    .io_outs_8(StickySelects_12_io_outs_8)
  );
  StickySelects StickySelects_13 ( // @[MemPrimitives.scala 121:29:@17644.4]
    .clock(StickySelects_13_clock),
    .reset(StickySelects_13_reset),
    .io_ins_0(StickySelects_13_io_ins_0),
    .io_ins_1(StickySelects_13_io_ins_1),
    .io_ins_2(StickySelects_13_io_ins_2),
    .io_ins_3(StickySelects_13_io_ins_3),
    .io_ins_4(StickySelects_13_io_ins_4),
    .io_ins_5(StickySelects_13_io_ins_5),
    .io_ins_6(StickySelects_13_io_ins_6),
    .io_ins_7(StickySelects_13_io_ins_7),
    .io_ins_8(StickySelects_13_io_ins_8),
    .io_outs_0(StickySelects_13_io_outs_0),
    .io_outs_1(StickySelects_13_io_outs_1),
    .io_outs_2(StickySelects_13_io_outs_2),
    .io_outs_3(StickySelects_13_io_outs_3),
    .io_outs_4(StickySelects_13_io_outs_4),
    .io_outs_5(StickySelects_13_io_outs_5),
    .io_outs_6(StickySelects_13_io_outs_6),
    .io_outs_7(StickySelects_13_io_outs_7),
    .io_outs_8(StickySelects_13_io_outs_8)
  );
  StickySelects StickySelects_14 ( // @[MemPrimitives.scala 121:29:@17733.4]
    .clock(StickySelects_14_clock),
    .reset(StickySelects_14_reset),
    .io_ins_0(StickySelects_14_io_ins_0),
    .io_ins_1(StickySelects_14_io_ins_1),
    .io_ins_2(StickySelects_14_io_ins_2),
    .io_ins_3(StickySelects_14_io_ins_3),
    .io_ins_4(StickySelects_14_io_ins_4),
    .io_ins_5(StickySelects_14_io_ins_5),
    .io_ins_6(StickySelects_14_io_ins_6),
    .io_ins_7(StickySelects_14_io_ins_7),
    .io_ins_8(StickySelects_14_io_ins_8),
    .io_outs_0(StickySelects_14_io_outs_0),
    .io_outs_1(StickySelects_14_io_outs_1),
    .io_outs_2(StickySelects_14_io_outs_2),
    .io_outs_3(StickySelects_14_io_outs_3),
    .io_outs_4(StickySelects_14_io_outs_4),
    .io_outs_5(StickySelects_14_io_outs_5),
    .io_outs_6(StickySelects_14_io_outs_6),
    .io_outs_7(StickySelects_14_io_outs_7),
    .io_outs_8(StickySelects_14_io_outs_8)
  );
  StickySelects StickySelects_15 ( // @[MemPrimitives.scala 121:29:@17822.4]
    .clock(StickySelects_15_clock),
    .reset(StickySelects_15_reset),
    .io_ins_0(StickySelects_15_io_ins_0),
    .io_ins_1(StickySelects_15_io_ins_1),
    .io_ins_2(StickySelects_15_io_ins_2),
    .io_ins_3(StickySelects_15_io_ins_3),
    .io_ins_4(StickySelects_15_io_ins_4),
    .io_ins_5(StickySelects_15_io_ins_5),
    .io_ins_6(StickySelects_15_io_ins_6),
    .io_ins_7(StickySelects_15_io_ins_7),
    .io_ins_8(StickySelects_15_io_ins_8),
    .io_outs_0(StickySelects_15_io_outs_0),
    .io_outs_1(StickySelects_15_io_outs_1),
    .io_outs_2(StickySelects_15_io_outs_2),
    .io_outs_3(StickySelects_15_io_outs_3),
    .io_outs_4(StickySelects_15_io_outs_4),
    .io_outs_5(StickySelects_15_io_outs_5),
    .io_outs_6(StickySelects_15_io_outs_6),
    .io_outs_7(StickySelects_15_io_outs_7),
    .io_outs_8(StickySelects_15_io_outs_8)
  );
  StickySelects StickySelects_16 ( // @[MemPrimitives.scala 121:29:@17911.4]
    .clock(StickySelects_16_clock),
    .reset(StickySelects_16_reset),
    .io_ins_0(StickySelects_16_io_ins_0),
    .io_ins_1(StickySelects_16_io_ins_1),
    .io_ins_2(StickySelects_16_io_ins_2),
    .io_ins_3(StickySelects_16_io_ins_3),
    .io_ins_4(StickySelects_16_io_ins_4),
    .io_ins_5(StickySelects_16_io_ins_5),
    .io_ins_6(StickySelects_16_io_ins_6),
    .io_ins_7(StickySelects_16_io_ins_7),
    .io_ins_8(StickySelects_16_io_ins_8),
    .io_outs_0(StickySelects_16_io_outs_0),
    .io_outs_1(StickySelects_16_io_outs_1),
    .io_outs_2(StickySelects_16_io_outs_2),
    .io_outs_3(StickySelects_16_io_outs_3),
    .io_outs_4(StickySelects_16_io_outs_4),
    .io_outs_5(StickySelects_16_io_outs_5),
    .io_outs_6(StickySelects_16_io_outs_6),
    .io_outs_7(StickySelects_16_io_outs_7),
    .io_outs_8(StickySelects_16_io_outs_8)
  );
  StickySelects StickySelects_17 ( // @[MemPrimitives.scala 121:29:@18000.4]
    .clock(StickySelects_17_clock),
    .reset(StickySelects_17_reset),
    .io_ins_0(StickySelects_17_io_ins_0),
    .io_ins_1(StickySelects_17_io_ins_1),
    .io_ins_2(StickySelects_17_io_ins_2),
    .io_ins_3(StickySelects_17_io_ins_3),
    .io_ins_4(StickySelects_17_io_ins_4),
    .io_ins_5(StickySelects_17_io_ins_5),
    .io_ins_6(StickySelects_17_io_ins_6),
    .io_ins_7(StickySelects_17_io_ins_7),
    .io_ins_8(StickySelects_17_io_ins_8),
    .io_outs_0(StickySelects_17_io_outs_0),
    .io_outs_1(StickySelects_17_io_outs_1),
    .io_outs_2(StickySelects_17_io_outs_2),
    .io_outs_3(StickySelects_17_io_outs_3),
    .io_outs_4(StickySelects_17_io_outs_4),
    .io_outs_5(StickySelects_17_io_outs_5),
    .io_outs_6(StickySelects_17_io_outs_6),
    .io_outs_7(StickySelects_17_io_outs_7),
    .io_outs_8(StickySelects_17_io_outs_8)
  );
  StickySelects StickySelects_18 ( // @[MemPrimitives.scala 121:29:@18089.4]
    .clock(StickySelects_18_clock),
    .reset(StickySelects_18_reset),
    .io_ins_0(StickySelects_18_io_ins_0),
    .io_ins_1(StickySelects_18_io_ins_1),
    .io_ins_2(StickySelects_18_io_ins_2),
    .io_ins_3(StickySelects_18_io_ins_3),
    .io_ins_4(StickySelects_18_io_ins_4),
    .io_ins_5(StickySelects_18_io_ins_5),
    .io_ins_6(StickySelects_18_io_ins_6),
    .io_ins_7(StickySelects_18_io_ins_7),
    .io_ins_8(StickySelects_18_io_ins_8),
    .io_outs_0(StickySelects_18_io_outs_0),
    .io_outs_1(StickySelects_18_io_outs_1),
    .io_outs_2(StickySelects_18_io_outs_2),
    .io_outs_3(StickySelects_18_io_outs_3),
    .io_outs_4(StickySelects_18_io_outs_4),
    .io_outs_5(StickySelects_18_io_outs_5),
    .io_outs_6(StickySelects_18_io_outs_6),
    .io_outs_7(StickySelects_18_io_outs_7),
    .io_outs_8(StickySelects_18_io_outs_8)
  );
  StickySelects StickySelects_19 ( // @[MemPrimitives.scala 121:29:@18178.4]
    .clock(StickySelects_19_clock),
    .reset(StickySelects_19_reset),
    .io_ins_0(StickySelects_19_io_ins_0),
    .io_ins_1(StickySelects_19_io_ins_1),
    .io_ins_2(StickySelects_19_io_ins_2),
    .io_ins_3(StickySelects_19_io_ins_3),
    .io_ins_4(StickySelects_19_io_ins_4),
    .io_ins_5(StickySelects_19_io_ins_5),
    .io_ins_6(StickySelects_19_io_ins_6),
    .io_ins_7(StickySelects_19_io_ins_7),
    .io_ins_8(StickySelects_19_io_ins_8),
    .io_outs_0(StickySelects_19_io_outs_0),
    .io_outs_1(StickySelects_19_io_outs_1),
    .io_outs_2(StickySelects_19_io_outs_2),
    .io_outs_3(StickySelects_19_io_outs_3),
    .io_outs_4(StickySelects_19_io_outs_4),
    .io_outs_5(StickySelects_19_io_outs_5),
    .io_outs_6(StickySelects_19_io_outs_6),
    .io_outs_7(StickySelects_19_io_outs_7),
    .io_outs_8(StickySelects_19_io_outs_8)
  );
  StickySelects StickySelects_20 ( // @[MemPrimitives.scala 121:29:@18267.4]
    .clock(StickySelects_20_clock),
    .reset(StickySelects_20_reset),
    .io_ins_0(StickySelects_20_io_ins_0),
    .io_ins_1(StickySelects_20_io_ins_1),
    .io_ins_2(StickySelects_20_io_ins_2),
    .io_ins_3(StickySelects_20_io_ins_3),
    .io_ins_4(StickySelects_20_io_ins_4),
    .io_ins_5(StickySelects_20_io_ins_5),
    .io_ins_6(StickySelects_20_io_ins_6),
    .io_ins_7(StickySelects_20_io_ins_7),
    .io_ins_8(StickySelects_20_io_ins_8),
    .io_outs_0(StickySelects_20_io_outs_0),
    .io_outs_1(StickySelects_20_io_outs_1),
    .io_outs_2(StickySelects_20_io_outs_2),
    .io_outs_3(StickySelects_20_io_outs_3),
    .io_outs_4(StickySelects_20_io_outs_4),
    .io_outs_5(StickySelects_20_io_outs_5),
    .io_outs_6(StickySelects_20_io_outs_6),
    .io_outs_7(StickySelects_20_io_outs_7),
    .io_outs_8(StickySelects_20_io_outs_8)
  );
  StickySelects StickySelects_21 ( // @[MemPrimitives.scala 121:29:@18356.4]
    .clock(StickySelects_21_clock),
    .reset(StickySelects_21_reset),
    .io_ins_0(StickySelects_21_io_ins_0),
    .io_ins_1(StickySelects_21_io_ins_1),
    .io_ins_2(StickySelects_21_io_ins_2),
    .io_ins_3(StickySelects_21_io_ins_3),
    .io_ins_4(StickySelects_21_io_ins_4),
    .io_ins_5(StickySelects_21_io_ins_5),
    .io_ins_6(StickySelects_21_io_ins_6),
    .io_ins_7(StickySelects_21_io_ins_7),
    .io_ins_8(StickySelects_21_io_ins_8),
    .io_outs_0(StickySelects_21_io_outs_0),
    .io_outs_1(StickySelects_21_io_outs_1),
    .io_outs_2(StickySelects_21_io_outs_2),
    .io_outs_3(StickySelects_21_io_outs_3),
    .io_outs_4(StickySelects_21_io_outs_4),
    .io_outs_5(StickySelects_21_io_outs_5),
    .io_outs_6(StickySelects_21_io_outs_6),
    .io_outs_7(StickySelects_21_io_outs_7),
    .io_outs_8(StickySelects_21_io_outs_8)
  );
  StickySelects StickySelects_22 ( // @[MemPrimitives.scala 121:29:@18445.4]
    .clock(StickySelects_22_clock),
    .reset(StickySelects_22_reset),
    .io_ins_0(StickySelects_22_io_ins_0),
    .io_ins_1(StickySelects_22_io_ins_1),
    .io_ins_2(StickySelects_22_io_ins_2),
    .io_ins_3(StickySelects_22_io_ins_3),
    .io_ins_4(StickySelects_22_io_ins_4),
    .io_ins_5(StickySelects_22_io_ins_5),
    .io_ins_6(StickySelects_22_io_ins_6),
    .io_ins_7(StickySelects_22_io_ins_7),
    .io_ins_8(StickySelects_22_io_ins_8),
    .io_outs_0(StickySelects_22_io_outs_0),
    .io_outs_1(StickySelects_22_io_outs_1),
    .io_outs_2(StickySelects_22_io_outs_2),
    .io_outs_3(StickySelects_22_io_outs_3),
    .io_outs_4(StickySelects_22_io_outs_4),
    .io_outs_5(StickySelects_22_io_outs_5),
    .io_outs_6(StickySelects_22_io_outs_6),
    .io_outs_7(StickySelects_22_io_outs_7),
    .io_outs_8(StickySelects_22_io_outs_8)
  );
  StickySelects StickySelects_23 ( // @[MemPrimitives.scala 121:29:@18534.4]
    .clock(StickySelects_23_clock),
    .reset(StickySelects_23_reset),
    .io_ins_0(StickySelects_23_io_ins_0),
    .io_ins_1(StickySelects_23_io_ins_1),
    .io_ins_2(StickySelects_23_io_ins_2),
    .io_ins_3(StickySelects_23_io_ins_3),
    .io_ins_4(StickySelects_23_io_ins_4),
    .io_ins_5(StickySelects_23_io_ins_5),
    .io_ins_6(StickySelects_23_io_ins_6),
    .io_ins_7(StickySelects_23_io_ins_7),
    .io_ins_8(StickySelects_23_io_ins_8),
    .io_outs_0(StickySelects_23_io_outs_0),
    .io_outs_1(StickySelects_23_io_outs_1),
    .io_outs_2(StickySelects_23_io_outs_2),
    .io_outs_3(StickySelects_23_io_outs_3),
    .io_outs_4(StickySelects_23_io_outs_4),
    .io_outs_5(StickySelects_23_io_outs_5),
    .io_outs_6(StickySelects_23_io_outs_6),
    .io_outs_7(StickySelects_23_io_outs_7),
    .io_outs_8(StickySelects_23_io_outs_8)
  );
  RetimeWrapper_44 RetimeWrapper ( // @[package.scala 93:22:@18624.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_1 ( // @[package.scala 93:22:@18632.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_2 ( // @[package.scala 93:22:@18640.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_3 ( // @[package.scala 93:22:@18648.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_4 ( // @[package.scala 93:22:@18656.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_5 ( // @[package.scala 93:22:@18664.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_6 ( // @[package.scala 93:22:@18672.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_7 ( // @[package.scala 93:22:@18680.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_8 ( // @[package.scala 93:22:@18688.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_9 ( // @[package.scala 93:22:@18696.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_10 ( // @[package.scala 93:22:@18704.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_11 ( // @[package.scala 93:22:@18712.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_12 ( // @[package.scala 93:22:@18768.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_13 ( // @[package.scala 93:22:@18776.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_14 ( // @[package.scala 93:22:@18784.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_15 ( // @[package.scala 93:22:@18792.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_16 ( // @[package.scala 93:22:@18800.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_17 ( // @[package.scala 93:22:@18808.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_18 ( // @[package.scala 93:22:@18816.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_19 ( // @[package.scala 93:22:@18824.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_20 ( // @[package.scala 93:22:@18832.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_21 ( // @[package.scala 93:22:@18840.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_22 ( // @[package.scala 93:22:@18848.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_23 ( // @[package.scala 93:22:@18856.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_24 ( // @[package.scala 93:22:@18912.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_25 ( // @[package.scala 93:22:@18920.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_26 ( // @[package.scala 93:22:@18928.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_27 ( // @[package.scala 93:22:@18936.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_28 ( // @[package.scala 93:22:@18944.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_29 ( // @[package.scala 93:22:@18952.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_30 ( // @[package.scala 93:22:@18960.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_31 ( // @[package.scala 93:22:@18968.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_32 ( // @[package.scala 93:22:@18976.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_33 ( // @[package.scala 93:22:@18984.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_34 ( // @[package.scala 93:22:@18992.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_35 ( // @[package.scala 93:22:@19000.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_36 ( // @[package.scala 93:22:@19056.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_37 ( // @[package.scala 93:22:@19064.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_38 ( // @[package.scala 93:22:@19072.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_39 ( // @[package.scala 93:22:@19080.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_40 ( // @[package.scala 93:22:@19088.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_41 ( // @[package.scala 93:22:@19096.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_42 ( // @[package.scala 93:22:@19104.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_43 ( // @[package.scala 93:22:@19112.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_44 ( // @[package.scala 93:22:@19120.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_45 ( // @[package.scala 93:22:@19128.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_46 ( // @[package.scala 93:22:@19136.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_47 ( // @[package.scala 93:22:@19144.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_48 ( // @[package.scala 93:22:@19200.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_49 ( // @[package.scala 93:22:@19208.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_50 ( // @[package.scala 93:22:@19216.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_51 ( // @[package.scala 93:22:@19224.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_52 ( // @[package.scala 93:22:@19232.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_53 ( // @[package.scala 93:22:@19240.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_54 ( // @[package.scala 93:22:@19248.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_55 ( // @[package.scala 93:22:@19256.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_56 ( // @[package.scala 93:22:@19264.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_57 ( // @[package.scala 93:22:@19272.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_58 ( // @[package.scala 93:22:@19280.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_59 ( // @[package.scala 93:22:@19288.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_60 ( // @[package.scala 93:22:@19344.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_61 ( // @[package.scala 93:22:@19352.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_62 ( // @[package.scala 93:22:@19360.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_63 ( // @[package.scala 93:22:@19368.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_64 ( // @[package.scala 93:22:@19376.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_65 ( // @[package.scala 93:22:@19384.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_66 ( // @[package.scala 93:22:@19392.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_67 ( // @[package.scala 93:22:@19400.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_68 ( // @[package.scala 93:22:@19408.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_69 ( // @[package.scala 93:22:@19416.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_70 ( // @[package.scala 93:22:@19424.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_71 ( // @[package.scala 93:22:@19432.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_72 ( // @[package.scala 93:22:@19488.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_73 ( // @[package.scala 93:22:@19496.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_74 ( // @[package.scala 93:22:@19504.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_75 ( // @[package.scala 93:22:@19512.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_76 ( // @[package.scala 93:22:@19520.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_77 ( // @[package.scala 93:22:@19528.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_78 ( // @[package.scala 93:22:@19536.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_79 ( // @[package.scala 93:22:@19544.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_80 ( // @[package.scala 93:22:@19552.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_81 ( // @[package.scala 93:22:@19560.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_82 ( // @[package.scala 93:22:@19568.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_83 ( // @[package.scala 93:22:@19576.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_84 ( // @[package.scala 93:22:@19632.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_85 ( // @[package.scala 93:22:@19640.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_86 ( // @[package.scala 93:22:@19648.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_87 ( // @[package.scala 93:22:@19656.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_88 ( // @[package.scala 93:22:@19664.4]
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_89 ( // @[package.scala 93:22:@19672.4]
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_90 ( // @[package.scala 93:22:@19680.4]
    .clock(RetimeWrapper_90_clock),
    .reset(RetimeWrapper_90_reset),
    .io_flow(RetimeWrapper_90_io_flow),
    .io_in(RetimeWrapper_90_io_in),
    .io_out(RetimeWrapper_90_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_91 ( // @[package.scala 93:22:@19688.4]
    .clock(RetimeWrapper_91_clock),
    .reset(RetimeWrapper_91_reset),
    .io_flow(RetimeWrapper_91_io_flow),
    .io_in(RetimeWrapper_91_io_in),
    .io_out(RetimeWrapper_91_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_92 ( // @[package.scala 93:22:@19696.4]
    .clock(RetimeWrapper_92_clock),
    .reset(RetimeWrapper_92_reset),
    .io_flow(RetimeWrapper_92_io_flow),
    .io_in(RetimeWrapper_92_io_in),
    .io_out(RetimeWrapper_92_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_93 ( // @[package.scala 93:22:@19704.4]
    .clock(RetimeWrapper_93_clock),
    .reset(RetimeWrapper_93_reset),
    .io_flow(RetimeWrapper_93_io_flow),
    .io_in(RetimeWrapper_93_io_in),
    .io_out(RetimeWrapper_93_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_94 ( // @[package.scala 93:22:@19712.4]
    .clock(RetimeWrapper_94_clock),
    .reset(RetimeWrapper_94_reset),
    .io_flow(RetimeWrapper_94_io_flow),
    .io_in(RetimeWrapper_94_io_in),
    .io_out(RetimeWrapper_94_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_95 ( // @[package.scala 93:22:@19720.4]
    .clock(RetimeWrapper_95_clock),
    .reset(RetimeWrapper_95_reset),
    .io_flow(RetimeWrapper_95_io_flow),
    .io_in(RetimeWrapper_95_io_in),
    .io_out(RetimeWrapper_95_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_96 ( // @[package.scala 93:22:@19776.4]
    .clock(RetimeWrapper_96_clock),
    .reset(RetimeWrapper_96_reset),
    .io_flow(RetimeWrapper_96_io_flow),
    .io_in(RetimeWrapper_96_io_in),
    .io_out(RetimeWrapper_96_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_97 ( // @[package.scala 93:22:@19784.4]
    .clock(RetimeWrapper_97_clock),
    .reset(RetimeWrapper_97_reset),
    .io_flow(RetimeWrapper_97_io_flow),
    .io_in(RetimeWrapper_97_io_in),
    .io_out(RetimeWrapper_97_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_98 ( // @[package.scala 93:22:@19792.4]
    .clock(RetimeWrapper_98_clock),
    .reset(RetimeWrapper_98_reset),
    .io_flow(RetimeWrapper_98_io_flow),
    .io_in(RetimeWrapper_98_io_in),
    .io_out(RetimeWrapper_98_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_99 ( // @[package.scala 93:22:@19800.4]
    .clock(RetimeWrapper_99_clock),
    .reset(RetimeWrapper_99_reset),
    .io_flow(RetimeWrapper_99_io_flow),
    .io_in(RetimeWrapper_99_io_in),
    .io_out(RetimeWrapper_99_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_100 ( // @[package.scala 93:22:@19808.4]
    .clock(RetimeWrapper_100_clock),
    .reset(RetimeWrapper_100_reset),
    .io_flow(RetimeWrapper_100_io_flow),
    .io_in(RetimeWrapper_100_io_in),
    .io_out(RetimeWrapper_100_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_101 ( // @[package.scala 93:22:@19816.4]
    .clock(RetimeWrapper_101_clock),
    .reset(RetimeWrapper_101_reset),
    .io_flow(RetimeWrapper_101_io_flow),
    .io_in(RetimeWrapper_101_io_in),
    .io_out(RetimeWrapper_101_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_102 ( // @[package.scala 93:22:@19824.4]
    .clock(RetimeWrapper_102_clock),
    .reset(RetimeWrapper_102_reset),
    .io_flow(RetimeWrapper_102_io_flow),
    .io_in(RetimeWrapper_102_io_in),
    .io_out(RetimeWrapper_102_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_103 ( // @[package.scala 93:22:@19832.4]
    .clock(RetimeWrapper_103_clock),
    .reset(RetimeWrapper_103_reset),
    .io_flow(RetimeWrapper_103_io_flow),
    .io_in(RetimeWrapper_103_io_in),
    .io_out(RetimeWrapper_103_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_104 ( // @[package.scala 93:22:@19840.4]
    .clock(RetimeWrapper_104_clock),
    .reset(RetimeWrapper_104_reset),
    .io_flow(RetimeWrapper_104_io_flow),
    .io_in(RetimeWrapper_104_io_in),
    .io_out(RetimeWrapper_104_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_105 ( // @[package.scala 93:22:@19848.4]
    .clock(RetimeWrapper_105_clock),
    .reset(RetimeWrapper_105_reset),
    .io_flow(RetimeWrapper_105_io_flow),
    .io_in(RetimeWrapper_105_io_in),
    .io_out(RetimeWrapper_105_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_106 ( // @[package.scala 93:22:@19856.4]
    .clock(RetimeWrapper_106_clock),
    .reset(RetimeWrapper_106_reset),
    .io_flow(RetimeWrapper_106_io_flow),
    .io_in(RetimeWrapper_106_io_in),
    .io_out(RetimeWrapper_106_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_107 ( // @[package.scala 93:22:@19864.4]
    .clock(RetimeWrapper_107_clock),
    .reset(RetimeWrapper_107_reset),
    .io_flow(RetimeWrapper_107_io_flow),
    .io_in(RetimeWrapper_107_io_in),
    .io_out(RetimeWrapper_107_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_108 ( // @[package.scala 93:22:@19920.4]
    .clock(RetimeWrapper_108_clock),
    .reset(RetimeWrapper_108_reset),
    .io_flow(RetimeWrapper_108_io_flow),
    .io_in(RetimeWrapper_108_io_in),
    .io_out(RetimeWrapper_108_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_109 ( // @[package.scala 93:22:@19928.4]
    .clock(RetimeWrapper_109_clock),
    .reset(RetimeWrapper_109_reset),
    .io_flow(RetimeWrapper_109_io_flow),
    .io_in(RetimeWrapper_109_io_in),
    .io_out(RetimeWrapper_109_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_110 ( // @[package.scala 93:22:@19936.4]
    .clock(RetimeWrapper_110_clock),
    .reset(RetimeWrapper_110_reset),
    .io_flow(RetimeWrapper_110_io_flow),
    .io_in(RetimeWrapper_110_io_in),
    .io_out(RetimeWrapper_110_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_111 ( // @[package.scala 93:22:@19944.4]
    .clock(RetimeWrapper_111_clock),
    .reset(RetimeWrapper_111_reset),
    .io_flow(RetimeWrapper_111_io_flow),
    .io_in(RetimeWrapper_111_io_in),
    .io_out(RetimeWrapper_111_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_112 ( // @[package.scala 93:22:@19952.4]
    .clock(RetimeWrapper_112_clock),
    .reset(RetimeWrapper_112_reset),
    .io_flow(RetimeWrapper_112_io_flow),
    .io_in(RetimeWrapper_112_io_in),
    .io_out(RetimeWrapper_112_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_113 ( // @[package.scala 93:22:@19960.4]
    .clock(RetimeWrapper_113_clock),
    .reset(RetimeWrapper_113_reset),
    .io_flow(RetimeWrapper_113_io_flow),
    .io_in(RetimeWrapper_113_io_in),
    .io_out(RetimeWrapper_113_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_114 ( // @[package.scala 93:22:@19968.4]
    .clock(RetimeWrapper_114_clock),
    .reset(RetimeWrapper_114_reset),
    .io_flow(RetimeWrapper_114_io_flow),
    .io_in(RetimeWrapper_114_io_in),
    .io_out(RetimeWrapper_114_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_115 ( // @[package.scala 93:22:@19976.4]
    .clock(RetimeWrapper_115_clock),
    .reset(RetimeWrapper_115_reset),
    .io_flow(RetimeWrapper_115_io_flow),
    .io_in(RetimeWrapper_115_io_in),
    .io_out(RetimeWrapper_115_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_116 ( // @[package.scala 93:22:@19984.4]
    .clock(RetimeWrapper_116_clock),
    .reset(RetimeWrapper_116_reset),
    .io_flow(RetimeWrapper_116_io_flow),
    .io_in(RetimeWrapper_116_io_in),
    .io_out(RetimeWrapper_116_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_117 ( // @[package.scala 93:22:@19992.4]
    .clock(RetimeWrapper_117_clock),
    .reset(RetimeWrapper_117_reset),
    .io_flow(RetimeWrapper_117_io_flow),
    .io_in(RetimeWrapper_117_io_in),
    .io_out(RetimeWrapper_117_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_118 ( // @[package.scala 93:22:@20000.4]
    .clock(RetimeWrapper_118_clock),
    .reset(RetimeWrapper_118_reset),
    .io_flow(RetimeWrapper_118_io_flow),
    .io_in(RetimeWrapper_118_io_in),
    .io_out(RetimeWrapper_118_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_119 ( // @[package.scala 93:22:@20008.4]
    .clock(RetimeWrapper_119_clock),
    .reset(RetimeWrapper_119_reset),
    .io_flow(RetimeWrapper_119_io_flow),
    .io_in(RetimeWrapper_119_io_in),
    .io_out(RetimeWrapper_119_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_120 ( // @[package.scala 93:22:@20064.4]
    .clock(RetimeWrapper_120_clock),
    .reset(RetimeWrapper_120_reset),
    .io_flow(RetimeWrapper_120_io_flow),
    .io_in(RetimeWrapper_120_io_in),
    .io_out(RetimeWrapper_120_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_121 ( // @[package.scala 93:22:@20072.4]
    .clock(RetimeWrapper_121_clock),
    .reset(RetimeWrapper_121_reset),
    .io_flow(RetimeWrapper_121_io_flow),
    .io_in(RetimeWrapper_121_io_in),
    .io_out(RetimeWrapper_121_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_122 ( // @[package.scala 93:22:@20080.4]
    .clock(RetimeWrapper_122_clock),
    .reset(RetimeWrapper_122_reset),
    .io_flow(RetimeWrapper_122_io_flow),
    .io_in(RetimeWrapper_122_io_in),
    .io_out(RetimeWrapper_122_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_123 ( // @[package.scala 93:22:@20088.4]
    .clock(RetimeWrapper_123_clock),
    .reset(RetimeWrapper_123_reset),
    .io_flow(RetimeWrapper_123_io_flow),
    .io_in(RetimeWrapper_123_io_in),
    .io_out(RetimeWrapper_123_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_124 ( // @[package.scala 93:22:@20096.4]
    .clock(RetimeWrapper_124_clock),
    .reset(RetimeWrapper_124_reset),
    .io_flow(RetimeWrapper_124_io_flow),
    .io_in(RetimeWrapper_124_io_in),
    .io_out(RetimeWrapper_124_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_125 ( // @[package.scala 93:22:@20104.4]
    .clock(RetimeWrapper_125_clock),
    .reset(RetimeWrapper_125_reset),
    .io_flow(RetimeWrapper_125_io_flow),
    .io_in(RetimeWrapper_125_io_in),
    .io_out(RetimeWrapper_125_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_126 ( // @[package.scala 93:22:@20112.4]
    .clock(RetimeWrapper_126_clock),
    .reset(RetimeWrapper_126_reset),
    .io_flow(RetimeWrapper_126_io_flow),
    .io_in(RetimeWrapper_126_io_in),
    .io_out(RetimeWrapper_126_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_127 ( // @[package.scala 93:22:@20120.4]
    .clock(RetimeWrapper_127_clock),
    .reset(RetimeWrapper_127_reset),
    .io_flow(RetimeWrapper_127_io_flow),
    .io_in(RetimeWrapper_127_io_in),
    .io_out(RetimeWrapper_127_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_128 ( // @[package.scala 93:22:@20128.4]
    .clock(RetimeWrapper_128_clock),
    .reset(RetimeWrapper_128_reset),
    .io_flow(RetimeWrapper_128_io_flow),
    .io_in(RetimeWrapper_128_io_in),
    .io_out(RetimeWrapper_128_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_129 ( // @[package.scala 93:22:@20136.4]
    .clock(RetimeWrapper_129_clock),
    .reset(RetimeWrapper_129_reset),
    .io_flow(RetimeWrapper_129_io_flow),
    .io_in(RetimeWrapper_129_io_in),
    .io_out(RetimeWrapper_129_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_130 ( // @[package.scala 93:22:@20144.4]
    .clock(RetimeWrapper_130_clock),
    .reset(RetimeWrapper_130_reset),
    .io_flow(RetimeWrapper_130_io_flow),
    .io_in(RetimeWrapper_130_io_in),
    .io_out(RetimeWrapper_130_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_131 ( // @[package.scala 93:22:@20152.4]
    .clock(RetimeWrapper_131_clock),
    .reset(RetimeWrapper_131_reset),
    .io_flow(RetimeWrapper_131_io_flow),
    .io_in(RetimeWrapper_131_io_in),
    .io_out(RetimeWrapper_131_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_132 ( // @[package.scala 93:22:@20208.4]
    .clock(RetimeWrapper_132_clock),
    .reset(RetimeWrapper_132_reset),
    .io_flow(RetimeWrapper_132_io_flow),
    .io_in(RetimeWrapper_132_io_in),
    .io_out(RetimeWrapper_132_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_133 ( // @[package.scala 93:22:@20216.4]
    .clock(RetimeWrapper_133_clock),
    .reset(RetimeWrapper_133_reset),
    .io_flow(RetimeWrapper_133_io_flow),
    .io_in(RetimeWrapper_133_io_in),
    .io_out(RetimeWrapper_133_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_134 ( // @[package.scala 93:22:@20224.4]
    .clock(RetimeWrapper_134_clock),
    .reset(RetimeWrapper_134_reset),
    .io_flow(RetimeWrapper_134_io_flow),
    .io_in(RetimeWrapper_134_io_in),
    .io_out(RetimeWrapper_134_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_135 ( // @[package.scala 93:22:@20232.4]
    .clock(RetimeWrapper_135_clock),
    .reset(RetimeWrapper_135_reset),
    .io_flow(RetimeWrapper_135_io_flow),
    .io_in(RetimeWrapper_135_io_in),
    .io_out(RetimeWrapper_135_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_136 ( // @[package.scala 93:22:@20240.4]
    .clock(RetimeWrapper_136_clock),
    .reset(RetimeWrapper_136_reset),
    .io_flow(RetimeWrapper_136_io_flow),
    .io_in(RetimeWrapper_136_io_in),
    .io_out(RetimeWrapper_136_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_137 ( // @[package.scala 93:22:@20248.4]
    .clock(RetimeWrapper_137_clock),
    .reset(RetimeWrapper_137_reset),
    .io_flow(RetimeWrapper_137_io_flow),
    .io_in(RetimeWrapper_137_io_in),
    .io_out(RetimeWrapper_137_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_138 ( // @[package.scala 93:22:@20256.4]
    .clock(RetimeWrapper_138_clock),
    .reset(RetimeWrapper_138_reset),
    .io_flow(RetimeWrapper_138_io_flow),
    .io_in(RetimeWrapper_138_io_in),
    .io_out(RetimeWrapper_138_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_139 ( // @[package.scala 93:22:@20264.4]
    .clock(RetimeWrapper_139_clock),
    .reset(RetimeWrapper_139_reset),
    .io_flow(RetimeWrapper_139_io_flow),
    .io_in(RetimeWrapper_139_io_in),
    .io_out(RetimeWrapper_139_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_140 ( // @[package.scala 93:22:@20272.4]
    .clock(RetimeWrapper_140_clock),
    .reset(RetimeWrapper_140_reset),
    .io_flow(RetimeWrapper_140_io_flow),
    .io_in(RetimeWrapper_140_io_in),
    .io_out(RetimeWrapper_140_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_141 ( // @[package.scala 93:22:@20280.4]
    .clock(RetimeWrapper_141_clock),
    .reset(RetimeWrapper_141_reset),
    .io_flow(RetimeWrapper_141_io_flow),
    .io_in(RetimeWrapper_141_io_in),
    .io_out(RetimeWrapper_141_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_142 ( // @[package.scala 93:22:@20288.4]
    .clock(RetimeWrapper_142_clock),
    .reset(RetimeWrapper_142_reset),
    .io_flow(RetimeWrapper_142_io_flow),
    .io_in(RetimeWrapper_142_io_in),
    .io_out(RetimeWrapper_142_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_143 ( // @[package.scala 93:22:@20296.4]
    .clock(RetimeWrapper_143_clock),
    .reset(RetimeWrapper_143_reset),
    .io_flow(RetimeWrapper_143_io_flow),
    .io_in(RetimeWrapper_143_io_in),
    .io_out(RetimeWrapper_143_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_144 ( // @[package.scala 93:22:@20352.4]
    .clock(RetimeWrapper_144_clock),
    .reset(RetimeWrapper_144_reset),
    .io_flow(RetimeWrapper_144_io_flow),
    .io_in(RetimeWrapper_144_io_in),
    .io_out(RetimeWrapper_144_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_145 ( // @[package.scala 93:22:@20360.4]
    .clock(RetimeWrapper_145_clock),
    .reset(RetimeWrapper_145_reset),
    .io_flow(RetimeWrapper_145_io_flow),
    .io_in(RetimeWrapper_145_io_in),
    .io_out(RetimeWrapper_145_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_146 ( // @[package.scala 93:22:@20368.4]
    .clock(RetimeWrapper_146_clock),
    .reset(RetimeWrapper_146_reset),
    .io_flow(RetimeWrapper_146_io_flow),
    .io_in(RetimeWrapper_146_io_in),
    .io_out(RetimeWrapper_146_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_147 ( // @[package.scala 93:22:@20376.4]
    .clock(RetimeWrapper_147_clock),
    .reset(RetimeWrapper_147_reset),
    .io_flow(RetimeWrapper_147_io_flow),
    .io_in(RetimeWrapper_147_io_in),
    .io_out(RetimeWrapper_147_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_148 ( // @[package.scala 93:22:@20384.4]
    .clock(RetimeWrapper_148_clock),
    .reset(RetimeWrapper_148_reset),
    .io_flow(RetimeWrapper_148_io_flow),
    .io_in(RetimeWrapper_148_io_in),
    .io_out(RetimeWrapper_148_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_149 ( // @[package.scala 93:22:@20392.4]
    .clock(RetimeWrapper_149_clock),
    .reset(RetimeWrapper_149_reset),
    .io_flow(RetimeWrapper_149_io_flow),
    .io_in(RetimeWrapper_149_io_in),
    .io_out(RetimeWrapper_149_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_150 ( // @[package.scala 93:22:@20400.4]
    .clock(RetimeWrapper_150_clock),
    .reset(RetimeWrapper_150_reset),
    .io_flow(RetimeWrapper_150_io_flow),
    .io_in(RetimeWrapper_150_io_in),
    .io_out(RetimeWrapper_150_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_151 ( // @[package.scala 93:22:@20408.4]
    .clock(RetimeWrapper_151_clock),
    .reset(RetimeWrapper_151_reset),
    .io_flow(RetimeWrapper_151_io_flow),
    .io_in(RetimeWrapper_151_io_in),
    .io_out(RetimeWrapper_151_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_152 ( // @[package.scala 93:22:@20416.4]
    .clock(RetimeWrapper_152_clock),
    .reset(RetimeWrapper_152_reset),
    .io_flow(RetimeWrapper_152_io_flow),
    .io_in(RetimeWrapper_152_io_in),
    .io_out(RetimeWrapper_152_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_153 ( // @[package.scala 93:22:@20424.4]
    .clock(RetimeWrapper_153_clock),
    .reset(RetimeWrapper_153_reset),
    .io_flow(RetimeWrapper_153_io_flow),
    .io_in(RetimeWrapper_153_io_in),
    .io_out(RetimeWrapper_153_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_154 ( // @[package.scala 93:22:@20432.4]
    .clock(RetimeWrapper_154_clock),
    .reset(RetimeWrapper_154_reset),
    .io_flow(RetimeWrapper_154_io_flow),
    .io_in(RetimeWrapper_154_io_in),
    .io_out(RetimeWrapper_154_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_155 ( // @[package.scala 93:22:@20440.4]
    .clock(RetimeWrapper_155_clock),
    .reset(RetimeWrapper_155_reset),
    .io_flow(RetimeWrapper_155_io_flow),
    .io_in(RetimeWrapper_155_io_in),
    .io_out(RetimeWrapper_155_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_156 ( // @[package.scala 93:22:@20496.4]
    .clock(RetimeWrapper_156_clock),
    .reset(RetimeWrapper_156_reset),
    .io_flow(RetimeWrapper_156_io_flow),
    .io_in(RetimeWrapper_156_io_in),
    .io_out(RetimeWrapper_156_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_157 ( // @[package.scala 93:22:@20504.4]
    .clock(RetimeWrapper_157_clock),
    .reset(RetimeWrapper_157_reset),
    .io_flow(RetimeWrapper_157_io_flow),
    .io_in(RetimeWrapper_157_io_in),
    .io_out(RetimeWrapper_157_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_158 ( // @[package.scala 93:22:@20512.4]
    .clock(RetimeWrapper_158_clock),
    .reset(RetimeWrapper_158_reset),
    .io_flow(RetimeWrapper_158_io_flow),
    .io_in(RetimeWrapper_158_io_in),
    .io_out(RetimeWrapper_158_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_159 ( // @[package.scala 93:22:@20520.4]
    .clock(RetimeWrapper_159_clock),
    .reset(RetimeWrapper_159_reset),
    .io_flow(RetimeWrapper_159_io_flow),
    .io_in(RetimeWrapper_159_io_in),
    .io_out(RetimeWrapper_159_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_160 ( // @[package.scala 93:22:@20528.4]
    .clock(RetimeWrapper_160_clock),
    .reset(RetimeWrapper_160_reset),
    .io_flow(RetimeWrapper_160_io_flow),
    .io_in(RetimeWrapper_160_io_in),
    .io_out(RetimeWrapper_160_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_161 ( // @[package.scala 93:22:@20536.4]
    .clock(RetimeWrapper_161_clock),
    .reset(RetimeWrapper_161_reset),
    .io_flow(RetimeWrapper_161_io_flow),
    .io_in(RetimeWrapper_161_io_in),
    .io_out(RetimeWrapper_161_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_162 ( // @[package.scala 93:22:@20544.4]
    .clock(RetimeWrapper_162_clock),
    .reset(RetimeWrapper_162_reset),
    .io_flow(RetimeWrapper_162_io_flow),
    .io_in(RetimeWrapper_162_io_in),
    .io_out(RetimeWrapper_162_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_163 ( // @[package.scala 93:22:@20552.4]
    .clock(RetimeWrapper_163_clock),
    .reset(RetimeWrapper_163_reset),
    .io_flow(RetimeWrapper_163_io_flow),
    .io_in(RetimeWrapper_163_io_in),
    .io_out(RetimeWrapper_163_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_164 ( // @[package.scala 93:22:@20560.4]
    .clock(RetimeWrapper_164_clock),
    .reset(RetimeWrapper_164_reset),
    .io_flow(RetimeWrapper_164_io_flow),
    .io_in(RetimeWrapper_164_io_in),
    .io_out(RetimeWrapper_164_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_165 ( // @[package.scala 93:22:@20568.4]
    .clock(RetimeWrapper_165_clock),
    .reset(RetimeWrapper_165_reset),
    .io_flow(RetimeWrapper_165_io_flow),
    .io_in(RetimeWrapper_165_io_in),
    .io_out(RetimeWrapper_165_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_166 ( // @[package.scala 93:22:@20576.4]
    .clock(RetimeWrapper_166_clock),
    .reset(RetimeWrapper_166_reset),
    .io_flow(RetimeWrapper_166_io_flow),
    .io_in(RetimeWrapper_166_io_in),
    .io_out(RetimeWrapper_166_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_167 ( // @[package.scala 93:22:@20584.4]
    .clock(RetimeWrapper_167_clock),
    .reset(RetimeWrapper_167_reset),
    .io_flow(RetimeWrapper_167_io_flow),
    .io_in(RetimeWrapper_167_io_in),
    .io_out(RetimeWrapper_167_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_168 ( // @[package.scala 93:22:@20640.4]
    .clock(RetimeWrapper_168_clock),
    .reset(RetimeWrapper_168_reset),
    .io_flow(RetimeWrapper_168_io_flow),
    .io_in(RetimeWrapper_168_io_in),
    .io_out(RetimeWrapper_168_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_169 ( // @[package.scala 93:22:@20648.4]
    .clock(RetimeWrapper_169_clock),
    .reset(RetimeWrapper_169_reset),
    .io_flow(RetimeWrapper_169_io_flow),
    .io_in(RetimeWrapper_169_io_in),
    .io_out(RetimeWrapper_169_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_170 ( // @[package.scala 93:22:@20656.4]
    .clock(RetimeWrapper_170_clock),
    .reset(RetimeWrapper_170_reset),
    .io_flow(RetimeWrapper_170_io_flow),
    .io_in(RetimeWrapper_170_io_in),
    .io_out(RetimeWrapper_170_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_171 ( // @[package.scala 93:22:@20664.4]
    .clock(RetimeWrapper_171_clock),
    .reset(RetimeWrapper_171_reset),
    .io_flow(RetimeWrapper_171_io_flow),
    .io_in(RetimeWrapper_171_io_in),
    .io_out(RetimeWrapper_171_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_172 ( // @[package.scala 93:22:@20672.4]
    .clock(RetimeWrapper_172_clock),
    .reset(RetimeWrapper_172_reset),
    .io_flow(RetimeWrapper_172_io_flow),
    .io_in(RetimeWrapper_172_io_in),
    .io_out(RetimeWrapper_172_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_173 ( // @[package.scala 93:22:@20680.4]
    .clock(RetimeWrapper_173_clock),
    .reset(RetimeWrapper_173_reset),
    .io_flow(RetimeWrapper_173_io_flow),
    .io_in(RetimeWrapper_173_io_in),
    .io_out(RetimeWrapper_173_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_174 ( // @[package.scala 93:22:@20688.4]
    .clock(RetimeWrapper_174_clock),
    .reset(RetimeWrapper_174_reset),
    .io_flow(RetimeWrapper_174_io_flow),
    .io_in(RetimeWrapper_174_io_in),
    .io_out(RetimeWrapper_174_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_175 ( // @[package.scala 93:22:@20696.4]
    .clock(RetimeWrapper_175_clock),
    .reset(RetimeWrapper_175_reset),
    .io_flow(RetimeWrapper_175_io_flow),
    .io_in(RetimeWrapper_175_io_in),
    .io_out(RetimeWrapper_175_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_176 ( // @[package.scala 93:22:@20704.4]
    .clock(RetimeWrapper_176_clock),
    .reset(RetimeWrapper_176_reset),
    .io_flow(RetimeWrapper_176_io_flow),
    .io_in(RetimeWrapper_176_io_in),
    .io_out(RetimeWrapper_176_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_177 ( // @[package.scala 93:22:@20712.4]
    .clock(RetimeWrapper_177_clock),
    .reset(RetimeWrapper_177_reset),
    .io_flow(RetimeWrapper_177_io_flow),
    .io_in(RetimeWrapper_177_io_in),
    .io_out(RetimeWrapper_177_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_178 ( // @[package.scala 93:22:@20720.4]
    .clock(RetimeWrapper_178_clock),
    .reset(RetimeWrapper_178_reset),
    .io_flow(RetimeWrapper_178_io_flow),
    .io_in(RetimeWrapper_178_io_in),
    .io_out(RetimeWrapper_178_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_179 ( // @[package.scala 93:22:@20728.4]
    .clock(RetimeWrapper_179_clock),
    .reset(RetimeWrapper_179_reset),
    .io_flow(RetimeWrapper_179_io_flow),
    .io_in(RetimeWrapper_179_io_in),
    .io_out(RetimeWrapper_179_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_180 ( // @[package.scala 93:22:@20784.4]
    .clock(RetimeWrapper_180_clock),
    .reset(RetimeWrapper_180_reset),
    .io_flow(RetimeWrapper_180_io_flow),
    .io_in(RetimeWrapper_180_io_in),
    .io_out(RetimeWrapper_180_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_181 ( // @[package.scala 93:22:@20792.4]
    .clock(RetimeWrapper_181_clock),
    .reset(RetimeWrapper_181_reset),
    .io_flow(RetimeWrapper_181_io_flow),
    .io_in(RetimeWrapper_181_io_in),
    .io_out(RetimeWrapper_181_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_182 ( // @[package.scala 93:22:@20800.4]
    .clock(RetimeWrapper_182_clock),
    .reset(RetimeWrapper_182_reset),
    .io_flow(RetimeWrapper_182_io_flow),
    .io_in(RetimeWrapper_182_io_in),
    .io_out(RetimeWrapper_182_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_183 ( // @[package.scala 93:22:@20808.4]
    .clock(RetimeWrapper_183_clock),
    .reset(RetimeWrapper_183_reset),
    .io_flow(RetimeWrapper_183_io_flow),
    .io_in(RetimeWrapper_183_io_in),
    .io_out(RetimeWrapper_183_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_184 ( // @[package.scala 93:22:@20816.4]
    .clock(RetimeWrapper_184_clock),
    .reset(RetimeWrapper_184_reset),
    .io_flow(RetimeWrapper_184_io_flow),
    .io_in(RetimeWrapper_184_io_in),
    .io_out(RetimeWrapper_184_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_185 ( // @[package.scala 93:22:@20824.4]
    .clock(RetimeWrapper_185_clock),
    .reset(RetimeWrapper_185_reset),
    .io_flow(RetimeWrapper_185_io_flow),
    .io_in(RetimeWrapper_185_io_in),
    .io_out(RetimeWrapper_185_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_186 ( // @[package.scala 93:22:@20832.4]
    .clock(RetimeWrapper_186_clock),
    .reset(RetimeWrapper_186_reset),
    .io_flow(RetimeWrapper_186_io_flow),
    .io_in(RetimeWrapper_186_io_in),
    .io_out(RetimeWrapper_186_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_187 ( // @[package.scala 93:22:@20840.4]
    .clock(RetimeWrapper_187_clock),
    .reset(RetimeWrapper_187_reset),
    .io_flow(RetimeWrapper_187_io_flow),
    .io_in(RetimeWrapper_187_io_in),
    .io_out(RetimeWrapper_187_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_188 ( // @[package.scala 93:22:@20848.4]
    .clock(RetimeWrapper_188_clock),
    .reset(RetimeWrapper_188_reset),
    .io_flow(RetimeWrapper_188_io_flow),
    .io_in(RetimeWrapper_188_io_in),
    .io_out(RetimeWrapper_188_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_189 ( // @[package.scala 93:22:@20856.4]
    .clock(RetimeWrapper_189_clock),
    .reset(RetimeWrapper_189_reset),
    .io_flow(RetimeWrapper_189_io_flow),
    .io_in(RetimeWrapper_189_io_in),
    .io_out(RetimeWrapper_189_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_190 ( // @[package.scala 93:22:@20864.4]
    .clock(RetimeWrapper_190_clock),
    .reset(RetimeWrapper_190_reset),
    .io_flow(RetimeWrapper_190_io_flow),
    .io_in(RetimeWrapper_190_io_in),
    .io_out(RetimeWrapper_190_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_191 ( // @[package.scala 93:22:@20872.4]
    .clock(RetimeWrapper_191_clock),
    .reset(RetimeWrapper_191_reset),
    .io_flow(RetimeWrapper_191_io_flow),
    .io_in(RetimeWrapper_191_io_in),
    .io_out(RetimeWrapper_191_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_192 ( // @[package.scala 93:22:@20928.4]
    .clock(RetimeWrapper_192_clock),
    .reset(RetimeWrapper_192_reset),
    .io_flow(RetimeWrapper_192_io_flow),
    .io_in(RetimeWrapper_192_io_in),
    .io_out(RetimeWrapper_192_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_193 ( // @[package.scala 93:22:@20936.4]
    .clock(RetimeWrapper_193_clock),
    .reset(RetimeWrapper_193_reset),
    .io_flow(RetimeWrapper_193_io_flow),
    .io_in(RetimeWrapper_193_io_in),
    .io_out(RetimeWrapper_193_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_194 ( // @[package.scala 93:22:@20944.4]
    .clock(RetimeWrapper_194_clock),
    .reset(RetimeWrapper_194_reset),
    .io_flow(RetimeWrapper_194_io_flow),
    .io_in(RetimeWrapper_194_io_in),
    .io_out(RetimeWrapper_194_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_195 ( // @[package.scala 93:22:@20952.4]
    .clock(RetimeWrapper_195_clock),
    .reset(RetimeWrapper_195_reset),
    .io_flow(RetimeWrapper_195_io_flow),
    .io_in(RetimeWrapper_195_io_in),
    .io_out(RetimeWrapper_195_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_196 ( // @[package.scala 93:22:@20960.4]
    .clock(RetimeWrapper_196_clock),
    .reset(RetimeWrapper_196_reset),
    .io_flow(RetimeWrapper_196_io_flow),
    .io_in(RetimeWrapper_196_io_in),
    .io_out(RetimeWrapper_196_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_197 ( // @[package.scala 93:22:@20968.4]
    .clock(RetimeWrapper_197_clock),
    .reset(RetimeWrapper_197_reset),
    .io_flow(RetimeWrapper_197_io_flow),
    .io_in(RetimeWrapper_197_io_in),
    .io_out(RetimeWrapper_197_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_198 ( // @[package.scala 93:22:@20976.4]
    .clock(RetimeWrapper_198_clock),
    .reset(RetimeWrapper_198_reset),
    .io_flow(RetimeWrapper_198_io_flow),
    .io_in(RetimeWrapper_198_io_in),
    .io_out(RetimeWrapper_198_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_199 ( // @[package.scala 93:22:@20984.4]
    .clock(RetimeWrapper_199_clock),
    .reset(RetimeWrapper_199_reset),
    .io_flow(RetimeWrapper_199_io_flow),
    .io_in(RetimeWrapper_199_io_in),
    .io_out(RetimeWrapper_199_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_200 ( // @[package.scala 93:22:@20992.4]
    .clock(RetimeWrapper_200_clock),
    .reset(RetimeWrapper_200_reset),
    .io_flow(RetimeWrapper_200_io_flow),
    .io_in(RetimeWrapper_200_io_in),
    .io_out(RetimeWrapper_200_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_201 ( // @[package.scala 93:22:@21000.4]
    .clock(RetimeWrapper_201_clock),
    .reset(RetimeWrapper_201_reset),
    .io_flow(RetimeWrapper_201_io_flow),
    .io_in(RetimeWrapper_201_io_in),
    .io_out(RetimeWrapper_201_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_202 ( // @[package.scala 93:22:@21008.4]
    .clock(RetimeWrapper_202_clock),
    .reset(RetimeWrapper_202_reset),
    .io_flow(RetimeWrapper_202_io_flow),
    .io_in(RetimeWrapper_202_io_in),
    .io_out(RetimeWrapper_202_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_203 ( // @[package.scala 93:22:@21016.4]
    .clock(RetimeWrapper_203_clock),
    .reset(RetimeWrapper_203_reset),
    .io_flow(RetimeWrapper_203_io_flow),
    .io_in(RetimeWrapper_203_io_in),
    .io_out(RetimeWrapper_203_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_204 ( // @[package.scala 93:22:@21072.4]
    .clock(RetimeWrapper_204_clock),
    .reset(RetimeWrapper_204_reset),
    .io_flow(RetimeWrapper_204_io_flow),
    .io_in(RetimeWrapper_204_io_in),
    .io_out(RetimeWrapper_204_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_205 ( // @[package.scala 93:22:@21080.4]
    .clock(RetimeWrapper_205_clock),
    .reset(RetimeWrapper_205_reset),
    .io_flow(RetimeWrapper_205_io_flow),
    .io_in(RetimeWrapper_205_io_in),
    .io_out(RetimeWrapper_205_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_206 ( // @[package.scala 93:22:@21088.4]
    .clock(RetimeWrapper_206_clock),
    .reset(RetimeWrapper_206_reset),
    .io_flow(RetimeWrapper_206_io_flow),
    .io_in(RetimeWrapper_206_io_in),
    .io_out(RetimeWrapper_206_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_207 ( // @[package.scala 93:22:@21096.4]
    .clock(RetimeWrapper_207_clock),
    .reset(RetimeWrapper_207_reset),
    .io_flow(RetimeWrapper_207_io_flow),
    .io_in(RetimeWrapper_207_io_in),
    .io_out(RetimeWrapper_207_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_208 ( // @[package.scala 93:22:@21104.4]
    .clock(RetimeWrapper_208_clock),
    .reset(RetimeWrapper_208_reset),
    .io_flow(RetimeWrapper_208_io_flow),
    .io_in(RetimeWrapper_208_io_in),
    .io_out(RetimeWrapper_208_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_209 ( // @[package.scala 93:22:@21112.4]
    .clock(RetimeWrapper_209_clock),
    .reset(RetimeWrapper_209_reset),
    .io_flow(RetimeWrapper_209_io_flow),
    .io_in(RetimeWrapper_209_io_in),
    .io_out(RetimeWrapper_209_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_210 ( // @[package.scala 93:22:@21120.4]
    .clock(RetimeWrapper_210_clock),
    .reset(RetimeWrapper_210_reset),
    .io_flow(RetimeWrapper_210_io_flow),
    .io_in(RetimeWrapper_210_io_in),
    .io_out(RetimeWrapper_210_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_211 ( // @[package.scala 93:22:@21128.4]
    .clock(RetimeWrapper_211_clock),
    .reset(RetimeWrapper_211_reset),
    .io_flow(RetimeWrapper_211_io_flow),
    .io_in(RetimeWrapper_211_io_in),
    .io_out(RetimeWrapper_211_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_212 ( // @[package.scala 93:22:@21136.4]
    .clock(RetimeWrapper_212_clock),
    .reset(RetimeWrapper_212_reset),
    .io_flow(RetimeWrapper_212_io_flow),
    .io_in(RetimeWrapper_212_io_in),
    .io_out(RetimeWrapper_212_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_213 ( // @[package.scala 93:22:@21144.4]
    .clock(RetimeWrapper_213_clock),
    .reset(RetimeWrapper_213_reset),
    .io_flow(RetimeWrapper_213_io_flow),
    .io_in(RetimeWrapper_213_io_in),
    .io_out(RetimeWrapper_213_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_214 ( // @[package.scala 93:22:@21152.4]
    .clock(RetimeWrapper_214_clock),
    .reset(RetimeWrapper_214_reset),
    .io_flow(RetimeWrapper_214_io_flow),
    .io_in(RetimeWrapper_214_io_in),
    .io_out(RetimeWrapper_214_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_215 ( // @[package.scala 93:22:@21160.4]
    .clock(RetimeWrapper_215_clock),
    .reset(RetimeWrapper_215_reset),
    .io_flow(RetimeWrapper_215_io_flow),
    .io_in(RetimeWrapper_215_io_in),
    .io_out(RetimeWrapper_215_io_out)
  );
  assign _T_700 = io_wPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@15995.4]
  assign _T_702 = io_wPort_0_banks_1 == 3'h0; // @[MemPrimitives.scala 82:210:@15996.4]
  assign _T_703 = _T_700 & _T_702; // @[MemPrimitives.scala 82:228:@15997.4]
  assign _T_704 = io_wPort_0_en_0 & _T_703; // @[MemPrimitives.scala 83:102:@15998.4]
  assign _T_706 = io_wPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@15999.4]
  assign _T_708 = io_wPort_2_banks_1 == 3'h0; // @[MemPrimitives.scala 82:210:@16000.4]
  assign _T_709 = _T_706 & _T_708; // @[MemPrimitives.scala 82:228:@16001.4]
  assign _T_710 = io_wPort_2_en_0 & _T_709; // @[MemPrimitives.scala 83:102:@16002.4]
  assign _T_712 = {_T_704,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@16004.4]
  assign _T_714 = {_T_710,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@16006.4]
  assign _T_715 = _T_704 ? _T_712 : _T_714; // @[Mux.scala 31:69:@16007.4]
  assign _T_720 = io_wPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@16014.4]
  assign _T_722 = io_wPort_1_banks_1 == 3'h1; // @[MemPrimitives.scala 82:210:@16015.4]
  assign _T_723 = _T_720 & _T_722; // @[MemPrimitives.scala 82:228:@16016.4]
  assign _T_724 = io_wPort_1_en_0 & _T_723; // @[MemPrimitives.scala 83:102:@16017.4]
  assign _T_726 = io_wPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@16018.4]
  assign _T_728 = io_wPort_3_banks_1 == 3'h1; // @[MemPrimitives.scala 82:210:@16019.4]
  assign _T_729 = _T_726 & _T_728; // @[MemPrimitives.scala 82:228:@16020.4]
  assign _T_730 = io_wPort_3_en_0 & _T_729; // @[MemPrimitives.scala 83:102:@16021.4]
  assign _T_732 = {_T_724,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@16023.4]
  assign _T_734 = {_T_730,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@16025.4]
  assign _T_735 = _T_724 ? _T_732 : _T_734; // @[Mux.scala 31:69:@16026.4]
  assign _T_742 = io_wPort_0_banks_1 == 3'h2; // @[MemPrimitives.scala 82:210:@16034.4]
  assign _T_743 = _T_700 & _T_742; // @[MemPrimitives.scala 82:228:@16035.4]
  assign _T_744 = io_wPort_0_en_0 & _T_743; // @[MemPrimitives.scala 83:102:@16036.4]
  assign _T_748 = io_wPort_2_banks_1 == 3'h2; // @[MemPrimitives.scala 82:210:@16038.4]
  assign _T_749 = _T_706 & _T_748; // @[MemPrimitives.scala 82:228:@16039.4]
  assign _T_750 = io_wPort_2_en_0 & _T_749; // @[MemPrimitives.scala 83:102:@16040.4]
  assign _T_752 = {_T_744,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@16042.4]
  assign _T_754 = {_T_750,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@16044.4]
  assign _T_755 = _T_744 ? _T_752 : _T_754; // @[Mux.scala 31:69:@16045.4]
  assign _T_762 = io_wPort_1_banks_1 == 3'h3; // @[MemPrimitives.scala 82:210:@16053.4]
  assign _T_763 = _T_720 & _T_762; // @[MemPrimitives.scala 82:228:@16054.4]
  assign _T_764 = io_wPort_1_en_0 & _T_763; // @[MemPrimitives.scala 83:102:@16055.4]
  assign _T_768 = io_wPort_3_banks_1 == 3'h3; // @[MemPrimitives.scala 82:210:@16057.4]
  assign _T_769 = _T_726 & _T_768; // @[MemPrimitives.scala 82:228:@16058.4]
  assign _T_770 = io_wPort_3_en_0 & _T_769; // @[MemPrimitives.scala 83:102:@16059.4]
  assign _T_772 = {_T_764,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@16061.4]
  assign _T_774 = {_T_770,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@16063.4]
  assign _T_775 = _T_764 ? _T_772 : _T_774; // @[Mux.scala 31:69:@16064.4]
  assign _T_782 = io_wPort_0_banks_1 == 3'h4; // @[MemPrimitives.scala 82:210:@16072.4]
  assign _T_783 = _T_700 & _T_782; // @[MemPrimitives.scala 82:228:@16073.4]
  assign _T_784 = io_wPort_0_en_0 & _T_783; // @[MemPrimitives.scala 83:102:@16074.4]
  assign _T_788 = io_wPort_2_banks_1 == 3'h4; // @[MemPrimitives.scala 82:210:@16076.4]
  assign _T_789 = _T_706 & _T_788; // @[MemPrimitives.scala 82:228:@16077.4]
  assign _T_790 = io_wPort_2_en_0 & _T_789; // @[MemPrimitives.scala 83:102:@16078.4]
  assign _T_792 = {_T_784,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@16080.4]
  assign _T_794 = {_T_790,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@16082.4]
  assign _T_795 = _T_784 ? _T_792 : _T_794; // @[Mux.scala 31:69:@16083.4]
  assign _T_802 = io_wPort_1_banks_1 == 3'h5; // @[MemPrimitives.scala 82:210:@16091.4]
  assign _T_803 = _T_720 & _T_802; // @[MemPrimitives.scala 82:228:@16092.4]
  assign _T_804 = io_wPort_1_en_0 & _T_803; // @[MemPrimitives.scala 83:102:@16093.4]
  assign _T_808 = io_wPort_3_banks_1 == 3'h5; // @[MemPrimitives.scala 82:210:@16095.4]
  assign _T_809 = _T_726 & _T_808; // @[MemPrimitives.scala 82:228:@16096.4]
  assign _T_810 = io_wPort_3_en_0 & _T_809; // @[MemPrimitives.scala 83:102:@16097.4]
  assign _T_812 = {_T_804,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@16099.4]
  assign _T_814 = {_T_810,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@16101.4]
  assign _T_815 = _T_804 ? _T_812 : _T_814; // @[Mux.scala 31:69:@16102.4]
  assign _T_820 = io_wPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@16109.4]
  assign _T_823 = _T_820 & _T_702; // @[MemPrimitives.scala 82:228:@16111.4]
  assign _T_824 = io_wPort_0_en_0 & _T_823; // @[MemPrimitives.scala 83:102:@16112.4]
  assign _T_826 = io_wPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@16113.4]
  assign _T_829 = _T_826 & _T_708; // @[MemPrimitives.scala 82:228:@16115.4]
  assign _T_830 = io_wPort_2_en_0 & _T_829; // @[MemPrimitives.scala 83:102:@16116.4]
  assign _T_832 = {_T_824,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@16118.4]
  assign _T_834 = {_T_830,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@16120.4]
  assign _T_835 = _T_824 ? _T_832 : _T_834; // @[Mux.scala 31:69:@16121.4]
  assign _T_840 = io_wPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@16128.4]
  assign _T_843 = _T_840 & _T_722; // @[MemPrimitives.scala 82:228:@16130.4]
  assign _T_844 = io_wPort_1_en_0 & _T_843; // @[MemPrimitives.scala 83:102:@16131.4]
  assign _T_846 = io_wPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@16132.4]
  assign _T_849 = _T_846 & _T_728; // @[MemPrimitives.scala 82:228:@16134.4]
  assign _T_850 = io_wPort_3_en_0 & _T_849; // @[MemPrimitives.scala 83:102:@16135.4]
  assign _T_852 = {_T_844,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@16137.4]
  assign _T_854 = {_T_850,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@16139.4]
  assign _T_855 = _T_844 ? _T_852 : _T_854; // @[Mux.scala 31:69:@16140.4]
  assign _T_863 = _T_820 & _T_742; // @[MemPrimitives.scala 82:228:@16149.4]
  assign _T_864 = io_wPort_0_en_0 & _T_863; // @[MemPrimitives.scala 83:102:@16150.4]
  assign _T_869 = _T_826 & _T_748; // @[MemPrimitives.scala 82:228:@16153.4]
  assign _T_870 = io_wPort_2_en_0 & _T_869; // @[MemPrimitives.scala 83:102:@16154.4]
  assign _T_872 = {_T_864,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@16156.4]
  assign _T_874 = {_T_870,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@16158.4]
  assign _T_875 = _T_864 ? _T_872 : _T_874; // @[Mux.scala 31:69:@16159.4]
  assign _T_883 = _T_840 & _T_762; // @[MemPrimitives.scala 82:228:@16168.4]
  assign _T_884 = io_wPort_1_en_0 & _T_883; // @[MemPrimitives.scala 83:102:@16169.4]
  assign _T_889 = _T_846 & _T_768; // @[MemPrimitives.scala 82:228:@16172.4]
  assign _T_890 = io_wPort_3_en_0 & _T_889; // @[MemPrimitives.scala 83:102:@16173.4]
  assign _T_892 = {_T_884,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@16175.4]
  assign _T_894 = {_T_890,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@16177.4]
  assign _T_895 = _T_884 ? _T_892 : _T_894; // @[Mux.scala 31:69:@16178.4]
  assign _T_903 = _T_820 & _T_782; // @[MemPrimitives.scala 82:228:@16187.4]
  assign _T_904 = io_wPort_0_en_0 & _T_903; // @[MemPrimitives.scala 83:102:@16188.4]
  assign _T_909 = _T_826 & _T_788; // @[MemPrimitives.scala 82:228:@16191.4]
  assign _T_910 = io_wPort_2_en_0 & _T_909; // @[MemPrimitives.scala 83:102:@16192.4]
  assign _T_912 = {_T_904,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@16194.4]
  assign _T_914 = {_T_910,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@16196.4]
  assign _T_915 = _T_904 ? _T_912 : _T_914; // @[Mux.scala 31:69:@16197.4]
  assign _T_923 = _T_840 & _T_802; // @[MemPrimitives.scala 82:228:@16206.4]
  assign _T_924 = io_wPort_1_en_0 & _T_923; // @[MemPrimitives.scala 83:102:@16207.4]
  assign _T_929 = _T_846 & _T_808; // @[MemPrimitives.scala 82:228:@16210.4]
  assign _T_930 = io_wPort_3_en_0 & _T_929; // @[MemPrimitives.scala 83:102:@16211.4]
  assign _T_932 = {_T_924,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@16213.4]
  assign _T_934 = {_T_930,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@16215.4]
  assign _T_935 = _T_924 ? _T_932 : _T_934; // @[Mux.scala 31:69:@16216.4]
  assign _T_940 = io_wPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@16223.4]
  assign _T_943 = _T_940 & _T_702; // @[MemPrimitives.scala 82:228:@16225.4]
  assign _T_944 = io_wPort_0_en_0 & _T_943; // @[MemPrimitives.scala 83:102:@16226.4]
  assign _T_946 = io_wPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@16227.4]
  assign _T_949 = _T_946 & _T_708; // @[MemPrimitives.scala 82:228:@16229.4]
  assign _T_950 = io_wPort_2_en_0 & _T_949; // @[MemPrimitives.scala 83:102:@16230.4]
  assign _T_952 = {_T_944,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@16232.4]
  assign _T_954 = {_T_950,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@16234.4]
  assign _T_955 = _T_944 ? _T_952 : _T_954; // @[Mux.scala 31:69:@16235.4]
  assign _T_960 = io_wPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@16242.4]
  assign _T_963 = _T_960 & _T_722; // @[MemPrimitives.scala 82:228:@16244.4]
  assign _T_964 = io_wPort_1_en_0 & _T_963; // @[MemPrimitives.scala 83:102:@16245.4]
  assign _T_966 = io_wPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@16246.4]
  assign _T_969 = _T_966 & _T_728; // @[MemPrimitives.scala 82:228:@16248.4]
  assign _T_970 = io_wPort_3_en_0 & _T_969; // @[MemPrimitives.scala 83:102:@16249.4]
  assign _T_972 = {_T_964,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@16251.4]
  assign _T_974 = {_T_970,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@16253.4]
  assign _T_975 = _T_964 ? _T_972 : _T_974; // @[Mux.scala 31:69:@16254.4]
  assign _T_983 = _T_940 & _T_742; // @[MemPrimitives.scala 82:228:@16263.4]
  assign _T_984 = io_wPort_0_en_0 & _T_983; // @[MemPrimitives.scala 83:102:@16264.4]
  assign _T_989 = _T_946 & _T_748; // @[MemPrimitives.scala 82:228:@16267.4]
  assign _T_990 = io_wPort_2_en_0 & _T_989; // @[MemPrimitives.scala 83:102:@16268.4]
  assign _T_992 = {_T_984,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@16270.4]
  assign _T_994 = {_T_990,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@16272.4]
  assign _T_995 = _T_984 ? _T_992 : _T_994; // @[Mux.scala 31:69:@16273.4]
  assign _T_1003 = _T_960 & _T_762; // @[MemPrimitives.scala 82:228:@16282.4]
  assign _T_1004 = io_wPort_1_en_0 & _T_1003; // @[MemPrimitives.scala 83:102:@16283.4]
  assign _T_1009 = _T_966 & _T_768; // @[MemPrimitives.scala 82:228:@16286.4]
  assign _T_1010 = io_wPort_3_en_0 & _T_1009; // @[MemPrimitives.scala 83:102:@16287.4]
  assign _T_1012 = {_T_1004,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@16289.4]
  assign _T_1014 = {_T_1010,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@16291.4]
  assign _T_1015 = _T_1004 ? _T_1012 : _T_1014; // @[Mux.scala 31:69:@16292.4]
  assign _T_1023 = _T_940 & _T_782; // @[MemPrimitives.scala 82:228:@16301.4]
  assign _T_1024 = io_wPort_0_en_0 & _T_1023; // @[MemPrimitives.scala 83:102:@16302.4]
  assign _T_1029 = _T_946 & _T_788; // @[MemPrimitives.scala 82:228:@16305.4]
  assign _T_1030 = io_wPort_2_en_0 & _T_1029; // @[MemPrimitives.scala 83:102:@16306.4]
  assign _T_1032 = {_T_1024,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@16308.4]
  assign _T_1034 = {_T_1030,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@16310.4]
  assign _T_1035 = _T_1024 ? _T_1032 : _T_1034; // @[Mux.scala 31:69:@16311.4]
  assign _T_1043 = _T_960 & _T_802; // @[MemPrimitives.scala 82:228:@16320.4]
  assign _T_1044 = io_wPort_1_en_0 & _T_1043; // @[MemPrimitives.scala 83:102:@16321.4]
  assign _T_1049 = _T_966 & _T_808; // @[MemPrimitives.scala 82:228:@16324.4]
  assign _T_1050 = io_wPort_3_en_0 & _T_1049; // @[MemPrimitives.scala 83:102:@16325.4]
  assign _T_1052 = {_T_1044,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@16327.4]
  assign _T_1054 = {_T_1050,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@16329.4]
  assign _T_1055 = _T_1044 ? _T_1052 : _T_1054; // @[Mux.scala 31:69:@16330.4]
  assign _T_1060 = io_wPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@16337.4]
  assign _T_1063 = _T_1060 & _T_702; // @[MemPrimitives.scala 82:228:@16339.4]
  assign _T_1064 = io_wPort_0_en_0 & _T_1063; // @[MemPrimitives.scala 83:102:@16340.4]
  assign _T_1066 = io_wPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@16341.4]
  assign _T_1069 = _T_1066 & _T_708; // @[MemPrimitives.scala 82:228:@16343.4]
  assign _T_1070 = io_wPort_2_en_0 & _T_1069; // @[MemPrimitives.scala 83:102:@16344.4]
  assign _T_1072 = {_T_1064,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@16346.4]
  assign _T_1074 = {_T_1070,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@16348.4]
  assign _T_1075 = _T_1064 ? _T_1072 : _T_1074; // @[Mux.scala 31:69:@16349.4]
  assign _T_1080 = io_wPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@16356.4]
  assign _T_1083 = _T_1080 & _T_722; // @[MemPrimitives.scala 82:228:@16358.4]
  assign _T_1084 = io_wPort_1_en_0 & _T_1083; // @[MemPrimitives.scala 83:102:@16359.4]
  assign _T_1086 = io_wPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@16360.4]
  assign _T_1089 = _T_1086 & _T_728; // @[MemPrimitives.scala 82:228:@16362.4]
  assign _T_1090 = io_wPort_3_en_0 & _T_1089; // @[MemPrimitives.scala 83:102:@16363.4]
  assign _T_1092 = {_T_1084,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@16365.4]
  assign _T_1094 = {_T_1090,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@16367.4]
  assign _T_1095 = _T_1084 ? _T_1092 : _T_1094; // @[Mux.scala 31:69:@16368.4]
  assign _T_1103 = _T_1060 & _T_742; // @[MemPrimitives.scala 82:228:@16377.4]
  assign _T_1104 = io_wPort_0_en_0 & _T_1103; // @[MemPrimitives.scala 83:102:@16378.4]
  assign _T_1109 = _T_1066 & _T_748; // @[MemPrimitives.scala 82:228:@16381.4]
  assign _T_1110 = io_wPort_2_en_0 & _T_1109; // @[MemPrimitives.scala 83:102:@16382.4]
  assign _T_1112 = {_T_1104,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@16384.4]
  assign _T_1114 = {_T_1110,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@16386.4]
  assign _T_1115 = _T_1104 ? _T_1112 : _T_1114; // @[Mux.scala 31:69:@16387.4]
  assign _T_1123 = _T_1080 & _T_762; // @[MemPrimitives.scala 82:228:@16396.4]
  assign _T_1124 = io_wPort_1_en_0 & _T_1123; // @[MemPrimitives.scala 83:102:@16397.4]
  assign _T_1129 = _T_1086 & _T_768; // @[MemPrimitives.scala 82:228:@16400.4]
  assign _T_1130 = io_wPort_3_en_0 & _T_1129; // @[MemPrimitives.scala 83:102:@16401.4]
  assign _T_1132 = {_T_1124,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@16403.4]
  assign _T_1134 = {_T_1130,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@16405.4]
  assign _T_1135 = _T_1124 ? _T_1132 : _T_1134; // @[Mux.scala 31:69:@16406.4]
  assign _T_1143 = _T_1060 & _T_782; // @[MemPrimitives.scala 82:228:@16415.4]
  assign _T_1144 = io_wPort_0_en_0 & _T_1143; // @[MemPrimitives.scala 83:102:@16416.4]
  assign _T_1149 = _T_1066 & _T_788; // @[MemPrimitives.scala 82:228:@16419.4]
  assign _T_1150 = io_wPort_2_en_0 & _T_1149; // @[MemPrimitives.scala 83:102:@16420.4]
  assign _T_1152 = {_T_1144,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@16422.4]
  assign _T_1154 = {_T_1150,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@16424.4]
  assign _T_1155 = _T_1144 ? _T_1152 : _T_1154; // @[Mux.scala 31:69:@16425.4]
  assign _T_1163 = _T_1080 & _T_802; // @[MemPrimitives.scala 82:228:@16434.4]
  assign _T_1164 = io_wPort_1_en_0 & _T_1163; // @[MemPrimitives.scala 83:102:@16435.4]
  assign _T_1169 = _T_1086 & _T_808; // @[MemPrimitives.scala 82:228:@16438.4]
  assign _T_1170 = io_wPort_3_en_0 & _T_1169; // @[MemPrimitives.scala 83:102:@16439.4]
  assign _T_1172 = {_T_1164,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@16441.4]
  assign _T_1174 = {_T_1170,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@16443.4]
  assign _T_1175 = _T_1164 ? _T_1172 : _T_1174; // @[Mux.scala 31:69:@16444.4]
  assign _T_1180 = io_rPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@16451.4]
  assign _T_1182 = io_rPort_0_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@16452.4]
  assign _T_1183 = _T_1180 & _T_1182; // @[MemPrimitives.scala 110:228:@16453.4]
  assign _T_1186 = io_rPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@16455.4]
  assign _T_1188 = io_rPort_1_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@16456.4]
  assign _T_1189 = _T_1186 & _T_1188; // @[MemPrimitives.scala 110:228:@16457.4]
  assign _T_1192 = io_rPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@16459.4]
  assign _T_1194 = io_rPort_3_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@16460.4]
  assign _T_1195 = _T_1192 & _T_1194; // @[MemPrimitives.scala 110:228:@16461.4]
  assign _T_1198 = io_rPort_4_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@16463.4]
  assign _T_1200 = io_rPort_4_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@16464.4]
  assign _T_1201 = _T_1198 & _T_1200; // @[MemPrimitives.scala 110:228:@16465.4]
  assign _T_1204 = io_rPort_8_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@16467.4]
  assign _T_1206 = io_rPort_8_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@16468.4]
  assign _T_1207 = _T_1204 & _T_1206; // @[MemPrimitives.scala 110:228:@16469.4]
  assign _T_1210 = io_rPort_10_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@16471.4]
  assign _T_1212 = io_rPort_10_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@16472.4]
  assign _T_1213 = _T_1210 & _T_1212; // @[MemPrimitives.scala 110:228:@16473.4]
  assign _T_1216 = io_rPort_14_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@16475.4]
  assign _T_1218 = io_rPort_14_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@16476.4]
  assign _T_1219 = _T_1216 & _T_1218; // @[MemPrimitives.scala 110:228:@16477.4]
  assign _T_1222 = io_rPort_15_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@16479.4]
  assign _T_1224 = io_rPort_15_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@16480.4]
  assign _T_1225 = _T_1222 & _T_1224; // @[MemPrimitives.scala 110:228:@16481.4]
  assign _T_1228 = io_rPort_17_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@16483.4]
  assign _T_1230 = io_rPort_17_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@16484.4]
  assign _T_1231 = _T_1228 & _T_1230; // @[MemPrimitives.scala 110:228:@16485.4]
  assign _T_1233 = StickySelects_io_outs_0; // @[MemPrimitives.scala 123:41:@16499.4]
  assign _T_1234 = StickySelects_io_outs_1; // @[MemPrimitives.scala 123:41:@16500.4]
  assign _T_1235 = StickySelects_io_outs_2; // @[MemPrimitives.scala 123:41:@16501.4]
  assign _T_1236 = StickySelects_io_outs_3; // @[MemPrimitives.scala 123:41:@16502.4]
  assign _T_1237 = StickySelects_io_outs_4; // @[MemPrimitives.scala 123:41:@16503.4]
  assign _T_1238 = StickySelects_io_outs_5; // @[MemPrimitives.scala 123:41:@16504.4]
  assign _T_1239 = StickySelects_io_outs_6; // @[MemPrimitives.scala 123:41:@16505.4]
  assign _T_1240 = StickySelects_io_outs_7; // @[MemPrimitives.scala 123:41:@16506.4]
  assign _T_1241 = StickySelects_io_outs_8; // @[MemPrimitives.scala 123:41:@16507.4]
  assign _T_1243 = {_T_1233,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@16509.4]
  assign _T_1245 = {_T_1234,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@16511.4]
  assign _T_1247 = {_T_1235,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@16513.4]
  assign _T_1249 = {_T_1236,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@16515.4]
  assign _T_1251 = {_T_1237,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@16517.4]
  assign _T_1253 = {_T_1238,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@16519.4]
  assign _T_1255 = {_T_1239,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@16521.4]
  assign _T_1257 = {_T_1240,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@16523.4]
  assign _T_1259 = {_T_1241,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@16525.4]
  assign _T_1260 = _T_1240 ? _T_1257 : _T_1259; // @[Mux.scala 31:69:@16526.4]
  assign _T_1261 = _T_1239 ? _T_1255 : _T_1260; // @[Mux.scala 31:69:@16527.4]
  assign _T_1262 = _T_1238 ? _T_1253 : _T_1261; // @[Mux.scala 31:69:@16528.4]
  assign _T_1263 = _T_1237 ? _T_1251 : _T_1262; // @[Mux.scala 31:69:@16529.4]
  assign _T_1264 = _T_1236 ? _T_1249 : _T_1263; // @[Mux.scala 31:69:@16530.4]
  assign _T_1265 = _T_1235 ? _T_1247 : _T_1264; // @[Mux.scala 31:69:@16531.4]
  assign _T_1266 = _T_1234 ? _T_1245 : _T_1265; // @[Mux.scala 31:69:@16532.4]
  assign _T_1267 = _T_1233 ? _T_1243 : _T_1266; // @[Mux.scala 31:69:@16533.4]
  assign _T_1272 = io_rPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@16540.4]
  assign _T_1274 = io_rPort_2_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@16541.4]
  assign _T_1275 = _T_1272 & _T_1274; // @[MemPrimitives.scala 110:228:@16542.4]
  assign _T_1278 = io_rPort_5_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@16544.4]
  assign _T_1280 = io_rPort_5_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@16545.4]
  assign _T_1281 = _T_1278 & _T_1280; // @[MemPrimitives.scala 110:228:@16546.4]
  assign _T_1284 = io_rPort_6_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@16548.4]
  assign _T_1286 = io_rPort_6_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@16549.4]
  assign _T_1287 = _T_1284 & _T_1286; // @[MemPrimitives.scala 110:228:@16550.4]
  assign _T_1290 = io_rPort_7_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@16552.4]
  assign _T_1292 = io_rPort_7_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@16553.4]
  assign _T_1293 = _T_1290 & _T_1292; // @[MemPrimitives.scala 110:228:@16554.4]
  assign _T_1296 = io_rPort_9_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@16556.4]
  assign _T_1298 = io_rPort_9_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@16557.4]
  assign _T_1299 = _T_1296 & _T_1298; // @[MemPrimitives.scala 110:228:@16558.4]
  assign _T_1302 = io_rPort_11_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@16560.4]
  assign _T_1304 = io_rPort_11_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@16561.4]
  assign _T_1305 = _T_1302 & _T_1304; // @[MemPrimitives.scala 110:228:@16562.4]
  assign _T_1308 = io_rPort_12_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@16564.4]
  assign _T_1310 = io_rPort_12_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@16565.4]
  assign _T_1311 = _T_1308 & _T_1310; // @[MemPrimitives.scala 110:228:@16566.4]
  assign _T_1314 = io_rPort_13_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@16568.4]
  assign _T_1316 = io_rPort_13_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@16569.4]
  assign _T_1317 = _T_1314 & _T_1316; // @[MemPrimitives.scala 110:228:@16570.4]
  assign _T_1320 = io_rPort_16_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@16572.4]
  assign _T_1322 = io_rPort_16_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@16573.4]
  assign _T_1323 = _T_1320 & _T_1322; // @[MemPrimitives.scala 110:228:@16574.4]
  assign _T_1325 = StickySelects_1_io_outs_0; // @[MemPrimitives.scala 123:41:@16588.4]
  assign _T_1326 = StickySelects_1_io_outs_1; // @[MemPrimitives.scala 123:41:@16589.4]
  assign _T_1327 = StickySelects_1_io_outs_2; // @[MemPrimitives.scala 123:41:@16590.4]
  assign _T_1328 = StickySelects_1_io_outs_3; // @[MemPrimitives.scala 123:41:@16591.4]
  assign _T_1329 = StickySelects_1_io_outs_4; // @[MemPrimitives.scala 123:41:@16592.4]
  assign _T_1330 = StickySelects_1_io_outs_5; // @[MemPrimitives.scala 123:41:@16593.4]
  assign _T_1331 = StickySelects_1_io_outs_6; // @[MemPrimitives.scala 123:41:@16594.4]
  assign _T_1332 = StickySelects_1_io_outs_7; // @[MemPrimitives.scala 123:41:@16595.4]
  assign _T_1333 = StickySelects_1_io_outs_8; // @[MemPrimitives.scala 123:41:@16596.4]
  assign _T_1335 = {_T_1325,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@16598.4]
  assign _T_1337 = {_T_1326,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@16600.4]
  assign _T_1339 = {_T_1327,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@16602.4]
  assign _T_1341 = {_T_1328,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@16604.4]
  assign _T_1343 = {_T_1329,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@16606.4]
  assign _T_1345 = {_T_1330,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@16608.4]
  assign _T_1347 = {_T_1331,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@16610.4]
  assign _T_1349 = {_T_1332,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@16612.4]
  assign _T_1351 = {_T_1333,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@16614.4]
  assign _T_1352 = _T_1332 ? _T_1349 : _T_1351; // @[Mux.scala 31:69:@16615.4]
  assign _T_1353 = _T_1331 ? _T_1347 : _T_1352; // @[Mux.scala 31:69:@16616.4]
  assign _T_1354 = _T_1330 ? _T_1345 : _T_1353; // @[Mux.scala 31:69:@16617.4]
  assign _T_1355 = _T_1329 ? _T_1343 : _T_1354; // @[Mux.scala 31:69:@16618.4]
  assign _T_1356 = _T_1328 ? _T_1341 : _T_1355; // @[Mux.scala 31:69:@16619.4]
  assign _T_1357 = _T_1327 ? _T_1339 : _T_1356; // @[Mux.scala 31:69:@16620.4]
  assign _T_1358 = _T_1326 ? _T_1337 : _T_1357; // @[Mux.scala 31:69:@16621.4]
  assign _T_1359 = _T_1325 ? _T_1335 : _T_1358; // @[Mux.scala 31:69:@16622.4]
  assign _T_1366 = io_rPort_0_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@16630.4]
  assign _T_1367 = _T_1180 & _T_1366; // @[MemPrimitives.scala 110:228:@16631.4]
  assign _T_1372 = io_rPort_1_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@16634.4]
  assign _T_1373 = _T_1186 & _T_1372; // @[MemPrimitives.scala 110:228:@16635.4]
  assign _T_1378 = io_rPort_3_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@16638.4]
  assign _T_1379 = _T_1192 & _T_1378; // @[MemPrimitives.scala 110:228:@16639.4]
  assign _T_1384 = io_rPort_4_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@16642.4]
  assign _T_1385 = _T_1198 & _T_1384; // @[MemPrimitives.scala 110:228:@16643.4]
  assign _T_1390 = io_rPort_8_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@16646.4]
  assign _T_1391 = _T_1204 & _T_1390; // @[MemPrimitives.scala 110:228:@16647.4]
  assign _T_1396 = io_rPort_10_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@16650.4]
  assign _T_1397 = _T_1210 & _T_1396; // @[MemPrimitives.scala 110:228:@16651.4]
  assign _T_1402 = io_rPort_14_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@16654.4]
  assign _T_1403 = _T_1216 & _T_1402; // @[MemPrimitives.scala 110:228:@16655.4]
  assign _T_1408 = io_rPort_15_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@16658.4]
  assign _T_1409 = _T_1222 & _T_1408; // @[MemPrimitives.scala 110:228:@16659.4]
  assign _T_1414 = io_rPort_17_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@16662.4]
  assign _T_1415 = _T_1228 & _T_1414; // @[MemPrimitives.scala 110:228:@16663.4]
  assign _T_1417 = StickySelects_2_io_outs_0; // @[MemPrimitives.scala 123:41:@16677.4]
  assign _T_1418 = StickySelects_2_io_outs_1; // @[MemPrimitives.scala 123:41:@16678.4]
  assign _T_1419 = StickySelects_2_io_outs_2; // @[MemPrimitives.scala 123:41:@16679.4]
  assign _T_1420 = StickySelects_2_io_outs_3; // @[MemPrimitives.scala 123:41:@16680.4]
  assign _T_1421 = StickySelects_2_io_outs_4; // @[MemPrimitives.scala 123:41:@16681.4]
  assign _T_1422 = StickySelects_2_io_outs_5; // @[MemPrimitives.scala 123:41:@16682.4]
  assign _T_1423 = StickySelects_2_io_outs_6; // @[MemPrimitives.scala 123:41:@16683.4]
  assign _T_1424 = StickySelects_2_io_outs_7; // @[MemPrimitives.scala 123:41:@16684.4]
  assign _T_1425 = StickySelects_2_io_outs_8; // @[MemPrimitives.scala 123:41:@16685.4]
  assign _T_1427 = {_T_1417,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@16687.4]
  assign _T_1429 = {_T_1418,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@16689.4]
  assign _T_1431 = {_T_1419,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@16691.4]
  assign _T_1433 = {_T_1420,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@16693.4]
  assign _T_1435 = {_T_1421,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@16695.4]
  assign _T_1437 = {_T_1422,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@16697.4]
  assign _T_1439 = {_T_1423,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@16699.4]
  assign _T_1441 = {_T_1424,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@16701.4]
  assign _T_1443 = {_T_1425,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@16703.4]
  assign _T_1444 = _T_1424 ? _T_1441 : _T_1443; // @[Mux.scala 31:69:@16704.4]
  assign _T_1445 = _T_1423 ? _T_1439 : _T_1444; // @[Mux.scala 31:69:@16705.4]
  assign _T_1446 = _T_1422 ? _T_1437 : _T_1445; // @[Mux.scala 31:69:@16706.4]
  assign _T_1447 = _T_1421 ? _T_1435 : _T_1446; // @[Mux.scala 31:69:@16707.4]
  assign _T_1448 = _T_1420 ? _T_1433 : _T_1447; // @[Mux.scala 31:69:@16708.4]
  assign _T_1449 = _T_1419 ? _T_1431 : _T_1448; // @[Mux.scala 31:69:@16709.4]
  assign _T_1450 = _T_1418 ? _T_1429 : _T_1449; // @[Mux.scala 31:69:@16710.4]
  assign _T_1451 = _T_1417 ? _T_1427 : _T_1450; // @[Mux.scala 31:69:@16711.4]
  assign _T_1458 = io_rPort_2_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@16719.4]
  assign _T_1459 = _T_1272 & _T_1458; // @[MemPrimitives.scala 110:228:@16720.4]
  assign _T_1464 = io_rPort_5_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@16723.4]
  assign _T_1465 = _T_1278 & _T_1464; // @[MemPrimitives.scala 110:228:@16724.4]
  assign _T_1470 = io_rPort_6_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@16727.4]
  assign _T_1471 = _T_1284 & _T_1470; // @[MemPrimitives.scala 110:228:@16728.4]
  assign _T_1476 = io_rPort_7_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@16731.4]
  assign _T_1477 = _T_1290 & _T_1476; // @[MemPrimitives.scala 110:228:@16732.4]
  assign _T_1482 = io_rPort_9_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@16735.4]
  assign _T_1483 = _T_1296 & _T_1482; // @[MemPrimitives.scala 110:228:@16736.4]
  assign _T_1488 = io_rPort_11_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@16739.4]
  assign _T_1489 = _T_1302 & _T_1488; // @[MemPrimitives.scala 110:228:@16740.4]
  assign _T_1494 = io_rPort_12_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@16743.4]
  assign _T_1495 = _T_1308 & _T_1494; // @[MemPrimitives.scala 110:228:@16744.4]
  assign _T_1500 = io_rPort_13_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@16747.4]
  assign _T_1501 = _T_1314 & _T_1500; // @[MemPrimitives.scala 110:228:@16748.4]
  assign _T_1506 = io_rPort_16_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@16751.4]
  assign _T_1507 = _T_1320 & _T_1506; // @[MemPrimitives.scala 110:228:@16752.4]
  assign _T_1509 = StickySelects_3_io_outs_0; // @[MemPrimitives.scala 123:41:@16766.4]
  assign _T_1510 = StickySelects_3_io_outs_1; // @[MemPrimitives.scala 123:41:@16767.4]
  assign _T_1511 = StickySelects_3_io_outs_2; // @[MemPrimitives.scala 123:41:@16768.4]
  assign _T_1512 = StickySelects_3_io_outs_3; // @[MemPrimitives.scala 123:41:@16769.4]
  assign _T_1513 = StickySelects_3_io_outs_4; // @[MemPrimitives.scala 123:41:@16770.4]
  assign _T_1514 = StickySelects_3_io_outs_5; // @[MemPrimitives.scala 123:41:@16771.4]
  assign _T_1515 = StickySelects_3_io_outs_6; // @[MemPrimitives.scala 123:41:@16772.4]
  assign _T_1516 = StickySelects_3_io_outs_7; // @[MemPrimitives.scala 123:41:@16773.4]
  assign _T_1517 = StickySelects_3_io_outs_8; // @[MemPrimitives.scala 123:41:@16774.4]
  assign _T_1519 = {_T_1509,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@16776.4]
  assign _T_1521 = {_T_1510,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@16778.4]
  assign _T_1523 = {_T_1511,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@16780.4]
  assign _T_1525 = {_T_1512,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@16782.4]
  assign _T_1527 = {_T_1513,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@16784.4]
  assign _T_1529 = {_T_1514,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@16786.4]
  assign _T_1531 = {_T_1515,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@16788.4]
  assign _T_1533 = {_T_1516,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@16790.4]
  assign _T_1535 = {_T_1517,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@16792.4]
  assign _T_1536 = _T_1516 ? _T_1533 : _T_1535; // @[Mux.scala 31:69:@16793.4]
  assign _T_1537 = _T_1515 ? _T_1531 : _T_1536; // @[Mux.scala 31:69:@16794.4]
  assign _T_1538 = _T_1514 ? _T_1529 : _T_1537; // @[Mux.scala 31:69:@16795.4]
  assign _T_1539 = _T_1513 ? _T_1527 : _T_1538; // @[Mux.scala 31:69:@16796.4]
  assign _T_1540 = _T_1512 ? _T_1525 : _T_1539; // @[Mux.scala 31:69:@16797.4]
  assign _T_1541 = _T_1511 ? _T_1523 : _T_1540; // @[Mux.scala 31:69:@16798.4]
  assign _T_1542 = _T_1510 ? _T_1521 : _T_1541; // @[Mux.scala 31:69:@16799.4]
  assign _T_1543 = _T_1509 ? _T_1519 : _T_1542; // @[Mux.scala 31:69:@16800.4]
  assign _T_1550 = io_rPort_0_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@16808.4]
  assign _T_1551 = _T_1180 & _T_1550; // @[MemPrimitives.scala 110:228:@16809.4]
  assign _T_1556 = io_rPort_1_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@16812.4]
  assign _T_1557 = _T_1186 & _T_1556; // @[MemPrimitives.scala 110:228:@16813.4]
  assign _T_1562 = io_rPort_3_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@16816.4]
  assign _T_1563 = _T_1192 & _T_1562; // @[MemPrimitives.scala 110:228:@16817.4]
  assign _T_1568 = io_rPort_4_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@16820.4]
  assign _T_1569 = _T_1198 & _T_1568; // @[MemPrimitives.scala 110:228:@16821.4]
  assign _T_1574 = io_rPort_8_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@16824.4]
  assign _T_1575 = _T_1204 & _T_1574; // @[MemPrimitives.scala 110:228:@16825.4]
  assign _T_1580 = io_rPort_10_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@16828.4]
  assign _T_1581 = _T_1210 & _T_1580; // @[MemPrimitives.scala 110:228:@16829.4]
  assign _T_1586 = io_rPort_14_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@16832.4]
  assign _T_1587 = _T_1216 & _T_1586; // @[MemPrimitives.scala 110:228:@16833.4]
  assign _T_1592 = io_rPort_15_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@16836.4]
  assign _T_1593 = _T_1222 & _T_1592; // @[MemPrimitives.scala 110:228:@16837.4]
  assign _T_1598 = io_rPort_17_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@16840.4]
  assign _T_1599 = _T_1228 & _T_1598; // @[MemPrimitives.scala 110:228:@16841.4]
  assign _T_1601 = StickySelects_4_io_outs_0; // @[MemPrimitives.scala 123:41:@16855.4]
  assign _T_1602 = StickySelects_4_io_outs_1; // @[MemPrimitives.scala 123:41:@16856.4]
  assign _T_1603 = StickySelects_4_io_outs_2; // @[MemPrimitives.scala 123:41:@16857.4]
  assign _T_1604 = StickySelects_4_io_outs_3; // @[MemPrimitives.scala 123:41:@16858.4]
  assign _T_1605 = StickySelects_4_io_outs_4; // @[MemPrimitives.scala 123:41:@16859.4]
  assign _T_1606 = StickySelects_4_io_outs_5; // @[MemPrimitives.scala 123:41:@16860.4]
  assign _T_1607 = StickySelects_4_io_outs_6; // @[MemPrimitives.scala 123:41:@16861.4]
  assign _T_1608 = StickySelects_4_io_outs_7; // @[MemPrimitives.scala 123:41:@16862.4]
  assign _T_1609 = StickySelects_4_io_outs_8; // @[MemPrimitives.scala 123:41:@16863.4]
  assign _T_1611 = {_T_1601,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@16865.4]
  assign _T_1613 = {_T_1602,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@16867.4]
  assign _T_1615 = {_T_1603,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@16869.4]
  assign _T_1617 = {_T_1604,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@16871.4]
  assign _T_1619 = {_T_1605,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@16873.4]
  assign _T_1621 = {_T_1606,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@16875.4]
  assign _T_1623 = {_T_1607,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@16877.4]
  assign _T_1625 = {_T_1608,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@16879.4]
  assign _T_1627 = {_T_1609,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@16881.4]
  assign _T_1628 = _T_1608 ? _T_1625 : _T_1627; // @[Mux.scala 31:69:@16882.4]
  assign _T_1629 = _T_1607 ? _T_1623 : _T_1628; // @[Mux.scala 31:69:@16883.4]
  assign _T_1630 = _T_1606 ? _T_1621 : _T_1629; // @[Mux.scala 31:69:@16884.4]
  assign _T_1631 = _T_1605 ? _T_1619 : _T_1630; // @[Mux.scala 31:69:@16885.4]
  assign _T_1632 = _T_1604 ? _T_1617 : _T_1631; // @[Mux.scala 31:69:@16886.4]
  assign _T_1633 = _T_1603 ? _T_1615 : _T_1632; // @[Mux.scala 31:69:@16887.4]
  assign _T_1634 = _T_1602 ? _T_1613 : _T_1633; // @[Mux.scala 31:69:@16888.4]
  assign _T_1635 = _T_1601 ? _T_1611 : _T_1634; // @[Mux.scala 31:69:@16889.4]
  assign _T_1642 = io_rPort_2_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@16897.4]
  assign _T_1643 = _T_1272 & _T_1642; // @[MemPrimitives.scala 110:228:@16898.4]
  assign _T_1648 = io_rPort_5_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@16901.4]
  assign _T_1649 = _T_1278 & _T_1648; // @[MemPrimitives.scala 110:228:@16902.4]
  assign _T_1654 = io_rPort_6_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@16905.4]
  assign _T_1655 = _T_1284 & _T_1654; // @[MemPrimitives.scala 110:228:@16906.4]
  assign _T_1660 = io_rPort_7_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@16909.4]
  assign _T_1661 = _T_1290 & _T_1660; // @[MemPrimitives.scala 110:228:@16910.4]
  assign _T_1666 = io_rPort_9_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@16913.4]
  assign _T_1667 = _T_1296 & _T_1666; // @[MemPrimitives.scala 110:228:@16914.4]
  assign _T_1672 = io_rPort_11_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@16917.4]
  assign _T_1673 = _T_1302 & _T_1672; // @[MemPrimitives.scala 110:228:@16918.4]
  assign _T_1678 = io_rPort_12_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@16921.4]
  assign _T_1679 = _T_1308 & _T_1678; // @[MemPrimitives.scala 110:228:@16922.4]
  assign _T_1684 = io_rPort_13_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@16925.4]
  assign _T_1685 = _T_1314 & _T_1684; // @[MemPrimitives.scala 110:228:@16926.4]
  assign _T_1690 = io_rPort_16_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@16929.4]
  assign _T_1691 = _T_1320 & _T_1690; // @[MemPrimitives.scala 110:228:@16930.4]
  assign _T_1693 = StickySelects_5_io_outs_0; // @[MemPrimitives.scala 123:41:@16944.4]
  assign _T_1694 = StickySelects_5_io_outs_1; // @[MemPrimitives.scala 123:41:@16945.4]
  assign _T_1695 = StickySelects_5_io_outs_2; // @[MemPrimitives.scala 123:41:@16946.4]
  assign _T_1696 = StickySelects_5_io_outs_3; // @[MemPrimitives.scala 123:41:@16947.4]
  assign _T_1697 = StickySelects_5_io_outs_4; // @[MemPrimitives.scala 123:41:@16948.4]
  assign _T_1698 = StickySelects_5_io_outs_5; // @[MemPrimitives.scala 123:41:@16949.4]
  assign _T_1699 = StickySelects_5_io_outs_6; // @[MemPrimitives.scala 123:41:@16950.4]
  assign _T_1700 = StickySelects_5_io_outs_7; // @[MemPrimitives.scala 123:41:@16951.4]
  assign _T_1701 = StickySelects_5_io_outs_8; // @[MemPrimitives.scala 123:41:@16952.4]
  assign _T_1703 = {_T_1693,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@16954.4]
  assign _T_1705 = {_T_1694,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@16956.4]
  assign _T_1707 = {_T_1695,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@16958.4]
  assign _T_1709 = {_T_1696,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@16960.4]
  assign _T_1711 = {_T_1697,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@16962.4]
  assign _T_1713 = {_T_1698,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@16964.4]
  assign _T_1715 = {_T_1699,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@16966.4]
  assign _T_1717 = {_T_1700,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@16968.4]
  assign _T_1719 = {_T_1701,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@16970.4]
  assign _T_1720 = _T_1700 ? _T_1717 : _T_1719; // @[Mux.scala 31:69:@16971.4]
  assign _T_1721 = _T_1699 ? _T_1715 : _T_1720; // @[Mux.scala 31:69:@16972.4]
  assign _T_1722 = _T_1698 ? _T_1713 : _T_1721; // @[Mux.scala 31:69:@16973.4]
  assign _T_1723 = _T_1697 ? _T_1711 : _T_1722; // @[Mux.scala 31:69:@16974.4]
  assign _T_1724 = _T_1696 ? _T_1709 : _T_1723; // @[Mux.scala 31:69:@16975.4]
  assign _T_1725 = _T_1695 ? _T_1707 : _T_1724; // @[Mux.scala 31:69:@16976.4]
  assign _T_1726 = _T_1694 ? _T_1705 : _T_1725; // @[Mux.scala 31:69:@16977.4]
  assign _T_1727 = _T_1693 ? _T_1703 : _T_1726; // @[Mux.scala 31:69:@16978.4]
  assign _T_1732 = io_rPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@16985.4]
  assign _T_1735 = _T_1732 & _T_1182; // @[MemPrimitives.scala 110:228:@16987.4]
  assign _T_1738 = io_rPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@16989.4]
  assign _T_1741 = _T_1738 & _T_1188; // @[MemPrimitives.scala 110:228:@16991.4]
  assign _T_1744 = io_rPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@16993.4]
  assign _T_1747 = _T_1744 & _T_1194; // @[MemPrimitives.scala 110:228:@16995.4]
  assign _T_1750 = io_rPort_4_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@16997.4]
  assign _T_1753 = _T_1750 & _T_1200; // @[MemPrimitives.scala 110:228:@16999.4]
  assign _T_1756 = io_rPort_8_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@17001.4]
  assign _T_1759 = _T_1756 & _T_1206; // @[MemPrimitives.scala 110:228:@17003.4]
  assign _T_1762 = io_rPort_10_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@17005.4]
  assign _T_1765 = _T_1762 & _T_1212; // @[MemPrimitives.scala 110:228:@17007.4]
  assign _T_1768 = io_rPort_14_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@17009.4]
  assign _T_1771 = _T_1768 & _T_1218; // @[MemPrimitives.scala 110:228:@17011.4]
  assign _T_1774 = io_rPort_15_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@17013.4]
  assign _T_1777 = _T_1774 & _T_1224; // @[MemPrimitives.scala 110:228:@17015.4]
  assign _T_1780 = io_rPort_17_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@17017.4]
  assign _T_1783 = _T_1780 & _T_1230; // @[MemPrimitives.scala 110:228:@17019.4]
  assign _T_1785 = StickySelects_6_io_outs_0; // @[MemPrimitives.scala 123:41:@17033.4]
  assign _T_1786 = StickySelects_6_io_outs_1; // @[MemPrimitives.scala 123:41:@17034.4]
  assign _T_1787 = StickySelects_6_io_outs_2; // @[MemPrimitives.scala 123:41:@17035.4]
  assign _T_1788 = StickySelects_6_io_outs_3; // @[MemPrimitives.scala 123:41:@17036.4]
  assign _T_1789 = StickySelects_6_io_outs_4; // @[MemPrimitives.scala 123:41:@17037.4]
  assign _T_1790 = StickySelects_6_io_outs_5; // @[MemPrimitives.scala 123:41:@17038.4]
  assign _T_1791 = StickySelects_6_io_outs_6; // @[MemPrimitives.scala 123:41:@17039.4]
  assign _T_1792 = StickySelects_6_io_outs_7; // @[MemPrimitives.scala 123:41:@17040.4]
  assign _T_1793 = StickySelects_6_io_outs_8; // @[MemPrimitives.scala 123:41:@17041.4]
  assign _T_1795 = {_T_1785,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@17043.4]
  assign _T_1797 = {_T_1786,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@17045.4]
  assign _T_1799 = {_T_1787,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@17047.4]
  assign _T_1801 = {_T_1788,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@17049.4]
  assign _T_1803 = {_T_1789,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@17051.4]
  assign _T_1805 = {_T_1790,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@17053.4]
  assign _T_1807 = {_T_1791,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@17055.4]
  assign _T_1809 = {_T_1792,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@17057.4]
  assign _T_1811 = {_T_1793,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@17059.4]
  assign _T_1812 = _T_1792 ? _T_1809 : _T_1811; // @[Mux.scala 31:69:@17060.4]
  assign _T_1813 = _T_1791 ? _T_1807 : _T_1812; // @[Mux.scala 31:69:@17061.4]
  assign _T_1814 = _T_1790 ? _T_1805 : _T_1813; // @[Mux.scala 31:69:@17062.4]
  assign _T_1815 = _T_1789 ? _T_1803 : _T_1814; // @[Mux.scala 31:69:@17063.4]
  assign _T_1816 = _T_1788 ? _T_1801 : _T_1815; // @[Mux.scala 31:69:@17064.4]
  assign _T_1817 = _T_1787 ? _T_1799 : _T_1816; // @[Mux.scala 31:69:@17065.4]
  assign _T_1818 = _T_1786 ? _T_1797 : _T_1817; // @[Mux.scala 31:69:@17066.4]
  assign _T_1819 = _T_1785 ? _T_1795 : _T_1818; // @[Mux.scala 31:69:@17067.4]
  assign _T_1824 = io_rPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@17074.4]
  assign _T_1827 = _T_1824 & _T_1274; // @[MemPrimitives.scala 110:228:@17076.4]
  assign _T_1830 = io_rPort_5_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@17078.4]
  assign _T_1833 = _T_1830 & _T_1280; // @[MemPrimitives.scala 110:228:@17080.4]
  assign _T_1836 = io_rPort_6_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@17082.4]
  assign _T_1839 = _T_1836 & _T_1286; // @[MemPrimitives.scala 110:228:@17084.4]
  assign _T_1842 = io_rPort_7_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@17086.4]
  assign _T_1845 = _T_1842 & _T_1292; // @[MemPrimitives.scala 110:228:@17088.4]
  assign _T_1848 = io_rPort_9_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@17090.4]
  assign _T_1851 = _T_1848 & _T_1298; // @[MemPrimitives.scala 110:228:@17092.4]
  assign _T_1854 = io_rPort_11_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@17094.4]
  assign _T_1857 = _T_1854 & _T_1304; // @[MemPrimitives.scala 110:228:@17096.4]
  assign _T_1860 = io_rPort_12_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@17098.4]
  assign _T_1863 = _T_1860 & _T_1310; // @[MemPrimitives.scala 110:228:@17100.4]
  assign _T_1866 = io_rPort_13_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@17102.4]
  assign _T_1869 = _T_1866 & _T_1316; // @[MemPrimitives.scala 110:228:@17104.4]
  assign _T_1872 = io_rPort_16_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@17106.4]
  assign _T_1875 = _T_1872 & _T_1322; // @[MemPrimitives.scala 110:228:@17108.4]
  assign _T_1877 = StickySelects_7_io_outs_0; // @[MemPrimitives.scala 123:41:@17122.4]
  assign _T_1878 = StickySelects_7_io_outs_1; // @[MemPrimitives.scala 123:41:@17123.4]
  assign _T_1879 = StickySelects_7_io_outs_2; // @[MemPrimitives.scala 123:41:@17124.4]
  assign _T_1880 = StickySelects_7_io_outs_3; // @[MemPrimitives.scala 123:41:@17125.4]
  assign _T_1881 = StickySelects_7_io_outs_4; // @[MemPrimitives.scala 123:41:@17126.4]
  assign _T_1882 = StickySelects_7_io_outs_5; // @[MemPrimitives.scala 123:41:@17127.4]
  assign _T_1883 = StickySelects_7_io_outs_6; // @[MemPrimitives.scala 123:41:@17128.4]
  assign _T_1884 = StickySelects_7_io_outs_7; // @[MemPrimitives.scala 123:41:@17129.4]
  assign _T_1885 = StickySelects_7_io_outs_8; // @[MemPrimitives.scala 123:41:@17130.4]
  assign _T_1887 = {_T_1877,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@17132.4]
  assign _T_1889 = {_T_1878,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@17134.4]
  assign _T_1891 = {_T_1879,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@17136.4]
  assign _T_1893 = {_T_1880,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@17138.4]
  assign _T_1895 = {_T_1881,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@17140.4]
  assign _T_1897 = {_T_1882,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@17142.4]
  assign _T_1899 = {_T_1883,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@17144.4]
  assign _T_1901 = {_T_1884,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@17146.4]
  assign _T_1903 = {_T_1885,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@17148.4]
  assign _T_1904 = _T_1884 ? _T_1901 : _T_1903; // @[Mux.scala 31:69:@17149.4]
  assign _T_1905 = _T_1883 ? _T_1899 : _T_1904; // @[Mux.scala 31:69:@17150.4]
  assign _T_1906 = _T_1882 ? _T_1897 : _T_1905; // @[Mux.scala 31:69:@17151.4]
  assign _T_1907 = _T_1881 ? _T_1895 : _T_1906; // @[Mux.scala 31:69:@17152.4]
  assign _T_1908 = _T_1880 ? _T_1893 : _T_1907; // @[Mux.scala 31:69:@17153.4]
  assign _T_1909 = _T_1879 ? _T_1891 : _T_1908; // @[Mux.scala 31:69:@17154.4]
  assign _T_1910 = _T_1878 ? _T_1889 : _T_1909; // @[Mux.scala 31:69:@17155.4]
  assign _T_1911 = _T_1877 ? _T_1887 : _T_1910; // @[Mux.scala 31:69:@17156.4]
  assign _T_1919 = _T_1732 & _T_1366; // @[MemPrimitives.scala 110:228:@17165.4]
  assign _T_1925 = _T_1738 & _T_1372; // @[MemPrimitives.scala 110:228:@17169.4]
  assign _T_1931 = _T_1744 & _T_1378; // @[MemPrimitives.scala 110:228:@17173.4]
  assign _T_1937 = _T_1750 & _T_1384; // @[MemPrimitives.scala 110:228:@17177.4]
  assign _T_1943 = _T_1756 & _T_1390; // @[MemPrimitives.scala 110:228:@17181.4]
  assign _T_1949 = _T_1762 & _T_1396; // @[MemPrimitives.scala 110:228:@17185.4]
  assign _T_1955 = _T_1768 & _T_1402; // @[MemPrimitives.scala 110:228:@17189.4]
  assign _T_1961 = _T_1774 & _T_1408; // @[MemPrimitives.scala 110:228:@17193.4]
  assign _T_1967 = _T_1780 & _T_1414; // @[MemPrimitives.scala 110:228:@17197.4]
  assign _T_1969 = StickySelects_8_io_outs_0; // @[MemPrimitives.scala 123:41:@17211.4]
  assign _T_1970 = StickySelects_8_io_outs_1; // @[MemPrimitives.scala 123:41:@17212.4]
  assign _T_1971 = StickySelects_8_io_outs_2; // @[MemPrimitives.scala 123:41:@17213.4]
  assign _T_1972 = StickySelects_8_io_outs_3; // @[MemPrimitives.scala 123:41:@17214.4]
  assign _T_1973 = StickySelects_8_io_outs_4; // @[MemPrimitives.scala 123:41:@17215.4]
  assign _T_1974 = StickySelects_8_io_outs_5; // @[MemPrimitives.scala 123:41:@17216.4]
  assign _T_1975 = StickySelects_8_io_outs_6; // @[MemPrimitives.scala 123:41:@17217.4]
  assign _T_1976 = StickySelects_8_io_outs_7; // @[MemPrimitives.scala 123:41:@17218.4]
  assign _T_1977 = StickySelects_8_io_outs_8; // @[MemPrimitives.scala 123:41:@17219.4]
  assign _T_1979 = {_T_1969,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@17221.4]
  assign _T_1981 = {_T_1970,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@17223.4]
  assign _T_1983 = {_T_1971,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@17225.4]
  assign _T_1985 = {_T_1972,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@17227.4]
  assign _T_1987 = {_T_1973,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@17229.4]
  assign _T_1989 = {_T_1974,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@17231.4]
  assign _T_1991 = {_T_1975,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@17233.4]
  assign _T_1993 = {_T_1976,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@17235.4]
  assign _T_1995 = {_T_1977,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@17237.4]
  assign _T_1996 = _T_1976 ? _T_1993 : _T_1995; // @[Mux.scala 31:69:@17238.4]
  assign _T_1997 = _T_1975 ? _T_1991 : _T_1996; // @[Mux.scala 31:69:@17239.4]
  assign _T_1998 = _T_1974 ? _T_1989 : _T_1997; // @[Mux.scala 31:69:@17240.4]
  assign _T_1999 = _T_1973 ? _T_1987 : _T_1998; // @[Mux.scala 31:69:@17241.4]
  assign _T_2000 = _T_1972 ? _T_1985 : _T_1999; // @[Mux.scala 31:69:@17242.4]
  assign _T_2001 = _T_1971 ? _T_1983 : _T_2000; // @[Mux.scala 31:69:@17243.4]
  assign _T_2002 = _T_1970 ? _T_1981 : _T_2001; // @[Mux.scala 31:69:@17244.4]
  assign _T_2003 = _T_1969 ? _T_1979 : _T_2002; // @[Mux.scala 31:69:@17245.4]
  assign _T_2011 = _T_1824 & _T_1458; // @[MemPrimitives.scala 110:228:@17254.4]
  assign _T_2017 = _T_1830 & _T_1464; // @[MemPrimitives.scala 110:228:@17258.4]
  assign _T_2023 = _T_1836 & _T_1470; // @[MemPrimitives.scala 110:228:@17262.4]
  assign _T_2029 = _T_1842 & _T_1476; // @[MemPrimitives.scala 110:228:@17266.4]
  assign _T_2035 = _T_1848 & _T_1482; // @[MemPrimitives.scala 110:228:@17270.4]
  assign _T_2041 = _T_1854 & _T_1488; // @[MemPrimitives.scala 110:228:@17274.4]
  assign _T_2047 = _T_1860 & _T_1494; // @[MemPrimitives.scala 110:228:@17278.4]
  assign _T_2053 = _T_1866 & _T_1500; // @[MemPrimitives.scala 110:228:@17282.4]
  assign _T_2059 = _T_1872 & _T_1506; // @[MemPrimitives.scala 110:228:@17286.4]
  assign _T_2061 = StickySelects_9_io_outs_0; // @[MemPrimitives.scala 123:41:@17300.4]
  assign _T_2062 = StickySelects_9_io_outs_1; // @[MemPrimitives.scala 123:41:@17301.4]
  assign _T_2063 = StickySelects_9_io_outs_2; // @[MemPrimitives.scala 123:41:@17302.4]
  assign _T_2064 = StickySelects_9_io_outs_3; // @[MemPrimitives.scala 123:41:@17303.4]
  assign _T_2065 = StickySelects_9_io_outs_4; // @[MemPrimitives.scala 123:41:@17304.4]
  assign _T_2066 = StickySelects_9_io_outs_5; // @[MemPrimitives.scala 123:41:@17305.4]
  assign _T_2067 = StickySelects_9_io_outs_6; // @[MemPrimitives.scala 123:41:@17306.4]
  assign _T_2068 = StickySelects_9_io_outs_7; // @[MemPrimitives.scala 123:41:@17307.4]
  assign _T_2069 = StickySelects_9_io_outs_8; // @[MemPrimitives.scala 123:41:@17308.4]
  assign _T_2071 = {_T_2061,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@17310.4]
  assign _T_2073 = {_T_2062,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@17312.4]
  assign _T_2075 = {_T_2063,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@17314.4]
  assign _T_2077 = {_T_2064,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@17316.4]
  assign _T_2079 = {_T_2065,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@17318.4]
  assign _T_2081 = {_T_2066,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@17320.4]
  assign _T_2083 = {_T_2067,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@17322.4]
  assign _T_2085 = {_T_2068,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@17324.4]
  assign _T_2087 = {_T_2069,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@17326.4]
  assign _T_2088 = _T_2068 ? _T_2085 : _T_2087; // @[Mux.scala 31:69:@17327.4]
  assign _T_2089 = _T_2067 ? _T_2083 : _T_2088; // @[Mux.scala 31:69:@17328.4]
  assign _T_2090 = _T_2066 ? _T_2081 : _T_2089; // @[Mux.scala 31:69:@17329.4]
  assign _T_2091 = _T_2065 ? _T_2079 : _T_2090; // @[Mux.scala 31:69:@17330.4]
  assign _T_2092 = _T_2064 ? _T_2077 : _T_2091; // @[Mux.scala 31:69:@17331.4]
  assign _T_2093 = _T_2063 ? _T_2075 : _T_2092; // @[Mux.scala 31:69:@17332.4]
  assign _T_2094 = _T_2062 ? _T_2073 : _T_2093; // @[Mux.scala 31:69:@17333.4]
  assign _T_2095 = _T_2061 ? _T_2071 : _T_2094; // @[Mux.scala 31:69:@17334.4]
  assign _T_2103 = _T_1732 & _T_1550; // @[MemPrimitives.scala 110:228:@17343.4]
  assign _T_2109 = _T_1738 & _T_1556; // @[MemPrimitives.scala 110:228:@17347.4]
  assign _T_2115 = _T_1744 & _T_1562; // @[MemPrimitives.scala 110:228:@17351.4]
  assign _T_2121 = _T_1750 & _T_1568; // @[MemPrimitives.scala 110:228:@17355.4]
  assign _T_2127 = _T_1756 & _T_1574; // @[MemPrimitives.scala 110:228:@17359.4]
  assign _T_2133 = _T_1762 & _T_1580; // @[MemPrimitives.scala 110:228:@17363.4]
  assign _T_2139 = _T_1768 & _T_1586; // @[MemPrimitives.scala 110:228:@17367.4]
  assign _T_2145 = _T_1774 & _T_1592; // @[MemPrimitives.scala 110:228:@17371.4]
  assign _T_2151 = _T_1780 & _T_1598; // @[MemPrimitives.scala 110:228:@17375.4]
  assign _T_2153 = StickySelects_10_io_outs_0; // @[MemPrimitives.scala 123:41:@17389.4]
  assign _T_2154 = StickySelects_10_io_outs_1; // @[MemPrimitives.scala 123:41:@17390.4]
  assign _T_2155 = StickySelects_10_io_outs_2; // @[MemPrimitives.scala 123:41:@17391.4]
  assign _T_2156 = StickySelects_10_io_outs_3; // @[MemPrimitives.scala 123:41:@17392.4]
  assign _T_2157 = StickySelects_10_io_outs_4; // @[MemPrimitives.scala 123:41:@17393.4]
  assign _T_2158 = StickySelects_10_io_outs_5; // @[MemPrimitives.scala 123:41:@17394.4]
  assign _T_2159 = StickySelects_10_io_outs_6; // @[MemPrimitives.scala 123:41:@17395.4]
  assign _T_2160 = StickySelects_10_io_outs_7; // @[MemPrimitives.scala 123:41:@17396.4]
  assign _T_2161 = StickySelects_10_io_outs_8; // @[MemPrimitives.scala 123:41:@17397.4]
  assign _T_2163 = {_T_2153,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@17399.4]
  assign _T_2165 = {_T_2154,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@17401.4]
  assign _T_2167 = {_T_2155,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@17403.4]
  assign _T_2169 = {_T_2156,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@17405.4]
  assign _T_2171 = {_T_2157,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@17407.4]
  assign _T_2173 = {_T_2158,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@17409.4]
  assign _T_2175 = {_T_2159,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@17411.4]
  assign _T_2177 = {_T_2160,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@17413.4]
  assign _T_2179 = {_T_2161,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@17415.4]
  assign _T_2180 = _T_2160 ? _T_2177 : _T_2179; // @[Mux.scala 31:69:@17416.4]
  assign _T_2181 = _T_2159 ? _T_2175 : _T_2180; // @[Mux.scala 31:69:@17417.4]
  assign _T_2182 = _T_2158 ? _T_2173 : _T_2181; // @[Mux.scala 31:69:@17418.4]
  assign _T_2183 = _T_2157 ? _T_2171 : _T_2182; // @[Mux.scala 31:69:@17419.4]
  assign _T_2184 = _T_2156 ? _T_2169 : _T_2183; // @[Mux.scala 31:69:@17420.4]
  assign _T_2185 = _T_2155 ? _T_2167 : _T_2184; // @[Mux.scala 31:69:@17421.4]
  assign _T_2186 = _T_2154 ? _T_2165 : _T_2185; // @[Mux.scala 31:69:@17422.4]
  assign _T_2187 = _T_2153 ? _T_2163 : _T_2186; // @[Mux.scala 31:69:@17423.4]
  assign _T_2195 = _T_1824 & _T_1642; // @[MemPrimitives.scala 110:228:@17432.4]
  assign _T_2201 = _T_1830 & _T_1648; // @[MemPrimitives.scala 110:228:@17436.4]
  assign _T_2207 = _T_1836 & _T_1654; // @[MemPrimitives.scala 110:228:@17440.4]
  assign _T_2213 = _T_1842 & _T_1660; // @[MemPrimitives.scala 110:228:@17444.4]
  assign _T_2219 = _T_1848 & _T_1666; // @[MemPrimitives.scala 110:228:@17448.4]
  assign _T_2225 = _T_1854 & _T_1672; // @[MemPrimitives.scala 110:228:@17452.4]
  assign _T_2231 = _T_1860 & _T_1678; // @[MemPrimitives.scala 110:228:@17456.4]
  assign _T_2237 = _T_1866 & _T_1684; // @[MemPrimitives.scala 110:228:@17460.4]
  assign _T_2243 = _T_1872 & _T_1690; // @[MemPrimitives.scala 110:228:@17464.4]
  assign _T_2245 = StickySelects_11_io_outs_0; // @[MemPrimitives.scala 123:41:@17478.4]
  assign _T_2246 = StickySelects_11_io_outs_1; // @[MemPrimitives.scala 123:41:@17479.4]
  assign _T_2247 = StickySelects_11_io_outs_2; // @[MemPrimitives.scala 123:41:@17480.4]
  assign _T_2248 = StickySelects_11_io_outs_3; // @[MemPrimitives.scala 123:41:@17481.4]
  assign _T_2249 = StickySelects_11_io_outs_4; // @[MemPrimitives.scala 123:41:@17482.4]
  assign _T_2250 = StickySelects_11_io_outs_5; // @[MemPrimitives.scala 123:41:@17483.4]
  assign _T_2251 = StickySelects_11_io_outs_6; // @[MemPrimitives.scala 123:41:@17484.4]
  assign _T_2252 = StickySelects_11_io_outs_7; // @[MemPrimitives.scala 123:41:@17485.4]
  assign _T_2253 = StickySelects_11_io_outs_8; // @[MemPrimitives.scala 123:41:@17486.4]
  assign _T_2255 = {_T_2245,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@17488.4]
  assign _T_2257 = {_T_2246,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@17490.4]
  assign _T_2259 = {_T_2247,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@17492.4]
  assign _T_2261 = {_T_2248,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@17494.4]
  assign _T_2263 = {_T_2249,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@17496.4]
  assign _T_2265 = {_T_2250,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@17498.4]
  assign _T_2267 = {_T_2251,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@17500.4]
  assign _T_2269 = {_T_2252,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@17502.4]
  assign _T_2271 = {_T_2253,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@17504.4]
  assign _T_2272 = _T_2252 ? _T_2269 : _T_2271; // @[Mux.scala 31:69:@17505.4]
  assign _T_2273 = _T_2251 ? _T_2267 : _T_2272; // @[Mux.scala 31:69:@17506.4]
  assign _T_2274 = _T_2250 ? _T_2265 : _T_2273; // @[Mux.scala 31:69:@17507.4]
  assign _T_2275 = _T_2249 ? _T_2263 : _T_2274; // @[Mux.scala 31:69:@17508.4]
  assign _T_2276 = _T_2248 ? _T_2261 : _T_2275; // @[Mux.scala 31:69:@17509.4]
  assign _T_2277 = _T_2247 ? _T_2259 : _T_2276; // @[Mux.scala 31:69:@17510.4]
  assign _T_2278 = _T_2246 ? _T_2257 : _T_2277; // @[Mux.scala 31:69:@17511.4]
  assign _T_2279 = _T_2245 ? _T_2255 : _T_2278; // @[Mux.scala 31:69:@17512.4]
  assign _T_2284 = io_rPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@17519.4]
  assign _T_2287 = _T_2284 & _T_1182; // @[MemPrimitives.scala 110:228:@17521.4]
  assign _T_2290 = io_rPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@17523.4]
  assign _T_2293 = _T_2290 & _T_1188; // @[MemPrimitives.scala 110:228:@17525.4]
  assign _T_2296 = io_rPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@17527.4]
  assign _T_2299 = _T_2296 & _T_1194; // @[MemPrimitives.scala 110:228:@17529.4]
  assign _T_2302 = io_rPort_4_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@17531.4]
  assign _T_2305 = _T_2302 & _T_1200; // @[MemPrimitives.scala 110:228:@17533.4]
  assign _T_2308 = io_rPort_8_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@17535.4]
  assign _T_2311 = _T_2308 & _T_1206; // @[MemPrimitives.scala 110:228:@17537.4]
  assign _T_2314 = io_rPort_10_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@17539.4]
  assign _T_2317 = _T_2314 & _T_1212; // @[MemPrimitives.scala 110:228:@17541.4]
  assign _T_2320 = io_rPort_14_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@17543.4]
  assign _T_2323 = _T_2320 & _T_1218; // @[MemPrimitives.scala 110:228:@17545.4]
  assign _T_2326 = io_rPort_15_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@17547.4]
  assign _T_2329 = _T_2326 & _T_1224; // @[MemPrimitives.scala 110:228:@17549.4]
  assign _T_2332 = io_rPort_17_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@17551.4]
  assign _T_2335 = _T_2332 & _T_1230; // @[MemPrimitives.scala 110:228:@17553.4]
  assign _T_2337 = StickySelects_12_io_outs_0; // @[MemPrimitives.scala 123:41:@17567.4]
  assign _T_2338 = StickySelects_12_io_outs_1; // @[MemPrimitives.scala 123:41:@17568.4]
  assign _T_2339 = StickySelects_12_io_outs_2; // @[MemPrimitives.scala 123:41:@17569.4]
  assign _T_2340 = StickySelects_12_io_outs_3; // @[MemPrimitives.scala 123:41:@17570.4]
  assign _T_2341 = StickySelects_12_io_outs_4; // @[MemPrimitives.scala 123:41:@17571.4]
  assign _T_2342 = StickySelects_12_io_outs_5; // @[MemPrimitives.scala 123:41:@17572.4]
  assign _T_2343 = StickySelects_12_io_outs_6; // @[MemPrimitives.scala 123:41:@17573.4]
  assign _T_2344 = StickySelects_12_io_outs_7; // @[MemPrimitives.scala 123:41:@17574.4]
  assign _T_2345 = StickySelects_12_io_outs_8; // @[MemPrimitives.scala 123:41:@17575.4]
  assign _T_2347 = {_T_2337,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@17577.4]
  assign _T_2349 = {_T_2338,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@17579.4]
  assign _T_2351 = {_T_2339,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@17581.4]
  assign _T_2353 = {_T_2340,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@17583.4]
  assign _T_2355 = {_T_2341,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@17585.4]
  assign _T_2357 = {_T_2342,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@17587.4]
  assign _T_2359 = {_T_2343,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@17589.4]
  assign _T_2361 = {_T_2344,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@17591.4]
  assign _T_2363 = {_T_2345,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@17593.4]
  assign _T_2364 = _T_2344 ? _T_2361 : _T_2363; // @[Mux.scala 31:69:@17594.4]
  assign _T_2365 = _T_2343 ? _T_2359 : _T_2364; // @[Mux.scala 31:69:@17595.4]
  assign _T_2366 = _T_2342 ? _T_2357 : _T_2365; // @[Mux.scala 31:69:@17596.4]
  assign _T_2367 = _T_2341 ? _T_2355 : _T_2366; // @[Mux.scala 31:69:@17597.4]
  assign _T_2368 = _T_2340 ? _T_2353 : _T_2367; // @[Mux.scala 31:69:@17598.4]
  assign _T_2369 = _T_2339 ? _T_2351 : _T_2368; // @[Mux.scala 31:69:@17599.4]
  assign _T_2370 = _T_2338 ? _T_2349 : _T_2369; // @[Mux.scala 31:69:@17600.4]
  assign _T_2371 = _T_2337 ? _T_2347 : _T_2370; // @[Mux.scala 31:69:@17601.4]
  assign _T_2376 = io_rPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@17608.4]
  assign _T_2379 = _T_2376 & _T_1274; // @[MemPrimitives.scala 110:228:@17610.4]
  assign _T_2382 = io_rPort_5_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@17612.4]
  assign _T_2385 = _T_2382 & _T_1280; // @[MemPrimitives.scala 110:228:@17614.4]
  assign _T_2388 = io_rPort_6_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@17616.4]
  assign _T_2391 = _T_2388 & _T_1286; // @[MemPrimitives.scala 110:228:@17618.4]
  assign _T_2394 = io_rPort_7_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@17620.4]
  assign _T_2397 = _T_2394 & _T_1292; // @[MemPrimitives.scala 110:228:@17622.4]
  assign _T_2400 = io_rPort_9_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@17624.4]
  assign _T_2403 = _T_2400 & _T_1298; // @[MemPrimitives.scala 110:228:@17626.4]
  assign _T_2406 = io_rPort_11_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@17628.4]
  assign _T_2409 = _T_2406 & _T_1304; // @[MemPrimitives.scala 110:228:@17630.4]
  assign _T_2412 = io_rPort_12_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@17632.4]
  assign _T_2415 = _T_2412 & _T_1310; // @[MemPrimitives.scala 110:228:@17634.4]
  assign _T_2418 = io_rPort_13_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@17636.4]
  assign _T_2421 = _T_2418 & _T_1316; // @[MemPrimitives.scala 110:228:@17638.4]
  assign _T_2424 = io_rPort_16_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@17640.4]
  assign _T_2427 = _T_2424 & _T_1322; // @[MemPrimitives.scala 110:228:@17642.4]
  assign _T_2429 = StickySelects_13_io_outs_0; // @[MemPrimitives.scala 123:41:@17656.4]
  assign _T_2430 = StickySelects_13_io_outs_1; // @[MemPrimitives.scala 123:41:@17657.4]
  assign _T_2431 = StickySelects_13_io_outs_2; // @[MemPrimitives.scala 123:41:@17658.4]
  assign _T_2432 = StickySelects_13_io_outs_3; // @[MemPrimitives.scala 123:41:@17659.4]
  assign _T_2433 = StickySelects_13_io_outs_4; // @[MemPrimitives.scala 123:41:@17660.4]
  assign _T_2434 = StickySelects_13_io_outs_5; // @[MemPrimitives.scala 123:41:@17661.4]
  assign _T_2435 = StickySelects_13_io_outs_6; // @[MemPrimitives.scala 123:41:@17662.4]
  assign _T_2436 = StickySelects_13_io_outs_7; // @[MemPrimitives.scala 123:41:@17663.4]
  assign _T_2437 = StickySelects_13_io_outs_8; // @[MemPrimitives.scala 123:41:@17664.4]
  assign _T_2439 = {_T_2429,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@17666.4]
  assign _T_2441 = {_T_2430,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@17668.4]
  assign _T_2443 = {_T_2431,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@17670.4]
  assign _T_2445 = {_T_2432,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@17672.4]
  assign _T_2447 = {_T_2433,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@17674.4]
  assign _T_2449 = {_T_2434,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@17676.4]
  assign _T_2451 = {_T_2435,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@17678.4]
  assign _T_2453 = {_T_2436,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@17680.4]
  assign _T_2455 = {_T_2437,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@17682.4]
  assign _T_2456 = _T_2436 ? _T_2453 : _T_2455; // @[Mux.scala 31:69:@17683.4]
  assign _T_2457 = _T_2435 ? _T_2451 : _T_2456; // @[Mux.scala 31:69:@17684.4]
  assign _T_2458 = _T_2434 ? _T_2449 : _T_2457; // @[Mux.scala 31:69:@17685.4]
  assign _T_2459 = _T_2433 ? _T_2447 : _T_2458; // @[Mux.scala 31:69:@17686.4]
  assign _T_2460 = _T_2432 ? _T_2445 : _T_2459; // @[Mux.scala 31:69:@17687.4]
  assign _T_2461 = _T_2431 ? _T_2443 : _T_2460; // @[Mux.scala 31:69:@17688.4]
  assign _T_2462 = _T_2430 ? _T_2441 : _T_2461; // @[Mux.scala 31:69:@17689.4]
  assign _T_2463 = _T_2429 ? _T_2439 : _T_2462; // @[Mux.scala 31:69:@17690.4]
  assign _T_2471 = _T_2284 & _T_1366; // @[MemPrimitives.scala 110:228:@17699.4]
  assign _T_2477 = _T_2290 & _T_1372; // @[MemPrimitives.scala 110:228:@17703.4]
  assign _T_2483 = _T_2296 & _T_1378; // @[MemPrimitives.scala 110:228:@17707.4]
  assign _T_2489 = _T_2302 & _T_1384; // @[MemPrimitives.scala 110:228:@17711.4]
  assign _T_2495 = _T_2308 & _T_1390; // @[MemPrimitives.scala 110:228:@17715.4]
  assign _T_2501 = _T_2314 & _T_1396; // @[MemPrimitives.scala 110:228:@17719.4]
  assign _T_2507 = _T_2320 & _T_1402; // @[MemPrimitives.scala 110:228:@17723.4]
  assign _T_2513 = _T_2326 & _T_1408; // @[MemPrimitives.scala 110:228:@17727.4]
  assign _T_2519 = _T_2332 & _T_1414; // @[MemPrimitives.scala 110:228:@17731.4]
  assign _T_2521 = StickySelects_14_io_outs_0; // @[MemPrimitives.scala 123:41:@17745.4]
  assign _T_2522 = StickySelects_14_io_outs_1; // @[MemPrimitives.scala 123:41:@17746.4]
  assign _T_2523 = StickySelects_14_io_outs_2; // @[MemPrimitives.scala 123:41:@17747.4]
  assign _T_2524 = StickySelects_14_io_outs_3; // @[MemPrimitives.scala 123:41:@17748.4]
  assign _T_2525 = StickySelects_14_io_outs_4; // @[MemPrimitives.scala 123:41:@17749.4]
  assign _T_2526 = StickySelects_14_io_outs_5; // @[MemPrimitives.scala 123:41:@17750.4]
  assign _T_2527 = StickySelects_14_io_outs_6; // @[MemPrimitives.scala 123:41:@17751.4]
  assign _T_2528 = StickySelects_14_io_outs_7; // @[MemPrimitives.scala 123:41:@17752.4]
  assign _T_2529 = StickySelects_14_io_outs_8; // @[MemPrimitives.scala 123:41:@17753.4]
  assign _T_2531 = {_T_2521,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@17755.4]
  assign _T_2533 = {_T_2522,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@17757.4]
  assign _T_2535 = {_T_2523,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@17759.4]
  assign _T_2537 = {_T_2524,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@17761.4]
  assign _T_2539 = {_T_2525,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@17763.4]
  assign _T_2541 = {_T_2526,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@17765.4]
  assign _T_2543 = {_T_2527,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@17767.4]
  assign _T_2545 = {_T_2528,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@17769.4]
  assign _T_2547 = {_T_2529,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@17771.4]
  assign _T_2548 = _T_2528 ? _T_2545 : _T_2547; // @[Mux.scala 31:69:@17772.4]
  assign _T_2549 = _T_2527 ? _T_2543 : _T_2548; // @[Mux.scala 31:69:@17773.4]
  assign _T_2550 = _T_2526 ? _T_2541 : _T_2549; // @[Mux.scala 31:69:@17774.4]
  assign _T_2551 = _T_2525 ? _T_2539 : _T_2550; // @[Mux.scala 31:69:@17775.4]
  assign _T_2552 = _T_2524 ? _T_2537 : _T_2551; // @[Mux.scala 31:69:@17776.4]
  assign _T_2553 = _T_2523 ? _T_2535 : _T_2552; // @[Mux.scala 31:69:@17777.4]
  assign _T_2554 = _T_2522 ? _T_2533 : _T_2553; // @[Mux.scala 31:69:@17778.4]
  assign _T_2555 = _T_2521 ? _T_2531 : _T_2554; // @[Mux.scala 31:69:@17779.4]
  assign _T_2563 = _T_2376 & _T_1458; // @[MemPrimitives.scala 110:228:@17788.4]
  assign _T_2569 = _T_2382 & _T_1464; // @[MemPrimitives.scala 110:228:@17792.4]
  assign _T_2575 = _T_2388 & _T_1470; // @[MemPrimitives.scala 110:228:@17796.4]
  assign _T_2581 = _T_2394 & _T_1476; // @[MemPrimitives.scala 110:228:@17800.4]
  assign _T_2587 = _T_2400 & _T_1482; // @[MemPrimitives.scala 110:228:@17804.4]
  assign _T_2593 = _T_2406 & _T_1488; // @[MemPrimitives.scala 110:228:@17808.4]
  assign _T_2599 = _T_2412 & _T_1494; // @[MemPrimitives.scala 110:228:@17812.4]
  assign _T_2605 = _T_2418 & _T_1500; // @[MemPrimitives.scala 110:228:@17816.4]
  assign _T_2611 = _T_2424 & _T_1506; // @[MemPrimitives.scala 110:228:@17820.4]
  assign _T_2613 = StickySelects_15_io_outs_0; // @[MemPrimitives.scala 123:41:@17834.4]
  assign _T_2614 = StickySelects_15_io_outs_1; // @[MemPrimitives.scala 123:41:@17835.4]
  assign _T_2615 = StickySelects_15_io_outs_2; // @[MemPrimitives.scala 123:41:@17836.4]
  assign _T_2616 = StickySelects_15_io_outs_3; // @[MemPrimitives.scala 123:41:@17837.4]
  assign _T_2617 = StickySelects_15_io_outs_4; // @[MemPrimitives.scala 123:41:@17838.4]
  assign _T_2618 = StickySelects_15_io_outs_5; // @[MemPrimitives.scala 123:41:@17839.4]
  assign _T_2619 = StickySelects_15_io_outs_6; // @[MemPrimitives.scala 123:41:@17840.4]
  assign _T_2620 = StickySelects_15_io_outs_7; // @[MemPrimitives.scala 123:41:@17841.4]
  assign _T_2621 = StickySelects_15_io_outs_8; // @[MemPrimitives.scala 123:41:@17842.4]
  assign _T_2623 = {_T_2613,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@17844.4]
  assign _T_2625 = {_T_2614,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@17846.4]
  assign _T_2627 = {_T_2615,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@17848.4]
  assign _T_2629 = {_T_2616,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@17850.4]
  assign _T_2631 = {_T_2617,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@17852.4]
  assign _T_2633 = {_T_2618,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@17854.4]
  assign _T_2635 = {_T_2619,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@17856.4]
  assign _T_2637 = {_T_2620,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@17858.4]
  assign _T_2639 = {_T_2621,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@17860.4]
  assign _T_2640 = _T_2620 ? _T_2637 : _T_2639; // @[Mux.scala 31:69:@17861.4]
  assign _T_2641 = _T_2619 ? _T_2635 : _T_2640; // @[Mux.scala 31:69:@17862.4]
  assign _T_2642 = _T_2618 ? _T_2633 : _T_2641; // @[Mux.scala 31:69:@17863.4]
  assign _T_2643 = _T_2617 ? _T_2631 : _T_2642; // @[Mux.scala 31:69:@17864.4]
  assign _T_2644 = _T_2616 ? _T_2629 : _T_2643; // @[Mux.scala 31:69:@17865.4]
  assign _T_2645 = _T_2615 ? _T_2627 : _T_2644; // @[Mux.scala 31:69:@17866.4]
  assign _T_2646 = _T_2614 ? _T_2625 : _T_2645; // @[Mux.scala 31:69:@17867.4]
  assign _T_2647 = _T_2613 ? _T_2623 : _T_2646; // @[Mux.scala 31:69:@17868.4]
  assign _T_2655 = _T_2284 & _T_1550; // @[MemPrimitives.scala 110:228:@17877.4]
  assign _T_2661 = _T_2290 & _T_1556; // @[MemPrimitives.scala 110:228:@17881.4]
  assign _T_2667 = _T_2296 & _T_1562; // @[MemPrimitives.scala 110:228:@17885.4]
  assign _T_2673 = _T_2302 & _T_1568; // @[MemPrimitives.scala 110:228:@17889.4]
  assign _T_2679 = _T_2308 & _T_1574; // @[MemPrimitives.scala 110:228:@17893.4]
  assign _T_2685 = _T_2314 & _T_1580; // @[MemPrimitives.scala 110:228:@17897.4]
  assign _T_2691 = _T_2320 & _T_1586; // @[MemPrimitives.scala 110:228:@17901.4]
  assign _T_2697 = _T_2326 & _T_1592; // @[MemPrimitives.scala 110:228:@17905.4]
  assign _T_2703 = _T_2332 & _T_1598; // @[MemPrimitives.scala 110:228:@17909.4]
  assign _T_2705 = StickySelects_16_io_outs_0; // @[MemPrimitives.scala 123:41:@17923.4]
  assign _T_2706 = StickySelects_16_io_outs_1; // @[MemPrimitives.scala 123:41:@17924.4]
  assign _T_2707 = StickySelects_16_io_outs_2; // @[MemPrimitives.scala 123:41:@17925.4]
  assign _T_2708 = StickySelects_16_io_outs_3; // @[MemPrimitives.scala 123:41:@17926.4]
  assign _T_2709 = StickySelects_16_io_outs_4; // @[MemPrimitives.scala 123:41:@17927.4]
  assign _T_2710 = StickySelects_16_io_outs_5; // @[MemPrimitives.scala 123:41:@17928.4]
  assign _T_2711 = StickySelects_16_io_outs_6; // @[MemPrimitives.scala 123:41:@17929.4]
  assign _T_2712 = StickySelects_16_io_outs_7; // @[MemPrimitives.scala 123:41:@17930.4]
  assign _T_2713 = StickySelects_16_io_outs_8; // @[MemPrimitives.scala 123:41:@17931.4]
  assign _T_2715 = {_T_2705,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@17933.4]
  assign _T_2717 = {_T_2706,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@17935.4]
  assign _T_2719 = {_T_2707,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@17937.4]
  assign _T_2721 = {_T_2708,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@17939.4]
  assign _T_2723 = {_T_2709,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@17941.4]
  assign _T_2725 = {_T_2710,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@17943.4]
  assign _T_2727 = {_T_2711,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@17945.4]
  assign _T_2729 = {_T_2712,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@17947.4]
  assign _T_2731 = {_T_2713,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@17949.4]
  assign _T_2732 = _T_2712 ? _T_2729 : _T_2731; // @[Mux.scala 31:69:@17950.4]
  assign _T_2733 = _T_2711 ? _T_2727 : _T_2732; // @[Mux.scala 31:69:@17951.4]
  assign _T_2734 = _T_2710 ? _T_2725 : _T_2733; // @[Mux.scala 31:69:@17952.4]
  assign _T_2735 = _T_2709 ? _T_2723 : _T_2734; // @[Mux.scala 31:69:@17953.4]
  assign _T_2736 = _T_2708 ? _T_2721 : _T_2735; // @[Mux.scala 31:69:@17954.4]
  assign _T_2737 = _T_2707 ? _T_2719 : _T_2736; // @[Mux.scala 31:69:@17955.4]
  assign _T_2738 = _T_2706 ? _T_2717 : _T_2737; // @[Mux.scala 31:69:@17956.4]
  assign _T_2739 = _T_2705 ? _T_2715 : _T_2738; // @[Mux.scala 31:69:@17957.4]
  assign _T_2747 = _T_2376 & _T_1642; // @[MemPrimitives.scala 110:228:@17966.4]
  assign _T_2753 = _T_2382 & _T_1648; // @[MemPrimitives.scala 110:228:@17970.4]
  assign _T_2759 = _T_2388 & _T_1654; // @[MemPrimitives.scala 110:228:@17974.4]
  assign _T_2765 = _T_2394 & _T_1660; // @[MemPrimitives.scala 110:228:@17978.4]
  assign _T_2771 = _T_2400 & _T_1666; // @[MemPrimitives.scala 110:228:@17982.4]
  assign _T_2777 = _T_2406 & _T_1672; // @[MemPrimitives.scala 110:228:@17986.4]
  assign _T_2783 = _T_2412 & _T_1678; // @[MemPrimitives.scala 110:228:@17990.4]
  assign _T_2789 = _T_2418 & _T_1684; // @[MemPrimitives.scala 110:228:@17994.4]
  assign _T_2795 = _T_2424 & _T_1690; // @[MemPrimitives.scala 110:228:@17998.4]
  assign _T_2797 = StickySelects_17_io_outs_0; // @[MemPrimitives.scala 123:41:@18012.4]
  assign _T_2798 = StickySelects_17_io_outs_1; // @[MemPrimitives.scala 123:41:@18013.4]
  assign _T_2799 = StickySelects_17_io_outs_2; // @[MemPrimitives.scala 123:41:@18014.4]
  assign _T_2800 = StickySelects_17_io_outs_3; // @[MemPrimitives.scala 123:41:@18015.4]
  assign _T_2801 = StickySelects_17_io_outs_4; // @[MemPrimitives.scala 123:41:@18016.4]
  assign _T_2802 = StickySelects_17_io_outs_5; // @[MemPrimitives.scala 123:41:@18017.4]
  assign _T_2803 = StickySelects_17_io_outs_6; // @[MemPrimitives.scala 123:41:@18018.4]
  assign _T_2804 = StickySelects_17_io_outs_7; // @[MemPrimitives.scala 123:41:@18019.4]
  assign _T_2805 = StickySelects_17_io_outs_8; // @[MemPrimitives.scala 123:41:@18020.4]
  assign _T_2807 = {_T_2797,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@18022.4]
  assign _T_2809 = {_T_2798,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@18024.4]
  assign _T_2811 = {_T_2799,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@18026.4]
  assign _T_2813 = {_T_2800,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@18028.4]
  assign _T_2815 = {_T_2801,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@18030.4]
  assign _T_2817 = {_T_2802,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@18032.4]
  assign _T_2819 = {_T_2803,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@18034.4]
  assign _T_2821 = {_T_2804,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@18036.4]
  assign _T_2823 = {_T_2805,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@18038.4]
  assign _T_2824 = _T_2804 ? _T_2821 : _T_2823; // @[Mux.scala 31:69:@18039.4]
  assign _T_2825 = _T_2803 ? _T_2819 : _T_2824; // @[Mux.scala 31:69:@18040.4]
  assign _T_2826 = _T_2802 ? _T_2817 : _T_2825; // @[Mux.scala 31:69:@18041.4]
  assign _T_2827 = _T_2801 ? _T_2815 : _T_2826; // @[Mux.scala 31:69:@18042.4]
  assign _T_2828 = _T_2800 ? _T_2813 : _T_2827; // @[Mux.scala 31:69:@18043.4]
  assign _T_2829 = _T_2799 ? _T_2811 : _T_2828; // @[Mux.scala 31:69:@18044.4]
  assign _T_2830 = _T_2798 ? _T_2809 : _T_2829; // @[Mux.scala 31:69:@18045.4]
  assign _T_2831 = _T_2797 ? _T_2807 : _T_2830; // @[Mux.scala 31:69:@18046.4]
  assign _T_2836 = io_rPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@18053.4]
  assign _T_2839 = _T_2836 & _T_1182; // @[MemPrimitives.scala 110:228:@18055.4]
  assign _T_2842 = io_rPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@18057.4]
  assign _T_2845 = _T_2842 & _T_1188; // @[MemPrimitives.scala 110:228:@18059.4]
  assign _T_2848 = io_rPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@18061.4]
  assign _T_2851 = _T_2848 & _T_1194; // @[MemPrimitives.scala 110:228:@18063.4]
  assign _T_2854 = io_rPort_4_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@18065.4]
  assign _T_2857 = _T_2854 & _T_1200; // @[MemPrimitives.scala 110:228:@18067.4]
  assign _T_2860 = io_rPort_8_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@18069.4]
  assign _T_2863 = _T_2860 & _T_1206; // @[MemPrimitives.scala 110:228:@18071.4]
  assign _T_2866 = io_rPort_10_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@18073.4]
  assign _T_2869 = _T_2866 & _T_1212; // @[MemPrimitives.scala 110:228:@18075.4]
  assign _T_2872 = io_rPort_14_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@18077.4]
  assign _T_2875 = _T_2872 & _T_1218; // @[MemPrimitives.scala 110:228:@18079.4]
  assign _T_2878 = io_rPort_15_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@18081.4]
  assign _T_2881 = _T_2878 & _T_1224; // @[MemPrimitives.scala 110:228:@18083.4]
  assign _T_2884 = io_rPort_17_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@18085.4]
  assign _T_2887 = _T_2884 & _T_1230; // @[MemPrimitives.scala 110:228:@18087.4]
  assign _T_2889 = StickySelects_18_io_outs_0; // @[MemPrimitives.scala 123:41:@18101.4]
  assign _T_2890 = StickySelects_18_io_outs_1; // @[MemPrimitives.scala 123:41:@18102.4]
  assign _T_2891 = StickySelects_18_io_outs_2; // @[MemPrimitives.scala 123:41:@18103.4]
  assign _T_2892 = StickySelects_18_io_outs_3; // @[MemPrimitives.scala 123:41:@18104.4]
  assign _T_2893 = StickySelects_18_io_outs_4; // @[MemPrimitives.scala 123:41:@18105.4]
  assign _T_2894 = StickySelects_18_io_outs_5; // @[MemPrimitives.scala 123:41:@18106.4]
  assign _T_2895 = StickySelects_18_io_outs_6; // @[MemPrimitives.scala 123:41:@18107.4]
  assign _T_2896 = StickySelects_18_io_outs_7; // @[MemPrimitives.scala 123:41:@18108.4]
  assign _T_2897 = StickySelects_18_io_outs_8; // @[MemPrimitives.scala 123:41:@18109.4]
  assign _T_2899 = {_T_2889,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@18111.4]
  assign _T_2901 = {_T_2890,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@18113.4]
  assign _T_2903 = {_T_2891,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@18115.4]
  assign _T_2905 = {_T_2892,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@18117.4]
  assign _T_2907 = {_T_2893,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@18119.4]
  assign _T_2909 = {_T_2894,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@18121.4]
  assign _T_2911 = {_T_2895,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@18123.4]
  assign _T_2913 = {_T_2896,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@18125.4]
  assign _T_2915 = {_T_2897,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@18127.4]
  assign _T_2916 = _T_2896 ? _T_2913 : _T_2915; // @[Mux.scala 31:69:@18128.4]
  assign _T_2917 = _T_2895 ? _T_2911 : _T_2916; // @[Mux.scala 31:69:@18129.4]
  assign _T_2918 = _T_2894 ? _T_2909 : _T_2917; // @[Mux.scala 31:69:@18130.4]
  assign _T_2919 = _T_2893 ? _T_2907 : _T_2918; // @[Mux.scala 31:69:@18131.4]
  assign _T_2920 = _T_2892 ? _T_2905 : _T_2919; // @[Mux.scala 31:69:@18132.4]
  assign _T_2921 = _T_2891 ? _T_2903 : _T_2920; // @[Mux.scala 31:69:@18133.4]
  assign _T_2922 = _T_2890 ? _T_2901 : _T_2921; // @[Mux.scala 31:69:@18134.4]
  assign _T_2923 = _T_2889 ? _T_2899 : _T_2922; // @[Mux.scala 31:69:@18135.4]
  assign _T_2928 = io_rPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@18142.4]
  assign _T_2931 = _T_2928 & _T_1274; // @[MemPrimitives.scala 110:228:@18144.4]
  assign _T_2934 = io_rPort_5_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@18146.4]
  assign _T_2937 = _T_2934 & _T_1280; // @[MemPrimitives.scala 110:228:@18148.4]
  assign _T_2940 = io_rPort_6_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@18150.4]
  assign _T_2943 = _T_2940 & _T_1286; // @[MemPrimitives.scala 110:228:@18152.4]
  assign _T_2946 = io_rPort_7_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@18154.4]
  assign _T_2949 = _T_2946 & _T_1292; // @[MemPrimitives.scala 110:228:@18156.4]
  assign _T_2952 = io_rPort_9_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@18158.4]
  assign _T_2955 = _T_2952 & _T_1298; // @[MemPrimitives.scala 110:228:@18160.4]
  assign _T_2958 = io_rPort_11_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@18162.4]
  assign _T_2961 = _T_2958 & _T_1304; // @[MemPrimitives.scala 110:228:@18164.4]
  assign _T_2964 = io_rPort_12_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@18166.4]
  assign _T_2967 = _T_2964 & _T_1310; // @[MemPrimitives.scala 110:228:@18168.4]
  assign _T_2970 = io_rPort_13_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@18170.4]
  assign _T_2973 = _T_2970 & _T_1316; // @[MemPrimitives.scala 110:228:@18172.4]
  assign _T_2976 = io_rPort_16_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@18174.4]
  assign _T_2979 = _T_2976 & _T_1322; // @[MemPrimitives.scala 110:228:@18176.4]
  assign _T_2981 = StickySelects_19_io_outs_0; // @[MemPrimitives.scala 123:41:@18190.4]
  assign _T_2982 = StickySelects_19_io_outs_1; // @[MemPrimitives.scala 123:41:@18191.4]
  assign _T_2983 = StickySelects_19_io_outs_2; // @[MemPrimitives.scala 123:41:@18192.4]
  assign _T_2984 = StickySelects_19_io_outs_3; // @[MemPrimitives.scala 123:41:@18193.4]
  assign _T_2985 = StickySelects_19_io_outs_4; // @[MemPrimitives.scala 123:41:@18194.4]
  assign _T_2986 = StickySelects_19_io_outs_5; // @[MemPrimitives.scala 123:41:@18195.4]
  assign _T_2987 = StickySelects_19_io_outs_6; // @[MemPrimitives.scala 123:41:@18196.4]
  assign _T_2988 = StickySelects_19_io_outs_7; // @[MemPrimitives.scala 123:41:@18197.4]
  assign _T_2989 = StickySelects_19_io_outs_8; // @[MemPrimitives.scala 123:41:@18198.4]
  assign _T_2991 = {_T_2981,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@18200.4]
  assign _T_2993 = {_T_2982,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@18202.4]
  assign _T_2995 = {_T_2983,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@18204.4]
  assign _T_2997 = {_T_2984,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@18206.4]
  assign _T_2999 = {_T_2985,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@18208.4]
  assign _T_3001 = {_T_2986,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@18210.4]
  assign _T_3003 = {_T_2987,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@18212.4]
  assign _T_3005 = {_T_2988,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@18214.4]
  assign _T_3007 = {_T_2989,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@18216.4]
  assign _T_3008 = _T_2988 ? _T_3005 : _T_3007; // @[Mux.scala 31:69:@18217.4]
  assign _T_3009 = _T_2987 ? _T_3003 : _T_3008; // @[Mux.scala 31:69:@18218.4]
  assign _T_3010 = _T_2986 ? _T_3001 : _T_3009; // @[Mux.scala 31:69:@18219.4]
  assign _T_3011 = _T_2985 ? _T_2999 : _T_3010; // @[Mux.scala 31:69:@18220.4]
  assign _T_3012 = _T_2984 ? _T_2997 : _T_3011; // @[Mux.scala 31:69:@18221.4]
  assign _T_3013 = _T_2983 ? _T_2995 : _T_3012; // @[Mux.scala 31:69:@18222.4]
  assign _T_3014 = _T_2982 ? _T_2993 : _T_3013; // @[Mux.scala 31:69:@18223.4]
  assign _T_3015 = _T_2981 ? _T_2991 : _T_3014; // @[Mux.scala 31:69:@18224.4]
  assign _T_3023 = _T_2836 & _T_1366; // @[MemPrimitives.scala 110:228:@18233.4]
  assign _T_3029 = _T_2842 & _T_1372; // @[MemPrimitives.scala 110:228:@18237.4]
  assign _T_3035 = _T_2848 & _T_1378; // @[MemPrimitives.scala 110:228:@18241.4]
  assign _T_3041 = _T_2854 & _T_1384; // @[MemPrimitives.scala 110:228:@18245.4]
  assign _T_3047 = _T_2860 & _T_1390; // @[MemPrimitives.scala 110:228:@18249.4]
  assign _T_3053 = _T_2866 & _T_1396; // @[MemPrimitives.scala 110:228:@18253.4]
  assign _T_3059 = _T_2872 & _T_1402; // @[MemPrimitives.scala 110:228:@18257.4]
  assign _T_3065 = _T_2878 & _T_1408; // @[MemPrimitives.scala 110:228:@18261.4]
  assign _T_3071 = _T_2884 & _T_1414; // @[MemPrimitives.scala 110:228:@18265.4]
  assign _T_3073 = StickySelects_20_io_outs_0; // @[MemPrimitives.scala 123:41:@18279.4]
  assign _T_3074 = StickySelects_20_io_outs_1; // @[MemPrimitives.scala 123:41:@18280.4]
  assign _T_3075 = StickySelects_20_io_outs_2; // @[MemPrimitives.scala 123:41:@18281.4]
  assign _T_3076 = StickySelects_20_io_outs_3; // @[MemPrimitives.scala 123:41:@18282.4]
  assign _T_3077 = StickySelects_20_io_outs_4; // @[MemPrimitives.scala 123:41:@18283.4]
  assign _T_3078 = StickySelects_20_io_outs_5; // @[MemPrimitives.scala 123:41:@18284.4]
  assign _T_3079 = StickySelects_20_io_outs_6; // @[MemPrimitives.scala 123:41:@18285.4]
  assign _T_3080 = StickySelects_20_io_outs_7; // @[MemPrimitives.scala 123:41:@18286.4]
  assign _T_3081 = StickySelects_20_io_outs_8; // @[MemPrimitives.scala 123:41:@18287.4]
  assign _T_3083 = {_T_3073,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@18289.4]
  assign _T_3085 = {_T_3074,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@18291.4]
  assign _T_3087 = {_T_3075,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@18293.4]
  assign _T_3089 = {_T_3076,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@18295.4]
  assign _T_3091 = {_T_3077,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@18297.4]
  assign _T_3093 = {_T_3078,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@18299.4]
  assign _T_3095 = {_T_3079,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@18301.4]
  assign _T_3097 = {_T_3080,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@18303.4]
  assign _T_3099 = {_T_3081,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@18305.4]
  assign _T_3100 = _T_3080 ? _T_3097 : _T_3099; // @[Mux.scala 31:69:@18306.4]
  assign _T_3101 = _T_3079 ? _T_3095 : _T_3100; // @[Mux.scala 31:69:@18307.4]
  assign _T_3102 = _T_3078 ? _T_3093 : _T_3101; // @[Mux.scala 31:69:@18308.4]
  assign _T_3103 = _T_3077 ? _T_3091 : _T_3102; // @[Mux.scala 31:69:@18309.4]
  assign _T_3104 = _T_3076 ? _T_3089 : _T_3103; // @[Mux.scala 31:69:@18310.4]
  assign _T_3105 = _T_3075 ? _T_3087 : _T_3104; // @[Mux.scala 31:69:@18311.4]
  assign _T_3106 = _T_3074 ? _T_3085 : _T_3105; // @[Mux.scala 31:69:@18312.4]
  assign _T_3107 = _T_3073 ? _T_3083 : _T_3106; // @[Mux.scala 31:69:@18313.4]
  assign _T_3115 = _T_2928 & _T_1458; // @[MemPrimitives.scala 110:228:@18322.4]
  assign _T_3121 = _T_2934 & _T_1464; // @[MemPrimitives.scala 110:228:@18326.4]
  assign _T_3127 = _T_2940 & _T_1470; // @[MemPrimitives.scala 110:228:@18330.4]
  assign _T_3133 = _T_2946 & _T_1476; // @[MemPrimitives.scala 110:228:@18334.4]
  assign _T_3139 = _T_2952 & _T_1482; // @[MemPrimitives.scala 110:228:@18338.4]
  assign _T_3145 = _T_2958 & _T_1488; // @[MemPrimitives.scala 110:228:@18342.4]
  assign _T_3151 = _T_2964 & _T_1494; // @[MemPrimitives.scala 110:228:@18346.4]
  assign _T_3157 = _T_2970 & _T_1500; // @[MemPrimitives.scala 110:228:@18350.4]
  assign _T_3163 = _T_2976 & _T_1506; // @[MemPrimitives.scala 110:228:@18354.4]
  assign _T_3165 = StickySelects_21_io_outs_0; // @[MemPrimitives.scala 123:41:@18368.4]
  assign _T_3166 = StickySelects_21_io_outs_1; // @[MemPrimitives.scala 123:41:@18369.4]
  assign _T_3167 = StickySelects_21_io_outs_2; // @[MemPrimitives.scala 123:41:@18370.4]
  assign _T_3168 = StickySelects_21_io_outs_3; // @[MemPrimitives.scala 123:41:@18371.4]
  assign _T_3169 = StickySelects_21_io_outs_4; // @[MemPrimitives.scala 123:41:@18372.4]
  assign _T_3170 = StickySelects_21_io_outs_5; // @[MemPrimitives.scala 123:41:@18373.4]
  assign _T_3171 = StickySelects_21_io_outs_6; // @[MemPrimitives.scala 123:41:@18374.4]
  assign _T_3172 = StickySelects_21_io_outs_7; // @[MemPrimitives.scala 123:41:@18375.4]
  assign _T_3173 = StickySelects_21_io_outs_8; // @[MemPrimitives.scala 123:41:@18376.4]
  assign _T_3175 = {_T_3165,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@18378.4]
  assign _T_3177 = {_T_3166,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@18380.4]
  assign _T_3179 = {_T_3167,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@18382.4]
  assign _T_3181 = {_T_3168,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@18384.4]
  assign _T_3183 = {_T_3169,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@18386.4]
  assign _T_3185 = {_T_3170,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@18388.4]
  assign _T_3187 = {_T_3171,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@18390.4]
  assign _T_3189 = {_T_3172,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@18392.4]
  assign _T_3191 = {_T_3173,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@18394.4]
  assign _T_3192 = _T_3172 ? _T_3189 : _T_3191; // @[Mux.scala 31:69:@18395.4]
  assign _T_3193 = _T_3171 ? _T_3187 : _T_3192; // @[Mux.scala 31:69:@18396.4]
  assign _T_3194 = _T_3170 ? _T_3185 : _T_3193; // @[Mux.scala 31:69:@18397.4]
  assign _T_3195 = _T_3169 ? _T_3183 : _T_3194; // @[Mux.scala 31:69:@18398.4]
  assign _T_3196 = _T_3168 ? _T_3181 : _T_3195; // @[Mux.scala 31:69:@18399.4]
  assign _T_3197 = _T_3167 ? _T_3179 : _T_3196; // @[Mux.scala 31:69:@18400.4]
  assign _T_3198 = _T_3166 ? _T_3177 : _T_3197; // @[Mux.scala 31:69:@18401.4]
  assign _T_3199 = _T_3165 ? _T_3175 : _T_3198; // @[Mux.scala 31:69:@18402.4]
  assign _T_3207 = _T_2836 & _T_1550; // @[MemPrimitives.scala 110:228:@18411.4]
  assign _T_3213 = _T_2842 & _T_1556; // @[MemPrimitives.scala 110:228:@18415.4]
  assign _T_3219 = _T_2848 & _T_1562; // @[MemPrimitives.scala 110:228:@18419.4]
  assign _T_3225 = _T_2854 & _T_1568; // @[MemPrimitives.scala 110:228:@18423.4]
  assign _T_3231 = _T_2860 & _T_1574; // @[MemPrimitives.scala 110:228:@18427.4]
  assign _T_3237 = _T_2866 & _T_1580; // @[MemPrimitives.scala 110:228:@18431.4]
  assign _T_3243 = _T_2872 & _T_1586; // @[MemPrimitives.scala 110:228:@18435.4]
  assign _T_3249 = _T_2878 & _T_1592; // @[MemPrimitives.scala 110:228:@18439.4]
  assign _T_3255 = _T_2884 & _T_1598; // @[MemPrimitives.scala 110:228:@18443.4]
  assign _T_3257 = StickySelects_22_io_outs_0; // @[MemPrimitives.scala 123:41:@18457.4]
  assign _T_3258 = StickySelects_22_io_outs_1; // @[MemPrimitives.scala 123:41:@18458.4]
  assign _T_3259 = StickySelects_22_io_outs_2; // @[MemPrimitives.scala 123:41:@18459.4]
  assign _T_3260 = StickySelects_22_io_outs_3; // @[MemPrimitives.scala 123:41:@18460.4]
  assign _T_3261 = StickySelects_22_io_outs_4; // @[MemPrimitives.scala 123:41:@18461.4]
  assign _T_3262 = StickySelects_22_io_outs_5; // @[MemPrimitives.scala 123:41:@18462.4]
  assign _T_3263 = StickySelects_22_io_outs_6; // @[MemPrimitives.scala 123:41:@18463.4]
  assign _T_3264 = StickySelects_22_io_outs_7; // @[MemPrimitives.scala 123:41:@18464.4]
  assign _T_3265 = StickySelects_22_io_outs_8; // @[MemPrimitives.scala 123:41:@18465.4]
  assign _T_3267 = {_T_3257,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@18467.4]
  assign _T_3269 = {_T_3258,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@18469.4]
  assign _T_3271 = {_T_3259,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@18471.4]
  assign _T_3273 = {_T_3260,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@18473.4]
  assign _T_3275 = {_T_3261,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@18475.4]
  assign _T_3277 = {_T_3262,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@18477.4]
  assign _T_3279 = {_T_3263,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@18479.4]
  assign _T_3281 = {_T_3264,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@18481.4]
  assign _T_3283 = {_T_3265,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@18483.4]
  assign _T_3284 = _T_3264 ? _T_3281 : _T_3283; // @[Mux.scala 31:69:@18484.4]
  assign _T_3285 = _T_3263 ? _T_3279 : _T_3284; // @[Mux.scala 31:69:@18485.4]
  assign _T_3286 = _T_3262 ? _T_3277 : _T_3285; // @[Mux.scala 31:69:@18486.4]
  assign _T_3287 = _T_3261 ? _T_3275 : _T_3286; // @[Mux.scala 31:69:@18487.4]
  assign _T_3288 = _T_3260 ? _T_3273 : _T_3287; // @[Mux.scala 31:69:@18488.4]
  assign _T_3289 = _T_3259 ? _T_3271 : _T_3288; // @[Mux.scala 31:69:@18489.4]
  assign _T_3290 = _T_3258 ? _T_3269 : _T_3289; // @[Mux.scala 31:69:@18490.4]
  assign _T_3291 = _T_3257 ? _T_3267 : _T_3290; // @[Mux.scala 31:69:@18491.4]
  assign _T_3299 = _T_2928 & _T_1642; // @[MemPrimitives.scala 110:228:@18500.4]
  assign _T_3305 = _T_2934 & _T_1648; // @[MemPrimitives.scala 110:228:@18504.4]
  assign _T_3311 = _T_2940 & _T_1654; // @[MemPrimitives.scala 110:228:@18508.4]
  assign _T_3317 = _T_2946 & _T_1660; // @[MemPrimitives.scala 110:228:@18512.4]
  assign _T_3323 = _T_2952 & _T_1666; // @[MemPrimitives.scala 110:228:@18516.4]
  assign _T_3329 = _T_2958 & _T_1672; // @[MemPrimitives.scala 110:228:@18520.4]
  assign _T_3335 = _T_2964 & _T_1678; // @[MemPrimitives.scala 110:228:@18524.4]
  assign _T_3341 = _T_2970 & _T_1684; // @[MemPrimitives.scala 110:228:@18528.4]
  assign _T_3347 = _T_2976 & _T_1690; // @[MemPrimitives.scala 110:228:@18532.4]
  assign _T_3349 = StickySelects_23_io_outs_0; // @[MemPrimitives.scala 123:41:@18546.4]
  assign _T_3350 = StickySelects_23_io_outs_1; // @[MemPrimitives.scala 123:41:@18547.4]
  assign _T_3351 = StickySelects_23_io_outs_2; // @[MemPrimitives.scala 123:41:@18548.4]
  assign _T_3352 = StickySelects_23_io_outs_3; // @[MemPrimitives.scala 123:41:@18549.4]
  assign _T_3353 = StickySelects_23_io_outs_4; // @[MemPrimitives.scala 123:41:@18550.4]
  assign _T_3354 = StickySelects_23_io_outs_5; // @[MemPrimitives.scala 123:41:@18551.4]
  assign _T_3355 = StickySelects_23_io_outs_6; // @[MemPrimitives.scala 123:41:@18552.4]
  assign _T_3356 = StickySelects_23_io_outs_7; // @[MemPrimitives.scala 123:41:@18553.4]
  assign _T_3357 = StickySelects_23_io_outs_8; // @[MemPrimitives.scala 123:41:@18554.4]
  assign _T_3359 = {_T_3349,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@18556.4]
  assign _T_3361 = {_T_3350,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@18558.4]
  assign _T_3363 = {_T_3351,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@18560.4]
  assign _T_3365 = {_T_3352,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@18562.4]
  assign _T_3367 = {_T_3353,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@18564.4]
  assign _T_3369 = {_T_3354,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@18566.4]
  assign _T_3371 = {_T_3355,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@18568.4]
  assign _T_3373 = {_T_3356,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@18570.4]
  assign _T_3375 = {_T_3357,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@18572.4]
  assign _T_3376 = _T_3356 ? _T_3373 : _T_3375; // @[Mux.scala 31:69:@18573.4]
  assign _T_3377 = _T_3355 ? _T_3371 : _T_3376; // @[Mux.scala 31:69:@18574.4]
  assign _T_3378 = _T_3354 ? _T_3369 : _T_3377; // @[Mux.scala 31:69:@18575.4]
  assign _T_3379 = _T_3353 ? _T_3367 : _T_3378; // @[Mux.scala 31:69:@18576.4]
  assign _T_3380 = _T_3352 ? _T_3365 : _T_3379; // @[Mux.scala 31:69:@18577.4]
  assign _T_3381 = _T_3351 ? _T_3363 : _T_3380; // @[Mux.scala 31:69:@18578.4]
  assign _T_3382 = _T_3350 ? _T_3361 : _T_3381; // @[Mux.scala 31:69:@18579.4]
  assign _T_3383 = _T_3349 ? _T_3359 : _T_3382; // @[Mux.scala 31:69:@18580.4]
  assign _T_3479 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@18709.4 package.scala 96:25:@18710.4]
  assign _T_3483 = _T_3479 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@18719.4]
  assign _T_3476 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@18701.4 package.scala 96:25:@18702.4]
  assign _T_3484 = _T_3476 ? Mem1D_18_io_output : _T_3483; // @[Mux.scala 31:69:@18720.4]
  assign _T_3473 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@18693.4 package.scala 96:25:@18694.4]
  assign _T_3485 = _T_3473 ? Mem1D_16_io_output : _T_3484; // @[Mux.scala 31:69:@18721.4]
  assign _T_3470 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@18685.4 package.scala 96:25:@18686.4]
  assign _T_3486 = _T_3470 ? Mem1D_14_io_output : _T_3485; // @[Mux.scala 31:69:@18722.4]
  assign _T_3467 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@18677.4 package.scala 96:25:@18678.4]
  assign _T_3487 = _T_3467 ? Mem1D_12_io_output : _T_3486; // @[Mux.scala 31:69:@18723.4]
  assign _T_3464 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@18669.4 package.scala 96:25:@18670.4]
  assign _T_3488 = _T_3464 ? Mem1D_10_io_output : _T_3487; // @[Mux.scala 31:69:@18724.4]
  assign _T_3461 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@18661.4 package.scala 96:25:@18662.4]
  assign _T_3489 = _T_3461 ? Mem1D_8_io_output : _T_3488; // @[Mux.scala 31:69:@18725.4]
  assign _T_3458 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@18653.4 package.scala 96:25:@18654.4]
  assign _T_3490 = _T_3458 ? Mem1D_6_io_output : _T_3489; // @[Mux.scala 31:69:@18726.4]
  assign _T_3455 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@18645.4 package.scala 96:25:@18646.4]
  assign _T_3491 = _T_3455 ? Mem1D_4_io_output : _T_3490; // @[Mux.scala 31:69:@18727.4]
  assign _T_3452 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@18637.4 package.scala 96:25:@18638.4]
  assign _T_3492 = _T_3452 ? Mem1D_2_io_output : _T_3491; // @[Mux.scala 31:69:@18728.4]
  assign _T_3449 = RetimeWrapper_io_out; // @[package.scala 96:25:@18629.4 package.scala 96:25:@18630.4]
  assign _T_3586 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@18853.4 package.scala 96:25:@18854.4]
  assign _T_3590 = _T_3586 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@18863.4]
  assign _T_3583 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@18845.4 package.scala 96:25:@18846.4]
  assign _T_3591 = _T_3583 ? Mem1D_18_io_output : _T_3590; // @[Mux.scala 31:69:@18864.4]
  assign _T_3580 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@18837.4 package.scala 96:25:@18838.4]
  assign _T_3592 = _T_3580 ? Mem1D_16_io_output : _T_3591; // @[Mux.scala 31:69:@18865.4]
  assign _T_3577 = RetimeWrapper_19_io_out; // @[package.scala 96:25:@18829.4 package.scala 96:25:@18830.4]
  assign _T_3593 = _T_3577 ? Mem1D_14_io_output : _T_3592; // @[Mux.scala 31:69:@18866.4]
  assign _T_3574 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@18821.4 package.scala 96:25:@18822.4]
  assign _T_3594 = _T_3574 ? Mem1D_12_io_output : _T_3593; // @[Mux.scala 31:69:@18867.4]
  assign _T_3571 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@18813.4 package.scala 96:25:@18814.4]
  assign _T_3595 = _T_3571 ? Mem1D_10_io_output : _T_3594; // @[Mux.scala 31:69:@18868.4]
  assign _T_3568 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@18805.4 package.scala 96:25:@18806.4]
  assign _T_3596 = _T_3568 ? Mem1D_8_io_output : _T_3595; // @[Mux.scala 31:69:@18869.4]
  assign _T_3565 = RetimeWrapper_15_io_out; // @[package.scala 96:25:@18797.4 package.scala 96:25:@18798.4]
  assign _T_3597 = _T_3565 ? Mem1D_6_io_output : _T_3596; // @[Mux.scala 31:69:@18870.4]
  assign _T_3562 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@18789.4 package.scala 96:25:@18790.4]
  assign _T_3598 = _T_3562 ? Mem1D_4_io_output : _T_3597; // @[Mux.scala 31:69:@18871.4]
  assign _T_3559 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@18781.4 package.scala 96:25:@18782.4]
  assign _T_3599 = _T_3559 ? Mem1D_2_io_output : _T_3598; // @[Mux.scala 31:69:@18872.4]
  assign _T_3556 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@18773.4 package.scala 96:25:@18774.4]
  assign _T_3693 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@18997.4 package.scala 96:25:@18998.4]
  assign _T_3697 = _T_3693 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@19007.4]
  assign _T_3690 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@18989.4 package.scala 96:25:@18990.4]
  assign _T_3698 = _T_3690 ? Mem1D_19_io_output : _T_3697; // @[Mux.scala 31:69:@19008.4]
  assign _T_3687 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@18981.4 package.scala 96:25:@18982.4]
  assign _T_3699 = _T_3687 ? Mem1D_17_io_output : _T_3698; // @[Mux.scala 31:69:@19009.4]
  assign _T_3684 = RetimeWrapper_31_io_out; // @[package.scala 96:25:@18973.4 package.scala 96:25:@18974.4]
  assign _T_3700 = _T_3684 ? Mem1D_15_io_output : _T_3699; // @[Mux.scala 31:69:@19010.4]
  assign _T_3681 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@18965.4 package.scala 96:25:@18966.4]
  assign _T_3701 = _T_3681 ? Mem1D_13_io_output : _T_3700; // @[Mux.scala 31:69:@19011.4]
  assign _T_3678 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@18957.4 package.scala 96:25:@18958.4]
  assign _T_3702 = _T_3678 ? Mem1D_11_io_output : _T_3701; // @[Mux.scala 31:69:@19012.4]
  assign _T_3675 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@18949.4 package.scala 96:25:@18950.4]
  assign _T_3703 = _T_3675 ? Mem1D_9_io_output : _T_3702; // @[Mux.scala 31:69:@19013.4]
  assign _T_3672 = RetimeWrapper_27_io_out; // @[package.scala 96:25:@18941.4 package.scala 96:25:@18942.4]
  assign _T_3704 = _T_3672 ? Mem1D_7_io_output : _T_3703; // @[Mux.scala 31:69:@19014.4]
  assign _T_3669 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@18933.4 package.scala 96:25:@18934.4]
  assign _T_3705 = _T_3669 ? Mem1D_5_io_output : _T_3704; // @[Mux.scala 31:69:@19015.4]
  assign _T_3666 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@18925.4 package.scala 96:25:@18926.4]
  assign _T_3706 = _T_3666 ? Mem1D_3_io_output : _T_3705; // @[Mux.scala 31:69:@19016.4]
  assign _T_3663 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@18917.4 package.scala 96:25:@18918.4]
  assign _T_3800 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@19141.4 package.scala 96:25:@19142.4]
  assign _T_3804 = _T_3800 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@19151.4]
  assign _T_3797 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@19133.4 package.scala 96:25:@19134.4]
  assign _T_3805 = _T_3797 ? Mem1D_18_io_output : _T_3804; // @[Mux.scala 31:69:@19152.4]
  assign _T_3794 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@19125.4 package.scala 96:25:@19126.4]
  assign _T_3806 = _T_3794 ? Mem1D_16_io_output : _T_3805; // @[Mux.scala 31:69:@19153.4]
  assign _T_3791 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@19117.4 package.scala 96:25:@19118.4]
  assign _T_3807 = _T_3791 ? Mem1D_14_io_output : _T_3806; // @[Mux.scala 31:69:@19154.4]
  assign _T_3788 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@19109.4 package.scala 96:25:@19110.4]
  assign _T_3808 = _T_3788 ? Mem1D_12_io_output : _T_3807; // @[Mux.scala 31:69:@19155.4]
  assign _T_3785 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@19101.4 package.scala 96:25:@19102.4]
  assign _T_3809 = _T_3785 ? Mem1D_10_io_output : _T_3808; // @[Mux.scala 31:69:@19156.4]
  assign _T_3782 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@19093.4 package.scala 96:25:@19094.4]
  assign _T_3810 = _T_3782 ? Mem1D_8_io_output : _T_3809; // @[Mux.scala 31:69:@19157.4]
  assign _T_3779 = RetimeWrapper_39_io_out; // @[package.scala 96:25:@19085.4 package.scala 96:25:@19086.4]
  assign _T_3811 = _T_3779 ? Mem1D_6_io_output : _T_3810; // @[Mux.scala 31:69:@19158.4]
  assign _T_3776 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@19077.4 package.scala 96:25:@19078.4]
  assign _T_3812 = _T_3776 ? Mem1D_4_io_output : _T_3811; // @[Mux.scala 31:69:@19159.4]
  assign _T_3773 = RetimeWrapper_37_io_out; // @[package.scala 96:25:@19069.4 package.scala 96:25:@19070.4]
  assign _T_3813 = _T_3773 ? Mem1D_2_io_output : _T_3812; // @[Mux.scala 31:69:@19160.4]
  assign _T_3770 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@19061.4 package.scala 96:25:@19062.4]
  assign _T_3907 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@19285.4 package.scala 96:25:@19286.4]
  assign _T_3911 = _T_3907 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@19295.4]
  assign _T_3904 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@19277.4 package.scala 96:25:@19278.4]
  assign _T_3912 = _T_3904 ? Mem1D_18_io_output : _T_3911; // @[Mux.scala 31:69:@19296.4]
  assign _T_3901 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@19269.4 package.scala 96:25:@19270.4]
  assign _T_3913 = _T_3901 ? Mem1D_16_io_output : _T_3912; // @[Mux.scala 31:69:@19297.4]
  assign _T_3898 = RetimeWrapper_55_io_out; // @[package.scala 96:25:@19261.4 package.scala 96:25:@19262.4]
  assign _T_3914 = _T_3898 ? Mem1D_14_io_output : _T_3913; // @[Mux.scala 31:69:@19298.4]
  assign _T_3895 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@19253.4 package.scala 96:25:@19254.4]
  assign _T_3915 = _T_3895 ? Mem1D_12_io_output : _T_3914; // @[Mux.scala 31:69:@19299.4]
  assign _T_3892 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@19245.4 package.scala 96:25:@19246.4]
  assign _T_3916 = _T_3892 ? Mem1D_10_io_output : _T_3915; // @[Mux.scala 31:69:@19300.4]
  assign _T_3889 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@19237.4 package.scala 96:25:@19238.4]
  assign _T_3917 = _T_3889 ? Mem1D_8_io_output : _T_3916; // @[Mux.scala 31:69:@19301.4]
  assign _T_3886 = RetimeWrapper_51_io_out; // @[package.scala 96:25:@19229.4 package.scala 96:25:@19230.4]
  assign _T_3918 = _T_3886 ? Mem1D_6_io_output : _T_3917; // @[Mux.scala 31:69:@19302.4]
  assign _T_3883 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@19221.4 package.scala 96:25:@19222.4]
  assign _T_3919 = _T_3883 ? Mem1D_4_io_output : _T_3918; // @[Mux.scala 31:69:@19303.4]
  assign _T_3880 = RetimeWrapper_49_io_out; // @[package.scala 96:25:@19213.4 package.scala 96:25:@19214.4]
  assign _T_3920 = _T_3880 ? Mem1D_2_io_output : _T_3919; // @[Mux.scala 31:69:@19304.4]
  assign _T_3877 = RetimeWrapper_48_io_out; // @[package.scala 96:25:@19205.4 package.scala 96:25:@19206.4]
  assign _T_4014 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@19429.4 package.scala 96:25:@19430.4]
  assign _T_4018 = _T_4014 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@19439.4]
  assign _T_4011 = RetimeWrapper_69_io_out; // @[package.scala 96:25:@19421.4 package.scala 96:25:@19422.4]
  assign _T_4019 = _T_4011 ? Mem1D_19_io_output : _T_4018; // @[Mux.scala 31:69:@19440.4]
  assign _T_4008 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@19413.4 package.scala 96:25:@19414.4]
  assign _T_4020 = _T_4008 ? Mem1D_17_io_output : _T_4019; // @[Mux.scala 31:69:@19441.4]
  assign _T_4005 = RetimeWrapper_67_io_out; // @[package.scala 96:25:@19405.4 package.scala 96:25:@19406.4]
  assign _T_4021 = _T_4005 ? Mem1D_15_io_output : _T_4020; // @[Mux.scala 31:69:@19442.4]
  assign _T_4002 = RetimeWrapper_66_io_out; // @[package.scala 96:25:@19397.4 package.scala 96:25:@19398.4]
  assign _T_4022 = _T_4002 ? Mem1D_13_io_output : _T_4021; // @[Mux.scala 31:69:@19443.4]
  assign _T_3999 = RetimeWrapper_65_io_out; // @[package.scala 96:25:@19389.4 package.scala 96:25:@19390.4]
  assign _T_4023 = _T_3999 ? Mem1D_11_io_output : _T_4022; // @[Mux.scala 31:69:@19444.4]
  assign _T_3996 = RetimeWrapper_64_io_out; // @[package.scala 96:25:@19381.4 package.scala 96:25:@19382.4]
  assign _T_4024 = _T_3996 ? Mem1D_9_io_output : _T_4023; // @[Mux.scala 31:69:@19445.4]
  assign _T_3993 = RetimeWrapper_63_io_out; // @[package.scala 96:25:@19373.4 package.scala 96:25:@19374.4]
  assign _T_4025 = _T_3993 ? Mem1D_7_io_output : _T_4024; // @[Mux.scala 31:69:@19446.4]
  assign _T_3990 = RetimeWrapper_62_io_out; // @[package.scala 96:25:@19365.4 package.scala 96:25:@19366.4]
  assign _T_4026 = _T_3990 ? Mem1D_5_io_output : _T_4025; // @[Mux.scala 31:69:@19447.4]
  assign _T_3987 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@19357.4 package.scala 96:25:@19358.4]
  assign _T_4027 = _T_3987 ? Mem1D_3_io_output : _T_4026; // @[Mux.scala 31:69:@19448.4]
  assign _T_3984 = RetimeWrapper_60_io_out; // @[package.scala 96:25:@19349.4 package.scala 96:25:@19350.4]
  assign _T_4121 = RetimeWrapper_82_io_out; // @[package.scala 96:25:@19573.4 package.scala 96:25:@19574.4]
  assign _T_4125 = _T_4121 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@19583.4]
  assign _T_4118 = RetimeWrapper_81_io_out; // @[package.scala 96:25:@19565.4 package.scala 96:25:@19566.4]
  assign _T_4126 = _T_4118 ? Mem1D_19_io_output : _T_4125; // @[Mux.scala 31:69:@19584.4]
  assign _T_4115 = RetimeWrapper_80_io_out; // @[package.scala 96:25:@19557.4 package.scala 96:25:@19558.4]
  assign _T_4127 = _T_4115 ? Mem1D_17_io_output : _T_4126; // @[Mux.scala 31:69:@19585.4]
  assign _T_4112 = RetimeWrapper_79_io_out; // @[package.scala 96:25:@19549.4 package.scala 96:25:@19550.4]
  assign _T_4128 = _T_4112 ? Mem1D_15_io_output : _T_4127; // @[Mux.scala 31:69:@19586.4]
  assign _T_4109 = RetimeWrapper_78_io_out; // @[package.scala 96:25:@19541.4 package.scala 96:25:@19542.4]
  assign _T_4129 = _T_4109 ? Mem1D_13_io_output : _T_4128; // @[Mux.scala 31:69:@19587.4]
  assign _T_4106 = RetimeWrapper_77_io_out; // @[package.scala 96:25:@19533.4 package.scala 96:25:@19534.4]
  assign _T_4130 = _T_4106 ? Mem1D_11_io_output : _T_4129; // @[Mux.scala 31:69:@19588.4]
  assign _T_4103 = RetimeWrapper_76_io_out; // @[package.scala 96:25:@19525.4 package.scala 96:25:@19526.4]
  assign _T_4131 = _T_4103 ? Mem1D_9_io_output : _T_4130; // @[Mux.scala 31:69:@19589.4]
  assign _T_4100 = RetimeWrapper_75_io_out; // @[package.scala 96:25:@19517.4 package.scala 96:25:@19518.4]
  assign _T_4132 = _T_4100 ? Mem1D_7_io_output : _T_4131; // @[Mux.scala 31:69:@19590.4]
  assign _T_4097 = RetimeWrapper_74_io_out; // @[package.scala 96:25:@19509.4 package.scala 96:25:@19510.4]
  assign _T_4133 = _T_4097 ? Mem1D_5_io_output : _T_4132; // @[Mux.scala 31:69:@19591.4]
  assign _T_4094 = RetimeWrapper_73_io_out; // @[package.scala 96:25:@19501.4 package.scala 96:25:@19502.4]
  assign _T_4134 = _T_4094 ? Mem1D_3_io_output : _T_4133; // @[Mux.scala 31:69:@19592.4]
  assign _T_4091 = RetimeWrapper_72_io_out; // @[package.scala 96:25:@19493.4 package.scala 96:25:@19494.4]
  assign _T_4228 = RetimeWrapper_94_io_out; // @[package.scala 96:25:@19717.4 package.scala 96:25:@19718.4]
  assign _T_4232 = _T_4228 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@19727.4]
  assign _T_4225 = RetimeWrapper_93_io_out; // @[package.scala 96:25:@19709.4 package.scala 96:25:@19710.4]
  assign _T_4233 = _T_4225 ? Mem1D_19_io_output : _T_4232; // @[Mux.scala 31:69:@19728.4]
  assign _T_4222 = RetimeWrapper_92_io_out; // @[package.scala 96:25:@19701.4 package.scala 96:25:@19702.4]
  assign _T_4234 = _T_4222 ? Mem1D_17_io_output : _T_4233; // @[Mux.scala 31:69:@19729.4]
  assign _T_4219 = RetimeWrapper_91_io_out; // @[package.scala 96:25:@19693.4 package.scala 96:25:@19694.4]
  assign _T_4235 = _T_4219 ? Mem1D_15_io_output : _T_4234; // @[Mux.scala 31:69:@19730.4]
  assign _T_4216 = RetimeWrapper_90_io_out; // @[package.scala 96:25:@19685.4 package.scala 96:25:@19686.4]
  assign _T_4236 = _T_4216 ? Mem1D_13_io_output : _T_4235; // @[Mux.scala 31:69:@19731.4]
  assign _T_4213 = RetimeWrapper_89_io_out; // @[package.scala 96:25:@19677.4 package.scala 96:25:@19678.4]
  assign _T_4237 = _T_4213 ? Mem1D_11_io_output : _T_4236; // @[Mux.scala 31:69:@19732.4]
  assign _T_4210 = RetimeWrapper_88_io_out; // @[package.scala 96:25:@19669.4 package.scala 96:25:@19670.4]
  assign _T_4238 = _T_4210 ? Mem1D_9_io_output : _T_4237; // @[Mux.scala 31:69:@19733.4]
  assign _T_4207 = RetimeWrapper_87_io_out; // @[package.scala 96:25:@19661.4 package.scala 96:25:@19662.4]
  assign _T_4239 = _T_4207 ? Mem1D_7_io_output : _T_4238; // @[Mux.scala 31:69:@19734.4]
  assign _T_4204 = RetimeWrapper_86_io_out; // @[package.scala 96:25:@19653.4 package.scala 96:25:@19654.4]
  assign _T_4240 = _T_4204 ? Mem1D_5_io_output : _T_4239; // @[Mux.scala 31:69:@19735.4]
  assign _T_4201 = RetimeWrapper_85_io_out; // @[package.scala 96:25:@19645.4 package.scala 96:25:@19646.4]
  assign _T_4241 = _T_4201 ? Mem1D_3_io_output : _T_4240; // @[Mux.scala 31:69:@19736.4]
  assign _T_4198 = RetimeWrapper_84_io_out; // @[package.scala 96:25:@19637.4 package.scala 96:25:@19638.4]
  assign _T_4335 = RetimeWrapper_106_io_out; // @[package.scala 96:25:@19861.4 package.scala 96:25:@19862.4]
  assign _T_4339 = _T_4335 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@19871.4]
  assign _T_4332 = RetimeWrapper_105_io_out; // @[package.scala 96:25:@19853.4 package.scala 96:25:@19854.4]
  assign _T_4340 = _T_4332 ? Mem1D_18_io_output : _T_4339; // @[Mux.scala 31:69:@19872.4]
  assign _T_4329 = RetimeWrapper_104_io_out; // @[package.scala 96:25:@19845.4 package.scala 96:25:@19846.4]
  assign _T_4341 = _T_4329 ? Mem1D_16_io_output : _T_4340; // @[Mux.scala 31:69:@19873.4]
  assign _T_4326 = RetimeWrapper_103_io_out; // @[package.scala 96:25:@19837.4 package.scala 96:25:@19838.4]
  assign _T_4342 = _T_4326 ? Mem1D_14_io_output : _T_4341; // @[Mux.scala 31:69:@19874.4]
  assign _T_4323 = RetimeWrapper_102_io_out; // @[package.scala 96:25:@19829.4 package.scala 96:25:@19830.4]
  assign _T_4343 = _T_4323 ? Mem1D_12_io_output : _T_4342; // @[Mux.scala 31:69:@19875.4]
  assign _T_4320 = RetimeWrapper_101_io_out; // @[package.scala 96:25:@19821.4 package.scala 96:25:@19822.4]
  assign _T_4344 = _T_4320 ? Mem1D_10_io_output : _T_4343; // @[Mux.scala 31:69:@19876.4]
  assign _T_4317 = RetimeWrapper_100_io_out; // @[package.scala 96:25:@19813.4 package.scala 96:25:@19814.4]
  assign _T_4345 = _T_4317 ? Mem1D_8_io_output : _T_4344; // @[Mux.scala 31:69:@19877.4]
  assign _T_4314 = RetimeWrapper_99_io_out; // @[package.scala 96:25:@19805.4 package.scala 96:25:@19806.4]
  assign _T_4346 = _T_4314 ? Mem1D_6_io_output : _T_4345; // @[Mux.scala 31:69:@19878.4]
  assign _T_4311 = RetimeWrapper_98_io_out; // @[package.scala 96:25:@19797.4 package.scala 96:25:@19798.4]
  assign _T_4347 = _T_4311 ? Mem1D_4_io_output : _T_4346; // @[Mux.scala 31:69:@19879.4]
  assign _T_4308 = RetimeWrapper_97_io_out; // @[package.scala 96:25:@19789.4 package.scala 96:25:@19790.4]
  assign _T_4348 = _T_4308 ? Mem1D_2_io_output : _T_4347; // @[Mux.scala 31:69:@19880.4]
  assign _T_4305 = RetimeWrapper_96_io_out; // @[package.scala 96:25:@19781.4 package.scala 96:25:@19782.4]
  assign _T_4442 = RetimeWrapper_118_io_out; // @[package.scala 96:25:@20005.4 package.scala 96:25:@20006.4]
  assign _T_4446 = _T_4442 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@20015.4]
  assign _T_4439 = RetimeWrapper_117_io_out; // @[package.scala 96:25:@19997.4 package.scala 96:25:@19998.4]
  assign _T_4447 = _T_4439 ? Mem1D_19_io_output : _T_4446; // @[Mux.scala 31:69:@20016.4]
  assign _T_4436 = RetimeWrapper_116_io_out; // @[package.scala 96:25:@19989.4 package.scala 96:25:@19990.4]
  assign _T_4448 = _T_4436 ? Mem1D_17_io_output : _T_4447; // @[Mux.scala 31:69:@20017.4]
  assign _T_4433 = RetimeWrapper_115_io_out; // @[package.scala 96:25:@19981.4 package.scala 96:25:@19982.4]
  assign _T_4449 = _T_4433 ? Mem1D_15_io_output : _T_4448; // @[Mux.scala 31:69:@20018.4]
  assign _T_4430 = RetimeWrapper_114_io_out; // @[package.scala 96:25:@19973.4 package.scala 96:25:@19974.4]
  assign _T_4450 = _T_4430 ? Mem1D_13_io_output : _T_4449; // @[Mux.scala 31:69:@20019.4]
  assign _T_4427 = RetimeWrapper_113_io_out; // @[package.scala 96:25:@19965.4 package.scala 96:25:@19966.4]
  assign _T_4451 = _T_4427 ? Mem1D_11_io_output : _T_4450; // @[Mux.scala 31:69:@20020.4]
  assign _T_4424 = RetimeWrapper_112_io_out; // @[package.scala 96:25:@19957.4 package.scala 96:25:@19958.4]
  assign _T_4452 = _T_4424 ? Mem1D_9_io_output : _T_4451; // @[Mux.scala 31:69:@20021.4]
  assign _T_4421 = RetimeWrapper_111_io_out; // @[package.scala 96:25:@19949.4 package.scala 96:25:@19950.4]
  assign _T_4453 = _T_4421 ? Mem1D_7_io_output : _T_4452; // @[Mux.scala 31:69:@20022.4]
  assign _T_4418 = RetimeWrapper_110_io_out; // @[package.scala 96:25:@19941.4 package.scala 96:25:@19942.4]
  assign _T_4454 = _T_4418 ? Mem1D_5_io_output : _T_4453; // @[Mux.scala 31:69:@20023.4]
  assign _T_4415 = RetimeWrapper_109_io_out; // @[package.scala 96:25:@19933.4 package.scala 96:25:@19934.4]
  assign _T_4455 = _T_4415 ? Mem1D_3_io_output : _T_4454; // @[Mux.scala 31:69:@20024.4]
  assign _T_4412 = RetimeWrapper_108_io_out; // @[package.scala 96:25:@19925.4 package.scala 96:25:@19926.4]
  assign _T_4549 = RetimeWrapper_130_io_out; // @[package.scala 96:25:@20149.4 package.scala 96:25:@20150.4]
  assign _T_4553 = _T_4549 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@20159.4]
  assign _T_4546 = RetimeWrapper_129_io_out; // @[package.scala 96:25:@20141.4 package.scala 96:25:@20142.4]
  assign _T_4554 = _T_4546 ? Mem1D_18_io_output : _T_4553; // @[Mux.scala 31:69:@20160.4]
  assign _T_4543 = RetimeWrapper_128_io_out; // @[package.scala 96:25:@20133.4 package.scala 96:25:@20134.4]
  assign _T_4555 = _T_4543 ? Mem1D_16_io_output : _T_4554; // @[Mux.scala 31:69:@20161.4]
  assign _T_4540 = RetimeWrapper_127_io_out; // @[package.scala 96:25:@20125.4 package.scala 96:25:@20126.4]
  assign _T_4556 = _T_4540 ? Mem1D_14_io_output : _T_4555; // @[Mux.scala 31:69:@20162.4]
  assign _T_4537 = RetimeWrapper_126_io_out; // @[package.scala 96:25:@20117.4 package.scala 96:25:@20118.4]
  assign _T_4557 = _T_4537 ? Mem1D_12_io_output : _T_4556; // @[Mux.scala 31:69:@20163.4]
  assign _T_4534 = RetimeWrapper_125_io_out; // @[package.scala 96:25:@20109.4 package.scala 96:25:@20110.4]
  assign _T_4558 = _T_4534 ? Mem1D_10_io_output : _T_4557; // @[Mux.scala 31:69:@20164.4]
  assign _T_4531 = RetimeWrapper_124_io_out; // @[package.scala 96:25:@20101.4 package.scala 96:25:@20102.4]
  assign _T_4559 = _T_4531 ? Mem1D_8_io_output : _T_4558; // @[Mux.scala 31:69:@20165.4]
  assign _T_4528 = RetimeWrapper_123_io_out; // @[package.scala 96:25:@20093.4 package.scala 96:25:@20094.4]
  assign _T_4560 = _T_4528 ? Mem1D_6_io_output : _T_4559; // @[Mux.scala 31:69:@20166.4]
  assign _T_4525 = RetimeWrapper_122_io_out; // @[package.scala 96:25:@20085.4 package.scala 96:25:@20086.4]
  assign _T_4561 = _T_4525 ? Mem1D_4_io_output : _T_4560; // @[Mux.scala 31:69:@20167.4]
  assign _T_4522 = RetimeWrapper_121_io_out; // @[package.scala 96:25:@20077.4 package.scala 96:25:@20078.4]
  assign _T_4562 = _T_4522 ? Mem1D_2_io_output : _T_4561; // @[Mux.scala 31:69:@20168.4]
  assign _T_4519 = RetimeWrapper_120_io_out; // @[package.scala 96:25:@20069.4 package.scala 96:25:@20070.4]
  assign _T_4656 = RetimeWrapper_142_io_out; // @[package.scala 96:25:@20293.4 package.scala 96:25:@20294.4]
  assign _T_4660 = _T_4656 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@20303.4]
  assign _T_4653 = RetimeWrapper_141_io_out; // @[package.scala 96:25:@20285.4 package.scala 96:25:@20286.4]
  assign _T_4661 = _T_4653 ? Mem1D_19_io_output : _T_4660; // @[Mux.scala 31:69:@20304.4]
  assign _T_4650 = RetimeWrapper_140_io_out; // @[package.scala 96:25:@20277.4 package.scala 96:25:@20278.4]
  assign _T_4662 = _T_4650 ? Mem1D_17_io_output : _T_4661; // @[Mux.scala 31:69:@20305.4]
  assign _T_4647 = RetimeWrapper_139_io_out; // @[package.scala 96:25:@20269.4 package.scala 96:25:@20270.4]
  assign _T_4663 = _T_4647 ? Mem1D_15_io_output : _T_4662; // @[Mux.scala 31:69:@20306.4]
  assign _T_4644 = RetimeWrapper_138_io_out; // @[package.scala 96:25:@20261.4 package.scala 96:25:@20262.4]
  assign _T_4664 = _T_4644 ? Mem1D_13_io_output : _T_4663; // @[Mux.scala 31:69:@20307.4]
  assign _T_4641 = RetimeWrapper_137_io_out; // @[package.scala 96:25:@20253.4 package.scala 96:25:@20254.4]
  assign _T_4665 = _T_4641 ? Mem1D_11_io_output : _T_4664; // @[Mux.scala 31:69:@20308.4]
  assign _T_4638 = RetimeWrapper_136_io_out; // @[package.scala 96:25:@20245.4 package.scala 96:25:@20246.4]
  assign _T_4666 = _T_4638 ? Mem1D_9_io_output : _T_4665; // @[Mux.scala 31:69:@20309.4]
  assign _T_4635 = RetimeWrapper_135_io_out; // @[package.scala 96:25:@20237.4 package.scala 96:25:@20238.4]
  assign _T_4667 = _T_4635 ? Mem1D_7_io_output : _T_4666; // @[Mux.scala 31:69:@20310.4]
  assign _T_4632 = RetimeWrapper_134_io_out; // @[package.scala 96:25:@20229.4 package.scala 96:25:@20230.4]
  assign _T_4668 = _T_4632 ? Mem1D_5_io_output : _T_4667; // @[Mux.scala 31:69:@20311.4]
  assign _T_4629 = RetimeWrapper_133_io_out; // @[package.scala 96:25:@20221.4 package.scala 96:25:@20222.4]
  assign _T_4669 = _T_4629 ? Mem1D_3_io_output : _T_4668; // @[Mux.scala 31:69:@20312.4]
  assign _T_4626 = RetimeWrapper_132_io_out; // @[package.scala 96:25:@20213.4 package.scala 96:25:@20214.4]
  assign _T_4763 = RetimeWrapper_154_io_out; // @[package.scala 96:25:@20437.4 package.scala 96:25:@20438.4]
  assign _T_4767 = _T_4763 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@20447.4]
  assign _T_4760 = RetimeWrapper_153_io_out; // @[package.scala 96:25:@20429.4 package.scala 96:25:@20430.4]
  assign _T_4768 = _T_4760 ? Mem1D_19_io_output : _T_4767; // @[Mux.scala 31:69:@20448.4]
  assign _T_4757 = RetimeWrapper_152_io_out; // @[package.scala 96:25:@20421.4 package.scala 96:25:@20422.4]
  assign _T_4769 = _T_4757 ? Mem1D_17_io_output : _T_4768; // @[Mux.scala 31:69:@20449.4]
  assign _T_4754 = RetimeWrapper_151_io_out; // @[package.scala 96:25:@20413.4 package.scala 96:25:@20414.4]
  assign _T_4770 = _T_4754 ? Mem1D_15_io_output : _T_4769; // @[Mux.scala 31:69:@20450.4]
  assign _T_4751 = RetimeWrapper_150_io_out; // @[package.scala 96:25:@20405.4 package.scala 96:25:@20406.4]
  assign _T_4771 = _T_4751 ? Mem1D_13_io_output : _T_4770; // @[Mux.scala 31:69:@20451.4]
  assign _T_4748 = RetimeWrapper_149_io_out; // @[package.scala 96:25:@20397.4 package.scala 96:25:@20398.4]
  assign _T_4772 = _T_4748 ? Mem1D_11_io_output : _T_4771; // @[Mux.scala 31:69:@20452.4]
  assign _T_4745 = RetimeWrapper_148_io_out; // @[package.scala 96:25:@20389.4 package.scala 96:25:@20390.4]
  assign _T_4773 = _T_4745 ? Mem1D_9_io_output : _T_4772; // @[Mux.scala 31:69:@20453.4]
  assign _T_4742 = RetimeWrapper_147_io_out; // @[package.scala 96:25:@20381.4 package.scala 96:25:@20382.4]
  assign _T_4774 = _T_4742 ? Mem1D_7_io_output : _T_4773; // @[Mux.scala 31:69:@20454.4]
  assign _T_4739 = RetimeWrapper_146_io_out; // @[package.scala 96:25:@20373.4 package.scala 96:25:@20374.4]
  assign _T_4775 = _T_4739 ? Mem1D_5_io_output : _T_4774; // @[Mux.scala 31:69:@20455.4]
  assign _T_4736 = RetimeWrapper_145_io_out; // @[package.scala 96:25:@20365.4 package.scala 96:25:@20366.4]
  assign _T_4776 = _T_4736 ? Mem1D_3_io_output : _T_4775; // @[Mux.scala 31:69:@20456.4]
  assign _T_4733 = RetimeWrapper_144_io_out; // @[package.scala 96:25:@20357.4 package.scala 96:25:@20358.4]
  assign _T_4870 = RetimeWrapper_166_io_out; // @[package.scala 96:25:@20581.4 package.scala 96:25:@20582.4]
  assign _T_4874 = _T_4870 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@20591.4]
  assign _T_4867 = RetimeWrapper_165_io_out; // @[package.scala 96:25:@20573.4 package.scala 96:25:@20574.4]
  assign _T_4875 = _T_4867 ? Mem1D_19_io_output : _T_4874; // @[Mux.scala 31:69:@20592.4]
  assign _T_4864 = RetimeWrapper_164_io_out; // @[package.scala 96:25:@20565.4 package.scala 96:25:@20566.4]
  assign _T_4876 = _T_4864 ? Mem1D_17_io_output : _T_4875; // @[Mux.scala 31:69:@20593.4]
  assign _T_4861 = RetimeWrapper_163_io_out; // @[package.scala 96:25:@20557.4 package.scala 96:25:@20558.4]
  assign _T_4877 = _T_4861 ? Mem1D_15_io_output : _T_4876; // @[Mux.scala 31:69:@20594.4]
  assign _T_4858 = RetimeWrapper_162_io_out; // @[package.scala 96:25:@20549.4 package.scala 96:25:@20550.4]
  assign _T_4878 = _T_4858 ? Mem1D_13_io_output : _T_4877; // @[Mux.scala 31:69:@20595.4]
  assign _T_4855 = RetimeWrapper_161_io_out; // @[package.scala 96:25:@20541.4 package.scala 96:25:@20542.4]
  assign _T_4879 = _T_4855 ? Mem1D_11_io_output : _T_4878; // @[Mux.scala 31:69:@20596.4]
  assign _T_4852 = RetimeWrapper_160_io_out; // @[package.scala 96:25:@20533.4 package.scala 96:25:@20534.4]
  assign _T_4880 = _T_4852 ? Mem1D_9_io_output : _T_4879; // @[Mux.scala 31:69:@20597.4]
  assign _T_4849 = RetimeWrapper_159_io_out; // @[package.scala 96:25:@20525.4 package.scala 96:25:@20526.4]
  assign _T_4881 = _T_4849 ? Mem1D_7_io_output : _T_4880; // @[Mux.scala 31:69:@20598.4]
  assign _T_4846 = RetimeWrapper_158_io_out; // @[package.scala 96:25:@20517.4 package.scala 96:25:@20518.4]
  assign _T_4882 = _T_4846 ? Mem1D_5_io_output : _T_4881; // @[Mux.scala 31:69:@20599.4]
  assign _T_4843 = RetimeWrapper_157_io_out; // @[package.scala 96:25:@20509.4 package.scala 96:25:@20510.4]
  assign _T_4883 = _T_4843 ? Mem1D_3_io_output : _T_4882; // @[Mux.scala 31:69:@20600.4]
  assign _T_4840 = RetimeWrapper_156_io_out; // @[package.scala 96:25:@20501.4 package.scala 96:25:@20502.4]
  assign _T_4977 = RetimeWrapper_178_io_out; // @[package.scala 96:25:@20725.4 package.scala 96:25:@20726.4]
  assign _T_4981 = _T_4977 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@20735.4]
  assign _T_4974 = RetimeWrapper_177_io_out; // @[package.scala 96:25:@20717.4 package.scala 96:25:@20718.4]
  assign _T_4982 = _T_4974 ? Mem1D_18_io_output : _T_4981; // @[Mux.scala 31:69:@20736.4]
  assign _T_4971 = RetimeWrapper_176_io_out; // @[package.scala 96:25:@20709.4 package.scala 96:25:@20710.4]
  assign _T_4983 = _T_4971 ? Mem1D_16_io_output : _T_4982; // @[Mux.scala 31:69:@20737.4]
  assign _T_4968 = RetimeWrapper_175_io_out; // @[package.scala 96:25:@20701.4 package.scala 96:25:@20702.4]
  assign _T_4984 = _T_4968 ? Mem1D_14_io_output : _T_4983; // @[Mux.scala 31:69:@20738.4]
  assign _T_4965 = RetimeWrapper_174_io_out; // @[package.scala 96:25:@20693.4 package.scala 96:25:@20694.4]
  assign _T_4985 = _T_4965 ? Mem1D_12_io_output : _T_4984; // @[Mux.scala 31:69:@20739.4]
  assign _T_4962 = RetimeWrapper_173_io_out; // @[package.scala 96:25:@20685.4 package.scala 96:25:@20686.4]
  assign _T_4986 = _T_4962 ? Mem1D_10_io_output : _T_4985; // @[Mux.scala 31:69:@20740.4]
  assign _T_4959 = RetimeWrapper_172_io_out; // @[package.scala 96:25:@20677.4 package.scala 96:25:@20678.4]
  assign _T_4987 = _T_4959 ? Mem1D_8_io_output : _T_4986; // @[Mux.scala 31:69:@20741.4]
  assign _T_4956 = RetimeWrapper_171_io_out; // @[package.scala 96:25:@20669.4 package.scala 96:25:@20670.4]
  assign _T_4988 = _T_4956 ? Mem1D_6_io_output : _T_4987; // @[Mux.scala 31:69:@20742.4]
  assign _T_4953 = RetimeWrapper_170_io_out; // @[package.scala 96:25:@20661.4 package.scala 96:25:@20662.4]
  assign _T_4989 = _T_4953 ? Mem1D_4_io_output : _T_4988; // @[Mux.scala 31:69:@20743.4]
  assign _T_4950 = RetimeWrapper_169_io_out; // @[package.scala 96:25:@20653.4 package.scala 96:25:@20654.4]
  assign _T_4990 = _T_4950 ? Mem1D_2_io_output : _T_4989; // @[Mux.scala 31:69:@20744.4]
  assign _T_4947 = RetimeWrapper_168_io_out; // @[package.scala 96:25:@20645.4 package.scala 96:25:@20646.4]
  assign _T_5084 = RetimeWrapper_190_io_out; // @[package.scala 96:25:@20869.4 package.scala 96:25:@20870.4]
  assign _T_5088 = _T_5084 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@20879.4]
  assign _T_5081 = RetimeWrapper_189_io_out; // @[package.scala 96:25:@20861.4 package.scala 96:25:@20862.4]
  assign _T_5089 = _T_5081 ? Mem1D_18_io_output : _T_5088; // @[Mux.scala 31:69:@20880.4]
  assign _T_5078 = RetimeWrapper_188_io_out; // @[package.scala 96:25:@20853.4 package.scala 96:25:@20854.4]
  assign _T_5090 = _T_5078 ? Mem1D_16_io_output : _T_5089; // @[Mux.scala 31:69:@20881.4]
  assign _T_5075 = RetimeWrapper_187_io_out; // @[package.scala 96:25:@20845.4 package.scala 96:25:@20846.4]
  assign _T_5091 = _T_5075 ? Mem1D_14_io_output : _T_5090; // @[Mux.scala 31:69:@20882.4]
  assign _T_5072 = RetimeWrapper_186_io_out; // @[package.scala 96:25:@20837.4 package.scala 96:25:@20838.4]
  assign _T_5092 = _T_5072 ? Mem1D_12_io_output : _T_5091; // @[Mux.scala 31:69:@20883.4]
  assign _T_5069 = RetimeWrapper_185_io_out; // @[package.scala 96:25:@20829.4 package.scala 96:25:@20830.4]
  assign _T_5093 = _T_5069 ? Mem1D_10_io_output : _T_5092; // @[Mux.scala 31:69:@20884.4]
  assign _T_5066 = RetimeWrapper_184_io_out; // @[package.scala 96:25:@20821.4 package.scala 96:25:@20822.4]
  assign _T_5094 = _T_5066 ? Mem1D_8_io_output : _T_5093; // @[Mux.scala 31:69:@20885.4]
  assign _T_5063 = RetimeWrapper_183_io_out; // @[package.scala 96:25:@20813.4 package.scala 96:25:@20814.4]
  assign _T_5095 = _T_5063 ? Mem1D_6_io_output : _T_5094; // @[Mux.scala 31:69:@20886.4]
  assign _T_5060 = RetimeWrapper_182_io_out; // @[package.scala 96:25:@20805.4 package.scala 96:25:@20806.4]
  assign _T_5096 = _T_5060 ? Mem1D_4_io_output : _T_5095; // @[Mux.scala 31:69:@20887.4]
  assign _T_5057 = RetimeWrapper_181_io_out; // @[package.scala 96:25:@20797.4 package.scala 96:25:@20798.4]
  assign _T_5097 = _T_5057 ? Mem1D_2_io_output : _T_5096; // @[Mux.scala 31:69:@20888.4]
  assign _T_5054 = RetimeWrapper_180_io_out; // @[package.scala 96:25:@20789.4 package.scala 96:25:@20790.4]
  assign _T_5191 = RetimeWrapper_202_io_out; // @[package.scala 96:25:@21013.4 package.scala 96:25:@21014.4]
  assign _T_5195 = _T_5191 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@21023.4]
  assign _T_5188 = RetimeWrapper_201_io_out; // @[package.scala 96:25:@21005.4 package.scala 96:25:@21006.4]
  assign _T_5196 = _T_5188 ? Mem1D_19_io_output : _T_5195; // @[Mux.scala 31:69:@21024.4]
  assign _T_5185 = RetimeWrapper_200_io_out; // @[package.scala 96:25:@20997.4 package.scala 96:25:@20998.4]
  assign _T_5197 = _T_5185 ? Mem1D_17_io_output : _T_5196; // @[Mux.scala 31:69:@21025.4]
  assign _T_5182 = RetimeWrapper_199_io_out; // @[package.scala 96:25:@20989.4 package.scala 96:25:@20990.4]
  assign _T_5198 = _T_5182 ? Mem1D_15_io_output : _T_5197; // @[Mux.scala 31:69:@21026.4]
  assign _T_5179 = RetimeWrapper_198_io_out; // @[package.scala 96:25:@20981.4 package.scala 96:25:@20982.4]
  assign _T_5199 = _T_5179 ? Mem1D_13_io_output : _T_5198; // @[Mux.scala 31:69:@21027.4]
  assign _T_5176 = RetimeWrapper_197_io_out; // @[package.scala 96:25:@20973.4 package.scala 96:25:@20974.4]
  assign _T_5200 = _T_5176 ? Mem1D_11_io_output : _T_5199; // @[Mux.scala 31:69:@21028.4]
  assign _T_5173 = RetimeWrapper_196_io_out; // @[package.scala 96:25:@20965.4 package.scala 96:25:@20966.4]
  assign _T_5201 = _T_5173 ? Mem1D_9_io_output : _T_5200; // @[Mux.scala 31:69:@21029.4]
  assign _T_5170 = RetimeWrapper_195_io_out; // @[package.scala 96:25:@20957.4 package.scala 96:25:@20958.4]
  assign _T_5202 = _T_5170 ? Mem1D_7_io_output : _T_5201; // @[Mux.scala 31:69:@21030.4]
  assign _T_5167 = RetimeWrapper_194_io_out; // @[package.scala 96:25:@20949.4 package.scala 96:25:@20950.4]
  assign _T_5203 = _T_5167 ? Mem1D_5_io_output : _T_5202; // @[Mux.scala 31:69:@21031.4]
  assign _T_5164 = RetimeWrapper_193_io_out; // @[package.scala 96:25:@20941.4 package.scala 96:25:@20942.4]
  assign _T_5204 = _T_5164 ? Mem1D_3_io_output : _T_5203; // @[Mux.scala 31:69:@21032.4]
  assign _T_5161 = RetimeWrapper_192_io_out; // @[package.scala 96:25:@20933.4 package.scala 96:25:@20934.4]
  assign _T_5298 = RetimeWrapper_214_io_out; // @[package.scala 96:25:@21157.4 package.scala 96:25:@21158.4]
  assign _T_5302 = _T_5298 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@21167.4]
  assign _T_5295 = RetimeWrapper_213_io_out; // @[package.scala 96:25:@21149.4 package.scala 96:25:@21150.4]
  assign _T_5303 = _T_5295 ? Mem1D_18_io_output : _T_5302; // @[Mux.scala 31:69:@21168.4]
  assign _T_5292 = RetimeWrapper_212_io_out; // @[package.scala 96:25:@21141.4 package.scala 96:25:@21142.4]
  assign _T_5304 = _T_5292 ? Mem1D_16_io_output : _T_5303; // @[Mux.scala 31:69:@21169.4]
  assign _T_5289 = RetimeWrapper_211_io_out; // @[package.scala 96:25:@21133.4 package.scala 96:25:@21134.4]
  assign _T_5305 = _T_5289 ? Mem1D_14_io_output : _T_5304; // @[Mux.scala 31:69:@21170.4]
  assign _T_5286 = RetimeWrapper_210_io_out; // @[package.scala 96:25:@21125.4 package.scala 96:25:@21126.4]
  assign _T_5306 = _T_5286 ? Mem1D_12_io_output : _T_5305; // @[Mux.scala 31:69:@21171.4]
  assign _T_5283 = RetimeWrapper_209_io_out; // @[package.scala 96:25:@21117.4 package.scala 96:25:@21118.4]
  assign _T_5307 = _T_5283 ? Mem1D_10_io_output : _T_5306; // @[Mux.scala 31:69:@21172.4]
  assign _T_5280 = RetimeWrapper_208_io_out; // @[package.scala 96:25:@21109.4 package.scala 96:25:@21110.4]
  assign _T_5308 = _T_5280 ? Mem1D_8_io_output : _T_5307; // @[Mux.scala 31:69:@21173.4]
  assign _T_5277 = RetimeWrapper_207_io_out; // @[package.scala 96:25:@21101.4 package.scala 96:25:@21102.4]
  assign _T_5309 = _T_5277 ? Mem1D_6_io_output : _T_5308; // @[Mux.scala 31:69:@21174.4]
  assign _T_5274 = RetimeWrapper_206_io_out; // @[package.scala 96:25:@21093.4 package.scala 96:25:@21094.4]
  assign _T_5310 = _T_5274 ? Mem1D_4_io_output : _T_5309; // @[Mux.scala 31:69:@21175.4]
  assign _T_5271 = RetimeWrapper_205_io_out; // @[package.scala 96:25:@21085.4 package.scala 96:25:@21086.4]
  assign _T_5311 = _T_5271 ? Mem1D_2_io_output : _T_5310; // @[Mux.scala 31:69:@21176.4]
  assign _T_5268 = RetimeWrapper_204_io_out; // @[package.scala 96:25:@21077.4 package.scala 96:25:@21078.4]
  assign io_rPort_17_output_0 = _T_5268 ? Mem1D_io_output : _T_5311; // @[MemPrimitives.scala 148:13:@21178.4]
  assign io_rPort_16_output_0 = _T_5161 ? Mem1D_1_io_output : _T_5204; // @[MemPrimitives.scala 148:13:@21034.4]
  assign io_rPort_15_output_0 = _T_5054 ? Mem1D_io_output : _T_5097; // @[MemPrimitives.scala 148:13:@20890.4]
  assign io_rPort_14_output_0 = _T_4947 ? Mem1D_io_output : _T_4990; // @[MemPrimitives.scala 148:13:@20746.4]
  assign io_rPort_13_output_0 = _T_4840 ? Mem1D_1_io_output : _T_4883; // @[MemPrimitives.scala 148:13:@20602.4]
  assign io_rPort_12_output_0 = _T_4733 ? Mem1D_1_io_output : _T_4776; // @[MemPrimitives.scala 148:13:@20458.4]
  assign io_rPort_11_output_0 = _T_4626 ? Mem1D_1_io_output : _T_4669; // @[MemPrimitives.scala 148:13:@20314.4]
  assign io_rPort_10_output_0 = _T_4519 ? Mem1D_io_output : _T_4562; // @[MemPrimitives.scala 148:13:@20170.4]
  assign io_rPort_9_output_0 = _T_4412 ? Mem1D_1_io_output : _T_4455; // @[MemPrimitives.scala 148:13:@20026.4]
  assign io_rPort_8_output_0 = _T_4305 ? Mem1D_io_output : _T_4348; // @[MemPrimitives.scala 148:13:@19882.4]
  assign io_rPort_7_output_0 = _T_4198 ? Mem1D_1_io_output : _T_4241; // @[MemPrimitives.scala 148:13:@19738.4]
  assign io_rPort_6_output_0 = _T_4091 ? Mem1D_1_io_output : _T_4134; // @[MemPrimitives.scala 148:13:@19594.4]
  assign io_rPort_5_output_0 = _T_3984 ? Mem1D_1_io_output : _T_4027; // @[MemPrimitives.scala 148:13:@19450.4]
  assign io_rPort_4_output_0 = _T_3877 ? Mem1D_io_output : _T_3920; // @[MemPrimitives.scala 148:13:@19306.4]
  assign io_rPort_3_output_0 = _T_3770 ? Mem1D_io_output : _T_3813; // @[MemPrimitives.scala 148:13:@19162.4]
  assign io_rPort_2_output_0 = _T_3663 ? Mem1D_1_io_output : _T_3706; // @[MemPrimitives.scala 148:13:@19018.4]
  assign io_rPort_1_output_0 = _T_3556 ? Mem1D_io_output : _T_3599; // @[MemPrimitives.scala 148:13:@18874.4]
  assign io_rPort_0_output_0 = _T_3449 ? Mem1D_io_output : _T_3492; // @[MemPrimitives.scala 148:13:@18730.4]
  assign Mem1D_clock = clock; // @[:@15612.4]
  assign Mem1D_reset = reset; // @[:@15613.4]
  assign Mem1D_io_r_ofs_0 = _T_1267[7:0]; // @[MemPrimitives.scala 127:28:@16537.4]
  assign Mem1D_io_r_backpressure = _T_1267[8]; // @[MemPrimitives.scala 128:32:@16538.4]
  assign Mem1D_io_w_ofs_0 = _T_715[7:0]; // @[MemPrimitives.scala 94:28:@16011.4]
  assign Mem1D_io_w_data_0 = _T_715[15:8]; // @[MemPrimitives.scala 95:29:@16012.4]
  assign Mem1D_io_w_en_0 = _T_715[16]; // @[MemPrimitives.scala 96:27:@16013.4]
  assign Mem1D_1_clock = clock; // @[:@15628.4]
  assign Mem1D_1_reset = reset; // @[:@15629.4]
  assign Mem1D_1_io_r_ofs_0 = _T_1359[7:0]; // @[MemPrimitives.scala 127:28:@16626.4]
  assign Mem1D_1_io_r_backpressure = _T_1359[8]; // @[MemPrimitives.scala 128:32:@16627.4]
  assign Mem1D_1_io_w_ofs_0 = _T_735[7:0]; // @[MemPrimitives.scala 94:28:@16030.4]
  assign Mem1D_1_io_w_data_0 = _T_735[15:8]; // @[MemPrimitives.scala 95:29:@16031.4]
  assign Mem1D_1_io_w_en_0 = _T_735[16]; // @[MemPrimitives.scala 96:27:@16032.4]
  assign Mem1D_2_clock = clock; // @[:@15644.4]
  assign Mem1D_2_reset = reset; // @[:@15645.4]
  assign Mem1D_2_io_r_ofs_0 = _T_1451[7:0]; // @[MemPrimitives.scala 127:28:@16715.4]
  assign Mem1D_2_io_r_backpressure = _T_1451[8]; // @[MemPrimitives.scala 128:32:@16716.4]
  assign Mem1D_2_io_w_ofs_0 = _T_755[7:0]; // @[MemPrimitives.scala 94:28:@16049.4]
  assign Mem1D_2_io_w_data_0 = _T_755[15:8]; // @[MemPrimitives.scala 95:29:@16050.4]
  assign Mem1D_2_io_w_en_0 = _T_755[16]; // @[MemPrimitives.scala 96:27:@16051.4]
  assign Mem1D_3_clock = clock; // @[:@15660.4]
  assign Mem1D_3_reset = reset; // @[:@15661.4]
  assign Mem1D_3_io_r_ofs_0 = _T_1543[7:0]; // @[MemPrimitives.scala 127:28:@16804.4]
  assign Mem1D_3_io_r_backpressure = _T_1543[8]; // @[MemPrimitives.scala 128:32:@16805.4]
  assign Mem1D_3_io_w_ofs_0 = _T_775[7:0]; // @[MemPrimitives.scala 94:28:@16068.4]
  assign Mem1D_3_io_w_data_0 = _T_775[15:8]; // @[MemPrimitives.scala 95:29:@16069.4]
  assign Mem1D_3_io_w_en_0 = _T_775[16]; // @[MemPrimitives.scala 96:27:@16070.4]
  assign Mem1D_4_clock = clock; // @[:@15676.4]
  assign Mem1D_4_reset = reset; // @[:@15677.4]
  assign Mem1D_4_io_r_ofs_0 = _T_1635[7:0]; // @[MemPrimitives.scala 127:28:@16893.4]
  assign Mem1D_4_io_r_backpressure = _T_1635[8]; // @[MemPrimitives.scala 128:32:@16894.4]
  assign Mem1D_4_io_w_ofs_0 = _T_795[7:0]; // @[MemPrimitives.scala 94:28:@16087.4]
  assign Mem1D_4_io_w_data_0 = _T_795[15:8]; // @[MemPrimitives.scala 95:29:@16088.4]
  assign Mem1D_4_io_w_en_0 = _T_795[16]; // @[MemPrimitives.scala 96:27:@16089.4]
  assign Mem1D_5_clock = clock; // @[:@15692.4]
  assign Mem1D_5_reset = reset; // @[:@15693.4]
  assign Mem1D_5_io_r_ofs_0 = _T_1727[7:0]; // @[MemPrimitives.scala 127:28:@16982.4]
  assign Mem1D_5_io_r_backpressure = _T_1727[8]; // @[MemPrimitives.scala 128:32:@16983.4]
  assign Mem1D_5_io_w_ofs_0 = _T_815[7:0]; // @[MemPrimitives.scala 94:28:@16106.4]
  assign Mem1D_5_io_w_data_0 = _T_815[15:8]; // @[MemPrimitives.scala 95:29:@16107.4]
  assign Mem1D_5_io_w_en_0 = _T_815[16]; // @[MemPrimitives.scala 96:27:@16108.4]
  assign Mem1D_6_clock = clock; // @[:@15708.4]
  assign Mem1D_6_reset = reset; // @[:@15709.4]
  assign Mem1D_6_io_r_ofs_0 = _T_1819[7:0]; // @[MemPrimitives.scala 127:28:@17071.4]
  assign Mem1D_6_io_r_backpressure = _T_1819[8]; // @[MemPrimitives.scala 128:32:@17072.4]
  assign Mem1D_6_io_w_ofs_0 = _T_835[7:0]; // @[MemPrimitives.scala 94:28:@16125.4]
  assign Mem1D_6_io_w_data_0 = _T_835[15:8]; // @[MemPrimitives.scala 95:29:@16126.4]
  assign Mem1D_6_io_w_en_0 = _T_835[16]; // @[MemPrimitives.scala 96:27:@16127.4]
  assign Mem1D_7_clock = clock; // @[:@15724.4]
  assign Mem1D_7_reset = reset; // @[:@15725.4]
  assign Mem1D_7_io_r_ofs_0 = _T_1911[7:0]; // @[MemPrimitives.scala 127:28:@17160.4]
  assign Mem1D_7_io_r_backpressure = _T_1911[8]; // @[MemPrimitives.scala 128:32:@17161.4]
  assign Mem1D_7_io_w_ofs_0 = _T_855[7:0]; // @[MemPrimitives.scala 94:28:@16144.4]
  assign Mem1D_7_io_w_data_0 = _T_855[15:8]; // @[MemPrimitives.scala 95:29:@16145.4]
  assign Mem1D_7_io_w_en_0 = _T_855[16]; // @[MemPrimitives.scala 96:27:@16146.4]
  assign Mem1D_8_clock = clock; // @[:@15740.4]
  assign Mem1D_8_reset = reset; // @[:@15741.4]
  assign Mem1D_8_io_r_ofs_0 = _T_2003[7:0]; // @[MemPrimitives.scala 127:28:@17249.4]
  assign Mem1D_8_io_r_backpressure = _T_2003[8]; // @[MemPrimitives.scala 128:32:@17250.4]
  assign Mem1D_8_io_w_ofs_0 = _T_875[7:0]; // @[MemPrimitives.scala 94:28:@16163.4]
  assign Mem1D_8_io_w_data_0 = _T_875[15:8]; // @[MemPrimitives.scala 95:29:@16164.4]
  assign Mem1D_8_io_w_en_0 = _T_875[16]; // @[MemPrimitives.scala 96:27:@16165.4]
  assign Mem1D_9_clock = clock; // @[:@15756.4]
  assign Mem1D_9_reset = reset; // @[:@15757.4]
  assign Mem1D_9_io_r_ofs_0 = _T_2095[7:0]; // @[MemPrimitives.scala 127:28:@17338.4]
  assign Mem1D_9_io_r_backpressure = _T_2095[8]; // @[MemPrimitives.scala 128:32:@17339.4]
  assign Mem1D_9_io_w_ofs_0 = _T_895[7:0]; // @[MemPrimitives.scala 94:28:@16182.4]
  assign Mem1D_9_io_w_data_0 = _T_895[15:8]; // @[MemPrimitives.scala 95:29:@16183.4]
  assign Mem1D_9_io_w_en_0 = _T_895[16]; // @[MemPrimitives.scala 96:27:@16184.4]
  assign Mem1D_10_clock = clock; // @[:@15772.4]
  assign Mem1D_10_reset = reset; // @[:@15773.4]
  assign Mem1D_10_io_r_ofs_0 = _T_2187[7:0]; // @[MemPrimitives.scala 127:28:@17427.4]
  assign Mem1D_10_io_r_backpressure = _T_2187[8]; // @[MemPrimitives.scala 128:32:@17428.4]
  assign Mem1D_10_io_w_ofs_0 = _T_915[7:0]; // @[MemPrimitives.scala 94:28:@16201.4]
  assign Mem1D_10_io_w_data_0 = _T_915[15:8]; // @[MemPrimitives.scala 95:29:@16202.4]
  assign Mem1D_10_io_w_en_0 = _T_915[16]; // @[MemPrimitives.scala 96:27:@16203.4]
  assign Mem1D_11_clock = clock; // @[:@15788.4]
  assign Mem1D_11_reset = reset; // @[:@15789.4]
  assign Mem1D_11_io_r_ofs_0 = _T_2279[7:0]; // @[MemPrimitives.scala 127:28:@17516.4]
  assign Mem1D_11_io_r_backpressure = _T_2279[8]; // @[MemPrimitives.scala 128:32:@17517.4]
  assign Mem1D_11_io_w_ofs_0 = _T_935[7:0]; // @[MemPrimitives.scala 94:28:@16220.4]
  assign Mem1D_11_io_w_data_0 = _T_935[15:8]; // @[MemPrimitives.scala 95:29:@16221.4]
  assign Mem1D_11_io_w_en_0 = _T_935[16]; // @[MemPrimitives.scala 96:27:@16222.4]
  assign Mem1D_12_clock = clock; // @[:@15804.4]
  assign Mem1D_12_reset = reset; // @[:@15805.4]
  assign Mem1D_12_io_r_ofs_0 = _T_2371[7:0]; // @[MemPrimitives.scala 127:28:@17605.4]
  assign Mem1D_12_io_r_backpressure = _T_2371[8]; // @[MemPrimitives.scala 128:32:@17606.4]
  assign Mem1D_12_io_w_ofs_0 = _T_955[7:0]; // @[MemPrimitives.scala 94:28:@16239.4]
  assign Mem1D_12_io_w_data_0 = _T_955[15:8]; // @[MemPrimitives.scala 95:29:@16240.4]
  assign Mem1D_12_io_w_en_0 = _T_955[16]; // @[MemPrimitives.scala 96:27:@16241.4]
  assign Mem1D_13_clock = clock; // @[:@15820.4]
  assign Mem1D_13_reset = reset; // @[:@15821.4]
  assign Mem1D_13_io_r_ofs_0 = _T_2463[7:0]; // @[MemPrimitives.scala 127:28:@17694.4]
  assign Mem1D_13_io_r_backpressure = _T_2463[8]; // @[MemPrimitives.scala 128:32:@17695.4]
  assign Mem1D_13_io_w_ofs_0 = _T_975[7:0]; // @[MemPrimitives.scala 94:28:@16258.4]
  assign Mem1D_13_io_w_data_0 = _T_975[15:8]; // @[MemPrimitives.scala 95:29:@16259.4]
  assign Mem1D_13_io_w_en_0 = _T_975[16]; // @[MemPrimitives.scala 96:27:@16260.4]
  assign Mem1D_14_clock = clock; // @[:@15836.4]
  assign Mem1D_14_reset = reset; // @[:@15837.4]
  assign Mem1D_14_io_r_ofs_0 = _T_2555[7:0]; // @[MemPrimitives.scala 127:28:@17783.4]
  assign Mem1D_14_io_r_backpressure = _T_2555[8]; // @[MemPrimitives.scala 128:32:@17784.4]
  assign Mem1D_14_io_w_ofs_0 = _T_995[7:0]; // @[MemPrimitives.scala 94:28:@16277.4]
  assign Mem1D_14_io_w_data_0 = _T_995[15:8]; // @[MemPrimitives.scala 95:29:@16278.4]
  assign Mem1D_14_io_w_en_0 = _T_995[16]; // @[MemPrimitives.scala 96:27:@16279.4]
  assign Mem1D_15_clock = clock; // @[:@15852.4]
  assign Mem1D_15_reset = reset; // @[:@15853.4]
  assign Mem1D_15_io_r_ofs_0 = _T_2647[7:0]; // @[MemPrimitives.scala 127:28:@17872.4]
  assign Mem1D_15_io_r_backpressure = _T_2647[8]; // @[MemPrimitives.scala 128:32:@17873.4]
  assign Mem1D_15_io_w_ofs_0 = _T_1015[7:0]; // @[MemPrimitives.scala 94:28:@16296.4]
  assign Mem1D_15_io_w_data_0 = _T_1015[15:8]; // @[MemPrimitives.scala 95:29:@16297.4]
  assign Mem1D_15_io_w_en_0 = _T_1015[16]; // @[MemPrimitives.scala 96:27:@16298.4]
  assign Mem1D_16_clock = clock; // @[:@15868.4]
  assign Mem1D_16_reset = reset; // @[:@15869.4]
  assign Mem1D_16_io_r_ofs_0 = _T_2739[7:0]; // @[MemPrimitives.scala 127:28:@17961.4]
  assign Mem1D_16_io_r_backpressure = _T_2739[8]; // @[MemPrimitives.scala 128:32:@17962.4]
  assign Mem1D_16_io_w_ofs_0 = _T_1035[7:0]; // @[MemPrimitives.scala 94:28:@16315.4]
  assign Mem1D_16_io_w_data_0 = _T_1035[15:8]; // @[MemPrimitives.scala 95:29:@16316.4]
  assign Mem1D_16_io_w_en_0 = _T_1035[16]; // @[MemPrimitives.scala 96:27:@16317.4]
  assign Mem1D_17_clock = clock; // @[:@15884.4]
  assign Mem1D_17_reset = reset; // @[:@15885.4]
  assign Mem1D_17_io_r_ofs_0 = _T_2831[7:0]; // @[MemPrimitives.scala 127:28:@18050.4]
  assign Mem1D_17_io_r_backpressure = _T_2831[8]; // @[MemPrimitives.scala 128:32:@18051.4]
  assign Mem1D_17_io_w_ofs_0 = _T_1055[7:0]; // @[MemPrimitives.scala 94:28:@16334.4]
  assign Mem1D_17_io_w_data_0 = _T_1055[15:8]; // @[MemPrimitives.scala 95:29:@16335.4]
  assign Mem1D_17_io_w_en_0 = _T_1055[16]; // @[MemPrimitives.scala 96:27:@16336.4]
  assign Mem1D_18_clock = clock; // @[:@15900.4]
  assign Mem1D_18_reset = reset; // @[:@15901.4]
  assign Mem1D_18_io_r_ofs_0 = _T_2923[7:0]; // @[MemPrimitives.scala 127:28:@18139.4]
  assign Mem1D_18_io_r_backpressure = _T_2923[8]; // @[MemPrimitives.scala 128:32:@18140.4]
  assign Mem1D_18_io_w_ofs_0 = _T_1075[7:0]; // @[MemPrimitives.scala 94:28:@16353.4]
  assign Mem1D_18_io_w_data_0 = _T_1075[15:8]; // @[MemPrimitives.scala 95:29:@16354.4]
  assign Mem1D_18_io_w_en_0 = _T_1075[16]; // @[MemPrimitives.scala 96:27:@16355.4]
  assign Mem1D_19_clock = clock; // @[:@15916.4]
  assign Mem1D_19_reset = reset; // @[:@15917.4]
  assign Mem1D_19_io_r_ofs_0 = _T_3015[7:0]; // @[MemPrimitives.scala 127:28:@18228.4]
  assign Mem1D_19_io_r_backpressure = _T_3015[8]; // @[MemPrimitives.scala 128:32:@18229.4]
  assign Mem1D_19_io_w_ofs_0 = _T_1095[7:0]; // @[MemPrimitives.scala 94:28:@16372.4]
  assign Mem1D_19_io_w_data_0 = _T_1095[15:8]; // @[MemPrimitives.scala 95:29:@16373.4]
  assign Mem1D_19_io_w_en_0 = _T_1095[16]; // @[MemPrimitives.scala 96:27:@16374.4]
  assign Mem1D_20_clock = clock; // @[:@15932.4]
  assign Mem1D_20_reset = reset; // @[:@15933.4]
  assign Mem1D_20_io_r_ofs_0 = _T_3107[7:0]; // @[MemPrimitives.scala 127:28:@18317.4]
  assign Mem1D_20_io_r_backpressure = _T_3107[8]; // @[MemPrimitives.scala 128:32:@18318.4]
  assign Mem1D_20_io_w_ofs_0 = _T_1115[7:0]; // @[MemPrimitives.scala 94:28:@16391.4]
  assign Mem1D_20_io_w_data_0 = _T_1115[15:8]; // @[MemPrimitives.scala 95:29:@16392.4]
  assign Mem1D_20_io_w_en_0 = _T_1115[16]; // @[MemPrimitives.scala 96:27:@16393.4]
  assign Mem1D_21_clock = clock; // @[:@15948.4]
  assign Mem1D_21_reset = reset; // @[:@15949.4]
  assign Mem1D_21_io_r_ofs_0 = _T_3199[7:0]; // @[MemPrimitives.scala 127:28:@18406.4]
  assign Mem1D_21_io_r_backpressure = _T_3199[8]; // @[MemPrimitives.scala 128:32:@18407.4]
  assign Mem1D_21_io_w_ofs_0 = _T_1135[7:0]; // @[MemPrimitives.scala 94:28:@16410.4]
  assign Mem1D_21_io_w_data_0 = _T_1135[15:8]; // @[MemPrimitives.scala 95:29:@16411.4]
  assign Mem1D_21_io_w_en_0 = _T_1135[16]; // @[MemPrimitives.scala 96:27:@16412.4]
  assign Mem1D_22_clock = clock; // @[:@15964.4]
  assign Mem1D_22_reset = reset; // @[:@15965.4]
  assign Mem1D_22_io_r_ofs_0 = _T_3291[7:0]; // @[MemPrimitives.scala 127:28:@18495.4]
  assign Mem1D_22_io_r_backpressure = _T_3291[8]; // @[MemPrimitives.scala 128:32:@18496.4]
  assign Mem1D_22_io_w_ofs_0 = _T_1155[7:0]; // @[MemPrimitives.scala 94:28:@16429.4]
  assign Mem1D_22_io_w_data_0 = _T_1155[15:8]; // @[MemPrimitives.scala 95:29:@16430.4]
  assign Mem1D_22_io_w_en_0 = _T_1155[16]; // @[MemPrimitives.scala 96:27:@16431.4]
  assign Mem1D_23_clock = clock; // @[:@15980.4]
  assign Mem1D_23_reset = reset; // @[:@15981.4]
  assign Mem1D_23_io_r_ofs_0 = _T_3383[7:0]; // @[MemPrimitives.scala 127:28:@18584.4]
  assign Mem1D_23_io_r_backpressure = _T_3383[8]; // @[MemPrimitives.scala 128:32:@18585.4]
  assign Mem1D_23_io_w_ofs_0 = _T_1175[7:0]; // @[MemPrimitives.scala 94:28:@16448.4]
  assign Mem1D_23_io_w_data_0 = _T_1175[15:8]; // @[MemPrimitives.scala 95:29:@16449.4]
  assign Mem1D_23_io_w_en_0 = _T_1175[16]; // @[MemPrimitives.scala 96:27:@16450.4]
  assign StickySelects_clock = clock; // @[:@16488.4]
  assign StickySelects_reset = reset; // @[:@16489.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0 & _T_1183; // @[MemPrimitives.scala 122:60:@16490.4]
  assign StickySelects_io_ins_1 = io_rPort_1_en_0 & _T_1189; // @[MemPrimitives.scala 122:60:@16491.4]
  assign StickySelects_io_ins_2 = io_rPort_3_en_0 & _T_1195; // @[MemPrimitives.scala 122:60:@16492.4]
  assign StickySelects_io_ins_3 = io_rPort_4_en_0 & _T_1201; // @[MemPrimitives.scala 122:60:@16493.4]
  assign StickySelects_io_ins_4 = io_rPort_8_en_0 & _T_1207; // @[MemPrimitives.scala 122:60:@16494.4]
  assign StickySelects_io_ins_5 = io_rPort_10_en_0 & _T_1213; // @[MemPrimitives.scala 122:60:@16495.4]
  assign StickySelects_io_ins_6 = io_rPort_14_en_0 & _T_1219; // @[MemPrimitives.scala 122:60:@16496.4]
  assign StickySelects_io_ins_7 = io_rPort_15_en_0 & _T_1225; // @[MemPrimitives.scala 122:60:@16497.4]
  assign StickySelects_io_ins_8 = io_rPort_17_en_0 & _T_1231; // @[MemPrimitives.scala 122:60:@16498.4]
  assign StickySelects_1_clock = clock; // @[:@16577.4]
  assign StickySelects_1_reset = reset; // @[:@16578.4]
  assign StickySelects_1_io_ins_0 = io_rPort_2_en_0 & _T_1275; // @[MemPrimitives.scala 122:60:@16579.4]
  assign StickySelects_1_io_ins_1 = io_rPort_5_en_0 & _T_1281; // @[MemPrimitives.scala 122:60:@16580.4]
  assign StickySelects_1_io_ins_2 = io_rPort_6_en_0 & _T_1287; // @[MemPrimitives.scala 122:60:@16581.4]
  assign StickySelects_1_io_ins_3 = io_rPort_7_en_0 & _T_1293; // @[MemPrimitives.scala 122:60:@16582.4]
  assign StickySelects_1_io_ins_4 = io_rPort_9_en_0 & _T_1299; // @[MemPrimitives.scala 122:60:@16583.4]
  assign StickySelects_1_io_ins_5 = io_rPort_11_en_0 & _T_1305; // @[MemPrimitives.scala 122:60:@16584.4]
  assign StickySelects_1_io_ins_6 = io_rPort_12_en_0 & _T_1311; // @[MemPrimitives.scala 122:60:@16585.4]
  assign StickySelects_1_io_ins_7 = io_rPort_13_en_0 & _T_1317; // @[MemPrimitives.scala 122:60:@16586.4]
  assign StickySelects_1_io_ins_8 = io_rPort_16_en_0 & _T_1323; // @[MemPrimitives.scala 122:60:@16587.4]
  assign StickySelects_2_clock = clock; // @[:@16666.4]
  assign StickySelects_2_reset = reset; // @[:@16667.4]
  assign StickySelects_2_io_ins_0 = io_rPort_0_en_0 & _T_1367; // @[MemPrimitives.scala 122:60:@16668.4]
  assign StickySelects_2_io_ins_1 = io_rPort_1_en_0 & _T_1373; // @[MemPrimitives.scala 122:60:@16669.4]
  assign StickySelects_2_io_ins_2 = io_rPort_3_en_0 & _T_1379; // @[MemPrimitives.scala 122:60:@16670.4]
  assign StickySelects_2_io_ins_3 = io_rPort_4_en_0 & _T_1385; // @[MemPrimitives.scala 122:60:@16671.4]
  assign StickySelects_2_io_ins_4 = io_rPort_8_en_0 & _T_1391; // @[MemPrimitives.scala 122:60:@16672.4]
  assign StickySelects_2_io_ins_5 = io_rPort_10_en_0 & _T_1397; // @[MemPrimitives.scala 122:60:@16673.4]
  assign StickySelects_2_io_ins_6 = io_rPort_14_en_0 & _T_1403; // @[MemPrimitives.scala 122:60:@16674.4]
  assign StickySelects_2_io_ins_7 = io_rPort_15_en_0 & _T_1409; // @[MemPrimitives.scala 122:60:@16675.4]
  assign StickySelects_2_io_ins_8 = io_rPort_17_en_0 & _T_1415; // @[MemPrimitives.scala 122:60:@16676.4]
  assign StickySelects_3_clock = clock; // @[:@16755.4]
  assign StickySelects_3_reset = reset; // @[:@16756.4]
  assign StickySelects_3_io_ins_0 = io_rPort_2_en_0 & _T_1459; // @[MemPrimitives.scala 122:60:@16757.4]
  assign StickySelects_3_io_ins_1 = io_rPort_5_en_0 & _T_1465; // @[MemPrimitives.scala 122:60:@16758.4]
  assign StickySelects_3_io_ins_2 = io_rPort_6_en_0 & _T_1471; // @[MemPrimitives.scala 122:60:@16759.4]
  assign StickySelects_3_io_ins_3 = io_rPort_7_en_0 & _T_1477; // @[MemPrimitives.scala 122:60:@16760.4]
  assign StickySelects_3_io_ins_4 = io_rPort_9_en_0 & _T_1483; // @[MemPrimitives.scala 122:60:@16761.4]
  assign StickySelects_3_io_ins_5 = io_rPort_11_en_0 & _T_1489; // @[MemPrimitives.scala 122:60:@16762.4]
  assign StickySelects_3_io_ins_6 = io_rPort_12_en_0 & _T_1495; // @[MemPrimitives.scala 122:60:@16763.4]
  assign StickySelects_3_io_ins_7 = io_rPort_13_en_0 & _T_1501; // @[MemPrimitives.scala 122:60:@16764.4]
  assign StickySelects_3_io_ins_8 = io_rPort_16_en_0 & _T_1507; // @[MemPrimitives.scala 122:60:@16765.4]
  assign StickySelects_4_clock = clock; // @[:@16844.4]
  assign StickySelects_4_reset = reset; // @[:@16845.4]
  assign StickySelects_4_io_ins_0 = io_rPort_0_en_0 & _T_1551; // @[MemPrimitives.scala 122:60:@16846.4]
  assign StickySelects_4_io_ins_1 = io_rPort_1_en_0 & _T_1557; // @[MemPrimitives.scala 122:60:@16847.4]
  assign StickySelects_4_io_ins_2 = io_rPort_3_en_0 & _T_1563; // @[MemPrimitives.scala 122:60:@16848.4]
  assign StickySelects_4_io_ins_3 = io_rPort_4_en_0 & _T_1569; // @[MemPrimitives.scala 122:60:@16849.4]
  assign StickySelects_4_io_ins_4 = io_rPort_8_en_0 & _T_1575; // @[MemPrimitives.scala 122:60:@16850.4]
  assign StickySelects_4_io_ins_5 = io_rPort_10_en_0 & _T_1581; // @[MemPrimitives.scala 122:60:@16851.4]
  assign StickySelects_4_io_ins_6 = io_rPort_14_en_0 & _T_1587; // @[MemPrimitives.scala 122:60:@16852.4]
  assign StickySelects_4_io_ins_7 = io_rPort_15_en_0 & _T_1593; // @[MemPrimitives.scala 122:60:@16853.4]
  assign StickySelects_4_io_ins_8 = io_rPort_17_en_0 & _T_1599; // @[MemPrimitives.scala 122:60:@16854.4]
  assign StickySelects_5_clock = clock; // @[:@16933.4]
  assign StickySelects_5_reset = reset; // @[:@16934.4]
  assign StickySelects_5_io_ins_0 = io_rPort_2_en_0 & _T_1643; // @[MemPrimitives.scala 122:60:@16935.4]
  assign StickySelects_5_io_ins_1 = io_rPort_5_en_0 & _T_1649; // @[MemPrimitives.scala 122:60:@16936.4]
  assign StickySelects_5_io_ins_2 = io_rPort_6_en_0 & _T_1655; // @[MemPrimitives.scala 122:60:@16937.4]
  assign StickySelects_5_io_ins_3 = io_rPort_7_en_0 & _T_1661; // @[MemPrimitives.scala 122:60:@16938.4]
  assign StickySelects_5_io_ins_4 = io_rPort_9_en_0 & _T_1667; // @[MemPrimitives.scala 122:60:@16939.4]
  assign StickySelects_5_io_ins_5 = io_rPort_11_en_0 & _T_1673; // @[MemPrimitives.scala 122:60:@16940.4]
  assign StickySelects_5_io_ins_6 = io_rPort_12_en_0 & _T_1679; // @[MemPrimitives.scala 122:60:@16941.4]
  assign StickySelects_5_io_ins_7 = io_rPort_13_en_0 & _T_1685; // @[MemPrimitives.scala 122:60:@16942.4]
  assign StickySelects_5_io_ins_8 = io_rPort_16_en_0 & _T_1691; // @[MemPrimitives.scala 122:60:@16943.4]
  assign StickySelects_6_clock = clock; // @[:@17022.4]
  assign StickySelects_6_reset = reset; // @[:@17023.4]
  assign StickySelects_6_io_ins_0 = io_rPort_0_en_0 & _T_1735; // @[MemPrimitives.scala 122:60:@17024.4]
  assign StickySelects_6_io_ins_1 = io_rPort_1_en_0 & _T_1741; // @[MemPrimitives.scala 122:60:@17025.4]
  assign StickySelects_6_io_ins_2 = io_rPort_3_en_0 & _T_1747; // @[MemPrimitives.scala 122:60:@17026.4]
  assign StickySelects_6_io_ins_3 = io_rPort_4_en_0 & _T_1753; // @[MemPrimitives.scala 122:60:@17027.4]
  assign StickySelects_6_io_ins_4 = io_rPort_8_en_0 & _T_1759; // @[MemPrimitives.scala 122:60:@17028.4]
  assign StickySelects_6_io_ins_5 = io_rPort_10_en_0 & _T_1765; // @[MemPrimitives.scala 122:60:@17029.4]
  assign StickySelects_6_io_ins_6 = io_rPort_14_en_0 & _T_1771; // @[MemPrimitives.scala 122:60:@17030.4]
  assign StickySelects_6_io_ins_7 = io_rPort_15_en_0 & _T_1777; // @[MemPrimitives.scala 122:60:@17031.4]
  assign StickySelects_6_io_ins_8 = io_rPort_17_en_0 & _T_1783; // @[MemPrimitives.scala 122:60:@17032.4]
  assign StickySelects_7_clock = clock; // @[:@17111.4]
  assign StickySelects_7_reset = reset; // @[:@17112.4]
  assign StickySelects_7_io_ins_0 = io_rPort_2_en_0 & _T_1827; // @[MemPrimitives.scala 122:60:@17113.4]
  assign StickySelects_7_io_ins_1 = io_rPort_5_en_0 & _T_1833; // @[MemPrimitives.scala 122:60:@17114.4]
  assign StickySelects_7_io_ins_2 = io_rPort_6_en_0 & _T_1839; // @[MemPrimitives.scala 122:60:@17115.4]
  assign StickySelects_7_io_ins_3 = io_rPort_7_en_0 & _T_1845; // @[MemPrimitives.scala 122:60:@17116.4]
  assign StickySelects_7_io_ins_4 = io_rPort_9_en_0 & _T_1851; // @[MemPrimitives.scala 122:60:@17117.4]
  assign StickySelects_7_io_ins_5 = io_rPort_11_en_0 & _T_1857; // @[MemPrimitives.scala 122:60:@17118.4]
  assign StickySelects_7_io_ins_6 = io_rPort_12_en_0 & _T_1863; // @[MemPrimitives.scala 122:60:@17119.4]
  assign StickySelects_7_io_ins_7 = io_rPort_13_en_0 & _T_1869; // @[MemPrimitives.scala 122:60:@17120.4]
  assign StickySelects_7_io_ins_8 = io_rPort_16_en_0 & _T_1875; // @[MemPrimitives.scala 122:60:@17121.4]
  assign StickySelects_8_clock = clock; // @[:@17200.4]
  assign StickySelects_8_reset = reset; // @[:@17201.4]
  assign StickySelects_8_io_ins_0 = io_rPort_0_en_0 & _T_1919; // @[MemPrimitives.scala 122:60:@17202.4]
  assign StickySelects_8_io_ins_1 = io_rPort_1_en_0 & _T_1925; // @[MemPrimitives.scala 122:60:@17203.4]
  assign StickySelects_8_io_ins_2 = io_rPort_3_en_0 & _T_1931; // @[MemPrimitives.scala 122:60:@17204.4]
  assign StickySelects_8_io_ins_3 = io_rPort_4_en_0 & _T_1937; // @[MemPrimitives.scala 122:60:@17205.4]
  assign StickySelects_8_io_ins_4 = io_rPort_8_en_0 & _T_1943; // @[MemPrimitives.scala 122:60:@17206.4]
  assign StickySelects_8_io_ins_5 = io_rPort_10_en_0 & _T_1949; // @[MemPrimitives.scala 122:60:@17207.4]
  assign StickySelects_8_io_ins_6 = io_rPort_14_en_0 & _T_1955; // @[MemPrimitives.scala 122:60:@17208.4]
  assign StickySelects_8_io_ins_7 = io_rPort_15_en_0 & _T_1961; // @[MemPrimitives.scala 122:60:@17209.4]
  assign StickySelects_8_io_ins_8 = io_rPort_17_en_0 & _T_1967; // @[MemPrimitives.scala 122:60:@17210.4]
  assign StickySelects_9_clock = clock; // @[:@17289.4]
  assign StickySelects_9_reset = reset; // @[:@17290.4]
  assign StickySelects_9_io_ins_0 = io_rPort_2_en_0 & _T_2011; // @[MemPrimitives.scala 122:60:@17291.4]
  assign StickySelects_9_io_ins_1 = io_rPort_5_en_0 & _T_2017; // @[MemPrimitives.scala 122:60:@17292.4]
  assign StickySelects_9_io_ins_2 = io_rPort_6_en_0 & _T_2023; // @[MemPrimitives.scala 122:60:@17293.4]
  assign StickySelects_9_io_ins_3 = io_rPort_7_en_0 & _T_2029; // @[MemPrimitives.scala 122:60:@17294.4]
  assign StickySelects_9_io_ins_4 = io_rPort_9_en_0 & _T_2035; // @[MemPrimitives.scala 122:60:@17295.4]
  assign StickySelects_9_io_ins_5 = io_rPort_11_en_0 & _T_2041; // @[MemPrimitives.scala 122:60:@17296.4]
  assign StickySelects_9_io_ins_6 = io_rPort_12_en_0 & _T_2047; // @[MemPrimitives.scala 122:60:@17297.4]
  assign StickySelects_9_io_ins_7 = io_rPort_13_en_0 & _T_2053; // @[MemPrimitives.scala 122:60:@17298.4]
  assign StickySelects_9_io_ins_8 = io_rPort_16_en_0 & _T_2059; // @[MemPrimitives.scala 122:60:@17299.4]
  assign StickySelects_10_clock = clock; // @[:@17378.4]
  assign StickySelects_10_reset = reset; // @[:@17379.4]
  assign StickySelects_10_io_ins_0 = io_rPort_0_en_0 & _T_2103; // @[MemPrimitives.scala 122:60:@17380.4]
  assign StickySelects_10_io_ins_1 = io_rPort_1_en_0 & _T_2109; // @[MemPrimitives.scala 122:60:@17381.4]
  assign StickySelects_10_io_ins_2 = io_rPort_3_en_0 & _T_2115; // @[MemPrimitives.scala 122:60:@17382.4]
  assign StickySelects_10_io_ins_3 = io_rPort_4_en_0 & _T_2121; // @[MemPrimitives.scala 122:60:@17383.4]
  assign StickySelects_10_io_ins_4 = io_rPort_8_en_0 & _T_2127; // @[MemPrimitives.scala 122:60:@17384.4]
  assign StickySelects_10_io_ins_5 = io_rPort_10_en_0 & _T_2133; // @[MemPrimitives.scala 122:60:@17385.4]
  assign StickySelects_10_io_ins_6 = io_rPort_14_en_0 & _T_2139; // @[MemPrimitives.scala 122:60:@17386.4]
  assign StickySelects_10_io_ins_7 = io_rPort_15_en_0 & _T_2145; // @[MemPrimitives.scala 122:60:@17387.4]
  assign StickySelects_10_io_ins_8 = io_rPort_17_en_0 & _T_2151; // @[MemPrimitives.scala 122:60:@17388.4]
  assign StickySelects_11_clock = clock; // @[:@17467.4]
  assign StickySelects_11_reset = reset; // @[:@17468.4]
  assign StickySelects_11_io_ins_0 = io_rPort_2_en_0 & _T_2195; // @[MemPrimitives.scala 122:60:@17469.4]
  assign StickySelects_11_io_ins_1 = io_rPort_5_en_0 & _T_2201; // @[MemPrimitives.scala 122:60:@17470.4]
  assign StickySelects_11_io_ins_2 = io_rPort_6_en_0 & _T_2207; // @[MemPrimitives.scala 122:60:@17471.4]
  assign StickySelects_11_io_ins_3 = io_rPort_7_en_0 & _T_2213; // @[MemPrimitives.scala 122:60:@17472.4]
  assign StickySelects_11_io_ins_4 = io_rPort_9_en_0 & _T_2219; // @[MemPrimitives.scala 122:60:@17473.4]
  assign StickySelects_11_io_ins_5 = io_rPort_11_en_0 & _T_2225; // @[MemPrimitives.scala 122:60:@17474.4]
  assign StickySelects_11_io_ins_6 = io_rPort_12_en_0 & _T_2231; // @[MemPrimitives.scala 122:60:@17475.4]
  assign StickySelects_11_io_ins_7 = io_rPort_13_en_0 & _T_2237; // @[MemPrimitives.scala 122:60:@17476.4]
  assign StickySelects_11_io_ins_8 = io_rPort_16_en_0 & _T_2243; // @[MemPrimitives.scala 122:60:@17477.4]
  assign StickySelects_12_clock = clock; // @[:@17556.4]
  assign StickySelects_12_reset = reset; // @[:@17557.4]
  assign StickySelects_12_io_ins_0 = io_rPort_0_en_0 & _T_2287; // @[MemPrimitives.scala 122:60:@17558.4]
  assign StickySelects_12_io_ins_1 = io_rPort_1_en_0 & _T_2293; // @[MemPrimitives.scala 122:60:@17559.4]
  assign StickySelects_12_io_ins_2 = io_rPort_3_en_0 & _T_2299; // @[MemPrimitives.scala 122:60:@17560.4]
  assign StickySelects_12_io_ins_3 = io_rPort_4_en_0 & _T_2305; // @[MemPrimitives.scala 122:60:@17561.4]
  assign StickySelects_12_io_ins_4 = io_rPort_8_en_0 & _T_2311; // @[MemPrimitives.scala 122:60:@17562.4]
  assign StickySelects_12_io_ins_5 = io_rPort_10_en_0 & _T_2317; // @[MemPrimitives.scala 122:60:@17563.4]
  assign StickySelects_12_io_ins_6 = io_rPort_14_en_0 & _T_2323; // @[MemPrimitives.scala 122:60:@17564.4]
  assign StickySelects_12_io_ins_7 = io_rPort_15_en_0 & _T_2329; // @[MemPrimitives.scala 122:60:@17565.4]
  assign StickySelects_12_io_ins_8 = io_rPort_17_en_0 & _T_2335; // @[MemPrimitives.scala 122:60:@17566.4]
  assign StickySelects_13_clock = clock; // @[:@17645.4]
  assign StickySelects_13_reset = reset; // @[:@17646.4]
  assign StickySelects_13_io_ins_0 = io_rPort_2_en_0 & _T_2379; // @[MemPrimitives.scala 122:60:@17647.4]
  assign StickySelects_13_io_ins_1 = io_rPort_5_en_0 & _T_2385; // @[MemPrimitives.scala 122:60:@17648.4]
  assign StickySelects_13_io_ins_2 = io_rPort_6_en_0 & _T_2391; // @[MemPrimitives.scala 122:60:@17649.4]
  assign StickySelects_13_io_ins_3 = io_rPort_7_en_0 & _T_2397; // @[MemPrimitives.scala 122:60:@17650.4]
  assign StickySelects_13_io_ins_4 = io_rPort_9_en_0 & _T_2403; // @[MemPrimitives.scala 122:60:@17651.4]
  assign StickySelects_13_io_ins_5 = io_rPort_11_en_0 & _T_2409; // @[MemPrimitives.scala 122:60:@17652.4]
  assign StickySelects_13_io_ins_6 = io_rPort_12_en_0 & _T_2415; // @[MemPrimitives.scala 122:60:@17653.4]
  assign StickySelects_13_io_ins_7 = io_rPort_13_en_0 & _T_2421; // @[MemPrimitives.scala 122:60:@17654.4]
  assign StickySelects_13_io_ins_8 = io_rPort_16_en_0 & _T_2427; // @[MemPrimitives.scala 122:60:@17655.4]
  assign StickySelects_14_clock = clock; // @[:@17734.4]
  assign StickySelects_14_reset = reset; // @[:@17735.4]
  assign StickySelects_14_io_ins_0 = io_rPort_0_en_0 & _T_2471; // @[MemPrimitives.scala 122:60:@17736.4]
  assign StickySelects_14_io_ins_1 = io_rPort_1_en_0 & _T_2477; // @[MemPrimitives.scala 122:60:@17737.4]
  assign StickySelects_14_io_ins_2 = io_rPort_3_en_0 & _T_2483; // @[MemPrimitives.scala 122:60:@17738.4]
  assign StickySelects_14_io_ins_3 = io_rPort_4_en_0 & _T_2489; // @[MemPrimitives.scala 122:60:@17739.4]
  assign StickySelects_14_io_ins_4 = io_rPort_8_en_0 & _T_2495; // @[MemPrimitives.scala 122:60:@17740.4]
  assign StickySelects_14_io_ins_5 = io_rPort_10_en_0 & _T_2501; // @[MemPrimitives.scala 122:60:@17741.4]
  assign StickySelects_14_io_ins_6 = io_rPort_14_en_0 & _T_2507; // @[MemPrimitives.scala 122:60:@17742.4]
  assign StickySelects_14_io_ins_7 = io_rPort_15_en_0 & _T_2513; // @[MemPrimitives.scala 122:60:@17743.4]
  assign StickySelects_14_io_ins_8 = io_rPort_17_en_0 & _T_2519; // @[MemPrimitives.scala 122:60:@17744.4]
  assign StickySelects_15_clock = clock; // @[:@17823.4]
  assign StickySelects_15_reset = reset; // @[:@17824.4]
  assign StickySelects_15_io_ins_0 = io_rPort_2_en_0 & _T_2563; // @[MemPrimitives.scala 122:60:@17825.4]
  assign StickySelects_15_io_ins_1 = io_rPort_5_en_0 & _T_2569; // @[MemPrimitives.scala 122:60:@17826.4]
  assign StickySelects_15_io_ins_2 = io_rPort_6_en_0 & _T_2575; // @[MemPrimitives.scala 122:60:@17827.4]
  assign StickySelects_15_io_ins_3 = io_rPort_7_en_0 & _T_2581; // @[MemPrimitives.scala 122:60:@17828.4]
  assign StickySelects_15_io_ins_4 = io_rPort_9_en_0 & _T_2587; // @[MemPrimitives.scala 122:60:@17829.4]
  assign StickySelects_15_io_ins_5 = io_rPort_11_en_0 & _T_2593; // @[MemPrimitives.scala 122:60:@17830.4]
  assign StickySelects_15_io_ins_6 = io_rPort_12_en_0 & _T_2599; // @[MemPrimitives.scala 122:60:@17831.4]
  assign StickySelects_15_io_ins_7 = io_rPort_13_en_0 & _T_2605; // @[MemPrimitives.scala 122:60:@17832.4]
  assign StickySelects_15_io_ins_8 = io_rPort_16_en_0 & _T_2611; // @[MemPrimitives.scala 122:60:@17833.4]
  assign StickySelects_16_clock = clock; // @[:@17912.4]
  assign StickySelects_16_reset = reset; // @[:@17913.4]
  assign StickySelects_16_io_ins_0 = io_rPort_0_en_0 & _T_2655; // @[MemPrimitives.scala 122:60:@17914.4]
  assign StickySelects_16_io_ins_1 = io_rPort_1_en_0 & _T_2661; // @[MemPrimitives.scala 122:60:@17915.4]
  assign StickySelects_16_io_ins_2 = io_rPort_3_en_0 & _T_2667; // @[MemPrimitives.scala 122:60:@17916.4]
  assign StickySelects_16_io_ins_3 = io_rPort_4_en_0 & _T_2673; // @[MemPrimitives.scala 122:60:@17917.4]
  assign StickySelects_16_io_ins_4 = io_rPort_8_en_0 & _T_2679; // @[MemPrimitives.scala 122:60:@17918.4]
  assign StickySelects_16_io_ins_5 = io_rPort_10_en_0 & _T_2685; // @[MemPrimitives.scala 122:60:@17919.4]
  assign StickySelects_16_io_ins_6 = io_rPort_14_en_0 & _T_2691; // @[MemPrimitives.scala 122:60:@17920.4]
  assign StickySelects_16_io_ins_7 = io_rPort_15_en_0 & _T_2697; // @[MemPrimitives.scala 122:60:@17921.4]
  assign StickySelects_16_io_ins_8 = io_rPort_17_en_0 & _T_2703; // @[MemPrimitives.scala 122:60:@17922.4]
  assign StickySelects_17_clock = clock; // @[:@18001.4]
  assign StickySelects_17_reset = reset; // @[:@18002.4]
  assign StickySelects_17_io_ins_0 = io_rPort_2_en_0 & _T_2747; // @[MemPrimitives.scala 122:60:@18003.4]
  assign StickySelects_17_io_ins_1 = io_rPort_5_en_0 & _T_2753; // @[MemPrimitives.scala 122:60:@18004.4]
  assign StickySelects_17_io_ins_2 = io_rPort_6_en_0 & _T_2759; // @[MemPrimitives.scala 122:60:@18005.4]
  assign StickySelects_17_io_ins_3 = io_rPort_7_en_0 & _T_2765; // @[MemPrimitives.scala 122:60:@18006.4]
  assign StickySelects_17_io_ins_4 = io_rPort_9_en_0 & _T_2771; // @[MemPrimitives.scala 122:60:@18007.4]
  assign StickySelects_17_io_ins_5 = io_rPort_11_en_0 & _T_2777; // @[MemPrimitives.scala 122:60:@18008.4]
  assign StickySelects_17_io_ins_6 = io_rPort_12_en_0 & _T_2783; // @[MemPrimitives.scala 122:60:@18009.4]
  assign StickySelects_17_io_ins_7 = io_rPort_13_en_0 & _T_2789; // @[MemPrimitives.scala 122:60:@18010.4]
  assign StickySelects_17_io_ins_8 = io_rPort_16_en_0 & _T_2795; // @[MemPrimitives.scala 122:60:@18011.4]
  assign StickySelects_18_clock = clock; // @[:@18090.4]
  assign StickySelects_18_reset = reset; // @[:@18091.4]
  assign StickySelects_18_io_ins_0 = io_rPort_0_en_0 & _T_2839; // @[MemPrimitives.scala 122:60:@18092.4]
  assign StickySelects_18_io_ins_1 = io_rPort_1_en_0 & _T_2845; // @[MemPrimitives.scala 122:60:@18093.4]
  assign StickySelects_18_io_ins_2 = io_rPort_3_en_0 & _T_2851; // @[MemPrimitives.scala 122:60:@18094.4]
  assign StickySelects_18_io_ins_3 = io_rPort_4_en_0 & _T_2857; // @[MemPrimitives.scala 122:60:@18095.4]
  assign StickySelects_18_io_ins_4 = io_rPort_8_en_0 & _T_2863; // @[MemPrimitives.scala 122:60:@18096.4]
  assign StickySelects_18_io_ins_5 = io_rPort_10_en_0 & _T_2869; // @[MemPrimitives.scala 122:60:@18097.4]
  assign StickySelects_18_io_ins_6 = io_rPort_14_en_0 & _T_2875; // @[MemPrimitives.scala 122:60:@18098.4]
  assign StickySelects_18_io_ins_7 = io_rPort_15_en_0 & _T_2881; // @[MemPrimitives.scala 122:60:@18099.4]
  assign StickySelects_18_io_ins_8 = io_rPort_17_en_0 & _T_2887; // @[MemPrimitives.scala 122:60:@18100.4]
  assign StickySelects_19_clock = clock; // @[:@18179.4]
  assign StickySelects_19_reset = reset; // @[:@18180.4]
  assign StickySelects_19_io_ins_0 = io_rPort_2_en_0 & _T_2931; // @[MemPrimitives.scala 122:60:@18181.4]
  assign StickySelects_19_io_ins_1 = io_rPort_5_en_0 & _T_2937; // @[MemPrimitives.scala 122:60:@18182.4]
  assign StickySelects_19_io_ins_2 = io_rPort_6_en_0 & _T_2943; // @[MemPrimitives.scala 122:60:@18183.4]
  assign StickySelects_19_io_ins_3 = io_rPort_7_en_0 & _T_2949; // @[MemPrimitives.scala 122:60:@18184.4]
  assign StickySelects_19_io_ins_4 = io_rPort_9_en_0 & _T_2955; // @[MemPrimitives.scala 122:60:@18185.4]
  assign StickySelects_19_io_ins_5 = io_rPort_11_en_0 & _T_2961; // @[MemPrimitives.scala 122:60:@18186.4]
  assign StickySelects_19_io_ins_6 = io_rPort_12_en_0 & _T_2967; // @[MemPrimitives.scala 122:60:@18187.4]
  assign StickySelects_19_io_ins_7 = io_rPort_13_en_0 & _T_2973; // @[MemPrimitives.scala 122:60:@18188.4]
  assign StickySelects_19_io_ins_8 = io_rPort_16_en_0 & _T_2979; // @[MemPrimitives.scala 122:60:@18189.4]
  assign StickySelects_20_clock = clock; // @[:@18268.4]
  assign StickySelects_20_reset = reset; // @[:@18269.4]
  assign StickySelects_20_io_ins_0 = io_rPort_0_en_0 & _T_3023; // @[MemPrimitives.scala 122:60:@18270.4]
  assign StickySelects_20_io_ins_1 = io_rPort_1_en_0 & _T_3029; // @[MemPrimitives.scala 122:60:@18271.4]
  assign StickySelects_20_io_ins_2 = io_rPort_3_en_0 & _T_3035; // @[MemPrimitives.scala 122:60:@18272.4]
  assign StickySelects_20_io_ins_3 = io_rPort_4_en_0 & _T_3041; // @[MemPrimitives.scala 122:60:@18273.4]
  assign StickySelects_20_io_ins_4 = io_rPort_8_en_0 & _T_3047; // @[MemPrimitives.scala 122:60:@18274.4]
  assign StickySelects_20_io_ins_5 = io_rPort_10_en_0 & _T_3053; // @[MemPrimitives.scala 122:60:@18275.4]
  assign StickySelects_20_io_ins_6 = io_rPort_14_en_0 & _T_3059; // @[MemPrimitives.scala 122:60:@18276.4]
  assign StickySelects_20_io_ins_7 = io_rPort_15_en_0 & _T_3065; // @[MemPrimitives.scala 122:60:@18277.4]
  assign StickySelects_20_io_ins_8 = io_rPort_17_en_0 & _T_3071; // @[MemPrimitives.scala 122:60:@18278.4]
  assign StickySelects_21_clock = clock; // @[:@18357.4]
  assign StickySelects_21_reset = reset; // @[:@18358.4]
  assign StickySelects_21_io_ins_0 = io_rPort_2_en_0 & _T_3115; // @[MemPrimitives.scala 122:60:@18359.4]
  assign StickySelects_21_io_ins_1 = io_rPort_5_en_0 & _T_3121; // @[MemPrimitives.scala 122:60:@18360.4]
  assign StickySelects_21_io_ins_2 = io_rPort_6_en_0 & _T_3127; // @[MemPrimitives.scala 122:60:@18361.4]
  assign StickySelects_21_io_ins_3 = io_rPort_7_en_0 & _T_3133; // @[MemPrimitives.scala 122:60:@18362.4]
  assign StickySelects_21_io_ins_4 = io_rPort_9_en_0 & _T_3139; // @[MemPrimitives.scala 122:60:@18363.4]
  assign StickySelects_21_io_ins_5 = io_rPort_11_en_0 & _T_3145; // @[MemPrimitives.scala 122:60:@18364.4]
  assign StickySelects_21_io_ins_6 = io_rPort_12_en_0 & _T_3151; // @[MemPrimitives.scala 122:60:@18365.4]
  assign StickySelects_21_io_ins_7 = io_rPort_13_en_0 & _T_3157; // @[MemPrimitives.scala 122:60:@18366.4]
  assign StickySelects_21_io_ins_8 = io_rPort_16_en_0 & _T_3163; // @[MemPrimitives.scala 122:60:@18367.4]
  assign StickySelects_22_clock = clock; // @[:@18446.4]
  assign StickySelects_22_reset = reset; // @[:@18447.4]
  assign StickySelects_22_io_ins_0 = io_rPort_0_en_0 & _T_3207; // @[MemPrimitives.scala 122:60:@18448.4]
  assign StickySelects_22_io_ins_1 = io_rPort_1_en_0 & _T_3213; // @[MemPrimitives.scala 122:60:@18449.4]
  assign StickySelects_22_io_ins_2 = io_rPort_3_en_0 & _T_3219; // @[MemPrimitives.scala 122:60:@18450.4]
  assign StickySelects_22_io_ins_3 = io_rPort_4_en_0 & _T_3225; // @[MemPrimitives.scala 122:60:@18451.4]
  assign StickySelects_22_io_ins_4 = io_rPort_8_en_0 & _T_3231; // @[MemPrimitives.scala 122:60:@18452.4]
  assign StickySelects_22_io_ins_5 = io_rPort_10_en_0 & _T_3237; // @[MemPrimitives.scala 122:60:@18453.4]
  assign StickySelects_22_io_ins_6 = io_rPort_14_en_0 & _T_3243; // @[MemPrimitives.scala 122:60:@18454.4]
  assign StickySelects_22_io_ins_7 = io_rPort_15_en_0 & _T_3249; // @[MemPrimitives.scala 122:60:@18455.4]
  assign StickySelects_22_io_ins_8 = io_rPort_17_en_0 & _T_3255; // @[MemPrimitives.scala 122:60:@18456.4]
  assign StickySelects_23_clock = clock; // @[:@18535.4]
  assign StickySelects_23_reset = reset; // @[:@18536.4]
  assign StickySelects_23_io_ins_0 = io_rPort_2_en_0 & _T_3299; // @[MemPrimitives.scala 122:60:@18537.4]
  assign StickySelects_23_io_ins_1 = io_rPort_5_en_0 & _T_3305; // @[MemPrimitives.scala 122:60:@18538.4]
  assign StickySelects_23_io_ins_2 = io_rPort_6_en_0 & _T_3311; // @[MemPrimitives.scala 122:60:@18539.4]
  assign StickySelects_23_io_ins_3 = io_rPort_7_en_0 & _T_3317; // @[MemPrimitives.scala 122:60:@18540.4]
  assign StickySelects_23_io_ins_4 = io_rPort_9_en_0 & _T_3323; // @[MemPrimitives.scala 122:60:@18541.4]
  assign StickySelects_23_io_ins_5 = io_rPort_11_en_0 & _T_3329; // @[MemPrimitives.scala 122:60:@18542.4]
  assign StickySelects_23_io_ins_6 = io_rPort_12_en_0 & _T_3335; // @[MemPrimitives.scala 122:60:@18543.4]
  assign StickySelects_23_io_ins_7 = io_rPort_13_en_0 & _T_3341; // @[MemPrimitives.scala 122:60:@18544.4]
  assign StickySelects_23_io_ins_8 = io_rPort_16_en_0 & _T_3347; // @[MemPrimitives.scala 122:60:@18545.4]
  assign RetimeWrapper_clock = clock; // @[:@18625.4]
  assign RetimeWrapper_reset = reset; // @[:@18626.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@18628.4]
  assign RetimeWrapper_io_in = _T_1183 & io_rPort_0_en_0; // @[package.scala 94:16:@18627.4]
  assign RetimeWrapper_1_clock = clock; // @[:@18633.4]
  assign RetimeWrapper_1_reset = reset; // @[:@18634.4]
  assign RetimeWrapper_1_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@18636.4]
  assign RetimeWrapper_1_io_in = _T_1367 & io_rPort_0_en_0; // @[package.scala 94:16:@18635.4]
  assign RetimeWrapper_2_clock = clock; // @[:@18641.4]
  assign RetimeWrapper_2_reset = reset; // @[:@18642.4]
  assign RetimeWrapper_2_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@18644.4]
  assign RetimeWrapper_2_io_in = _T_1551 & io_rPort_0_en_0; // @[package.scala 94:16:@18643.4]
  assign RetimeWrapper_3_clock = clock; // @[:@18649.4]
  assign RetimeWrapper_3_reset = reset; // @[:@18650.4]
  assign RetimeWrapper_3_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@18652.4]
  assign RetimeWrapper_3_io_in = _T_1735 & io_rPort_0_en_0; // @[package.scala 94:16:@18651.4]
  assign RetimeWrapper_4_clock = clock; // @[:@18657.4]
  assign RetimeWrapper_4_reset = reset; // @[:@18658.4]
  assign RetimeWrapper_4_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@18660.4]
  assign RetimeWrapper_4_io_in = _T_1919 & io_rPort_0_en_0; // @[package.scala 94:16:@18659.4]
  assign RetimeWrapper_5_clock = clock; // @[:@18665.4]
  assign RetimeWrapper_5_reset = reset; // @[:@18666.4]
  assign RetimeWrapper_5_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@18668.4]
  assign RetimeWrapper_5_io_in = _T_2103 & io_rPort_0_en_0; // @[package.scala 94:16:@18667.4]
  assign RetimeWrapper_6_clock = clock; // @[:@18673.4]
  assign RetimeWrapper_6_reset = reset; // @[:@18674.4]
  assign RetimeWrapper_6_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@18676.4]
  assign RetimeWrapper_6_io_in = _T_2287 & io_rPort_0_en_0; // @[package.scala 94:16:@18675.4]
  assign RetimeWrapper_7_clock = clock; // @[:@18681.4]
  assign RetimeWrapper_7_reset = reset; // @[:@18682.4]
  assign RetimeWrapper_7_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@18684.4]
  assign RetimeWrapper_7_io_in = _T_2471 & io_rPort_0_en_0; // @[package.scala 94:16:@18683.4]
  assign RetimeWrapper_8_clock = clock; // @[:@18689.4]
  assign RetimeWrapper_8_reset = reset; // @[:@18690.4]
  assign RetimeWrapper_8_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@18692.4]
  assign RetimeWrapper_8_io_in = _T_2655 & io_rPort_0_en_0; // @[package.scala 94:16:@18691.4]
  assign RetimeWrapper_9_clock = clock; // @[:@18697.4]
  assign RetimeWrapper_9_reset = reset; // @[:@18698.4]
  assign RetimeWrapper_9_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@18700.4]
  assign RetimeWrapper_9_io_in = _T_2839 & io_rPort_0_en_0; // @[package.scala 94:16:@18699.4]
  assign RetimeWrapper_10_clock = clock; // @[:@18705.4]
  assign RetimeWrapper_10_reset = reset; // @[:@18706.4]
  assign RetimeWrapper_10_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@18708.4]
  assign RetimeWrapper_10_io_in = _T_3023 & io_rPort_0_en_0; // @[package.scala 94:16:@18707.4]
  assign RetimeWrapper_11_clock = clock; // @[:@18713.4]
  assign RetimeWrapper_11_reset = reset; // @[:@18714.4]
  assign RetimeWrapper_11_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@18716.4]
  assign RetimeWrapper_11_io_in = _T_3207 & io_rPort_0_en_0; // @[package.scala 94:16:@18715.4]
  assign RetimeWrapper_12_clock = clock; // @[:@18769.4]
  assign RetimeWrapper_12_reset = reset; // @[:@18770.4]
  assign RetimeWrapper_12_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@18772.4]
  assign RetimeWrapper_12_io_in = _T_1189 & io_rPort_1_en_0; // @[package.scala 94:16:@18771.4]
  assign RetimeWrapper_13_clock = clock; // @[:@18777.4]
  assign RetimeWrapper_13_reset = reset; // @[:@18778.4]
  assign RetimeWrapper_13_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@18780.4]
  assign RetimeWrapper_13_io_in = _T_1373 & io_rPort_1_en_0; // @[package.scala 94:16:@18779.4]
  assign RetimeWrapper_14_clock = clock; // @[:@18785.4]
  assign RetimeWrapper_14_reset = reset; // @[:@18786.4]
  assign RetimeWrapper_14_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@18788.4]
  assign RetimeWrapper_14_io_in = _T_1557 & io_rPort_1_en_0; // @[package.scala 94:16:@18787.4]
  assign RetimeWrapper_15_clock = clock; // @[:@18793.4]
  assign RetimeWrapper_15_reset = reset; // @[:@18794.4]
  assign RetimeWrapper_15_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@18796.4]
  assign RetimeWrapper_15_io_in = _T_1741 & io_rPort_1_en_0; // @[package.scala 94:16:@18795.4]
  assign RetimeWrapper_16_clock = clock; // @[:@18801.4]
  assign RetimeWrapper_16_reset = reset; // @[:@18802.4]
  assign RetimeWrapper_16_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@18804.4]
  assign RetimeWrapper_16_io_in = _T_1925 & io_rPort_1_en_0; // @[package.scala 94:16:@18803.4]
  assign RetimeWrapper_17_clock = clock; // @[:@18809.4]
  assign RetimeWrapper_17_reset = reset; // @[:@18810.4]
  assign RetimeWrapper_17_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@18812.4]
  assign RetimeWrapper_17_io_in = _T_2109 & io_rPort_1_en_0; // @[package.scala 94:16:@18811.4]
  assign RetimeWrapper_18_clock = clock; // @[:@18817.4]
  assign RetimeWrapper_18_reset = reset; // @[:@18818.4]
  assign RetimeWrapper_18_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@18820.4]
  assign RetimeWrapper_18_io_in = _T_2293 & io_rPort_1_en_0; // @[package.scala 94:16:@18819.4]
  assign RetimeWrapper_19_clock = clock; // @[:@18825.4]
  assign RetimeWrapper_19_reset = reset; // @[:@18826.4]
  assign RetimeWrapper_19_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@18828.4]
  assign RetimeWrapper_19_io_in = _T_2477 & io_rPort_1_en_0; // @[package.scala 94:16:@18827.4]
  assign RetimeWrapper_20_clock = clock; // @[:@18833.4]
  assign RetimeWrapper_20_reset = reset; // @[:@18834.4]
  assign RetimeWrapper_20_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@18836.4]
  assign RetimeWrapper_20_io_in = _T_2661 & io_rPort_1_en_0; // @[package.scala 94:16:@18835.4]
  assign RetimeWrapper_21_clock = clock; // @[:@18841.4]
  assign RetimeWrapper_21_reset = reset; // @[:@18842.4]
  assign RetimeWrapper_21_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@18844.4]
  assign RetimeWrapper_21_io_in = _T_2845 & io_rPort_1_en_0; // @[package.scala 94:16:@18843.4]
  assign RetimeWrapper_22_clock = clock; // @[:@18849.4]
  assign RetimeWrapper_22_reset = reset; // @[:@18850.4]
  assign RetimeWrapper_22_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@18852.4]
  assign RetimeWrapper_22_io_in = _T_3029 & io_rPort_1_en_0; // @[package.scala 94:16:@18851.4]
  assign RetimeWrapper_23_clock = clock; // @[:@18857.4]
  assign RetimeWrapper_23_reset = reset; // @[:@18858.4]
  assign RetimeWrapper_23_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@18860.4]
  assign RetimeWrapper_23_io_in = _T_3213 & io_rPort_1_en_0; // @[package.scala 94:16:@18859.4]
  assign RetimeWrapper_24_clock = clock; // @[:@18913.4]
  assign RetimeWrapper_24_reset = reset; // @[:@18914.4]
  assign RetimeWrapper_24_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@18916.4]
  assign RetimeWrapper_24_io_in = _T_1275 & io_rPort_2_en_0; // @[package.scala 94:16:@18915.4]
  assign RetimeWrapper_25_clock = clock; // @[:@18921.4]
  assign RetimeWrapper_25_reset = reset; // @[:@18922.4]
  assign RetimeWrapper_25_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@18924.4]
  assign RetimeWrapper_25_io_in = _T_1459 & io_rPort_2_en_0; // @[package.scala 94:16:@18923.4]
  assign RetimeWrapper_26_clock = clock; // @[:@18929.4]
  assign RetimeWrapper_26_reset = reset; // @[:@18930.4]
  assign RetimeWrapper_26_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@18932.4]
  assign RetimeWrapper_26_io_in = _T_1643 & io_rPort_2_en_0; // @[package.scala 94:16:@18931.4]
  assign RetimeWrapper_27_clock = clock; // @[:@18937.4]
  assign RetimeWrapper_27_reset = reset; // @[:@18938.4]
  assign RetimeWrapper_27_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@18940.4]
  assign RetimeWrapper_27_io_in = _T_1827 & io_rPort_2_en_0; // @[package.scala 94:16:@18939.4]
  assign RetimeWrapper_28_clock = clock; // @[:@18945.4]
  assign RetimeWrapper_28_reset = reset; // @[:@18946.4]
  assign RetimeWrapper_28_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@18948.4]
  assign RetimeWrapper_28_io_in = _T_2011 & io_rPort_2_en_0; // @[package.scala 94:16:@18947.4]
  assign RetimeWrapper_29_clock = clock; // @[:@18953.4]
  assign RetimeWrapper_29_reset = reset; // @[:@18954.4]
  assign RetimeWrapper_29_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@18956.4]
  assign RetimeWrapper_29_io_in = _T_2195 & io_rPort_2_en_0; // @[package.scala 94:16:@18955.4]
  assign RetimeWrapper_30_clock = clock; // @[:@18961.4]
  assign RetimeWrapper_30_reset = reset; // @[:@18962.4]
  assign RetimeWrapper_30_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@18964.4]
  assign RetimeWrapper_30_io_in = _T_2379 & io_rPort_2_en_0; // @[package.scala 94:16:@18963.4]
  assign RetimeWrapper_31_clock = clock; // @[:@18969.4]
  assign RetimeWrapper_31_reset = reset; // @[:@18970.4]
  assign RetimeWrapper_31_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@18972.4]
  assign RetimeWrapper_31_io_in = _T_2563 & io_rPort_2_en_0; // @[package.scala 94:16:@18971.4]
  assign RetimeWrapper_32_clock = clock; // @[:@18977.4]
  assign RetimeWrapper_32_reset = reset; // @[:@18978.4]
  assign RetimeWrapper_32_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@18980.4]
  assign RetimeWrapper_32_io_in = _T_2747 & io_rPort_2_en_0; // @[package.scala 94:16:@18979.4]
  assign RetimeWrapper_33_clock = clock; // @[:@18985.4]
  assign RetimeWrapper_33_reset = reset; // @[:@18986.4]
  assign RetimeWrapper_33_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@18988.4]
  assign RetimeWrapper_33_io_in = _T_2931 & io_rPort_2_en_0; // @[package.scala 94:16:@18987.4]
  assign RetimeWrapper_34_clock = clock; // @[:@18993.4]
  assign RetimeWrapper_34_reset = reset; // @[:@18994.4]
  assign RetimeWrapper_34_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@18996.4]
  assign RetimeWrapper_34_io_in = _T_3115 & io_rPort_2_en_0; // @[package.scala 94:16:@18995.4]
  assign RetimeWrapper_35_clock = clock; // @[:@19001.4]
  assign RetimeWrapper_35_reset = reset; // @[:@19002.4]
  assign RetimeWrapper_35_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@19004.4]
  assign RetimeWrapper_35_io_in = _T_3299 & io_rPort_2_en_0; // @[package.scala 94:16:@19003.4]
  assign RetimeWrapper_36_clock = clock; // @[:@19057.4]
  assign RetimeWrapper_36_reset = reset; // @[:@19058.4]
  assign RetimeWrapper_36_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@19060.4]
  assign RetimeWrapper_36_io_in = _T_1195 & io_rPort_3_en_0; // @[package.scala 94:16:@19059.4]
  assign RetimeWrapper_37_clock = clock; // @[:@19065.4]
  assign RetimeWrapper_37_reset = reset; // @[:@19066.4]
  assign RetimeWrapper_37_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@19068.4]
  assign RetimeWrapper_37_io_in = _T_1379 & io_rPort_3_en_0; // @[package.scala 94:16:@19067.4]
  assign RetimeWrapper_38_clock = clock; // @[:@19073.4]
  assign RetimeWrapper_38_reset = reset; // @[:@19074.4]
  assign RetimeWrapper_38_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@19076.4]
  assign RetimeWrapper_38_io_in = _T_1563 & io_rPort_3_en_0; // @[package.scala 94:16:@19075.4]
  assign RetimeWrapper_39_clock = clock; // @[:@19081.4]
  assign RetimeWrapper_39_reset = reset; // @[:@19082.4]
  assign RetimeWrapper_39_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@19084.4]
  assign RetimeWrapper_39_io_in = _T_1747 & io_rPort_3_en_0; // @[package.scala 94:16:@19083.4]
  assign RetimeWrapper_40_clock = clock; // @[:@19089.4]
  assign RetimeWrapper_40_reset = reset; // @[:@19090.4]
  assign RetimeWrapper_40_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@19092.4]
  assign RetimeWrapper_40_io_in = _T_1931 & io_rPort_3_en_0; // @[package.scala 94:16:@19091.4]
  assign RetimeWrapper_41_clock = clock; // @[:@19097.4]
  assign RetimeWrapper_41_reset = reset; // @[:@19098.4]
  assign RetimeWrapper_41_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@19100.4]
  assign RetimeWrapper_41_io_in = _T_2115 & io_rPort_3_en_0; // @[package.scala 94:16:@19099.4]
  assign RetimeWrapper_42_clock = clock; // @[:@19105.4]
  assign RetimeWrapper_42_reset = reset; // @[:@19106.4]
  assign RetimeWrapper_42_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@19108.4]
  assign RetimeWrapper_42_io_in = _T_2299 & io_rPort_3_en_0; // @[package.scala 94:16:@19107.4]
  assign RetimeWrapper_43_clock = clock; // @[:@19113.4]
  assign RetimeWrapper_43_reset = reset; // @[:@19114.4]
  assign RetimeWrapper_43_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@19116.4]
  assign RetimeWrapper_43_io_in = _T_2483 & io_rPort_3_en_0; // @[package.scala 94:16:@19115.4]
  assign RetimeWrapper_44_clock = clock; // @[:@19121.4]
  assign RetimeWrapper_44_reset = reset; // @[:@19122.4]
  assign RetimeWrapper_44_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@19124.4]
  assign RetimeWrapper_44_io_in = _T_2667 & io_rPort_3_en_0; // @[package.scala 94:16:@19123.4]
  assign RetimeWrapper_45_clock = clock; // @[:@19129.4]
  assign RetimeWrapper_45_reset = reset; // @[:@19130.4]
  assign RetimeWrapper_45_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@19132.4]
  assign RetimeWrapper_45_io_in = _T_2851 & io_rPort_3_en_0; // @[package.scala 94:16:@19131.4]
  assign RetimeWrapper_46_clock = clock; // @[:@19137.4]
  assign RetimeWrapper_46_reset = reset; // @[:@19138.4]
  assign RetimeWrapper_46_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@19140.4]
  assign RetimeWrapper_46_io_in = _T_3035 & io_rPort_3_en_0; // @[package.scala 94:16:@19139.4]
  assign RetimeWrapper_47_clock = clock; // @[:@19145.4]
  assign RetimeWrapper_47_reset = reset; // @[:@19146.4]
  assign RetimeWrapper_47_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@19148.4]
  assign RetimeWrapper_47_io_in = _T_3219 & io_rPort_3_en_0; // @[package.scala 94:16:@19147.4]
  assign RetimeWrapper_48_clock = clock; // @[:@19201.4]
  assign RetimeWrapper_48_reset = reset; // @[:@19202.4]
  assign RetimeWrapper_48_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@19204.4]
  assign RetimeWrapper_48_io_in = _T_1201 & io_rPort_4_en_0; // @[package.scala 94:16:@19203.4]
  assign RetimeWrapper_49_clock = clock; // @[:@19209.4]
  assign RetimeWrapper_49_reset = reset; // @[:@19210.4]
  assign RetimeWrapper_49_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@19212.4]
  assign RetimeWrapper_49_io_in = _T_1385 & io_rPort_4_en_0; // @[package.scala 94:16:@19211.4]
  assign RetimeWrapper_50_clock = clock; // @[:@19217.4]
  assign RetimeWrapper_50_reset = reset; // @[:@19218.4]
  assign RetimeWrapper_50_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@19220.4]
  assign RetimeWrapper_50_io_in = _T_1569 & io_rPort_4_en_0; // @[package.scala 94:16:@19219.4]
  assign RetimeWrapper_51_clock = clock; // @[:@19225.4]
  assign RetimeWrapper_51_reset = reset; // @[:@19226.4]
  assign RetimeWrapper_51_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@19228.4]
  assign RetimeWrapper_51_io_in = _T_1753 & io_rPort_4_en_0; // @[package.scala 94:16:@19227.4]
  assign RetimeWrapper_52_clock = clock; // @[:@19233.4]
  assign RetimeWrapper_52_reset = reset; // @[:@19234.4]
  assign RetimeWrapper_52_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@19236.4]
  assign RetimeWrapper_52_io_in = _T_1937 & io_rPort_4_en_0; // @[package.scala 94:16:@19235.4]
  assign RetimeWrapper_53_clock = clock; // @[:@19241.4]
  assign RetimeWrapper_53_reset = reset; // @[:@19242.4]
  assign RetimeWrapper_53_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@19244.4]
  assign RetimeWrapper_53_io_in = _T_2121 & io_rPort_4_en_0; // @[package.scala 94:16:@19243.4]
  assign RetimeWrapper_54_clock = clock; // @[:@19249.4]
  assign RetimeWrapper_54_reset = reset; // @[:@19250.4]
  assign RetimeWrapper_54_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@19252.4]
  assign RetimeWrapper_54_io_in = _T_2305 & io_rPort_4_en_0; // @[package.scala 94:16:@19251.4]
  assign RetimeWrapper_55_clock = clock; // @[:@19257.4]
  assign RetimeWrapper_55_reset = reset; // @[:@19258.4]
  assign RetimeWrapper_55_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@19260.4]
  assign RetimeWrapper_55_io_in = _T_2489 & io_rPort_4_en_0; // @[package.scala 94:16:@19259.4]
  assign RetimeWrapper_56_clock = clock; // @[:@19265.4]
  assign RetimeWrapper_56_reset = reset; // @[:@19266.4]
  assign RetimeWrapper_56_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@19268.4]
  assign RetimeWrapper_56_io_in = _T_2673 & io_rPort_4_en_0; // @[package.scala 94:16:@19267.4]
  assign RetimeWrapper_57_clock = clock; // @[:@19273.4]
  assign RetimeWrapper_57_reset = reset; // @[:@19274.4]
  assign RetimeWrapper_57_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@19276.4]
  assign RetimeWrapper_57_io_in = _T_2857 & io_rPort_4_en_0; // @[package.scala 94:16:@19275.4]
  assign RetimeWrapper_58_clock = clock; // @[:@19281.4]
  assign RetimeWrapper_58_reset = reset; // @[:@19282.4]
  assign RetimeWrapper_58_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@19284.4]
  assign RetimeWrapper_58_io_in = _T_3041 & io_rPort_4_en_0; // @[package.scala 94:16:@19283.4]
  assign RetimeWrapper_59_clock = clock; // @[:@19289.4]
  assign RetimeWrapper_59_reset = reset; // @[:@19290.4]
  assign RetimeWrapper_59_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@19292.4]
  assign RetimeWrapper_59_io_in = _T_3225 & io_rPort_4_en_0; // @[package.scala 94:16:@19291.4]
  assign RetimeWrapper_60_clock = clock; // @[:@19345.4]
  assign RetimeWrapper_60_reset = reset; // @[:@19346.4]
  assign RetimeWrapper_60_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@19348.4]
  assign RetimeWrapper_60_io_in = _T_1281 & io_rPort_5_en_0; // @[package.scala 94:16:@19347.4]
  assign RetimeWrapper_61_clock = clock; // @[:@19353.4]
  assign RetimeWrapper_61_reset = reset; // @[:@19354.4]
  assign RetimeWrapper_61_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@19356.4]
  assign RetimeWrapper_61_io_in = _T_1465 & io_rPort_5_en_0; // @[package.scala 94:16:@19355.4]
  assign RetimeWrapper_62_clock = clock; // @[:@19361.4]
  assign RetimeWrapper_62_reset = reset; // @[:@19362.4]
  assign RetimeWrapper_62_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@19364.4]
  assign RetimeWrapper_62_io_in = _T_1649 & io_rPort_5_en_0; // @[package.scala 94:16:@19363.4]
  assign RetimeWrapper_63_clock = clock; // @[:@19369.4]
  assign RetimeWrapper_63_reset = reset; // @[:@19370.4]
  assign RetimeWrapper_63_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@19372.4]
  assign RetimeWrapper_63_io_in = _T_1833 & io_rPort_5_en_0; // @[package.scala 94:16:@19371.4]
  assign RetimeWrapper_64_clock = clock; // @[:@19377.4]
  assign RetimeWrapper_64_reset = reset; // @[:@19378.4]
  assign RetimeWrapper_64_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@19380.4]
  assign RetimeWrapper_64_io_in = _T_2017 & io_rPort_5_en_0; // @[package.scala 94:16:@19379.4]
  assign RetimeWrapper_65_clock = clock; // @[:@19385.4]
  assign RetimeWrapper_65_reset = reset; // @[:@19386.4]
  assign RetimeWrapper_65_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@19388.4]
  assign RetimeWrapper_65_io_in = _T_2201 & io_rPort_5_en_0; // @[package.scala 94:16:@19387.4]
  assign RetimeWrapper_66_clock = clock; // @[:@19393.4]
  assign RetimeWrapper_66_reset = reset; // @[:@19394.4]
  assign RetimeWrapper_66_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@19396.4]
  assign RetimeWrapper_66_io_in = _T_2385 & io_rPort_5_en_0; // @[package.scala 94:16:@19395.4]
  assign RetimeWrapper_67_clock = clock; // @[:@19401.4]
  assign RetimeWrapper_67_reset = reset; // @[:@19402.4]
  assign RetimeWrapper_67_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@19404.4]
  assign RetimeWrapper_67_io_in = _T_2569 & io_rPort_5_en_0; // @[package.scala 94:16:@19403.4]
  assign RetimeWrapper_68_clock = clock; // @[:@19409.4]
  assign RetimeWrapper_68_reset = reset; // @[:@19410.4]
  assign RetimeWrapper_68_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@19412.4]
  assign RetimeWrapper_68_io_in = _T_2753 & io_rPort_5_en_0; // @[package.scala 94:16:@19411.4]
  assign RetimeWrapper_69_clock = clock; // @[:@19417.4]
  assign RetimeWrapper_69_reset = reset; // @[:@19418.4]
  assign RetimeWrapper_69_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@19420.4]
  assign RetimeWrapper_69_io_in = _T_2937 & io_rPort_5_en_0; // @[package.scala 94:16:@19419.4]
  assign RetimeWrapper_70_clock = clock; // @[:@19425.4]
  assign RetimeWrapper_70_reset = reset; // @[:@19426.4]
  assign RetimeWrapper_70_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@19428.4]
  assign RetimeWrapper_70_io_in = _T_3121 & io_rPort_5_en_0; // @[package.scala 94:16:@19427.4]
  assign RetimeWrapper_71_clock = clock; // @[:@19433.4]
  assign RetimeWrapper_71_reset = reset; // @[:@19434.4]
  assign RetimeWrapper_71_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@19436.4]
  assign RetimeWrapper_71_io_in = _T_3305 & io_rPort_5_en_0; // @[package.scala 94:16:@19435.4]
  assign RetimeWrapper_72_clock = clock; // @[:@19489.4]
  assign RetimeWrapper_72_reset = reset; // @[:@19490.4]
  assign RetimeWrapper_72_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@19492.4]
  assign RetimeWrapper_72_io_in = _T_1287 & io_rPort_6_en_0; // @[package.scala 94:16:@19491.4]
  assign RetimeWrapper_73_clock = clock; // @[:@19497.4]
  assign RetimeWrapper_73_reset = reset; // @[:@19498.4]
  assign RetimeWrapper_73_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@19500.4]
  assign RetimeWrapper_73_io_in = _T_1471 & io_rPort_6_en_0; // @[package.scala 94:16:@19499.4]
  assign RetimeWrapper_74_clock = clock; // @[:@19505.4]
  assign RetimeWrapper_74_reset = reset; // @[:@19506.4]
  assign RetimeWrapper_74_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@19508.4]
  assign RetimeWrapper_74_io_in = _T_1655 & io_rPort_6_en_0; // @[package.scala 94:16:@19507.4]
  assign RetimeWrapper_75_clock = clock; // @[:@19513.4]
  assign RetimeWrapper_75_reset = reset; // @[:@19514.4]
  assign RetimeWrapper_75_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@19516.4]
  assign RetimeWrapper_75_io_in = _T_1839 & io_rPort_6_en_0; // @[package.scala 94:16:@19515.4]
  assign RetimeWrapper_76_clock = clock; // @[:@19521.4]
  assign RetimeWrapper_76_reset = reset; // @[:@19522.4]
  assign RetimeWrapper_76_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@19524.4]
  assign RetimeWrapper_76_io_in = _T_2023 & io_rPort_6_en_0; // @[package.scala 94:16:@19523.4]
  assign RetimeWrapper_77_clock = clock; // @[:@19529.4]
  assign RetimeWrapper_77_reset = reset; // @[:@19530.4]
  assign RetimeWrapper_77_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@19532.4]
  assign RetimeWrapper_77_io_in = _T_2207 & io_rPort_6_en_0; // @[package.scala 94:16:@19531.4]
  assign RetimeWrapper_78_clock = clock; // @[:@19537.4]
  assign RetimeWrapper_78_reset = reset; // @[:@19538.4]
  assign RetimeWrapper_78_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@19540.4]
  assign RetimeWrapper_78_io_in = _T_2391 & io_rPort_6_en_0; // @[package.scala 94:16:@19539.4]
  assign RetimeWrapper_79_clock = clock; // @[:@19545.4]
  assign RetimeWrapper_79_reset = reset; // @[:@19546.4]
  assign RetimeWrapper_79_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@19548.4]
  assign RetimeWrapper_79_io_in = _T_2575 & io_rPort_6_en_0; // @[package.scala 94:16:@19547.4]
  assign RetimeWrapper_80_clock = clock; // @[:@19553.4]
  assign RetimeWrapper_80_reset = reset; // @[:@19554.4]
  assign RetimeWrapper_80_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@19556.4]
  assign RetimeWrapper_80_io_in = _T_2759 & io_rPort_6_en_0; // @[package.scala 94:16:@19555.4]
  assign RetimeWrapper_81_clock = clock; // @[:@19561.4]
  assign RetimeWrapper_81_reset = reset; // @[:@19562.4]
  assign RetimeWrapper_81_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@19564.4]
  assign RetimeWrapper_81_io_in = _T_2943 & io_rPort_6_en_0; // @[package.scala 94:16:@19563.4]
  assign RetimeWrapper_82_clock = clock; // @[:@19569.4]
  assign RetimeWrapper_82_reset = reset; // @[:@19570.4]
  assign RetimeWrapper_82_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@19572.4]
  assign RetimeWrapper_82_io_in = _T_3127 & io_rPort_6_en_0; // @[package.scala 94:16:@19571.4]
  assign RetimeWrapper_83_clock = clock; // @[:@19577.4]
  assign RetimeWrapper_83_reset = reset; // @[:@19578.4]
  assign RetimeWrapper_83_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@19580.4]
  assign RetimeWrapper_83_io_in = _T_3311 & io_rPort_6_en_0; // @[package.scala 94:16:@19579.4]
  assign RetimeWrapper_84_clock = clock; // @[:@19633.4]
  assign RetimeWrapper_84_reset = reset; // @[:@19634.4]
  assign RetimeWrapper_84_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@19636.4]
  assign RetimeWrapper_84_io_in = _T_1293 & io_rPort_7_en_0; // @[package.scala 94:16:@19635.4]
  assign RetimeWrapper_85_clock = clock; // @[:@19641.4]
  assign RetimeWrapper_85_reset = reset; // @[:@19642.4]
  assign RetimeWrapper_85_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@19644.4]
  assign RetimeWrapper_85_io_in = _T_1477 & io_rPort_7_en_0; // @[package.scala 94:16:@19643.4]
  assign RetimeWrapper_86_clock = clock; // @[:@19649.4]
  assign RetimeWrapper_86_reset = reset; // @[:@19650.4]
  assign RetimeWrapper_86_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@19652.4]
  assign RetimeWrapper_86_io_in = _T_1661 & io_rPort_7_en_0; // @[package.scala 94:16:@19651.4]
  assign RetimeWrapper_87_clock = clock; // @[:@19657.4]
  assign RetimeWrapper_87_reset = reset; // @[:@19658.4]
  assign RetimeWrapper_87_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@19660.4]
  assign RetimeWrapper_87_io_in = _T_1845 & io_rPort_7_en_0; // @[package.scala 94:16:@19659.4]
  assign RetimeWrapper_88_clock = clock; // @[:@19665.4]
  assign RetimeWrapper_88_reset = reset; // @[:@19666.4]
  assign RetimeWrapper_88_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@19668.4]
  assign RetimeWrapper_88_io_in = _T_2029 & io_rPort_7_en_0; // @[package.scala 94:16:@19667.4]
  assign RetimeWrapper_89_clock = clock; // @[:@19673.4]
  assign RetimeWrapper_89_reset = reset; // @[:@19674.4]
  assign RetimeWrapper_89_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@19676.4]
  assign RetimeWrapper_89_io_in = _T_2213 & io_rPort_7_en_0; // @[package.scala 94:16:@19675.4]
  assign RetimeWrapper_90_clock = clock; // @[:@19681.4]
  assign RetimeWrapper_90_reset = reset; // @[:@19682.4]
  assign RetimeWrapper_90_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@19684.4]
  assign RetimeWrapper_90_io_in = _T_2397 & io_rPort_7_en_0; // @[package.scala 94:16:@19683.4]
  assign RetimeWrapper_91_clock = clock; // @[:@19689.4]
  assign RetimeWrapper_91_reset = reset; // @[:@19690.4]
  assign RetimeWrapper_91_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@19692.4]
  assign RetimeWrapper_91_io_in = _T_2581 & io_rPort_7_en_0; // @[package.scala 94:16:@19691.4]
  assign RetimeWrapper_92_clock = clock; // @[:@19697.4]
  assign RetimeWrapper_92_reset = reset; // @[:@19698.4]
  assign RetimeWrapper_92_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@19700.4]
  assign RetimeWrapper_92_io_in = _T_2765 & io_rPort_7_en_0; // @[package.scala 94:16:@19699.4]
  assign RetimeWrapper_93_clock = clock; // @[:@19705.4]
  assign RetimeWrapper_93_reset = reset; // @[:@19706.4]
  assign RetimeWrapper_93_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@19708.4]
  assign RetimeWrapper_93_io_in = _T_2949 & io_rPort_7_en_0; // @[package.scala 94:16:@19707.4]
  assign RetimeWrapper_94_clock = clock; // @[:@19713.4]
  assign RetimeWrapper_94_reset = reset; // @[:@19714.4]
  assign RetimeWrapper_94_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@19716.4]
  assign RetimeWrapper_94_io_in = _T_3133 & io_rPort_7_en_0; // @[package.scala 94:16:@19715.4]
  assign RetimeWrapper_95_clock = clock; // @[:@19721.4]
  assign RetimeWrapper_95_reset = reset; // @[:@19722.4]
  assign RetimeWrapper_95_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@19724.4]
  assign RetimeWrapper_95_io_in = _T_3317 & io_rPort_7_en_0; // @[package.scala 94:16:@19723.4]
  assign RetimeWrapper_96_clock = clock; // @[:@19777.4]
  assign RetimeWrapper_96_reset = reset; // @[:@19778.4]
  assign RetimeWrapper_96_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@19780.4]
  assign RetimeWrapper_96_io_in = _T_1207 & io_rPort_8_en_0; // @[package.scala 94:16:@19779.4]
  assign RetimeWrapper_97_clock = clock; // @[:@19785.4]
  assign RetimeWrapper_97_reset = reset; // @[:@19786.4]
  assign RetimeWrapper_97_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@19788.4]
  assign RetimeWrapper_97_io_in = _T_1391 & io_rPort_8_en_0; // @[package.scala 94:16:@19787.4]
  assign RetimeWrapper_98_clock = clock; // @[:@19793.4]
  assign RetimeWrapper_98_reset = reset; // @[:@19794.4]
  assign RetimeWrapper_98_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@19796.4]
  assign RetimeWrapper_98_io_in = _T_1575 & io_rPort_8_en_0; // @[package.scala 94:16:@19795.4]
  assign RetimeWrapper_99_clock = clock; // @[:@19801.4]
  assign RetimeWrapper_99_reset = reset; // @[:@19802.4]
  assign RetimeWrapper_99_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@19804.4]
  assign RetimeWrapper_99_io_in = _T_1759 & io_rPort_8_en_0; // @[package.scala 94:16:@19803.4]
  assign RetimeWrapper_100_clock = clock; // @[:@19809.4]
  assign RetimeWrapper_100_reset = reset; // @[:@19810.4]
  assign RetimeWrapper_100_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@19812.4]
  assign RetimeWrapper_100_io_in = _T_1943 & io_rPort_8_en_0; // @[package.scala 94:16:@19811.4]
  assign RetimeWrapper_101_clock = clock; // @[:@19817.4]
  assign RetimeWrapper_101_reset = reset; // @[:@19818.4]
  assign RetimeWrapper_101_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@19820.4]
  assign RetimeWrapper_101_io_in = _T_2127 & io_rPort_8_en_0; // @[package.scala 94:16:@19819.4]
  assign RetimeWrapper_102_clock = clock; // @[:@19825.4]
  assign RetimeWrapper_102_reset = reset; // @[:@19826.4]
  assign RetimeWrapper_102_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@19828.4]
  assign RetimeWrapper_102_io_in = _T_2311 & io_rPort_8_en_0; // @[package.scala 94:16:@19827.4]
  assign RetimeWrapper_103_clock = clock; // @[:@19833.4]
  assign RetimeWrapper_103_reset = reset; // @[:@19834.4]
  assign RetimeWrapper_103_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@19836.4]
  assign RetimeWrapper_103_io_in = _T_2495 & io_rPort_8_en_0; // @[package.scala 94:16:@19835.4]
  assign RetimeWrapper_104_clock = clock; // @[:@19841.4]
  assign RetimeWrapper_104_reset = reset; // @[:@19842.4]
  assign RetimeWrapper_104_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@19844.4]
  assign RetimeWrapper_104_io_in = _T_2679 & io_rPort_8_en_0; // @[package.scala 94:16:@19843.4]
  assign RetimeWrapper_105_clock = clock; // @[:@19849.4]
  assign RetimeWrapper_105_reset = reset; // @[:@19850.4]
  assign RetimeWrapper_105_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@19852.4]
  assign RetimeWrapper_105_io_in = _T_2863 & io_rPort_8_en_0; // @[package.scala 94:16:@19851.4]
  assign RetimeWrapper_106_clock = clock; // @[:@19857.4]
  assign RetimeWrapper_106_reset = reset; // @[:@19858.4]
  assign RetimeWrapper_106_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@19860.4]
  assign RetimeWrapper_106_io_in = _T_3047 & io_rPort_8_en_0; // @[package.scala 94:16:@19859.4]
  assign RetimeWrapper_107_clock = clock; // @[:@19865.4]
  assign RetimeWrapper_107_reset = reset; // @[:@19866.4]
  assign RetimeWrapper_107_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@19868.4]
  assign RetimeWrapper_107_io_in = _T_3231 & io_rPort_8_en_0; // @[package.scala 94:16:@19867.4]
  assign RetimeWrapper_108_clock = clock; // @[:@19921.4]
  assign RetimeWrapper_108_reset = reset; // @[:@19922.4]
  assign RetimeWrapper_108_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@19924.4]
  assign RetimeWrapper_108_io_in = _T_1299 & io_rPort_9_en_0; // @[package.scala 94:16:@19923.4]
  assign RetimeWrapper_109_clock = clock; // @[:@19929.4]
  assign RetimeWrapper_109_reset = reset; // @[:@19930.4]
  assign RetimeWrapper_109_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@19932.4]
  assign RetimeWrapper_109_io_in = _T_1483 & io_rPort_9_en_0; // @[package.scala 94:16:@19931.4]
  assign RetimeWrapper_110_clock = clock; // @[:@19937.4]
  assign RetimeWrapper_110_reset = reset; // @[:@19938.4]
  assign RetimeWrapper_110_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@19940.4]
  assign RetimeWrapper_110_io_in = _T_1667 & io_rPort_9_en_0; // @[package.scala 94:16:@19939.4]
  assign RetimeWrapper_111_clock = clock; // @[:@19945.4]
  assign RetimeWrapper_111_reset = reset; // @[:@19946.4]
  assign RetimeWrapper_111_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@19948.4]
  assign RetimeWrapper_111_io_in = _T_1851 & io_rPort_9_en_0; // @[package.scala 94:16:@19947.4]
  assign RetimeWrapper_112_clock = clock; // @[:@19953.4]
  assign RetimeWrapper_112_reset = reset; // @[:@19954.4]
  assign RetimeWrapper_112_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@19956.4]
  assign RetimeWrapper_112_io_in = _T_2035 & io_rPort_9_en_0; // @[package.scala 94:16:@19955.4]
  assign RetimeWrapper_113_clock = clock; // @[:@19961.4]
  assign RetimeWrapper_113_reset = reset; // @[:@19962.4]
  assign RetimeWrapper_113_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@19964.4]
  assign RetimeWrapper_113_io_in = _T_2219 & io_rPort_9_en_0; // @[package.scala 94:16:@19963.4]
  assign RetimeWrapper_114_clock = clock; // @[:@19969.4]
  assign RetimeWrapper_114_reset = reset; // @[:@19970.4]
  assign RetimeWrapper_114_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@19972.4]
  assign RetimeWrapper_114_io_in = _T_2403 & io_rPort_9_en_0; // @[package.scala 94:16:@19971.4]
  assign RetimeWrapper_115_clock = clock; // @[:@19977.4]
  assign RetimeWrapper_115_reset = reset; // @[:@19978.4]
  assign RetimeWrapper_115_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@19980.4]
  assign RetimeWrapper_115_io_in = _T_2587 & io_rPort_9_en_0; // @[package.scala 94:16:@19979.4]
  assign RetimeWrapper_116_clock = clock; // @[:@19985.4]
  assign RetimeWrapper_116_reset = reset; // @[:@19986.4]
  assign RetimeWrapper_116_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@19988.4]
  assign RetimeWrapper_116_io_in = _T_2771 & io_rPort_9_en_0; // @[package.scala 94:16:@19987.4]
  assign RetimeWrapper_117_clock = clock; // @[:@19993.4]
  assign RetimeWrapper_117_reset = reset; // @[:@19994.4]
  assign RetimeWrapper_117_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@19996.4]
  assign RetimeWrapper_117_io_in = _T_2955 & io_rPort_9_en_0; // @[package.scala 94:16:@19995.4]
  assign RetimeWrapper_118_clock = clock; // @[:@20001.4]
  assign RetimeWrapper_118_reset = reset; // @[:@20002.4]
  assign RetimeWrapper_118_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@20004.4]
  assign RetimeWrapper_118_io_in = _T_3139 & io_rPort_9_en_0; // @[package.scala 94:16:@20003.4]
  assign RetimeWrapper_119_clock = clock; // @[:@20009.4]
  assign RetimeWrapper_119_reset = reset; // @[:@20010.4]
  assign RetimeWrapper_119_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@20012.4]
  assign RetimeWrapper_119_io_in = _T_3323 & io_rPort_9_en_0; // @[package.scala 94:16:@20011.4]
  assign RetimeWrapper_120_clock = clock; // @[:@20065.4]
  assign RetimeWrapper_120_reset = reset; // @[:@20066.4]
  assign RetimeWrapper_120_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@20068.4]
  assign RetimeWrapper_120_io_in = _T_1213 & io_rPort_10_en_0; // @[package.scala 94:16:@20067.4]
  assign RetimeWrapper_121_clock = clock; // @[:@20073.4]
  assign RetimeWrapper_121_reset = reset; // @[:@20074.4]
  assign RetimeWrapper_121_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@20076.4]
  assign RetimeWrapper_121_io_in = _T_1397 & io_rPort_10_en_0; // @[package.scala 94:16:@20075.4]
  assign RetimeWrapper_122_clock = clock; // @[:@20081.4]
  assign RetimeWrapper_122_reset = reset; // @[:@20082.4]
  assign RetimeWrapper_122_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@20084.4]
  assign RetimeWrapper_122_io_in = _T_1581 & io_rPort_10_en_0; // @[package.scala 94:16:@20083.4]
  assign RetimeWrapper_123_clock = clock; // @[:@20089.4]
  assign RetimeWrapper_123_reset = reset; // @[:@20090.4]
  assign RetimeWrapper_123_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@20092.4]
  assign RetimeWrapper_123_io_in = _T_1765 & io_rPort_10_en_0; // @[package.scala 94:16:@20091.4]
  assign RetimeWrapper_124_clock = clock; // @[:@20097.4]
  assign RetimeWrapper_124_reset = reset; // @[:@20098.4]
  assign RetimeWrapper_124_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@20100.4]
  assign RetimeWrapper_124_io_in = _T_1949 & io_rPort_10_en_0; // @[package.scala 94:16:@20099.4]
  assign RetimeWrapper_125_clock = clock; // @[:@20105.4]
  assign RetimeWrapper_125_reset = reset; // @[:@20106.4]
  assign RetimeWrapper_125_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@20108.4]
  assign RetimeWrapper_125_io_in = _T_2133 & io_rPort_10_en_0; // @[package.scala 94:16:@20107.4]
  assign RetimeWrapper_126_clock = clock; // @[:@20113.4]
  assign RetimeWrapper_126_reset = reset; // @[:@20114.4]
  assign RetimeWrapper_126_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@20116.4]
  assign RetimeWrapper_126_io_in = _T_2317 & io_rPort_10_en_0; // @[package.scala 94:16:@20115.4]
  assign RetimeWrapper_127_clock = clock; // @[:@20121.4]
  assign RetimeWrapper_127_reset = reset; // @[:@20122.4]
  assign RetimeWrapper_127_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@20124.4]
  assign RetimeWrapper_127_io_in = _T_2501 & io_rPort_10_en_0; // @[package.scala 94:16:@20123.4]
  assign RetimeWrapper_128_clock = clock; // @[:@20129.4]
  assign RetimeWrapper_128_reset = reset; // @[:@20130.4]
  assign RetimeWrapper_128_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@20132.4]
  assign RetimeWrapper_128_io_in = _T_2685 & io_rPort_10_en_0; // @[package.scala 94:16:@20131.4]
  assign RetimeWrapper_129_clock = clock; // @[:@20137.4]
  assign RetimeWrapper_129_reset = reset; // @[:@20138.4]
  assign RetimeWrapper_129_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@20140.4]
  assign RetimeWrapper_129_io_in = _T_2869 & io_rPort_10_en_0; // @[package.scala 94:16:@20139.4]
  assign RetimeWrapper_130_clock = clock; // @[:@20145.4]
  assign RetimeWrapper_130_reset = reset; // @[:@20146.4]
  assign RetimeWrapper_130_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@20148.4]
  assign RetimeWrapper_130_io_in = _T_3053 & io_rPort_10_en_0; // @[package.scala 94:16:@20147.4]
  assign RetimeWrapper_131_clock = clock; // @[:@20153.4]
  assign RetimeWrapper_131_reset = reset; // @[:@20154.4]
  assign RetimeWrapper_131_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@20156.4]
  assign RetimeWrapper_131_io_in = _T_3237 & io_rPort_10_en_0; // @[package.scala 94:16:@20155.4]
  assign RetimeWrapper_132_clock = clock; // @[:@20209.4]
  assign RetimeWrapper_132_reset = reset; // @[:@20210.4]
  assign RetimeWrapper_132_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@20212.4]
  assign RetimeWrapper_132_io_in = _T_1305 & io_rPort_11_en_0; // @[package.scala 94:16:@20211.4]
  assign RetimeWrapper_133_clock = clock; // @[:@20217.4]
  assign RetimeWrapper_133_reset = reset; // @[:@20218.4]
  assign RetimeWrapper_133_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@20220.4]
  assign RetimeWrapper_133_io_in = _T_1489 & io_rPort_11_en_0; // @[package.scala 94:16:@20219.4]
  assign RetimeWrapper_134_clock = clock; // @[:@20225.4]
  assign RetimeWrapper_134_reset = reset; // @[:@20226.4]
  assign RetimeWrapper_134_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@20228.4]
  assign RetimeWrapper_134_io_in = _T_1673 & io_rPort_11_en_0; // @[package.scala 94:16:@20227.4]
  assign RetimeWrapper_135_clock = clock; // @[:@20233.4]
  assign RetimeWrapper_135_reset = reset; // @[:@20234.4]
  assign RetimeWrapper_135_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@20236.4]
  assign RetimeWrapper_135_io_in = _T_1857 & io_rPort_11_en_0; // @[package.scala 94:16:@20235.4]
  assign RetimeWrapper_136_clock = clock; // @[:@20241.4]
  assign RetimeWrapper_136_reset = reset; // @[:@20242.4]
  assign RetimeWrapper_136_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@20244.4]
  assign RetimeWrapper_136_io_in = _T_2041 & io_rPort_11_en_0; // @[package.scala 94:16:@20243.4]
  assign RetimeWrapper_137_clock = clock; // @[:@20249.4]
  assign RetimeWrapper_137_reset = reset; // @[:@20250.4]
  assign RetimeWrapper_137_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@20252.4]
  assign RetimeWrapper_137_io_in = _T_2225 & io_rPort_11_en_0; // @[package.scala 94:16:@20251.4]
  assign RetimeWrapper_138_clock = clock; // @[:@20257.4]
  assign RetimeWrapper_138_reset = reset; // @[:@20258.4]
  assign RetimeWrapper_138_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@20260.4]
  assign RetimeWrapper_138_io_in = _T_2409 & io_rPort_11_en_0; // @[package.scala 94:16:@20259.4]
  assign RetimeWrapper_139_clock = clock; // @[:@20265.4]
  assign RetimeWrapper_139_reset = reset; // @[:@20266.4]
  assign RetimeWrapper_139_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@20268.4]
  assign RetimeWrapper_139_io_in = _T_2593 & io_rPort_11_en_0; // @[package.scala 94:16:@20267.4]
  assign RetimeWrapper_140_clock = clock; // @[:@20273.4]
  assign RetimeWrapper_140_reset = reset; // @[:@20274.4]
  assign RetimeWrapper_140_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@20276.4]
  assign RetimeWrapper_140_io_in = _T_2777 & io_rPort_11_en_0; // @[package.scala 94:16:@20275.4]
  assign RetimeWrapper_141_clock = clock; // @[:@20281.4]
  assign RetimeWrapper_141_reset = reset; // @[:@20282.4]
  assign RetimeWrapper_141_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@20284.4]
  assign RetimeWrapper_141_io_in = _T_2961 & io_rPort_11_en_0; // @[package.scala 94:16:@20283.4]
  assign RetimeWrapper_142_clock = clock; // @[:@20289.4]
  assign RetimeWrapper_142_reset = reset; // @[:@20290.4]
  assign RetimeWrapper_142_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@20292.4]
  assign RetimeWrapper_142_io_in = _T_3145 & io_rPort_11_en_0; // @[package.scala 94:16:@20291.4]
  assign RetimeWrapper_143_clock = clock; // @[:@20297.4]
  assign RetimeWrapper_143_reset = reset; // @[:@20298.4]
  assign RetimeWrapper_143_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@20300.4]
  assign RetimeWrapper_143_io_in = _T_3329 & io_rPort_11_en_0; // @[package.scala 94:16:@20299.4]
  assign RetimeWrapper_144_clock = clock; // @[:@20353.4]
  assign RetimeWrapper_144_reset = reset; // @[:@20354.4]
  assign RetimeWrapper_144_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@20356.4]
  assign RetimeWrapper_144_io_in = _T_1311 & io_rPort_12_en_0; // @[package.scala 94:16:@20355.4]
  assign RetimeWrapper_145_clock = clock; // @[:@20361.4]
  assign RetimeWrapper_145_reset = reset; // @[:@20362.4]
  assign RetimeWrapper_145_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@20364.4]
  assign RetimeWrapper_145_io_in = _T_1495 & io_rPort_12_en_0; // @[package.scala 94:16:@20363.4]
  assign RetimeWrapper_146_clock = clock; // @[:@20369.4]
  assign RetimeWrapper_146_reset = reset; // @[:@20370.4]
  assign RetimeWrapper_146_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@20372.4]
  assign RetimeWrapper_146_io_in = _T_1679 & io_rPort_12_en_0; // @[package.scala 94:16:@20371.4]
  assign RetimeWrapper_147_clock = clock; // @[:@20377.4]
  assign RetimeWrapper_147_reset = reset; // @[:@20378.4]
  assign RetimeWrapper_147_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@20380.4]
  assign RetimeWrapper_147_io_in = _T_1863 & io_rPort_12_en_0; // @[package.scala 94:16:@20379.4]
  assign RetimeWrapper_148_clock = clock; // @[:@20385.4]
  assign RetimeWrapper_148_reset = reset; // @[:@20386.4]
  assign RetimeWrapper_148_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@20388.4]
  assign RetimeWrapper_148_io_in = _T_2047 & io_rPort_12_en_0; // @[package.scala 94:16:@20387.4]
  assign RetimeWrapper_149_clock = clock; // @[:@20393.4]
  assign RetimeWrapper_149_reset = reset; // @[:@20394.4]
  assign RetimeWrapper_149_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@20396.4]
  assign RetimeWrapper_149_io_in = _T_2231 & io_rPort_12_en_0; // @[package.scala 94:16:@20395.4]
  assign RetimeWrapper_150_clock = clock; // @[:@20401.4]
  assign RetimeWrapper_150_reset = reset; // @[:@20402.4]
  assign RetimeWrapper_150_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@20404.4]
  assign RetimeWrapper_150_io_in = _T_2415 & io_rPort_12_en_0; // @[package.scala 94:16:@20403.4]
  assign RetimeWrapper_151_clock = clock; // @[:@20409.4]
  assign RetimeWrapper_151_reset = reset; // @[:@20410.4]
  assign RetimeWrapper_151_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@20412.4]
  assign RetimeWrapper_151_io_in = _T_2599 & io_rPort_12_en_0; // @[package.scala 94:16:@20411.4]
  assign RetimeWrapper_152_clock = clock; // @[:@20417.4]
  assign RetimeWrapper_152_reset = reset; // @[:@20418.4]
  assign RetimeWrapper_152_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@20420.4]
  assign RetimeWrapper_152_io_in = _T_2783 & io_rPort_12_en_0; // @[package.scala 94:16:@20419.4]
  assign RetimeWrapper_153_clock = clock; // @[:@20425.4]
  assign RetimeWrapper_153_reset = reset; // @[:@20426.4]
  assign RetimeWrapper_153_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@20428.4]
  assign RetimeWrapper_153_io_in = _T_2967 & io_rPort_12_en_0; // @[package.scala 94:16:@20427.4]
  assign RetimeWrapper_154_clock = clock; // @[:@20433.4]
  assign RetimeWrapper_154_reset = reset; // @[:@20434.4]
  assign RetimeWrapper_154_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@20436.4]
  assign RetimeWrapper_154_io_in = _T_3151 & io_rPort_12_en_0; // @[package.scala 94:16:@20435.4]
  assign RetimeWrapper_155_clock = clock; // @[:@20441.4]
  assign RetimeWrapper_155_reset = reset; // @[:@20442.4]
  assign RetimeWrapper_155_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@20444.4]
  assign RetimeWrapper_155_io_in = _T_3335 & io_rPort_12_en_0; // @[package.scala 94:16:@20443.4]
  assign RetimeWrapper_156_clock = clock; // @[:@20497.4]
  assign RetimeWrapper_156_reset = reset; // @[:@20498.4]
  assign RetimeWrapper_156_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@20500.4]
  assign RetimeWrapper_156_io_in = _T_1317 & io_rPort_13_en_0; // @[package.scala 94:16:@20499.4]
  assign RetimeWrapper_157_clock = clock; // @[:@20505.4]
  assign RetimeWrapper_157_reset = reset; // @[:@20506.4]
  assign RetimeWrapper_157_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@20508.4]
  assign RetimeWrapper_157_io_in = _T_1501 & io_rPort_13_en_0; // @[package.scala 94:16:@20507.4]
  assign RetimeWrapper_158_clock = clock; // @[:@20513.4]
  assign RetimeWrapper_158_reset = reset; // @[:@20514.4]
  assign RetimeWrapper_158_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@20516.4]
  assign RetimeWrapper_158_io_in = _T_1685 & io_rPort_13_en_0; // @[package.scala 94:16:@20515.4]
  assign RetimeWrapper_159_clock = clock; // @[:@20521.4]
  assign RetimeWrapper_159_reset = reset; // @[:@20522.4]
  assign RetimeWrapper_159_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@20524.4]
  assign RetimeWrapper_159_io_in = _T_1869 & io_rPort_13_en_0; // @[package.scala 94:16:@20523.4]
  assign RetimeWrapper_160_clock = clock; // @[:@20529.4]
  assign RetimeWrapper_160_reset = reset; // @[:@20530.4]
  assign RetimeWrapper_160_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@20532.4]
  assign RetimeWrapper_160_io_in = _T_2053 & io_rPort_13_en_0; // @[package.scala 94:16:@20531.4]
  assign RetimeWrapper_161_clock = clock; // @[:@20537.4]
  assign RetimeWrapper_161_reset = reset; // @[:@20538.4]
  assign RetimeWrapper_161_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@20540.4]
  assign RetimeWrapper_161_io_in = _T_2237 & io_rPort_13_en_0; // @[package.scala 94:16:@20539.4]
  assign RetimeWrapper_162_clock = clock; // @[:@20545.4]
  assign RetimeWrapper_162_reset = reset; // @[:@20546.4]
  assign RetimeWrapper_162_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@20548.4]
  assign RetimeWrapper_162_io_in = _T_2421 & io_rPort_13_en_0; // @[package.scala 94:16:@20547.4]
  assign RetimeWrapper_163_clock = clock; // @[:@20553.4]
  assign RetimeWrapper_163_reset = reset; // @[:@20554.4]
  assign RetimeWrapper_163_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@20556.4]
  assign RetimeWrapper_163_io_in = _T_2605 & io_rPort_13_en_0; // @[package.scala 94:16:@20555.4]
  assign RetimeWrapper_164_clock = clock; // @[:@20561.4]
  assign RetimeWrapper_164_reset = reset; // @[:@20562.4]
  assign RetimeWrapper_164_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@20564.4]
  assign RetimeWrapper_164_io_in = _T_2789 & io_rPort_13_en_0; // @[package.scala 94:16:@20563.4]
  assign RetimeWrapper_165_clock = clock; // @[:@20569.4]
  assign RetimeWrapper_165_reset = reset; // @[:@20570.4]
  assign RetimeWrapper_165_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@20572.4]
  assign RetimeWrapper_165_io_in = _T_2973 & io_rPort_13_en_0; // @[package.scala 94:16:@20571.4]
  assign RetimeWrapper_166_clock = clock; // @[:@20577.4]
  assign RetimeWrapper_166_reset = reset; // @[:@20578.4]
  assign RetimeWrapper_166_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@20580.4]
  assign RetimeWrapper_166_io_in = _T_3157 & io_rPort_13_en_0; // @[package.scala 94:16:@20579.4]
  assign RetimeWrapper_167_clock = clock; // @[:@20585.4]
  assign RetimeWrapper_167_reset = reset; // @[:@20586.4]
  assign RetimeWrapper_167_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@20588.4]
  assign RetimeWrapper_167_io_in = _T_3341 & io_rPort_13_en_0; // @[package.scala 94:16:@20587.4]
  assign RetimeWrapper_168_clock = clock; // @[:@20641.4]
  assign RetimeWrapper_168_reset = reset; // @[:@20642.4]
  assign RetimeWrapper_168_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@20644.4]
  assign RetimeWrapper_168_io_in = _T_1219 & io_rPort_14_en_0; // @[package.scala 94:16:@20643.4]
  assign RetimeWrapper_169_clock = clock; // @[:@20649.4]
  assign RetimeWrapper_169_reset = reset; // @[:@20650.4]
  assign RetimeWrapper_169_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@20652.4]
  assign RetimeWrapper_169_io_in = _T_1403 & io_rPort_14_en_0; // @[package.scala 94:16:@20651.4]
  assign RetimeWrapper_170_clock = clock; // @[:@20657.4]
  assign RetimeWrapper_170_reset = reset; // @[:@20658.4]
  assign RetimeWrapper_170_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@20660.4]
  assign RetimeWrapper_170_io_in = _T_1587 & io_rPort_14_en_0; // @[package.scala 94:16:@20659.4]
  assign RetimeWrapper_171_clock = clock; // @[:@20665.4]
  assign RetimeWrapper_171_reset = reset; // @[:@20666.4]
  assign RetimeWrapper_171_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@20668.4]
  assign RetimeWrapper_171_io_in = _T_1771 & io_rPort_14_en_0; // @[package.scala 94:16:@20667.4]
  assign RetimeWrapper_172_clock = clock; // @[:@20673.4]
  assign RetimeWrapper_172_reset = reset; // @[:@20674.4]
  assign RetimeWrapper_172_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@20676.4]
  assign RetimeWrapper_172_io_in = _T_1955 & io_rPort_14_en_0; // @[package.scala 94:16:@20675.4]
  assign RetimeWrapper_173_clock = clock; // @[:@20681.4]
  assign RetimeWrapper_173_reset = reset; // @[:@20682.4]
  assign RetimeWrapper_173_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@20684.4]
  assign RetimeWrapper_173_io_in = _T_2139 & io_rPort_14_en_0; // @[package.scala 94:16:@20683.4]
  assign RetimeWrapper_174_clock = clock; // @[:@20689.4]
  assign RetimeWrapper_174_reset = reset; // @[:@20690.4]
  assign RetimeWrapper_174_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@20692.4]
  assign RetimeWrapper_174_io_in = _T_2323 & io_rPort_14_en_0; // @[package.scala 94:16:@20691.4]
  assign RetimeWrapper_175_clock = clock; // @[:@20697.4]
  assign RetimeWrapper_175_reset = reset; // @[:@20698.4]
  assign RetimeWrapper_175_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@20700.4]
  assign RetimeWrapper_175_io_in = _T_2507 & io_rPort_14_en_0; // @[package.scala 94:16:@20699.4]
  assign RetimeWrapper_176_clock = clock; // @[:@20705.4]
  assign RetimeWrapper_176_reset = reset; // @[:@20706.4]
  assign RetimeWrapper_176_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@20708.4]
  assign RetimeWrapper_176_io_in = _T_2691 & io_rPort_14_en_0; // @[package.scala 94:16:@20707.4]
  assign RetimeWrapper_177_clock = clock; // @[:@20713.4]
  assign RetimeWrapper_177_reset = reset; // @[:@20714.4]
  assign RetimeWrapper_177_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@20716.4]
  assign RetimeWrapper_177_io_in = _T_2875 & io_rPort_14_en_0; // @[package.scala 94:16:@20715.4]
  assign RetimeWrapper_178_clock = clock; // @[:@20721.4]
  assign RetimeWrapper_178_reset = reset; // @[:@20722.4]
  assign RetimeWrapper_178_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@20724.4]
  assign RetimeWrapper_178_io_in = _T_3059 & io_rPort_14_en_0; // @[package.scala 94:16:@20723.4]
  assign RetimeWrapper_179_clock = clock; // @[:@20729.4]
  assign RetimeWrapper_179_reset = reset; // @[:@20730.4]
  assign RetimeWrapper_179_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@20732.4]
  assign RetimeWrapper_179_io_in = _T_3243 & io_rPort_14_en_0; // @[package.scala 94:16:@20731.4]
  assign RetimeWrapper_180_clock = clock; // @[:@20785.4]
  assign RetimeWrapper_180_reset = reset; // @[:@20786.4]
  assign RetimeWrapper_180_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@20788.4]
  assign RetimeWrapper_180_io_in = _T_1225 & io_rPort_15_en_0; // @[package.scala 94:16:@20787.4]
  assign RetimeWrapper_181_clock = clock; // @[:@20793.4]
  assign RetimeWrapper_181_reset = reset; // @[:@20794.4]
  assign RetimeWrapper_181_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@20796.4]
  assign RetimeWrapper_181_io_in = _T_1409 & io_rPort_15_en_0; // @[package.scala 94:16:@20795.4]
  assign RetimeWrapper_182_clock = clock; // @[:@20801.4]
  assign RetimeWrapper_182_reset = reset; // @[:@20802.4]
  assign RetimeWrapper_182_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@20804.4]
  assign RetimeWrapper_182_io_in = _T_1593 & io_rPort_15_en_0; // @[package.scala 94:16:@20803.4]
  assign RetimeWrapper_183_clock = clock; // @[:@20809.4]
  assign RetimeWrapper_183_reset = reset; // @[:@20810.4]
  assign RetimeWrapper_183_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@20812.4]
  assign RetimeWrapper_183_io_in = _T_1777 & io_rPort_15_en_0; // @[package.scala 94:16:@20811.4]
  assign RetimeWrapper_184_clock = clock; // @[:@20817.4]
  assign RetimeWrapper_184_reset = reset; // @[:@20818.4]
  assign RetimeWrapper_184_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@20820.4]
  assign RetimeWrapper_184_io_in = _T_1961 & io_rPort_15_en_0; // @[package.scala 94:16:@20819.4]
  assign RetimeWrapper_185_clock = clock; // @[:@20825.4]
  assign RetimeWrapper_185_reset = reset; // @[:@20826.4]
  assign RetimeWrapper_185_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@20828.4]
  assign RetimeWrapper_185_io_in = _T_2145 & io_rPort_15_en_0; // @[package.scala 94:16:@20827.4]
  assign RetimeWrapper_186_clock = clock; // @[:@20833.4]
  assign RetimeWrapper_186_reset = reset; // @[:@20834.4]
  assign RetimeWrapper_186_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@20836.4]
  assign RetimeWrapper_186_io_in = _T_2329 & io_rPort_15_en_0; // @[package.scala 94:16:@20835.4]
  assign RetimeWrapper_187_clock = clock; // @[:@20841.4]
  assign RetimeWrapper_187_reset = reset; // @[:@20842.4]
  assign RetimeWrapper_187_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@20844.4]
  assign RetimeWrapper_187_io_in = _T_2513 & io_rPort_15_en_0; // @[package.scala 94:16:@20843.4]
  assign RetimeWrapper_188_clock = clock; // @[:@20849.4]
  assign RetimeWrapper_188_reset = reset; // @[:@20850.4]
  assign RetimeWrapper_188_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@20852.4]
  assign RetimeWrapper_188_io_in = _T_2697 & io_rPort_15_en_0; // @[package.scala 94:16:@20851.4]
  assign RetimeWrapper_189_clock = clock; // @[:@20857.4]
  assign RetimeWrapper_189_reset = reset; // @[:@20858.4]
  assign RetimeWrapper_189_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@20860.4]
  assign RetimeWrapper_189_io_in = _T_2881 & io_rPort_15_en_0; // @[package.scala 94:16:@20859.4]
  assign RetimeWrapper_190_clock = clock; // @[:@20865.4]
  assign RetimeWrapper_190_reset = reset; // @[:@20866.4]
  assign RetimeWrapper_190_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@20868.4]
  assign RetimeWrapper_190_io_in = _T_3065 & io_rPort_15_en_0; // @[package.scala 94:16:@20867.4]
  assign RetimeWrapper_191_clock = clock; // @[:@20873.4]
  assign RetimeWrapper_191_reset = reset; // @[:@20874.4]
  assign RetimeWrapper_191_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@20876.4]
  assign RetimeWrapper_191_io_in = _T_3249 & io_rPort_15_en_0; // @[package.scala 94:16:@20875.4]
  assign RetimeWrapper_192_clock = clock; // @[:@20929.4]
  assign RetimeWrapper_192_reset = reset; // @[:@20930.4]
  assign RetimeWrapper_192_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@20932.4]
  assign RetimeWrapper_192_io_in = _T_1323 & io_rPort_16_en_0; // @[package.scala 94:16:@20931.4]
  assign RetimeWrapper_193_clock = clock; // @[:@20937.4]
  assign RetimeWrapper_193_reset = reset; // @[:@20938.4]
  assign RetimeWrapper_193_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@20940.4]
  assign RetimeWrapper_193_io_in = _T_1507 & io_rPort_16_en_0; // @[package.scala 94:16:@20939.4]
  assign RetimeWrapper_194_clock = clock; // @[:@20945.4]
  assign RetimeWrapper_194_reset = reset; // @[:@20946.4]
  assign RetimeWrapper_194_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@20948.4]
  assign RetimeWrapper_194_io_in = _T_1691 & io_rPort_16_en_0; // @[package.scala 94:16:@20947.4]
  assign RetimeWrapper_195_clock = clock; // @[:@20953.4]
  assign RetimeWrapper_195_reset = reset; // @[:@20954.4]
  assign RetimeWrapper_195_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@20956.4]
  assign RetimeWrapper_195_io_in = _T_1875 & io_rPort_16_en_0; // @[package.scala 94:16:@20955.4]
  assign RetimeWrapper_196_clock = clock; // @[:@20961.4]
  assign RetimeWrapper_196_reset = reset; // @[:@20962.4]
  assign RetimeWrapper_196_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@20964.4]
  assign RetimeWrapper_196_io_in = _T_2059 & io_rPort_16_en_0; // @[package.scala 94:16:@20963.4]
  assign RetimeWrapper_197_clock = clock; // @[:@20969.4]
  assign RetimeWrapper_197_reset = reset; // @[:@20970.4]
  assign RetimeWrapper_197_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@20972.4]
  assign RetimeWrapper_197_io_in = _T_2243 & io_rPort_16_en_0; // @[package.scala 94:16:@20971.4]
  assign RetimeWrapper_198_clock = clock; // @[:@20977.4]
  assign RetimeWrapper_198_reset = reset; // @[:@20978.4]
  assign RetimeWrapper_198_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@20980.4]
  assign RetimeWrapper_198_io_in = _T_2427 & io_rPort_16_en_0; // @[package.scala 94:16:@20979.4]
  assign RetimeWrapper_199_clock = clock; // @[:@20985.4]
  assign RetimeWrapper_199_reset = reset; // @[:@20986.4]
  assign RetimeWrapper_199_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@20988.4]
  assign RetimeWrapper_199_io_in = _T_2611 & io_rPort_16_en_0; // @[package.scala 94:16:@20987.4]
  assign RetimeWrapper_200_clock = clock; // @[:@20993.4]
  assign RetimeWrapper_200_reset = reset; // @[:@20994.4]
  assign RetimeWrapper_200_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@20996.4]
  assign RetimeWrapper_200_io_in = _T_2795 & io_rPort_16_en_0; // @[package.scala 94:16:@20995.4]
  assign RetimeWrapper_201_clock = clock; // @[:@21001.4]
  assign RetimeWrapper_201_reset = reset; // @[:@21002.4]
  assign RetimeWrapper_201_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@21004.4]
  assign RetimeWrapper_201_io_in = _T_2979 & io_rPort_16_en_0; // @[package.scala 94:16:@21003.4]
  assign RetimeWrapper_202_clock = clock; // @[:@21009.4]
  assign RetimeWrapper_202_reset = reset; // @[:@21010.4]
  assign RetimeWrapper_202_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@21012.4]
  assign RetimeWrapper_202_io_in = _T_3163 & io_rPort_16_en_0; // @[package.scala 94:16:@21011.4]
  assign RetimeWrapper_203_clock = clock; // @[:@21017.4]
  assign RetimeWrapper_203_reset = reset; // @[:@21018.4]
  assign RetimeWrapper_203_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@21020.4]
  assign RetimeWrapper_203_io_in = _T_3347 & io_rPort_16_en_0; // @[package.scala 94:16:@21019.4]
  assign RetimeWrapper_204_clock = clock; // @[:@21073.4]
  assign RetimeWrapper_204_reset = reset; // @[:@21074.4]
  assign RetimeWrapper_204_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@21076.4]
  assign RetimeWrapper_204_io_in = _T_1231 & io_rPort_17_en_0; // @[package.scala 94:16:@21075.4]
  assign RetimeWrapper_205_clock = clock; // @[:@21081.4]
  assign RetimeWrapper_205_reset = reset; // @[:@21082.4]
  assign RetimeWrapper_205_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@21084.4]
  assign RetimeWrapper_205_io_in = _T_1415 & io_rPort_17_en_0; // @[package.scala 94:16:@21083.4]
  assign RetimeWrapper_206_clock = clock; // @[:@21089.4]
  assign RetimeWrapper_206_reset = reset; // @[:@21090.4]
  assign RetimeWrapper_206_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@21092.4]
  assign RetimeWrapper_206_io_in = _T_1599 & io_rPort_17_en_0; // @[package.scala 94:16:@21091.4]
  assign RetimeWrapper_207_clock = clock; // @[:@21097.4]
  assign RetimeWrapper_207_reset = reset; // @[:@21098.4]
  assign RetimeWrapper_207_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@21100.4]
  assign RetimeWrapper_207_io_in = _T_1783 & io_rPort_17_en_0; // @[package.scala 94:16:@21099.4]
  assign RetimeWrapper_208_clock = clock; // @[:@21105.4]
  assign RetimeWrapper_208_reset = reset; // @[:@21106.4]
  assign RetimeWrapper_208_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@21108.4]
  assign RetimeWrapper_208_io_in = _T_1967 & io_rPort_17_en_0; // @[package.scala 94:16:@21107.4]
  assign RetimeWrapper_209_clock = clock; // @[:@21113.4]
  assign RetimeWrapper_209_reset = reset; // @[:@21114.4]
  assign RetimeWrapper_209_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@21116.4]
  assign RetimeWrapper_209_io_in = _T_2151 & io_rPort_17_en_0; // @[package.scala 94:16:@21115.4]
  assign RetimeWrapper_210_clock = clock; // @[:@21121.4]
  assign RetimeWrapper_210_reset = reset; // @[:@21122.4]
  assign RetimeWrapper_210_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@21124.4]
  assign RetimeWrapper_210_io_in = _T_2335 & io_rPort_17_en_0; // @[package.scala 94:16:@21123.4]
  assign RetimeWrapper_211_clock = clock; // @[:@21129.4]
  assign RetimeWrapper_211_reset = reset; // @[:@21130.4]
  assign RetimeWrapper_211_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@21132.4]
  assign RetimeWrapper_211_io_in = _T_2519 & io_rPort_17_en_0; // @[package.scala 94:16:@21131.4]
  assign RetimeWrapper_212_clock = clock; // @[:@21137.4]
  assign RetimeWrapper_212_reset = reset; // @[:@21138.4]
  assign RetimeWrapper_212_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@21140.4]
  assign RetimeWrapper_212_io_in = _T_2703 & io_rPort_17_en_0; // @[package.scala 94:16:@21139.4]
  assign RetimeWrapper_213_clock = clock; // @[:@21145.4]
  assign RetimeWrapper_213_reset = reset; // @[:@21146.4]
  assign RetimeWrapper_213_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@21148.4]
  assign RetimeWrapper_213_io_in = _T_2887 & io_rPort_17_en_0; // @[package.scala 94:16:@21147.4]
  assign RetimeWrapper_214_clock = clock; // @[:@21153.4]
  assign RetimeWrapper_214_reset = reset; // @[:@21154.4]
  assign RetimeWrapper_214_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@21156.4]
  assign RetimeWrapper_214_io_in = _T_3071 & io_rPort_17_en_0; // @[package.scala 94:16:@21155.4]
  assign RetimeWrapper_215_clock = clock; // @[:@21161.4]
  assign RetimeWrapper_215_reset = reset; // @[:@21162.4]
  assign RetimeWrapper_215_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@21164.4]
  assign RetimeWrapper_215_io_in = _T_3255 & io_rPort_17_en_0; // @[package.scala 94:16:@21163.4]
endmodule
module RetimeWrapper_260( // @[:@21192.2]
  input         clock, // @[:@21193.4]
  input         reset, // @[:@21194.4]
  input         io_flow, // @[:@21195.4]
  input  [31:0] io_in, // @[:@21195.4]
  output [31:0] io_out // @[:@21195.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@21197.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@21197.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@21197.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@21197.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@21197.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@21197.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@21197.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@21210.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@21209.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@21208.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@21207.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@21206.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@21204.4]
endmodule
module RetimeWrapper_261( // @[:@21224.2]
  input         clock, // @[:@21225.4]
  input         reset, // @[:@21226.4]
  input         io_flow, // @[:@21227.4]
  input  [31:0] io_in, // @[:@21227.4]
  output [31:0] io_out // @[:@21227.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@21229.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@21229.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@21229.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@21229.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@21229.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@21229.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(16)) sr ( // @[RetimeShiftRegister.scala 15:20:@21229.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@21242.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@21241.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@21240.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@21239.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@21238.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@21236.4]
endmodule
module fix2fixBox( // @[:@21244.2]
  input  [63:0] io_a, // @[:@21247.4]
  output [31:0] io_b // @[:@21247.4]
);
  assign io_b = io_a[31:0]; // @[Converter.scala 95:38:@21260.4]
endmodule
module x340( // @[:@21262.2]
  input         clock, // @[:@21263.4]
  input         reset, // @[:@21264.4]
  input  [31:0] io_a, // @[:@21265.4]
  input  [31:0] io_b, // @[:@21265.4]
  input         io_flow, // @[:@21265.4]
  output [31:0] io_result // @[:@21265.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@21274.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@21274.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@21274.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@21274.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@21274.4]
  wire [63:0] fix2fixBox_io_a; // @[Math.scala 357:30:@21282.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 357:30:@21282.4]
  wire [31:0] _T_19; // @[package.scala 96:25:@21279.4 package.scala 96:25:@21280.4]
  wire [31:0] _GEN_0; // @[package.scala 94:16:@21277.4]
  RetimeWrapper_261 RetimeWrapper ( // @[package.scala 93:22:@21274.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  fix2fixBox fix2fixBox ( // @[Math.scala 357:30:@21282.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign _T_19 = RetimeWrapper_io_out; // @[package.scala 96:25:@21279.4 package.scala 96:25:@21280.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 363:17:@21290.4]
  assign RetimeWrapper_clock = clock; // @[:@21275.4]
  assign RetimeWrapper_reset = reset; // @[:@21276.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@21278.4]
  assign _GEN_0 = io_a % io_b; // @[package.scala 94:16:@21277.4]
  assign RetimeWrapper_io_in = _GEN_0[31:0]; // @[package.scala 94:16:@21277.4]
  assign fix2fixBox_io_a = {{32'd0}, _T_19}; // @[Math.scala 358:23:@21285.4]
endmodule
module RetimeWrapper_262( // @[:@21304.2]
  input         clock, // @[:@21305.4]
  input         reset, // @[:@21306.4]
  input         io_flow, // @[:@21307.4]
  input  [63:0] io_in, // @[:@21307.4]
  output [63:0] io_out // @[:@21307.4]
);
  wire [63:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@21309.4]
  wire [63:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@21309.4]
  wire [63:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@21309.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@21309.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@21309.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@21309.4]
  RetimeShiftRegister #(.WIDTH(64), .STAGES(6)) sr ( // @[RetimeShiftRegister.scala 15:20:@21309.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@21322.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@21321.4]
  assign sr_init = 64'h0; // @[RetimeShiftRegister.scala 19:16:@21320.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@21319.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@21318.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@21316.4]
endmodule
module RetimeWrapper_263( // @[:@21336.2]
  input   clock, // @[:@21337.4]
  input   reset, // @[:@21338.4]
  input   io_flow, // @[:@21339.4]
  input   io_in // @[:@21339.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@21341.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@21341.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@21341.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@21341.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@21341.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@21341.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(6)) sr ( // @[RetimeShiftRegister.scala 15:20:@21341.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@21353.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@21352.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@21351.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@21350.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@21348.4]
endmodule
module x342_mul( // @[:@21406.2]
  input         clock, // @[:@21407.4]
  input         reset, // @[:@21408.4]
  input  [31:0] io_a, // @[:@21409.4]
  input         io_flow, // @[:@21409.4]
  output [31:0] io_result // @[:@21409.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@21417.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@21417.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@21417.4]
  wire [63:0] RetimeWrapper_io_in; // @[package.scala 93:22:@21417.4]
  wire [63:0] RetimeWrapper_io_out; // @[package.scala 93:22:@21417.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@21430.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@21430.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@21430.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@21430.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@21441.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@21441.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@21441.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@21441.4]
  wire [31:0] fix2fixBox_io_a; // @[Math.scala 253:30:@21448.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 253:30:@21448.4]
  wire [63:0] _T_18; // @[package.scala 96:25:@21422.4 package.scala 96:25:@21423.4]
  wire  _T_21; // @[FixedPoint.scala 50:25:@21427.4]
  RetimeWrapper_262 RetimeWrapper ( // @[package.scala 93:22:@21417.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_263 RetimeWrapper_1 ( // @[package.scala 93:22:@21430.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in)
  );
  RetimeWrapper_263 RetimeWrapper_2 ( // @[package.scala 93:22:@21441.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in)
  );
  SimBlackBoxesfix2fixBox fix2fixBox ( // @[Math.scala 253:30:@21448.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@21422.4 package.scala 96:25:@21423.4]
  assign _T_21 = io_a[31]; // @[FixedPoint.scala 50:25:@21427.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 259:17:@21456.4]
  assign RetimeWrapper_clock = clock; // @[:@21418.4]
  assign RetimeWrapper_reset = reset; // @[:@21419.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@21421.4]
  assign RetimeWrapper_io_in = io_a * 32'hab; // @[package.scala 94:16:@21420.4]
  assign RetimeWrapper_1_clock = clock; // @[:@21431.4]
  assign RetimeWrapper_1_reset = reset; // @[:@21432.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@21434.4]
  assign RetimeWrapper_1_io_in = io_a[31]; // @[package.scala 94:16:@21433.4]
  assign RetimeWrapper_2_clock = clock; // @[:@21442.4]
  assign RetimeWrapper_2_reset = reset; // @[:@21443.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@21445.4]
  assign RetimeWrapper_2_io_in = _T_21 == 1'h0; // @[package.scala 94:16:@21444.4]
  assign fix2fixBox_io_a = _T_18[31:0]; // @[Math.scala 254:23:@21451.4]
endmodule
module RetimeWrapper_265( // @[:@21470.2]
  input         clock, // @[:@21471.4]
  input         reset, // @[:@21472.4]
  input         io_flow, // @[:@21473.4]
  input  [31:0] io_in, // @[:@21473.4]
  output [31:0] io_out // @[:@21473.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@21475.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@21475.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@21475.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@21475.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@21475.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@21475.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(20)) sr ( // @[RetimeShiftRegister.scala 15:20:@21475.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@21488.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@21487.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@21486.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@21485.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@21484.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@21482.4]
endmodule
module x343_div( // @[:@21531.2]
  input         clock, // @[:@21532.4]
  input         reset, // @[:@21533.4]
  input  [31:0] io_a, // @[:@21534.4]
  input         io_flow, // @[:@21534.4]
  output [31:0] io_result // @[:@21534.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@21543.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@21543.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@21543.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@21543.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@21543.4]
  wire [31:0] __io_b; // @[Math.scala 709:24:@21556.4]
  wire [31:0] __io_result; // @[Math.scala 709:24:@21556.4]
  wire [31:0] _T_15; // @[FixedPoint.scala 24:59:@21540.4]
  wire [32:0] _T_17; // @[BigIPSim.scala 23:39:@21542.4]
  wire [32:0] _T_18; // @[package.scala 94:23:@21546.4]
  wire [31:0] _T_21; // @[package.scala 96:25:@21550.4]
  RetimeWrapper_265 RetimeWrapper ( // @[package.scala 93:22:@21543.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  _ _ ( // @[Math.scala 709:24:@21556.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  assign _T_15 = $signed(io_a); // @[FixedPoint.scala 24:59:@21540.4]
  assign _T_17 = $signed(_T_15) / $signed(32'sh6); // @[BigIPSim.scala 23:39:@21542.4]
  assign _T_18 = $unsigned(_T_17); // @[package.scala 94:23:@21546.4]
  assign _T_21 = $signed(RetimeWrapper_io_out); // @[package.scala 96:25:@21550.4]
  assign io_result = __io_result; // @[Math.scala 290:34:@21564.4]
  assign RetimeWrapper_clock = clock; // @[:@21544.4]
  assign RetimeWrapper_reset = reset; // @[:@21545.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@21548.4]
  assign RetimeWrapper_io_in = _T_18[31:0]; // @[package.scala 94:16:@21547.4]
  assign __io_b = $unsigned(_T_21); // @[Math.scala 710:17:@21559.4]
endmodule
module RetimeWrapper_266( // @[:@21578.2]
  input         clock, // @[:@21579.4]
  input         reset, // @[:@21580.4]
  input         io_flow, // @[:@21581.4]
  input  [31:0] io_in, // @[:@21581.4]
  output [31:0] io_out // @[:@21581.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@21583.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@21583.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@21583.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@21583.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@21583.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@21583.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(14)) sr ( // @[RetimeShiftRegister.scala 15:20:@21583.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@21596.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@21595.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@21594.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@21593.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@21592.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@21590.4]
endmodule
module SimBlackBoxesfix2fixBox_3( // @[:@21598.2]
  input  [31:0] io_a, // @[:@21601.4]
  output [32:0] io_b // @[:@21601.4]
);
  wire  _T_20; // @[implicits.scala 69:16:@21611.4]
  assign _T_20 = io_a[31]; // @[implicits.scala 69:16:@21611.4]
  assign io_b = {_T_20,io_a}; // @[SimBlackBoxes.scala 99:40:@21616.4]
endmodule
module __3( // @[:@21618.2]
  input  [31:0] io_b, // @[:@21621.4]
  output [32:0] io_result // @[:@21621.4]
);
  wire [31:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@21626.4]
  wire [32:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@21626.4]
  SimBlackBoxesfix2fixBox_3 SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@21626.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@21639.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@21634.4]
endmodule
module fix2fixBox_2( // @[:@21716.2]
  input         clock, // @[:@21717.4]
  input         reset, // @[:@21718.4]
  input  [32:0] io_a, // @[:@21719.4]
  input         io_flow, // @[:@21719.4]
  output [31:0] io_b // @[:@21719.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@21732.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@21732.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@21732.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@21732.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@21732.4]
  RetimeWrapper_260 RetimeWrapper ( // @[package.scala 93:22:@21732.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@21739.4]
  assign RetimeWrapper_clock = clock; // @[:@21733.4]
  assign RetimeWrapper_reset = reset; // @[:@21734.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@21736.4]
  assign RetimeWrapper_io_in = io_a[31:0]; // @[package.scala 94:16:@21735.4]
endmodule
module x344_sum( // @[:@21741.2]
  input         clock, // @[:@21742.4]
  input         reset, // @[:@21743.4]
  input  [31:0] io_a, // @[:@21744.4]
  input  [31:0] io_b, // @[:@21744.4]
  input         io_flow, // @[:@21744.4]
  output [31:0] io_result // @[:@21744.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@21752.4]
  wire [32:0] __io_result; // @[Math.scala 709:24:@21752.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@21759.4]
  wire [32:0] __1_io_result; // @[Math.scala 709:24:@21759.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@21777.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@21777.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@21777.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@21777.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@21777.4]
  wire [32:0] a_upcast_number; // @[Math.scala 712:22:@21757.4 Math.scala 713:14:@21758.4]
  wire [32:0] b_upcast_number; // @[Math.scala 712:22:@21764.4 Math.scala 713:14:@21765.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@21766.4]
  __3 _ ( // @[Math.scala 709:24:@21752.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __3 __1 ( // @[Math.scala 709:24:@21759.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_2 fix2fixBox ( // @[Math.scala 141:30:@21777.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@21757.4 Math.scala 713:14:@21758.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@21764.4 Math.scala 713:14:@21765.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@21766.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@21785.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@21755.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@21762.4]
  assign fix2fixBox_clock = clock; // @[:@21778.4]
  assign fix2fixBox_reset = reset; // @[:@21779.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@21780.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@21783.4]
endmodule
module RetimeWrapper_268( // @[:@21799.2]
  input         clock, // @[:@21800.4]
  input         reset, // @[:@21801.4]
  input         io_flow, // @[:@21802.4]
  input  [31:0] io_in, // @[:@21802.4]
  output [31:0] io_out // @[:@21802.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@21804.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@21804.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@21804.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@21804.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@21804.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@21804.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(8)) sr ( // @[RetimeShiftRegister.scala 15:20:@21804.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@21817.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@21816.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@21815.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@21814.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@21813.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@21811.4]
endmodule
module RetimeWrapper_269( // @[:@21831.2]
  input         clock, // @[:@21832.4]
  input         reset, // @[:@21833.4]
  input         io_flow, // @[:@21834.4]
  input  [31:0] io_in, // @[:@21834.4]
  output [31:0] io_out // @[:@21834.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@21836.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@21836.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@21836.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@21836.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@21836.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@21836.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@21836.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@21849.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@21848.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@21847.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@21846.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@21845.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@21843.4]
endmodule
module RetimeWrapper_270( // @[:@21863.2]
  input         clock, // @[:@21864.4]
  input         reset, // @[:@21865.4]
  input         io_flow, // @[:@21866.4]
  input  [31:0] io_in, // @[:@21866.4]
  output [31:0] io_out // @[:@21866.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@21868.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@21868.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@21868.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@21868.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@21868.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@21868.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(24)) sr ( // @[RetimeShiftRegister.scala 15:20:@21868.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@21881.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@21880.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@21879.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@21878.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@21877.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@21875.4]
endmodule
module RetimeWrapper_271( // @[:@21895.2]
  input   clock, // @[:@21896.4]
  input   reset, // @[:@21897.4]
  input   io_flow, // @[:@21898.4]
  input   io_in, // @[:@21898.4]
  output  io_out // @[:@21898.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@21900.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@21900.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@21900.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@21900.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@21900.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@21900.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(24)) sr ( // @[RetimeShiftRegister.scala 15:20:@21900.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@21913.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@21912.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@21911.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@21910.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@21909.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@21907.4]
endmodule
module RetimeWrapper_273( // @[:@21959.2]
  input        clock, // @[:@21960.4]
  input        reset, // @[:@21961.4]
  input        io_flow, // @[:@21962.4]
  input  [7:0] io_in, // @[:@21962.4]
  output [7:0] io_out // @[:@21962.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@21964.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@21964.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@21964.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@21964.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@21964.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@21964.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(23)) sr ( // @[RetimeShiftRegister.scala 15:20:@21964.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@21977.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@21976.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@21975.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@21974.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@21973.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@21971.4]
endmodule
module RetimeWrapper_278( // @[:@22400.2]
  input         clock, // @[:@22401.4]
  input         reset, // @[:@22402.4]
  input         io_flow, // @[:@22403.4]
  input  [31:0] io_in, // @[:@22403.4]
  output [31:0] io_out // @[:@22403.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@22405.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@22405.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@22405.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@22405.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@22405.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@22405.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(15)) sr ( // @[RetimeShiftRegister.scala 15:20:@22405.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@22418.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@22417.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@22416.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@22415.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@22414.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@22412.4]
endmodule
module RetimeWrapper_281( // @[:@22653.2]
  input         clock, // @[:@22654.4]
  input         reset, // @[:@22655.4]
  input         io_flow, // @[:@22656.4]
  input  [31:0] io_in, // @[:@22656.4]
  output [31:0] io_out // @[:@22656.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@22658.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@22658.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@22658.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@22658.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@22658.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@22658.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(7)) sr ( // @[RetimeShiftRegister.scala 15:20:@22658.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@22671.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@22670.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@22669.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@22668.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@22667.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@22665.4]
endmodule
module RetimeWrapper_282( // @[:@22685.2]
  input         clock, // @[:@22686.4]
  input         reset, // @[:@22687.4]
  input         io_flow, // @[:@22688.4]
  input  [31:0] io_in, // @[:@22688.4]
  output [31:0] io_out // @[:@22688.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@22690.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@22690.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@22690.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@22690.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@22690.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@22690.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@22690.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@22703.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@22702.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@22701.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@22700.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@22699.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@22697.4]
endmodule
module RetimeWrapper_300( // @[:@24137.2]
  input         clock, // @[:@24138.4]
  input         reset, // @[:@24139.4]
  input         io_flow, // @[:@24140.4]
  input  [31:0] io_in, // @[:@24140.4]
  output [31:0] io_out // @[:@24140.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@24142.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@24142.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@24142.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@24142.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@24142.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@24142.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(26)) sr ( // @[RetimeShiftRegister.scala 15:20:@24142.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@24155.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@24154.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@24153.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@24152.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@24151.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@24149.4]
endmodule
module RetimeWrapper_309( // @[:@24543.2]
  input         clock, // @[:@24544.4]
  input         reset, // @[:@24545.4]
  input         io_flow, // @[:@24546.4]
  input  [31:0] io_in, // @[:@24546.4]
  output [31:0] io_out // @[:@24546.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@24548.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@24548.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@24548.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@24548.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@24548.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@24548.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(27)) sr ( // @[RetimeShiftRegister.scala 15:20:@24548.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@24561.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@24560.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@24559.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@24558.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@24557.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@24555.4]
endmodule
module RetimeWrapper_311( // @[:@24764.2]
  input   clock, // @[:@24765.4]
  input   reset, // @[:@24766.4]
  input   io_flow, // @[:@24767.4]
  input   io_in, // @[:@24767.4]
  output  io_out // @[:@24767.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@24769.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@24769.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@24769.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@24769.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@24769.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@24769.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(50)) sr ( // @[RetimeShiftRegister.scala 15:20:@24769.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@24782.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@24781.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@24780.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@24779.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@24778.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@24776.4]
endmodule
module RetimeWrapper_312( // @[:@24796.2]
  input         clock, // @[:@24797.4]
  input         reset, // @[:@24798.4]
  input         io_flow, // @[:@24799.4]
  input  [31:0] io_in, // @[:@24799.4]
  output [31:0] io_out // @[:@24799.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@24801.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@24801.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@24801.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@24801.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@24801.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@24801.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(33)) sr ( // @[RetimeShiftRegister.scala 15:20:@24801.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@24814.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@24813.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@24812.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@24811.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@24810.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@24808.4]
endmodule
module RetimeWrapper_316( // @[:@24924.2]
  input   clock, // @[:@24925.4]
  input   reset, // @[:@24926.4]
  input   io_flow, // @[:@24927.4]
  input   io_in, // @[:@24927.4]
  output  io_out // @[:@24927.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@24929.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@24929.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@24929.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@24929.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@24929.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@24929.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(22)) sr ( // @[RetimeShiftRegister.scala 15:20:@24929.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@24942.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@24941.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@24940.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@24939.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@24938.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@24936.4]
endmodule
module RetimeWrapper_336( // @[:@25878.2]
  input         clock, // @[:@25879.4]
  input         reset, // @[:@25880.4]
  input         io_flow, // @[:@25881.4]
  input  [31:0] io_in, // @[:@25881.4]
  output [31:0] io_out // @[:@25881.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@25883.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@25883.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@25883.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@25883.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@25883.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@25883.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(28)) sr ( // @[RetimeShiftRegister.scala 15:20:@25883.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@25896.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@25895.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@25894.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@25893.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@25892.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@25890.4]
endmodule
module RetimeWrapper_338( // @[:@26099.2]
  input         clock, // @[:@26100.4]
  input         reset, // @[:@26101.4]
  input         io_flow, // @[:@26102.4]
  input  [31:0] io_in, // @[:@26102.4]
  output [31:0] io_out // @[:@26102.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@26104.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@26104.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@26104.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@26104.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@26104.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@26104.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(34)) sr ( // @[RetimeShiftRegister.scala 15:20:@26104.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@26117.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@26116.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@26115.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@26114.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@26113.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@26111.4]
endmodule
module RetimeWrapper_340( // @[:@26163.2]
  input   clock, // @[:@26164.4]
  input   reset, // @[:@26165.4]
  input   io_flow, // @[:@26166.4]
  input   io_in, // @[:@26166.4]
  output  io_out // @[:@26166.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@26168.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@26168.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@26168.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@26168.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@26168.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@26168.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(23)) sr ( // @[RetimeShiftRegister.scala 15:20:@26168.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@26181.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@26180.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@26179.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@26178.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@26177.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@26175.4]
endmodule
module x412_rdrow( // @[:@27874.2]
  input         clock, // @[:@27875.4]
  input         reset, // @[:@27876.4]
  input  [31:0] io_a, // @[:@27877.4]
  input  [31:0] io_b, // @[:@27877.4]
  input         io_flow, // @[:@27877.4]
  output [31:0] io_result // @[:@27877.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@27885.4]
  wire [32:0] __io_result; // @[Math.scala 709:24:@27885.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@27892.4]
  wire [32:0] __1_io_result; // @[Math.scala 709:24:@27892.4]
  wire  fix2fixBox_clock; // @[Math.scala 182:30:@27911.4]
  wire  fix2fixBox_reset; // @[Math.scala 182:30:@27911.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 182:30:@27911.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 182:30:@27911.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 182:30:@27911.4]
  wire [32:0] a_upcast_number; // @[Math.scala 712:22:@27890.4 Math.scala 713:14:@27891.4]
  wire [32:0] b_upcast_number; // @[Math.scala 712:22:@27897.4 Math.scala 713:14:@27898.4]
  wire [33:0] _T_21; // @[Math.scala 177:37:@27899.4]
  wire [33:0] _T_22; // @[Math.scala 177:37:@27900.4]
  __3 _ ( // @[Math.scala 709:24:@27885.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __3 __1 ( // @[Math.scala 709:24:@27892.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_2 fix2fixBox ( // @[Math.scala 182:30:@27911.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@27890.4 Math.scala 713:14:@27891.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@27897.4 Math.scala 713:14:@27898.4]
  assign _T_21 = a_upcast_number - b_upcast_number; // @[Math.scala 177:37:@27899.4]
  assign _T_22 = $unsigned(_T_21); // @[Math.scala 177:37:@27900.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 188:17:@27919.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@27888.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@27895.4]
  assign fix2fixBox_clock = clock; // @[:@27912.4]
  assign fix2fixBox_reset = reset; // @[:@27913.4]
  assign fix2fixBox_io_a = _T_22[32:0]; // @[Math.scala 183:23:@27914.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 186:26:@27917.4]
endmodule
module RetimeWrapper_382( // @[:@29130.2]
  input         clock, // @[:@29131.4]
  input         reset, // @[:@29132.4]
  input         io_flow, // @[:@29133.4]
  input  [31:0] io_in, // @[:@29133.4]
  output [31:0] io_out // @[:@29133.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@29135.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@29135.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@29135.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@29135.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@29135.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@29135.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(29)) sr ( // @[RetimeShiftRegister.scala 15:20:@29135.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@29148.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@29147.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@29146.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@29145.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@29144.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@29142.4]
endmodule
module RetimeWrapper_419( // @[:@32003.2]
  input        clock, // @[:@32004.4]
  input        reset, // @[:@32005.4]
  input        io_flow, // @[:@32006.4]
  input  [8:0] io_in, // @[:@32006.4]
  output [8:0] io_out // @[:@32006.4]
);
  wire [8:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@32008.4]
  wire [8:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@32008.4]
  wire [8:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@32008.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@32008.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@32008.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@32008.4]
  RetimeShiftRegister #(.WIDTH(9), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@32008.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@32021.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@32020.4]
  assign sr_init = 9'h0; // @[RetimeShiftRegister.scala 19:16:@32019.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@32018.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@32017.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@32015.4]
endmodule
module RetimeWrapper_421( // @[:@32067.2]
  input        clock, // @[:@32068.4]
  input        reset, // @[:@32069.4]
  input        io_flow, // @[:@32070.4]
  input  [9:0] io_in, // @[:@32070.4]
  output [9:0] io_out // @[:@32070.4]
);
  wire [9:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@32072.4]
  wire [9:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@32072.4]
  wire [9:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@32072.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@32072.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@32072.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@32072.4]
  RetimeShiftRegister #(.WIDTH(10), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@32072.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@32085.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@32084.4]
  assign sr_init = 10'h0; // @[RetimeShiftRegister.scala 19:16:@32083.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@32082.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@32081.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@32079.4]
endmodule
module RetimeWrapper_424( // @[:@32163.2]
  input        clock, // @[:@32164.4]
  input        reset, // @[:@32165.4]
  input        io_flow, // @[:@32166.4]
  input  [7:0] io_in, // @[:@32166.4]
  output [7:0] io_out // @[:@32166.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@32168.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@32168.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@32168.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@32168.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@32168.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@32168.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@32168.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@32181.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@32180.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@32179.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@32178.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@32177.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@32175.4]
endmodule
module SimBlackBoxesfix2fixBox_66( // @[:@32215.2]
  input  [7:0] io_a, // @[:@32218.4]
  output [8:0] io_b // @[:@32218.4]
);
  assign io_b = {1'h0,io_a}; // @[SimBlackBoxes.scala 99:40:@32232.4]
endmodule
module __66( // @[:@32234.2]
  input  [7:0] io_b, // @[:@32237.4]
  output [8:0] io_result // @[:@32237.4]
);
  wire [7:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@32242.4]
  wire [8:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@32242.4]
  SimBlackBoxesfix2fixBox_66 SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@32242.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@32255.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@32250.4]
endmodule
module fix2fixBox_42( // @[:@32299.2]
  input  [8:0] io_a, // @[:@32302.4]
  output [7:0] io_b // @[:@32302.4]
);
  assign io_b = io_a[7:0]; // @[Converter.scala 95:38:@32315.4]
endmodule
module x489_x11( // @[:@32317.2]
  input  [7:0] io_a, // @[:@32320.4]
  input  [7:0] io_b, // @[:@32320.4]
  output [7:0] io_result // @[:@32320.4]
);
  wire [7:0] __io_b; // @[Math.scala 709:24:@32328.4]
  wire [8:0] __io_result; // @[Math.scala 709:24:@32328.4]
  wire [7:0] __1_io_b; // @[Math.scala 709:24:@32335.4]
  wire [8:0] __1_io_result; // @[Math.scala 709:24:@32335.4]
  wire [8:0] fix2fixBox_io_a; // @[Math.scala 141:30:@32345.4]
  wire [7:0] fix2fixBox_io_b; // @[Math.scala 141:30:@32345.4]
  wire [8:0] a_upcast_number; // @[Math.scala 712:22:@32333.4 Math.scala 713:14:@32334.4]
  wire [8:0] b_upcast_number; // @[Math.scala 712:22:@32340.4 Math.scala 713:14:@32341.4]
  wire [9:0] _T_21; // @[Math.scala 136:37:@32342.4]
  __66 _ ( // @[Math.scala 709:24:@32328.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __66 __1 ( // @[Math.scala 709:24:@32335.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_42 fix2fixBox ( // @[Math.scala 141:30:@32345.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@32333.4 Math.scala 713:14:@32334.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@32340.4 Math.scala 713:14:@32341.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@32342.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@32353.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@32331.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@32338.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@32348.4]
endmodule
module RetimeWrapper_431( // @[:@33227.2]
  input        clock, // @[:@33228.4]
  input        reset, // @[:@33229.4]
  input        io_flow, // @[:@33230.4]
  input  [7:0] io_in, // @[:@33230.4]
  output [7:0] io_out // @[:@33230.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@33232.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@33232.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@33232.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@33232.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@33232.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@33232.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@33232.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@33245.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@33244.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@33243.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@33242.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@33241.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@33239.4]
endmodule
module RetimeWrapper_432( // @[:@33399.2]
  input        clock, // @[:@33400.4]
  input        reset, // @[:@33401.4]
  input        io_flow, // @[:@33402.4]
  input  [7:0] io_in, // @[:@33402.4]
  output [7:0] io_out // @[:@33402.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@33404.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@33404.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@33404.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@33404.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@33404.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@33404.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(4)) sr ( // @[RetimeShiftRegister.scala 15:20:@33404.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@33417.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@33416.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@33415.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@33414.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@33413.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@33411.4]
endmodule
module fix2fixBox_49( // @[:@33535.2]
  input        clock, // @[:@33536.4]
  input        reset, // @[:@33537.4]
  input  [8:0] io_a, // @[:@33538.4]
  input        io_flow, // @[:@33538.4]
  output [7:0] io_b // @[:@33538.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@33551.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@33551.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@33551.4]
  wire [7:0] RetimeWrapper_io_in; // @[package.scala 93:22:@33551.4]
  wire [7:0] RetimeWrapper_io_out; // @[package.scala 93:22:@33551.4]
  RetimeWrapper_20 RetimeWrapper ( // @[package.scala 93:22:@33551.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@33558.4]
  assign RetimeWrapper_clock = clock; // @[:@33552.4]
  assign RetimeWrapper_reset = reset; // @[:@33553.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@33555.4]
  assign RetimeWrapper_io_in = io_a[7:0]; // @[package.scala 94:16:@33554.4]
endmodule
module x496_sum( // @[:@33560.2]
  input        clock, // @[:@33561.4]
  input        reset, // @[:@33562.4]
  input  [7:0] io_a, // @[:@33563.4]
  input  [7:0] io_b, // @[:@33563.4]
  input        io_flow, // @[:@33563.4]
  output [7:0] io_result // @[:@33563.4]
);
  wire [7:0] __io_b; // @[Math.scala 709:24:@33571.4]
  wire [8:0] __io_result; // @[Math.scala 709:24:@33571.4]
  wire [7:0] __1_io_b; // @[Math.scala 709:24:@33578.4]
  wire [8:0] __1_io_result; // @[Math.scala 709:24:@33578.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@33588.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@33588.4]
  wire [8:0] fix2fixBox_io_a; // @[Math.scala 141:30:@33588.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@33588.4]
  wire [7:0] fix2fixBox_io_b; // @[Math.scala 141:30:@33588.4]
  wire [8:0] a_upcast_number; // @[Math.scala 712:22:@33576.4 Math.scala 713:14:@33577.4]
  wire [8:0] b_upcast_number; // @[Math.scala 712:22:@33583.4 Math.scala 713:14:@33584.4]
  wire [9:0] _T_21; // @[Math.scala 136:37:@33585.4]
  __66 _ ( // @[Math.scala 709:24:@33571.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __66 __1 ( // @[Math.scala 709:24:@33578.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_49 fix2fixBox ( // @[Math.scala 141:30:@33588.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@33576.4 Math.scala 713:14:@33577.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@33583.4 Math.scala 713:14:@33584.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@33585.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@33596.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@33574.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@33581.4]
  assign fix2fixBox_clock = clock; // @[:@33589.4]
  assign fix2fixBox_reset = reset; // @[:@33590.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@33591.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@33594.4]
endmodule
module x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1( // @[:@38547.2]
  input          clock, // @[:@38548.4]
  input          reset, // @[:@38549.4]
  output         io_in_x316_TREADY, // @[:@38550.4]
  input  [255:0] io_in_x316_TDATA, // @[:@38550.4]
  input  [7:0]   io_in_x316_TID, // @[:@38550.4]
  input  [7:0]   io_in_x316_TDEST, // @[:@38550.4]
  output         io_in_x317_TVALID, // @[:@38550.4]
  input          io_in_x317_TREADY, // @[:@38550.4]
  output [255:0] io_in_x317_TDATA, // @[:@38550.4]
  input          io_sigsIn_backpressure, // @[:@38550.4]
  input          io_sigsIn_datapathEn, // @[:@38550.4]
  input          io_sigsIn_break, // @[:@38550.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_1, // @[:@38550.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_0, // @[:@38550.4]
  input          io_sigsIn_cchainOutputs_0_oobs_0, // @[:@38550.4]
  input          io_sigsIn_cchainOutputs_0_oobs_1, // @[:@38550.4]
  input          io_rr // @[:@38550.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@38564.4]
  wire [31:0] __io_result; // @[Math.scala 709:24:@38564.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@38576.4]
  wire [31:0] __1_io_result; // @[Math.scala 709:24:@38576.4]
  wire  x329_lb_0_clock; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire  x329_lb_0_reset; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_rPort_17_banks_1; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_rPort_17_banks_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_rPort_17_ofs_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire  x329_lb_0_io_rPort_17_en_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire  x329_lb_0_io_rPort_17_backpressure; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_rPort_17_output_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_rPort_16_banks_1; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_rPort_16_banks_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_rPort_16_ofs_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire  x329_lb_0_io_rPort_16_en_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire  x329_lb_0_io_rPort_16_backpressure; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_rPort_16_output_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_rPort_15_banks_1; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_rPort_15_banks_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_rPort_15_ofs_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire  x329_lb_0_io_rPort_15_en_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire  x329_lb_0_io_rPort_15_backpressure; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_rPort_15_output_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_rPort_14_banks_1; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_rPort_14_banks_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_rPort_14_ofs_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire  x329_lb_0_io_rPort_14_en_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire  x329_lb_0_io_rPort_14_backpressure; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_rPort_14_output_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_rPort_13_banks_1; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_rPort_13_banks_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_rPort_13_ofs_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire  x329_lb_0_io_rPort_13_en_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire  x329_lb_0_io_rPort_13_backpressure; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_rPort_13_output_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_rPort_12_banks_1; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_rPort_12_banks_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_rPort_12_ofs_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire  x329_lb_0_io_rPort_12_en_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire  x329_lb_0_io_rPort_12_backpressure; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_rPort_12_output_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_rPort_11_banks_1; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_rPort_11_banks_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_rPort_11_ofs_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire  x329_lb_0_io_rPort_11_en_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire  x329_lb_0_io_rPort_11_backpressure; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_rPort_11_output_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_rPort_10_banks_1; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_rPort_10_banks_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_rPort_10_ofs_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire  x329_lb_0_io_rPort_10_en_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire  x329_lb_0_io_rPort_10_backpressure; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_rPort_10_output_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_rPort_9_banks_1; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_rPort_9_banks_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_rPort_9_ofs_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire  x329_lb_0_io_rPort_9_en_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire  x329_lb_0_io_rPort_9_backpressure; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_rPort_9_output_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_rPort_8_banks_1; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_rPort_8_banks_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_rPort_8_ofs_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire  x329_lb_0_io_rPort_8_en_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire  x329_lb_0_io_rPort_8_backpressure; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_rPort_8_output_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_rPort_7_banks_1; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_rPort_7_banks_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_rPort_7_ofs_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire  x329_lb_0_io_rPort_7_en_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire  x329_lb_0_io_rPort_7_backpressure; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_rPort_7_output_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_rPort_6_banks_1; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_rPort_6_banks_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_rPort_6_ofs_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire  x329_lb_0_io_rPort_6_en_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire  x329_lb_0_io_rPort_6_backpressure; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_rPort_6_output_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_rPort_5_banks_1; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_rPort_5_banks_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_rPort_5_ofs_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire  x329_lb_0_io_rPort_5_en_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire  x329_lb_0_io_rPort_5_backpressure; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_rPort_5_output_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_rPort_4_banks_1; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_rPort_4_banks_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_rPort_4_ofs_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire  x329_lb_0_io_rPort_4_en_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire  x329_lb_0_io_rPort_4_backpressure; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_rPort_4_output_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_rPort_3_banks_1; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_rPort_3_banks_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_rPort_3_ofs_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire  x329_lb_0_io_rPort_3_en_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire  x329_lb_0_io_rPort_3_backpressure; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_rPort_3_output_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_rPort_2_banks_1; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_rPort_2_banks_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_rPort_2_ofs_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire  x329_lb_0_io_rPort_2_en_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire  x329_lb_0_io_rPort_2_backpressure; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_rPort_2_output_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_rPort_1_banks_1; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_rPort_1_banks_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_rPort_1_ofs_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire  x329_lb_0_io_rPort_1_en_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire  x329_lb_0_io_rPort_1_backpressure; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_rPort_1_output_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_rPort_0_banks_1; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_rPort_0_banks_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_rPort_0_ofs_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire  x329_lb_0_io_rPort_0_en_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire  x329_lb_0_io_rPort_0_backpressure; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_rPort_0_output_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_wPort_3_banks_1; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_wPort_3_banks_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_wPort_3_ofs_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_wPort_3_data_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire  x329_lb_0_io_wPort_3_en_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_wPort_2_banks_1; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_wPort_2_banks_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_wPort_2_ofs_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_wPort_2_data_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire  x329_lb_0_io_wPort_2_en_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_wPort_1_banks_1; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_wPort_1_banks_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_wPort_1_ofs_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_wPort_1_data_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire  x329_lb_0_io_wPort_1_en_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_wPort_0_banks_1; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [2:0] x329_lb_0_io_wPort_0_banks_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_wPort_0_ofs_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire [7:0] x329_lb_0_io_wPort_0_data_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire  x329_lb_0_io_wPort_0_en_0; // @[m_x329_lb_0.scala 47:17:@38586.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@38744.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@38744.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@38744.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@38744.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@38744.4]
  wire  x340_1_clock; // @[Math.scala 366:24:@38828.4]
  wire  x340_1_reset; // @[Math.scala 366:24:@38828.4]
  wire [31:0] x340_1_io_a; // @[Math.scala 366:24:@38828.4]
  wire [31:0] x340_1_io_b; // @[Math.scala 366:24:@38828.4]
  wire  x340_1_io_flow; // @[Math.scala 366:24:@38828.4]
  wire [31:0] x340_1_io_result; // @[Math.scala 366:24:@38828.4]
  wire  x342_mul_1_clock; // @[Math.scala 262:24:@38849.4]
  wire  x342_mul_1_reset; // @[Math.scala 262:24:@38849.4]
  wire [31:0] x342_mul_1_io_a; // @[Math.scala 262:24:@38849.4]
  wire  x342_mul_1_io_flow; // @[Math.scala 262:24:@38849.4]
  wire [31:0] x342_mul_1_io_result; // @[Math.scala 262:24:@38849.4]
  wire  x343_div_1_clock; // @[Math.scala 327:24:@38861.4]
  wire  x343_div_1_reset; // @[Math.scala 327:24:@38861.4]
  wire [31:0] x343_div_1_io_a; // @[Math.scala 327:24:@38861.4]
  wire  x343_div_1_io_flow; // @[Math.scala 327:24:@38861.4]
  wire [31:0] x343_div_1_io_result; // @[Math.scala 327:24:@38861.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@38871.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@38871.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@38871.4]
  wire [31:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@38871.4]
  wire [31:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@38871.4]
  wire  x344_sum_1_clock; // @[Math.scala 150:24:@38880.4]
  wire  x344_sum_1_reset; // @[Math.scala 150:24:@38880.4]
  wire [31:0] x344_sum_1_io_a; // @[Math.scala 150:24:@38880.4]
  wire [31:0] x344_sum_1_io_b; // @[Math.scala 150:24:@38880.4]
  wire  x344_sum_1_io_flow; // @[Math.scala 150:24:@38880.4]
  wire [31:0] x344_sum_1_io_result; // @[Math.scala 150:24:@38880.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@38890.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@38890.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@38890.4]
  wire [31:0] RetimeWrapper_2_io_in; // @[package.scala 93:22:@38890.4]
  wire [31:0] RetimeWrapper_2_io_out; // @[package.scala 93:22:@38890.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@38899.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@38899.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@38899.4]
  wire [31:0] RetimeWrapper_3_io_in; // @[package.scala 93:22:@38899.4]
  wire [31:0] RetimeWrapper_3_io_out; // @[package.scala 93:22:@38899.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@38908.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@38908.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@38908.4]
  wire [31:0] RetimeWrapper_4_io_in; // @[package.scala 93:22:@38908.4]
  wire [31:0] RetimeWrapper_4_io_out; // @[package.scala 93:22:@38908.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@38917.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@38917.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@38917.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@38917.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@38917.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@38926.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@38926.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@38926.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@38926.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@38926.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@38935.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@38935.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@38935.4]
  wire [7:0] RetimeWrapper_7_io_in; // @[package.scala 93:22:@38935.4]
  wire [7:0] RetimeWrapper_7_io_out; // @[package.scala 93:22:@38935.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@38946.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@38946.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@38946.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@38946.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@38946.4]
  wire  x346_rdcol_1_clock; // @[Math.scala 150:24:@38969.4]
  wire  x346_rdcol_1_reset; // @[Math.scala 150:24:@38969.4]
  wire [31:0] x346_rdcol_1_io_a; // @[Math.scala 150:24:@38969.4]
  wire [31:0] x346_rdcol_1_io_b; // @[Math.scala 150:24:@38969.4]
  wire  x346_rdcol_1_io_flow; // @[Math.scala 150:24:@38969.4]
  wire [31:0] x346_rdcol_1_io_result; // @[Math.scala 150:24:@38969.4]
  wire  x348_1_clock; // @[Math.scala 366:24:@38983.4]
  wire  x348_1_reset; // @[Math.scala 366:24:@38983.4]
  wire [31:0] x348_1_io_a; // @[Math.scala 366:24:@38983.4]
  wire [31:0] x348_1_io_b; // @[Math.scala 366:24:@38983.4]
  wire  x348_1_io_flow; // @[Math.scala 366:24:@38983.4]
  wire [31:0] x348_1_io_result; // @[Math.scala 366:24:@38983.4]
  wire  x349_div_1_clock; // @[Math.scala 327:24:@38995.4]
  wire  x349_div_1_reset; // @[Math.scala 327:24:@38995.4]
  wire [31:0] x349_div_1_io_a; // @[Math.scala 327:24:@38995.4]
  wire  x349_div_1_io_flow; // @[Math.scala 327:24:@38995.4]
  wire [31:0] x349_div_1_io_result; // @[Math.scala 327:24:@38995.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@39005.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@39005.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@39005.4]
  wire [31:0] RetimeWrapper_9_io_in; // @[package.scala 93:22:@39005.4]
  wire [31:0] RetimeWrapper_9_io_out; // @[package.scala 93:22:@39005.4]
  wire  x350_sum_1_clock; // @[Math.scala 150:24:@39014.4]
  wire  x350_sum_1_reset; // @[Math.scala 150:24:@39014.4]
  wire [31:0] x350_sum_1_io_a; // @[Math.scala 150:24:@39014.4]
  wire [31:0] x350_sum_1_io_b; // @[Math.scala 150:24:@39014.4]
  wire  x350_sum_1_io_flow; // @[Math.scala 150:24:@39014.4]
  wire [31:0] x350_sum_1_io_result; // @[Math.scala 150:24:@39014.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@39024.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@39024.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@39024.4]
  wire [7:0] RetimeWrapper_10_io_in; // @[package.scala 93:22:@39024.4]
  wire [7:0] RetimeWrapper_10_io_out; // @[package.scala 93:22:@39024.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@39033.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@39033.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@39033.4]
  wire [31:0] RetimeWrapper_11_io_in; // @[package.scala 93:22:@39033.4]
  wire [31:0] RetimeWrapper_11_io_out; // @[package.scala 93:22:@39033.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@39042.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@39042.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@39042.4]
  wire [31:0] RetimeWrapper_12_io_in; // @[package.scala 93:22:@39042.4]
  wire [31:0] RetimeWrapper_12_io_out; // @[package.scala 93:22:@39042.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@39053.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@39053.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@39053.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@39053.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@39053.4]
  wire  x352_rdcol_1_clock; // @[Math.scala 150:24:@39076.4]
  wire  x352_rdcol_1_reset; // @[Math.scala 150:24:@39076.4]
  wire [31:0] x352_rdcol_1_io_a; // @[Math.scala 150:24:@39076.4]
  wire [31:0] x352_rdcol_1_io_b; // @[Math.scala 150:24:@39076.4]
  wire  x352_rdcol_1_io_flow; // @[Math.scala 150:24:@39076.4]
  wire [31:0] x352_rdcol_1_io_result; // @[Math.scala 150:24:@39076.4]
  wire  x354_1_clock; // @[Math.scala 366:24:@39090.4]
  wire  x354_1_reset; // @[Math.scala 366:24:@39090.4]
  wire [31:0] x354_1_io_a; // @[Math.scala 366:24:@39090.4]
  wire [31:0] x354_1_io_b; // @[Math.scala 366:24:@39090.4]
  wire  x354_1_io_flow; // @[Math.scala 366:24:@39090.4]
  wire [31:0] x354_1_io_result; // @[Math.scala 366:24:@39090.4]
  wire  x355_div_1_clock; // @[Math.scala 327:24:@39102.4]
  wire  x355_div_1_reset; // @[Math.scala 327:24:@39102.4]
  wire [31:0] x355_div_1_io_a; // @[Math.scala 327:24:@39102.4]
  wire  x355_div_1_io_flow; // @[Math.scala 327:24:@39102.4]
  wire [31:0] x355_div_1_io_result; // @[Math.scala 327:24:@39102.4]
  wire  x356_sum_1_clock; // @[Math.scala 150:24:@39112.4]
  wire  x356_sum_1_reset; // @[Math.scala 150:24:@39112.4]
  wire [31:0] x356_sum_1_io_a; // @[Math.scala 150:24:@39112.4]
  wire [31:0] x356_sum_1_io_b; // @[Math.scala 150:24:@39112.4]
  wire  x356_sum_1_io_flow; // @[Math.scala 150:24:@39112.4]
  wire [31:0] x356_sum_1_io_result; // @[Math.scala 150:24:@39112.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@39122.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@39122.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@39122.4]
  wire [7:0] RetimeWrapper_14_io_in; // @[package.scala 93:22:@39122.4]
  wire [7:0] RetimeWrapper_14_io_out; // @[package.scala 93:22:@39122.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@39131.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@39131.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@39131.4]
  wire [31:0] RetimeWrapper_15_io_in; // @[package.scala 93:22:@39131.4]
  wire [31:0] RetimeWrapper_15_io_out; // @[package.scala 93:22:@39131.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@39140.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@39140.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@39140.4]
  wire [31:0] RetimeWrapper_16_io_in; // @[package.scala 93:22:@39140.4]
  wire [31:0] RetimeWrapper_16_io_out; // @[package.scala 93:22:@39140.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@39151.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@39151.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@39151.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@39151.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@39151.4]
  wire  x358_rdcol_1_clock; // @[Math.scala 150:24:@39174.4]
  wire  x358_rdcol_1_reset; // @[Math.scala 150:24:@39174.4]
  wire [31:0] x358_rdcol_1_io_a; // @[Math.scala 150:24:@39174.4]
  wire [31:0] x358_rdcol_1_io_b; // @[Math.scala 150:24:@39174.4]
  wire  x358_rdcol_1_io_flow; // @[Math.scala 150:24:@39174.4]
  wire [31:0] x358_rdcol_1_io_result; // @[Math.scala 150:24:@39174.4]
  wire  x360_1_clock; // @[Math.scala 366:24:@39188.4]
  wire  x360_1_reset; // @[Math.scala 366:24:@39188.4]
  wire [31:0] x360_1_io_a; // @[Math.scala 366:24:@39188.4]
  wire [31:0] x360_1_io_b; // @[Math.scala 366:24:@39188.4]
  wire  x360_1_io_flow; // @[Math.scala 366:24:@39188.4]
  wire [31:0] x360_1_io_result; // @[Math.scala 366:24:@39188.4]
  wire  x361_div_1_clock; // @[Math.scala 327:24:@39200.4]
  wire  x361_div_1_reset; // @[Math.scala 327:24:@39200.4]
  wire [31:0] x361_div_1_io_a; // @[Math.scala 327:24:@39200.4]
  wire  x361_div_1_io_flow; // @[Math.scala 327:24:@39200.4]
  wire [31:0] x361_div_1_io_result; // @[Math.scala 327:24:@39200.4]
  wire  x362_sum_1_clock; // @[Math.scala 150:24:@39210.4]
  wire  x362_sum_1_reset; // @[Math.scala 150:24:@39210.4]
  wire [31:0] x362_sum_1_io_a; // @[Math.scala 150:24:@39210.4]
  wire [31:0] x362_sum_1_io_b; // @[Math.scala 150:24:@39210.4]
  wire  x362_sum_1_io_flow; // @[Math.scala 150:24:@39210.4]
  wire [31:0] x362_sum_1_io_result; // @[Math.scala 150:24:@39210.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@39220.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@39220.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@39220.4]
  wire [31:0] RetimeWrapper_18_io_in; // @[package.scala 93:22:@39220.4]
  wire [31:0] RetimeWrapper_18_io_out; // @[package.scala 93:22:@39220.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@39229.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@39229.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@39229.4]
  wire [31:0] RetimeWrapper_19_io_in; // @[package.scala 93:22:@39229.4]
  wire [31:0] RetimeWrapper_19_io_out; // @[package.scala 93:22:@39229.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@39238.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@39238.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@39238.4]
  wire [7:0] RetimeWrapper_20_io_in; // @[package.scala 93:22:@39238.4]
  wire [7:0] RetimeWrapper_20_io_out; // @[package.scala 93:22:@39238.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@39249.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@39249.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@39249.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@39249.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@39249.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@39270.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@39270.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@39270.4]
  wire [31:0] RetimeWrapper_22_io_in; // @[package.scala 93:22:@39270.4]
  wire [31:0] RetimeWrapper_22_io_out; // @[package.scala 93:22:@39270.4]
  wire  x365_1_clock; // @[Math.scala 366:24:@39283.4]
  wire  x365_1_reset; // @[Math.scala 366:24:@39283.4]
  wire [31:0] x365_1_io_a; // @[Math.scala 366:24:@39283.4]
  wire [31:0] x365_1_io_b; // @[Math.scala 366:24:@39283.4]
  wire  x365_1_io_flow; // @[Math.scala 366:24:@39283.4]
  wire [31:0] x365_1_io_result; // @[Math.scala 366:24:@39283.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@39298.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@39298.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@39298.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@39298.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@39298.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@39307.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@39307.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@39307.4]
  wire [31:0] RetimeWrapper_24_io_in; // @[package.scala 93:22:@39307.4]
  wire [31:0] RetimeWrapper_24_io_out; // @[package.scala 93:22:@39307.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@39321.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@39321.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@39321.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@39321.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@39321.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@39330.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@39330.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@39330.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@39330.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@39330.4]
  wire  x372_mul_1_clock; // @[Math.scala 262:24:@39367.4]
  wire  x372_mul_1_reset; // @[Math.scala 262:24:@39367.4]
  wire [31:0] x372_mul_1_io_a; // @[Math.scala 262:24:@39367.4]
  wire  x372_mul_1_io_flow; // @[Math.scala 262:24:@39367.4]
  wire [31:0] x372_mul_1_io_result; // @[Math.scala 262:24:@39367.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@39377.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@39377.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@39377.4]
  wire [31:0] RetimeWrapper_27_io_in; // @[package.scala 93:22:@39377.4]
  wire [31:0] RetimeWrapper_27_io_out; // @[package.scala 93:22:@39377.4]
  wire  x373_sum_1_clock; // @[Math.scala 150:24:@39386.4]
  wire  x373_sum_1_reset; // @[Math.scala 150:24:@39386.4]
  wire [31:0] x373_sum_1_io_a; // @[Math.scala 150:24:@39386.4]
  wire [31:0] x373_sum_1_io_b; // @[Math.scala 150:24:@39386.4]
  wire  x373_sum_1_io_flow; // @[Math.scala 150:24:@39386.4]
  wire [31:0] x373_sum_1_io_result; // @[Math.scala 150:24:@39386.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@39396.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@39396.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@39396.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@39396.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@39396.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@39405.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@39405.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@39405.4]
  wire [31:0] RetimeWrapper_29_io_in; // @[package.scala 93:22:@39405.4]
  wire [31:0] RetimeWrapper_29_io_out; // @[package.scala 93:22:@39405.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@39414.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@39414.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@39414.4]
  wire [31:0] RetimeWrapper_30_io_in; // @[package.scala 93:22:@39414.4]
  wire [31:0] RetimeWrapper_30_io_out; // @[package.scala 93:22:@39414.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@39423.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@39423.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@39423.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@39423.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@39423.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@39432.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@39432.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@39432.4]
  wire [31:0] RetimeWrapper_32_io_in; // @[package.scala 93:22:@39432.4]
  wire [31:0] RetimeWrapper_32_io_out; // @[package.scala 93:22:@39432.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@39441.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@39441.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@39441.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@39441.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@39441.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@39453.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@39453.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@39453.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@39453.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@39453.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@39474.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@39474.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@39474.4]
  wire [31:0] RetimeWrapper_35_io_in; // @[package.scala 93:22:@39474.4]
  wire [31:0] RetimeWrapper_35_io_out; // @[package.scala 93:22:@39474.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@39488.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@39488.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@39488.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@39488.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@39488.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@39503.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@39503.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@39503.4]
  wire [31:0] RetimeWrapper_37_io_in; // @[package.scala 93:22:@39503.4]
  wire [31:0] RetimeWrapper_37_io_out; // @[package.scala 93:22:@39503.4]
  wire  x379_sum_1_clock; // @[Math.scala 150:24:@39512.4]
  wire  x379_sum_1_reset; // @[Math.scala 150:24:@39512.4]
  wire [31:0] x379_sum_1_io_a; // @[Math.scala 150:24:@39512.4]
  wire [31:0] x379_sum_1_io_b; // @[Math.scala 150:24:@39512.4]
  wire  x379_sum_1_io_flow; // @[Math.scala 150:24:@39512.4]
  wire [31:0] x379_sum_1_io_result; // @[Math.scala 150:24:@39512.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@39522.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@39522.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@39522.4]
  wire [31:0] RetimeWrapper_38_io_in; // @[package.scala 93:22:@39522.4]
  wire [31:0] RetimeWrapper_38_io_out; // @[package.scala 93:22:@39522.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@39531.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@39531.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@39531.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@39531.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@39531.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@39540.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@39540.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@39540.4]
  wire [31:0] RetimeWrapper_40_io_in; // @[package.scala 93:22:@39540.4]
  wire [31:0] RetimeWrapper_40_io_out; // @[package.scala 93:22:@39540.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@39552.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@39552.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@39552.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@39552.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@39552.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@39573.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@39573.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@39573.4]
  wire [31:0] RetimeWrapper_42_io_in; // @[package.scala 93:22:@39573.4]
  wire [31:0] RetimeWrapper_42_io_out; // @[package.scala 93:22:@39573.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@39587.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@39587.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@39587.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@39587.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@39587.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@39602.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@39602.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@39602.4]
  wire [31:0] RetimeWrapper_44_io_in; // @[package.scala 93:22:@39602.4]
  wire [31:0] RetimeWrapper_44_io_out; // @[package.scala 93:22:@39602.4]
  wire  x385_sum_1_clock; // @[Math.scala 150:24:@39611.4]
  wire  x385_sum_1_reset; // @[Math.scala 150:24:@39611.4]
  wire [31:0] x385_sum_1_io_a; // @[Math.scala 150:24:@39611.4]
  wire [31:0] x385_sum_1_io_b; // @[Math.scala 150:24:@39611.4]
  wire  x385_sum_1_io_flow; // @[Math.scala 150:24:@39611.4]
  wire [31:0] x385_sum_1_io_result; // @[Math.scala 150:24:@39611.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@39621.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@39621.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@39621.4]
  wire [31:0] RetimeWrapper_45_io_in; // @[package.scala 93:22:@39621.4]
  wire [31:0] RetimeWrapper_45_io_out; // @[package.scala 93:22:@39621.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@39630.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@39630.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@39630.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@39630.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@39630.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@39639.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@39639.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@39639.4]
  wire [31:0] RetimeWrapper_47_io_in; // @[package.scala 93:22:@39639.4]
  wire [31:0] RetimeWrapper_47_io_out; // @[package.scala 93:22:@39639.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@39651.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@39651.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@39651.4]
  wire  RetimeWrapper_48_io_in; // @[package.scala 93:22:@39651.4]
  wire  RetimeWrapper_48_io_out; // @[package.scala 93:22:@39651.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@39672.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@39672.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@39672.4]
  wire [31:0] RetimeWrapper_49_io_in; // @[package.scala 93:22:@39672.4]
  wire [31:0] RetimeWrapper_49_io_out; // @[package.scala 93:22:@39672.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@39688.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@39688.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@39688.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@39688.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@39688.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@39703.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@39703.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@39703.4]
  wire [31:0] RetimeWrapper_51_io_in; // @[package.scala 93:22:@39703.4]
  wire [31:0] RetimeWrapper_51_io_out; // @[package.scala 93:22:@39703.4]
  wire  x391_sum_1_clock; // @[Math.scala 150:24:@39712.4]
  wire  x391_sum_1_reset; // @[Math.scala 150:24:@39712.4]
  wire [31:0] x391_sum_1_io_a; // @[Math.scala 150:24:@39712.4]
  wire [31:0] x391_sum_1_io_b; // @[Math.scala 150:24:@39712.4]
  wire  x391_sum_1_io_flow; // @[Math.scala 150:24:@39712.4]
  wire [31:0] x391_sum_1_io_result; // @[Math.scala 150:24:@39712.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@39722.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@39722.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@39722.4]
  wire [31:0] RetimeWrapper_52_io_in; // @[package.scala 93:22:@39722.4]
  wire [31:0] RetimeWrapper_52_io_out; // @[package.scala 93:22:@39722.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@39731.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@39731.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@39731.4]
  wire [31:0] RetimeWrapper_53_io_in; // @[package.scala 93:22:@39731.4]
  wire [31:0] RetimeWrapper_53_io_out; // @[package.scala 93:22:@39731.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@39740.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@39740.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@39740.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@39740.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@39740.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@39752.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@39752.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@39752.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@39752.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@39752.4]
  wire  x394_rdcol_1_clock; // @[Math.scala 150:24:@39775.4]
  wire  x394_rdcol_1_reset; // @[Math.scala 150:24:@39775.4]
  wire [31:0] x394_rdcol_1_io_a; // @[Math.scala 150:24:@39775.4]
  wire [31:0] x394_rdcol_1_io_b; // @[Math.scala 150:24:@39775.4]
  wire  x394_rdcol_1_io_flow; // @[Math.scala 150:24:@39775.4]
  wire [31:0] x394_rdcol_1_io_result; // @[Math.scala 150:24:@39775.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@39790.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@39790.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@39790.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@39790.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@39790.4]
  wire  x398_1_clock; // @[Math.scala 366:24:@39807.4]
  wire  x398_1_reset; // @[Math.scala 366:24:@39807.4]
  wire [31:0] x398_1_io_a; // @[Math.scala 366:24:@39807.4]
  wire [31:0] x398_1_io_b; // @[Math.scala 366:24:@39807.4]
  wire  x398_1_io_flow; // @[Math.scala 366:24:@39807.4]
  wire [31:0] x398_1_io_result; // @[Math.scala 366:24:@39807.4]
  wire  x399_div_1_clock; // @[Math.scala 327:24:@39819.4]
  wire  x399_div_1_reset; // @[Math.scala 327:24:@39819.4]
  wire [31:0] x399_div_1_io_a; // @[Math.scala 327:24:@39819.4]
  wire  x399_div_1_io_flow; // @[Math.scala 327:24:@39819.4]
  wire [31:0] x399_div_1_io_result; // @[Math.scala 327:24:@39819.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@39829.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@39829.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@39829.4]
  wire [31:0] RetimeWrapper_57_io_in; // @[package.scala 93:22:@39829.4]
  wire [31:0] RetimeWrapper_57_io_out; // @[package.scala 93:22:@39829.4]
  wire  x400_sum_1_clock; // @[Math.scala 150:24:@39838.4]
  wire  x400_sum_1_reset; // @[Math.scala 150:24:@39838.4]
  wire [31:0] x400_sum_1_io_a; // @[Math.scala 150:24:@39838.4]
  wire [31:0] x400_sum_1_io_b; // @[Math.scala 150:24:@39838.4]
  wire  x400_sum_1_io_flow; // @[Math.scala 150:24:@39838.4]
  wire [31:0] x400_sum_1_io_result; // @[Math.scala 150:24:@39838.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@39848.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@39848.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@39848.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@39848.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@39848.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@39857.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@39857.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@39857.4]
  wire [31:0] RetimeWrapper_59_io_in; // @[package.scala 93:22:@39857.4]
  wire [31:0] RetimeWrapper_59_io_out; // @[package.scala 93:22:@39857.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@39866.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@39866.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@39866.4]
  wire [31:0] RetimeWrapper_60_io_in; // @[package.scala 93:22:@39866.4]
  wire [31:0] RetimeWrapper_60_io_out; // @[package.scala 93:22:@39866.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@39878.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@39878.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@39878.4]
  wire  RetimeWrapper_61_io_in; // @[package.scala 93:22:@39878.4]
  wire  RetimeWrapper_61_io_out; // @[package.scala 93:22:@39878.4]
  wire  x403_rdcol_1_clock; // @[Math.scala 150:24:@39901.4]
  wire  x403_rdcol_1_reset; // @[Math.scala 150:24:@39901.4]
  wire [31:0] x403_rdcol_1_io_a; // @[Math.scala 150:24:@39901.4]
  wire [31:0] x403_rdcol_1_io_b; // @[Math.scala 150:24:@39901.4]
  wire  x403_rdcol_1_io_flow; // @[Math.scala 150:24:@39901.4]
  wire [31:0] x403_rdcol_1_io_result; // @[Math.scala 150:24:@39901.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@39916.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@39916.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@39916.4]
  wire  RetimeWrapper_62_io_in; // @[package.scala 93:22:@39916.4]
  wire  RetimeWrapper_62_io_out; // @[package.scala 93:22:@39916.4]
  wire  x407_1_clock; // @[Math.scala 366:24:@39933.4]
  wire  x407_1_reset; // @[Math.scala 366:24:@39933.4]
  wire [31:0] x407_1_io_a; // @[Math.scala 366:24:@39933.4]
  wire [31:0] x407_1_io_b; // @[Math.scala 366:24:@39933.4]
  wire  x407_1_io_flow; // @[Math.scala 366:24:@39933.4]
  wire [31:0] x407_1_io_result; // @[Math.scala 366:24:@39933.4]
  wire  x408_div_1_clock; // @[Math.scala 327:24:@39945.4]
  wire  x408_div_1_reset; // @[Math.scala 327:24:@39945.4]
  wire [31:0] x408_div_1_io_a; // @[Math.scala 327:24:@39945.4]
  wire  x408_div_1_io_flow; // @[Math.scala 327:24:@39945.4]
  wire [31:0] x408_div_1_io_result; // @[Math.scala 327:24:@39945.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@39955.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@39955.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@39955.4]
  wire [31:0] RetimeWrapper_63_io_in; // @[package.scala 93:22:@39955.4]
  wire [31:0] RetimeWrapper_63_io_out; // @[package.scala 93:22:@39955.4]
  wire  x409_sum_1_clock; // @[Math.scala 150:24:@39964.4]
  wire  x409_sum_1_reset; // @[Math.scala 150:24:@39964.4]
  wire [31:0] x409_sum_1_io_a; // @[Math.scala 150:24:@39964.4]
  wire [31:0] x409_sum_1_io_b; // @[Math.scala 150:24:@39964.4]
  wire  x409_sum_1_io_flow; // @[Math.scala 150:24:@39964.4]
  wire [31:0] x409_sum_1_io_result; // @[Math.scala 150:24:@39964.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@39974.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@39974.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@39974.4]
  wire [31:0] RetimeWrapper_64_io_in; // @[package.scala 93:22:@39974.4]
  wire [31:0] RetimeWrapper_64_io_out; // @[package.scala 93:22:@39974.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@39983.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@39983.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@39983.4]
  wire  RetimeWrapper_65_io_in; // @[package.scala 93:22:@39983.4]
  wire  RetimeWrapper_65_io_out; // @[package.scala 93:22:@39983.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@39992.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@39992.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@39992.4]
  wire [31:0] RetimeWrapper_66_io_in; // @[package.scala 93:22:@39992.4]
  wire [31:0] RetimeWrapper_66_io_out; // @[package.scala 93:22:@39992.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@40004.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@40004.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@40004.4]
  wire  RetimeWrapper_67_io_in; // @[package.scala 93:22:@40004.4]
  wire  RetimeWrapper_67_io_out; // @[package.scala 93:22:@40004.4]
  wire  x412_rdrow_1_clock; // @[Math.scala 191:24:@40027.4]
  wire  x412_rdrow_1_reset; // @[Math.scala 191:24:@40027.4]
  wire [31:0] x412_rdrow_1_io_a; // @[Math.scala 191:24:@40027.4]
  wire [31:0] x412_rdrow_1_io_b; // @[Math.scala 191:24:@40027.4]
  wire  x412_rdrow_1_io_flow; // @[Math.scala 191:24:@40027.4]
  wire [31:0] x412_rdrow_1_io_result; // @[Math.scala 191:24:@40027.4]
  wire  x413_1_clock; // @[Math.scala 366:24:@40039.4]
  wire  x413_1_reset; // @[Math.scala 366:24:@40039.4]
  wire [31:0] x413_1_io_a; // @[Math.scala 366:24:@40039.4]
  wire [31:0] x413_1_io_b; // @[Math.scala 366:24:@40039.4]
  wire  x413_1_io_flow; // @[Math.scala 366:24:@40039.4]
  wire [31:0] x413_1_io_result; // @[Math.scala 366:24:@40039.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@40054.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@40054.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@40054.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@40054.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@40054.4]
  wire  x419_mul_1_clock; // @[Math.scala 262:24:@40091.4]
  wire  x419_mul_1_reset; // @[Math.scala 262:24:@40091.4]
  wire [31:0] x419_mul_1_io_a; // @[Math.scala 262:24:@40091.4]
  wire  x419_mul_1_io_flow; // @[Math.scala 262:24:@40091.4]
  wire [31:0] x419_mul_1_io_result; // @[Math.scala 262:24:@40091.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@40101.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@40101.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@40101.4]
  wire [31:0] RetimeWrapper_69_io_in; // @[package.scala 93:22:@40101.4]
  wire [31:0] RetimeWrapper_69_io_out; // @[package.scala 93:22:@40101.4]
  wire  x420_sum_1_clock; // @[Math.scala 150:24:@40110.4]
  wire  x420_sum_1_reset; // @[Math.scala 150:24:@40110.4]
  wire [31:0] x420_sum_1_io_a; // @[Math.scala 150:24:@40110.4]
  wire [31:0] x420_sum_1_io_b; // @[Math.scala 150:24:@40110.4]
  wire  x420_sum_1_io_flow; // @[Math.scala 150:24:@40110.4]
  wire [31:0] x420_sum_1_io_result; // @[Math.scala 150:24:@40110.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@40120.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@40120.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@40120.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@40120.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@40120.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@40129.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@40129.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@40129.4]
  wire [31:0] RetimeWrapper_71_io_in; // @[package.scala 93:22:@40129.4]
  wire [31:0] RetimeWrapper_71_io_out; // @[package.scala 93:22:@40129.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@40141.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@40141.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@40141.4]
  wire  RetimeWrapper_72_io_in; // @[package.scala 93:22:@40141.4]
  wire  RetimeWrapper_72_io_out; // @[package.scala 93:22:@40141.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@40168.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@40168.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@40168.4]
  wire [31:0] RetimeWrapper_73_io_in; // @[package.scala 93:22:@40168.4]
  wire [31:0] RetimeWrapper_73_io_out; // @[package.scala 93:22:@40168.4]
  wire  x425_sum_1_clock; // @[Math.scala 150:24:@40179.4]
  wire  x425_sum_1_reset; // @[Math.scala 150:24:@40179.4]
  wire [31:0] x425_sum_1_io_a; // @[Math.scala 150:24:@40179.4]
  wire [31:0] x425_sum_1_io_b; // @[Math.scala 150:24:@40179.4]
  wire  x425_sum_1_io_flow; // @[Math.scala 150:24:@40179.4]
  wire [31:0] x425_sum_1_io_result; // @[Math.scala 150:24:@40179.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@40189.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@40189.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@40189.4]
  wire  RetimeWrapper_74_io_in; // @[package.scala 93:22:@40189.4]
  wire  RetimeWrapper_74_io_out; // @[package.scala 93:22:@40189.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@40201.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@40201.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@40201.4]
  wire  RetimeWrapper_75_io_in; // @[package.scala 93:22:@40201.4]
  wire  RetimeWrapper_75_io_out; // @[package.scala 93:22:@40201.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@40228.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@40228.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@40228.4]
  wire [31:0] RetimeWrapper_76_io_in; // @[package.scala 93:22:@40228.4]
  wire [31:0] RetimeWrapper_76_io_out; // @[package.scala 93:22:@40228.4]
  wire  x430_sum_1_clock; // @[Math.scala 150:24:@40237.4]
  wire  x430_sum_1_reset; // @[Math.scala 150:24:@40237.4]
  wire [31:0] x430_sum_1_io_a; // @[Math.scala 150:24:@40237.4]
  wire [31:0] x430_sum_1_io_b; // @[Math.scala 150:24:@40237.4]
  wire  x430_sum_1_io_flow; // @[Math.scala 150:24:@40237.4]
  wire [31:0] x430_sum_1_io_result; // @[Math.scala 150:24:@40237.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@40247.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@40247.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@40247.4]
  wire  RetimeWrapper_77_io_in; // @[package.scala 93:22:@40247.4]
  wire  RetimeWrapper_77_io_out; // @[package.scala 93:22:@40247.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@40259.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@40259.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@40259.4]
  wire  RetimeWrapper_78_io_in; // @[package.scala 93:22:@40259.4]
  wire  RetimeWrapper_78_io_out; // @[package.scala 93:22:@40259.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@40280.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@40280.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@40280.4]
  wire  RetimeWrapper_79_io_in; // @[package.scala 93:22:@40280.4]
  wire  RetimeWrapper_79_io_out; // @[package.scala 93:22:@40280.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@40295.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@40295.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@40295.4]
  wire [31:0] RetimeWrapper_80_io_in; // @[package.scala 93:22:@40295.4]
  wire [31:0] RetimeWrapper_80_io_out; // @[package.scala 93:22:@40295.4]
  wire  x435_sum_1_clock; // @[Math.scala 150:24:@40304.4]
  wire  x435_sum_1_reset; // @[Math.scala 150:24:@40304.4]
  wire [31:0] x435_sum_1_io_a; // @[Math.scala 150:24:@40304.4]
  wire [31:0] x435_sum_1_io_b; // @[Math.scala 150:24:@40304.4]
  wire  x435_sum_1_io_flow; // @[Math.scala 150:24:@40304.4]
  wire [31:0] x435_sum_1_io_result; // @[Math.scala 150:24:@40304.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@40314.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@40314.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@40314.4]
  wire  RetimeWrapper_81_io_in; // @[package.scala 93:22:@40314.4]
  wire  RetimeWrapper_81_io_out; // @[package.scala 93:22:@40314.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@40326.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@40326.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@40326.4]
  wire  RetimeWrapper_82_io_in; // @[package.scala 93:22:@40326.4]
  wire  RetimeWrapper_82_io_out; // @[package.scala 93:22:@40326.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@40353.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@40353.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@40353.4]
  wire [31:0] RetimeWrapper_83_io_in; // @[package.scala 93:22:@40353.4]
  wire [31:0] RetimeWrapper_83_io_out; // @[package.scala 93:22:@40353.4]
  wire  x440_sum_1_clock; // @[Math.scala 150:24:@40362.4]
  wire  x440_sum_1_reset; // @[Math.scala 150:24:@40362.4]
  wire [31:0] x440_sum_1_io_a; // @[Math.scala 150:24:@40362.4]
  wire [31:0] x440_sum_1_io_b; // @[Math.scala 150:24:@40362.4]
  wire  x440_sum_1_io_flow; // @[Math.scala 150:24:@40362.4]
  wire [31:0] x440_sum_1_io_result; // @[Math.scala 150:24:@40362.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@40372.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@40372.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@40372.4]
  wire  RetimeWrapper_84_io_in; // @[package.scala 93:22:@40372.4]
  wire  RetimeWrapper_84_io_out; // @[package.scala 93:22:@40372.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@40384.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@40384.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@40384.4]
  wire  RetimeWrapper_85_io_in; // @[package.scala 93:22:@40384.4]
  wire  RetimeWrapper_85_io_out; // @[package.scala 93:22:@40384.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@40411.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@40411.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@40411.4]
  wire [31:0] RetimeWrapper_86_io_in; // @[package.scala 93:22:@40411.4]
  wire [31:0] RetimeWrapper_86_io_out; // @[package.scala 93:22:@40411.4]
  wire  x445_sum_1_clock; // @[Math.scala 150:24:@40420.4]
  wire  x445_sum_1_reset; // @[Math.scala 150:24:@40420.4]
  wire [31:0] x445_sum_1_io_a; // @[Math.scala 150:24:@40420.4]
  wire [31:0] x445_sum_1_io_b; // @[Math.scala 150:24:@40420.4]
  wire  x445_sum_1_io_flow; // @[Math.scala 150:24:@40420.4]
  wire [31:0] x445_sum_1_io_result; // @[Math.scala 150:24:@40420.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@40430.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@40430.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@40430.4]
  wire  RetimeWrapper_87_io_in; // @[package.scala 93:22:@40430.4]
  wire  RetimeWrapper_87_io_out; // @[package.scala 93:22:@40430.4]
  wire  RetimeWrapper_88_clock; // @[package.scala 93:22:@40442.4]
  wire  RetimeWrapper_88_reset; // @[package.scala 93:22:@40442.4]
  wire  RetimeWrapper_88_io_flow; // @[package.scala 93:22:@40442.4]
  wire  RetimeWrapper_88_io_in; // @[package.scala 93:22:@40442.4]
  wire  RetimeWrapper_88_io_out; // @[package.scala 93:22:@40442.4]
  wire  x448_rdrow_1_clock; // @[Math.scala 191:24:@40465.4]
  wire  x448_rdrow_1_reset; // @[Math.scala 191:24:@40465.4]
  wire [31:0] x448_rdrow_1_io_a; // @[Math.scala 191:24:@40465.4]
  wire [31:0] x448_rdrow_1_io_b; // @[Math.scala 191:24:@40465.4]
  wire  x448_rdrow_1_io_flow; // @[Math.scala 191:24:@40465.4]
  wire [31:0] x448_rdrow_1_io_result; // @[Math.scala 191:24:@40465.4]
  wire  x449_1_clock; // @[Math.scala 366:24:@40477.4]
  wire  x449_1_reset; // @[Math.scala 366:24:@40477.4]
  wire [31:0] x449_1_io_a; // @[Math.scala 366:24:@40477.4]
  wire [31:0] x449_1_io_b; // @[Math.scala 366:24:@40477.4]
  wire  x449_1_io_flow; // @[Math.scala 366:24:@40477.4]
  wire [31:0] x449_1_io_result; // @[Math.scala 366:24:@40477.4]
  wire  RetimeWrapper_89_clock; // @[package.scala 93:22:@40492.4]
  wire  RetimeWrapper_89_reset; // @[package.scala 93:22:@40492.4]
  wire  RetimeWrapper_89_io_flow; // @[package.scala 93:22:@40492.4]
  wire  RetimeWrapper_89_io_in; // @[package.scala 93:22:@40492.4]
  wire  RetimeWrapper_89_io_out; // @[package.scala 93:22:@40492.4]
  wire  x455_mul_1_clock; // @[Math.scala 262:24:@40529.4]
  wire  x455_mul_1_reset; // @[Math.scala 262:24:@40529.4]
  wire [31:0] x455_mul_1_io_a; // @[Math.scala 262:24:@40529.4]
  wire  x455_mul_1_io_flow; // @[Math.scala 262:24:@40529.4]
  wire [31:0] x455_mul_1_io_result; // @[Math.scala 262:24:@40529.4]
  wire  x456_sum_1_clock; // @[Math.scala 150:24:@40539.4]
  wire  x456_sum_1_reset; // @[Math.scala 150:24:@40539.4]
  wire [31:0] x456_sum_1_io_a; // @[Math.scala 150:24:@40539.4]
  wire [31:0] x456_sum_1_io_b; // @[Math.scala 150:24:@40539.4]
  wire  x456_sum_1_io_flow; // @[Math.scala 150:24:@40539.4]
  wire [31:0] x456_sum_1_io_result; // @[Math.scala 150:24:@40539.4]
  wire  RetimeWrapper_90_clock; // @[package.scala 93:22:@40549.4]
  wire  RetimeWrapper_90_reset; // @[package.scala 93:22:@40549.4]
  wire  RetimeWrapper_90_io_flow; // @[package.scala 93:22:@40549.4]
  wire  RetimeWrapper_90_io_in; // @[package.scala 93:22:@40549.4]
  wire  RetimeWrapper_90_io_out; // @[package.scala 93:22:@40549.4]
  wire  RetimeWrapper_91_clock; // @[package.scala 93:22:@40558.4]
  wire  RetimeWrapper_91_reset; // @[package.scala 93:22:@40558.4]
  wire  RetimeWrapper_91_io_flow; // @[package.scala 93:22:@40558.4]
  wire [31:0] RetimeWrapper_91_io_in; // @[package.scala 93:22:@40558.4]
  wire [31:0] RetimeWrapper_91_io_out; // @[package.scala 93:22:@40558.4]
  wire  RetimeWrapper_92_clock; // @[package.scala 93:22:@40570.4]
  wire  RetimeWrapper_92_reset; // @[package.scala 93:22:@40570.4]
  wire  RetimeWrapper_92_io_flow; // @[package.scala 93:22:@40570.4]
  wire  RetimeWrapper_92_io_in; // @[package.scala 93:22:@40570.4]
  wire  RetimeWrapper_92_io_out; // @[package.scala 93:22:@40570.4]
  wire  x461_sum_1_clock; // @[Math.scala 150:24:@40599.4]
  wire  x461_sum_1_reset; // @[Math.scala 150:24:@40599.4]
  wire [31:0] x461_sum_1_io_a; // @[Math.scala 150:24:@40599.4]
  wire [31:0] x461_sum_1_io_b; // @[Math.scala 150:24:@40599.4]
  wire  x461_sum_1_io_flow; // @[Math.scala 150:24:@40599.4]
  wire [31:0] x461_sum_1_io_result; // @[Math.scala 150:24:@40599.4]
  wire  RetimeWrapper_93_clock; // @[package.scala 93:22:@40609.4]
  wire  RetimeWrapper_93_reset; // @[package.scala 93:22:@40609.4]
  wire  RetimeWrapper_93_io_flow; // @[package.scala 93:22:@40609.4]
  wire  RetimeWrapper_93_io_in; // @[package.scala 93:22:@40609.4]
  wire  RetimeWrapper_93_io_out; // @[package.scala 93:22:@40609.4]
  wire  RetimeWrapper_94_clock; // @[package.scala 93:22:@40621.4]
  wire  RetimeWrapper_94_reset; // @[package.scala 93:22:@40621.4]
  wire  RetimeWrapper_94_io_flow; // @[package.scala 93:22:@40621.4]
  wire  RetimeWrapper_94_io_in; // @[package.scala 93:22:@40621.4]
  wire  RetimeWrapper_94_io_out; // @[package.scala 93:22:@40621.4]
  wire  x466_sum_1_clock; // @[Math.scala 150:24:@40648.4]
  wire  x466_sum_1_reset; // @[Math.scala 150:24:@40648.4]
  wire [31:0] x466_sum_1_io_a; // @[Math.scala 150:24:@40648.4]
  wire [31:0] x466_sum_1_io_b; // @[Math.scala 150:24:@40648.4]
  wire  x466_sum_1_io_flow; // @[Math.scala 150:24:@40648.4]
  wire [31:0] x466_sum_1_io_result; // @[Math.scala 150:24:@40648.4]
  wire  RetimeWrapper_95_clock; // @[package.scala 93:22:@40658.4]
  wire  RetimeWrapper_95_reset; // @[package.scala 93:22:@40658.4]
  wire  RetimeWrapper_95_io_flow; // @[package.scala 93:22:@40658.4]
  wire  RetimeWrapper_95_io_in; // @[package.scala 93:22:@40658.4]
  wire  RetimeWrapper_95_io_out; // @[package.scala 93:22:@40658.4]
  wire  RetimeWrapper_96_clock; // @[package.scala 93:22:@40670.4]
  wire  RetimeWrapper_96_reset; // @[package.scala 93:22:@40670.4]
  wire  RetimeWrapper_96_io_flow; // @[package.scala 93:22:@40670.4]
  wire  RetimeWrapper_96_io_in; // @[package.scala 93:22:@40670.4]
  wire  RetimeWrapper_96_io_out; // @[package.scala 93:22:@40670.4]
  wire  x471_sum_1_clock; // @[Math.scala 150:24:@40697.4]
  wire  x471_sum_1_reset; // @[Math.scala 150:24:@40697.4]
  wire [31:0] x471_sum_1_io_a; // @[Math.scala 150:24:@40697.4]
  wire [31:0] x471_sum_1_io_b; // @[Math.scala 150:24:@40697.4]
  wire  x471_sum_1_io_flow; // @[Math.scala 150:24:@40697.4]
  wire [31:0] x471_sum_1_io_result; // @[Math.scala 150:24:@40697.4]
  wire  RetimeWrapper_97_clock; // @[package.scala 93:22:@40707.4]
  wire  RetimeWrapper_97_reset; // @[package.scala 93:22:@40707.4]
  wire  RetimeWrapper_97_io_flow; // @[package.scala 93:22:@40707.4]
  wire  RetimeWrapper_97_io_in; // @[package.scala 93:22:@40707.4]
  wire  RetimeWrapper_97_io_out; // @[package.scala 93:22:@40707.4]
  wire  RetimeWrapper_98_clock; // @[package.scala 93:22:@40719.4]
  wire  RetimeWrapper_98_reset; // @[package.scala 93:22:@40719.4]
  wire  RetimeWrapper_98_io_flow; // @[package.scala 93:22:@40719.4]
  wire  RetimeWrapper_98_io_in; // @[package.scala 93:22:@40719.4]
  wire  RetimeWrapper_98_io_out; // @[package.scala 93:22:@40719.4]
  wire  x476_sum_1_clock; // @[Math.scala 150:24:@40746.4]
  wire  x476_sum_1_reset; // @[Math.scala 150:24:@40746.4]
  wire [31:0] x476_sum_1_io_a; // @[Math.scala 150:24:@40746.4]
  wire [31:0] x476_sum_1_io_b; // @[Math.scala 150:24:@40746.4]
  wire  x476_sum_1_io_flow; // @[Math.scala 150:24:@40746.4]
  wire [31:0] x476_sum_1_io_result; // @[Math.scala 150:24:@40746.4]
  wire  RetimeWrapper_99_clock; // @[package.scala 93:22:@40756.4]
  wire  RetimeWrapper_99_reset; // @[package.scala 93:22:@40756.4]
  wire  RetimeWrapper_99_io_flow; // @[package.scala 93:22:@40756.4]
  wire  RetimeWrapper_99_io_in; // @[package.scala 93:22:@40756.4]
  wire  RetimeWrapper_99_io_out; // @[package.scala 93:22:@40756.4]
  wire  RetimeWrapper_100_clock; // @[package.scala 93:22:@40768.4]
  wire  RetimeWrapper_100_reset; // @[package.scala 93:22:@40768.4]
  wire  RetimeWrapper_100_io_flow; // @[package.scala 93:22:@40768.4]
  wire  RetimeWrapper_100_io_in; // @[package.scala 93:22:@40768.4]
  wire  RetimeWrapper_100_io_out; // @[package.scala 93:22:@40768.4]
  wire  x481_sum_1_clock; // @[Math.scala 150:24:@40795.4]
  wire  x481_sum_1_reset; // @[Math.scala 150:24:@40795.4]
  wire [31:0] x481_sum_1_io_a; // @[Math.scala 150:24:@40795.4]
  wire [31:0] x481_sum_1_io_b; // @[Math.scala 150:24:@40795.4]
  wire  x481_sum_1_io_flow; // @[Math.scala 150:24:@40795.4]
  wire [31:0] x481_sum_1_io_result; // @[Math.scala 150:24:@40795.4]
  wire  RetimeWrapper_101_clock; // @[package.scala 93:22:@40805.4]
  wire  RetimeWrapper_101_reset; // @[package.scala 93:22:@40805.4]
  wire  RetimeWrapper_101_io_flow; // @[package.scala 93:22:@40805.4]
  wire  RetimeWrapper_101_io_in; // @[package.scala 93:22:@40805.4]
  wire  RetimeWrapper_101_io_out; // @[package.scala 93:22:@40805.4]
  wire  RetimeWrapper_102_clock; // @[package.scala 93:22:@40817.4]
  wire  RetimeWrapper_102_reset; // @[package.scala 93:22:@40817.4]
  wire  RetimeWrapper_102_io_flow; // @[package.scala 93:22:@40817.4]
  wire  RetimeWrapper_102_io_in; // @[package.scala 93:22:@40817.4]
  wire  RetimeWrapper_102_io_out; // @[package.scala 93:22:@40817.4]
  wire  RetimeWrapper_103_clock; // @[package.scala 93:22:@40840.4]
  wire  RetimeWrapper_103_reset; // @[package.scala 93:22:@40840.4]
  wire  RetimeWrapper_103_io_flow; // @[package.scala 93:22:@40840.4]
  wire [8:0] RetimeWrapper_103_io_in; // @[package.scala 93:22:@40840.4]
  wire [8:0] RetimeWrapper_103_io_out; // @[package.scala 93:22:@40840.4]
  wire  RetimeWrapper_104_clock; // @[package.scala 93:22:@40852.4]
  wire  RetimeWrapper_104_reset; // @[package.scala 93:22:@40852.4]
  wire  RetimeWrapper_104_io_flow; // @[package.scala 93:22:@40852.4]
  wire [8:0] RetimeWrapper_104_io_in; // @[package.scala 93:22:@40852.4]
  wire [8:0] RetimeWrapper_104_io_out; // @[package.scala 93:22:@40852.4]
  wire  RetimeWrapper_105_clock; // @[package.scala 93:22:@40864.4]
  wire  RetimeWrapper_105_reset; // @[package.scala 93:22:@40864.4]
  wire  RetimeWrapper_105_io_flow; // @[package.scala 93:22:@40864.4]
  wire [9:0] RetimeWrapper_105_io_in; // @[package.scala 93:22:@40864.4]
  wire [9:0] RetimeWrapper_105_io_out; // @[package.scala 93:22:@40864.4]
  wire  RetimeWrapper_106_clock; // @[package.scala 93:22:@40876.4]
  wire  RetimeWrapper_106_reset; // @[package.scala 93:22:@40876.4]
  wire  RetimeWrapper_106_io_flow; // @[package.scala 93:22:@40876.4]
  wire [8:0] RetimeWrapper_106_io_in; // @[package.scala 93:22:@40876.4]
  wire [8:0] RetimeWrapper_106_io_out; // @[package.scala 93:22:@40876.4]
  wire  RetimeWrapper_107_clock; // @[package.scala 93:22:@40888.4]
  wire  RetimeWrapper_107_reset; // @[package.scala 93:22:@40888.4]
  wire  RetimeWrapper_107_io_flow; // @[package.scala 93:22:@40888.4]
  wire [8:0] RetimeWrapper_107_io_in; // @[package.scala 93:22:@40888.4]
  wire [8:0] RetimeWrapper_107_io_out; // @[package.scala 93:22:@40888.4]
  wire  RetimeWrapper_108_clock; // @[package.scala 93:22:@40898.4]
  wire  RetimeWrapper_108_reset; // @[package.scala 93:22:@40898.4]
  wire  RetimeWrapper_108_io_flow; // @[package.scala 93:22:@40898.4]
  wire [7:0] RetimeWrapper_108_io_in; // @[package.scala 93:22:@40898.4]
  wire [7:0] RetimeWrapper_108_io_out; // @[package.scala 93:22:@40898.4]
  wire  RetimeWrapper_109_clock; // @[package.scala 93:22:@40907.4]
  wire  RetimeWrapper_109_reset; // @[package.scala 93:22:@40907.4]
  wire  RetimeWrapper_109_io_flow; // @[package.scala 93:22:@40907.4]
  wire [7:0] RetimeWrapper_109_io_in; // @[package.scala 93:22:@40907.4]
  wire [7:0] RetimeWrapper_109_io_out; // @[package.scala 93:22:@40907.4]
  wire [7:0] x489_x11_1_io_a; // @[Math.scala 150:24:@40916.4]
  wire [7:0] x489_x11_1_io_b; // @[Math.scala 150:24:@40916.4]
  wire [7:0] x489_x11_1_io_result; // @[Math.scala 150:24:@40916.4]
  wire  RetimeWrapper_110_clock; // @[package.scala 93:22:@40926.4]
  wire  RetimeWrapper_110_reset; // @[package.scala 93:22:@40926.4]
  wire  RetimeWrapper_110_io_flow; // @[package.scala 93:22:@40926.4]
  wire [7:0] RetimeWrapper_110_io_in; // @[package.scala 93:22:@40926.4]
  wire [7:0] RetimeWrapper_110_io_out; // @[package.scala 93:22:@40926.4]
  wire  RetimeWrapper_111_clock; // @[package.scala 93:22:@40935.4]
  wire  RetimeWrapper_111_reset; // @[package.scala 93:22:@40935.4]
  wire  RetimeWrapper_111_io_flow; // @[package.scala 93:22:@40935.4]
  wire [7:0] RetimeWrapper_111_io_in; // @[package.scala 93:22:@40935.4]
  wire [7:0] RetimeWrapper_111_io_out; // @[package.scala 93:22:@40935.4]
  wire [7:0] x490_x12_1_io_a; // @[Math.scala 150:24:@40944.4]
  wire [7:0] x490_x12_1_io_b; // @[Math.scala 150:24:@40944.4]
  wire [7:0] x490_x12_1_io_result; // @[Math.scala 150:24:@40944.4]
  wire [7:0] x491_x11_1_io_a; // @[Math.scala 150:24:@40954.4]
  wire [7:0] x491_x11_1_io_b; // @[Math.scala 150:24:@40954.4]
  wire [7:0] x491_x11_1_io_result; // @[Math.scala 150:24:@40954.4]
  wire  RetimeWrapper_112_clock; // @[package.scala 93:22:@40964.4]
  wire  RetimeWrapper_112_reset; // @[package.scala 93:22:@40964.4]
  wire  RetimeWrapper_112_io_flow; // @[package.scala 93:22:@40964.4]
  wire [7:0] RetimeWrapper_112_io_in; // @[package.scala 93:22:@40964.4]
  wire [7:0] RetimeWrapper_112_io_out; // @[package.scala 93:22:@40964.4]
  wire [7:0] x492_x12_1_io_a; // @[Math.scala 150:24:@40973.4]
  wire [7:0] x492_x12_1_io_b; // @[Math.scala 150:24:@40973.4]
  wire [7:0] x492_x12_1_io_result; // @[Math.scala 150:24:@40973.4]
  wire  RetimeWrapper_113_clock; // @[package.scala 93:22:@40983.4]
  wire  RetimeWrapper_113_reset; // @[package.scala 93:22:@40983.4]
  wire  RetimeWrapper_113_io_flow; // @[package.scala 93:22:@40983.4]
  wire [7:0] RetimeWrapper_113_io_in; // @[package.scala 93:22:@40983.4]
  wire [7:0] RetimeWrapper_113_io_out; // @[package.scala 93:22:@40983.4]
  wire  RetimeWrapper_114_clock; // @[package.scala 93:22:@40992.4]
  wire  RetimeWrapper_114_reset; // @[package.scala 93:22:@40992.4]
  wire  RetimeWrapper_114_io_flow; // @[package.scala 93:22:@40992.4]
  wire [7:0] RetimeWrapper_114_io_in; // @[package.scala 93:22:@40992.4]
  wire [7:0] RetimeWrapper_114_io_out; // @[package.scala 93:22:@40992.4]
  wire [7:0] x493_x11_1_io_a; // @[Math.scala 150:24:@41001.4]
  wire [7:0] x493_x11_1_io_b; // @[Math.scala 150:24:@41001.4]
  wire [7:0] x493_x11_1_io_result; // @[Math.scala 150:24:@41001.4]
  wire [7:0] x494_x12_1_io_a; // @[Math.scala 150:24:@41011.4]
  wire [7:0] x494_x12_1_io_b; // @[Math.scala 150:24:@41011.4]
  wire [7:0] x494_x12_1_io_result; // @[Math.scala 150:24:@41011.4]
  wire  RetimeWrapper_115_clock; // @[package.scala 93:22:@41021.4]
  wire  RetimeWrapper_115_reset; // @[package.scala 93:22:@41021.4]
  wire  RetimeWrapper_115_io_flow; // @[package.scala 93:22:@41021.4]
  wire [7:0] RetimeWrapper_115_io_in; // @[package.scala 93:22:@41021.4]
  wire [7:0] RetimeWrapper_115_io_out; // @[package.scala 93:22:@41021.4]
  wire [7:0] x495_x11_1_io_a; // @[Math.scala 150:24:@41032.4]
  wire [7:0] x495_x11_1_io_b; // @[Math.scala 150:24:@41032.4]
  wire [7:0] x495_x11_1_io_result; // @[Math.scala 150:24:@41032.4]
  wire  RetimeWrapper_116_clock; // @[package.scala 93:22:@41042.4]
  wire  RetimeWrapper_116_reset; // @[package.scala 93:22:@41042.4]
  wire  RetimeWrapper_116_io_flow; // @[package.scala 93:22:@41042.4]
  wire [7:0] RetimeWrapper_116_io_in; // @[package.scala 93:22:@41042.4]
  wire [7:0] RetimeWrapper_116_io_out; // @[package.scala 93:22:@41042.4]
  wire  x496_sum_1_clock; // @[Math.scala 150:24:@41051.4]
  wire  x496_sum_1_reset; // @[Math.scala 150:24:@41051.4]
  wire [7:0] x496_sum_1_io_a; // @[Math.scala 150:24:@41051.4]
  wire [7:0] x496_sum_1_io_b; // @[Math.scala 150:24:@41051.4]
  wire  x496_sum_1_io_flow; // @[Math.scala 150:24:@41051.4]
  wire [7:0] x496_sum_1_io_result; // @[Math.scala 150:24:@41051.4]
  wire  RetimeWrapper_117_clock; // @[package.scala 93:22:@41070.4]
  wire  RetimeWrapper_117_reset; // @[package.scala 93:22:@41070.4]
  wire  RetimeWrapper_117_io_flow; // @[package.scala 93:22:@41070.4]
  wire [8:0] RetimeWrapper_117_io_in; // @[package.scala 93:22:@41070.4]
  wire [8:0] RetimeWrapper_117_io_out; // @[package.scala 93:22:@41070.4]
  wire  RetimeWrapper_118_clock; // @[package.scala 93:22:@41082.4]
  wire  RetimeWrapper_118_reset; // @[package.scala 93:22:@41082.4]
  wire  RetimeWrapper_118_io_flow; // @[package.scala 93:22:@41082.4]
  wire [8:0] RetimeWrapper_118_io_in; // @[package.scala 93:22:@41082.4]
  wire [8:0] RetimeWrapper_118_io_out; // @[package.scala 93:22:@41082.4]
  wire  RetimeWrapper_119_clock; // @[package.scala 93:22:@41094.4]
  wire  RetimeWrapper_119_reset; // @[package.scala 93:22:@41094.4]
  wire  RetimeWrapper_119_io_flow; // @[package.scala 93:22:@41094.4]
  wire [9:0] RetimeWrapper_119_io_in; // @[package.scala 93:22:@41094.4]
  wire [9:0] RetimeWrapper_119_io_out; // @[package.scala 93:22:@41094.4]
  wire  RetimeWrapper_120_clock; // @[package.scala 93:22:@41106.4]
  wire  RetimeWrapper_120_reset; // @[package.scala 93:22:@41106.4]
  wire  RetimeWrapper_120_io_flow; // @[package.scala 93:22:@41106.4]
  wire [8:0] RetimeWrapper_120_io_in; // @[package.scala 93:22:@41106.4]
  wire [8:0] RetimeWrapper_120_io_out; // @[package.scala 93:22:@41106.4]
  wire  RetimeWrapper_121_clock; // @[package.scala 93:22:@41118.4]
  wire  RetimeWrapper_121_reset; // @[package.scala 93:22:@41118.4]
  wire  RetimeWrapper_121_io_flow; // @[package.scala 93:22:@41118.4]
  wire [8:0] RetimeWrapper_121_io_in; // @[package.scala 93:22:@41118.4]
  wire [8:0] RetimeWrapper_121_io_out; // @[package.scala 93:22:@41118.4]
  wire  RetimeWrapper_122_clock; // @[package.scala 93:22:@41128.4]
  wire  RetimeWrapper_122_reset; // @[package.scala 93:22:@41128.4]
  wire  RetimeWrapper_122_io_flow; // @[package.scala 93:22:@41128.4]
  wire [7:0] RetimeWrapper_122_io_in; // @[package.scala 93:22:@41128.4]
  wire [7:0] RetimeWrapper_122_io_out; // @[package.scala 93:22:@41128.4]
  wire  RetimeWrapper_123_clock; // @[package.scala 93:22:@41137.4]
  wire  RetimeWrapper_123_reset; // @[package.scala 93:22:@41137.4]
  wire  RetimeWrapper_123_io_flow; // @[package.scala 93:22:@41137.4]
  wire [7:0] RetimeWrapper_123_io_in; // @[package.scala 93:22:@41137.4]
  wire [7:0] RetimeWrapper_123_io_out; // @[package.scala 93:22:@41137.4]
  wire [7:0] x503_x11_1_io_a; // @[Math.scala 150:24:@41146.4]
  wire [7:0] x503_x11_1_io_b; // @[Math.scala 150:24:@41146.4]
  wire [7:0] x503_x11_1_io_result; // @[Math.scala 150:24:@41146.4]
  wire  RetimeWrapper_124_clock; // @[package.scala 93:22:@41156.4]
  wire  RetimeWrapper_124_reset; // @[package.scala 93:22:@41156.4]
  wire  RetimeWrapper_124_io_flow; // @[package.scala 93:22:@41156.4]
  wire [7:0] RetimeWrapper_124_io_in; // @[package.scala 93:22:@41156.4]
  wire [7:0] RetimeWrapper_124_io_out; // @[package.scala 93:22:@41156.4]
  wire  RetimeWrapper_125_clock; // @[package.scala 93:22:@41165.4]
  wire  RetimeWrapper_125_reset; // @[package.scala 93:22:@41165.4]
  wire  RetimeWrapper_125_io_flow; // @[package.scala 93:22:@41165.4]
  wire [7:0] RetimeWrapper_125_io_in; // @[package.scala 93:22:@41165.4]
  wire [7:0] RetimeWrapper_125_io_out; // @[package.scala 93:22:@41165.4]
  wire [7:0] x504_x12_1_io_a; // @[Math.scala 150:24:@41174.4]
  wire [7:0] x504_x12_1_io_b; // @[Math.scala 150:24:@41174.4]
  wire [7:0] x504_x12_1_io_result; // @[Math.scala 150:24:@41174.4]
  wire [7:0] x505_x11_1_io_a; // @[Math.scala 150:24:@41184.4]
  wire [7:0] x505_x11_1_io_b; // @[Math.scala 150:24:@41184.4]
  wire [7:0] x505_x11_1_io_result; // @[Math.scala 150:24:@41184.4]
  wire  RetimeWrapper_126_clock; // @[package.scala 93:22:@41194.4]
  wire  RetimeWrapper_126_reset; // @[package.scala 93:22:@41194.4]
  wire  RetimeWrapper_126_io_flow; // @[package.scala 93:22:@41194.4]
  wire [7:0] RetimeWrapper_126_io_in; // @[package.scala 93:22:@41194.4]
  wire [7:0] RetimeWrapper_126_io_out; // @[package.scala 93:22:@41194.4]
  wire [7:0] x506_x12_1_io_a; // @[Math.scala 150:24:@41203.4]
  wire [7:0] x506_x12_1_io_b; // @[Math.scala 150:24:@41203.4]
  wire [7:0] x506_x12_1_io_result; // @[Math.scala 150:24:@41203.4]
  wire  RetimeWrapper_127_clock; // @[package.scala 93:22:@41213.4]
  wire  RetimeWrapper_127_reset; // @[package.scala 93:22:@41213.4]
  wire  RetimeWrapper_127_io_flow; // @[package.scala 93:22:@41213.4]
  wire [7:0] RetimeWrapper_127_io_in; // @[package.scala 93:22:@41213.4]
  wire [7:0] RetimeWrapper_127_io_out; // @[package.scala 93:22:@41213.4]
  wire  RetimeWrapper_128_clock; // @[package.scala 93:22:@41222.4]
  wire  RetimeWrapper_128_reset; // @[package.scala 93:22:@41222.4]
  wire  RetimeWrapper_128_io_flow; // @[package.scala 93:22:@41222.4]
  wire [7:0] RetimeWrapper_128_io_in; // @[package.scala 93:22:@41222.4]
  wire [7:0] RetimeWrapper_128_io_out; // @[package.scala 93:22:@41222.4]
  wire [7:0] x507_x11_1_io_a; // @[Math.scala 150:24:@41231.4]
  wire [7:0] x507_x11_1_io_b; // @[Math.scala 150:24:@41231.4]
  wire [7:0] x507_x11_1_io_result; // @[Math.scala 150:24:@41231.4]
  wire [7:0] x508_x12_1_io_a; // @[Math.scala 150:24:@41241.4]
  wire [7:0] x508_x12_1_io_b; // @[Math.scala 150:24:@41241.4]
  wire [7:0] x508_x12_1_io_result; // @[Math.scala 150:24:@41241.4]
  wire  RetimeWrapper_129_clock; // @[package.scala 93:22:@41251.4]
  wire  RetimeWrapper_129_reset; // @[package.scala 93:22:@41251.4]
  wire  RetimeWrapper_129_io_flow; // @[package.scala 93:22:@41251.4]
  wire [7:0] RetimeWrapper_129_io_in; // @[package.scala 93:22:@41251.4]
  wire [7:0] RetimeWrapper_129_io_out; // @[package.scala 93:22:@41251.4]
  wire [7:0] x509_x11_1_io_a; // @[Math.scala 150:24:@41260.4]
  wire [7:0] x509_x11_1_io_b; // @[Math.scala 150:24:@41260.4]
  wire [7:0] x509_x11_1_io_result; // @[Math.scala 150:24:@41260.4]
  wire  RetimeWrapper_130_clock; // @[package.scala 93:22:@41270.4]
  wire  RetimeWrapper_130_reset; // @[package.scala 93:22:@41270.4]
  wire  RetimeWrapper_130_io_flow; // @[package.scala 93:22:@41270.4]
  wire [7:0] RetimeWrapper_130_io_in; // @[package.scala 93:22:@41270.4]
  wire [7:0] RetimeWrapper_130_io_out; // @[package.scala 93:22:@41270.4]
  wire  x510_sum_1_clock; // @[Math.scala 150:24:@41279.4]
  wire  x510_sum_1_reset; // @[Math.scala 150:24:@41279.4]
  wire [7:0] x510_sum_1_io_a; // @[Math.scala 150:24:@41279.4]
  wire [7:0] x510_sum_1_io_b; // @[Math.scala 150:24:@41279.4]
  wire  x510_sum_1_io_flow; // @[Math.scala 150:24:@41279.4]
  wire [7:0] x510_sum_1_io_result; // @[Math.scala 150:24:@41279.4]
  wire  RetimeWrapper_131_clock; // @[package.scala 93:22:@41298.4]
  wire  RetimeWrapper_131_reset; // @[package.scala 93:22:@41298.4]
  wire  RetimeWrapper_131_io_flow; // @[package.scala 93:22:@41298.4]
  wire [8:0] RetimeWrapper_131_io_in; // @[package.scala 93:22:@41298.4]
  wire [8:0] RetimeWrapper_131_io_out; // @[package.scala 93:22:@41298.4]
  wire  RetimeWrapper_132_clock; // @[package.scala 93:22:@41310.4]
  wire  RetimeWrapper_132_reset; // @[package.scala 93:22:@41310.4]
  wire  RetimeWrapper_132_io_flow; // @[package.scala 93:22:@41310.4]
  wire [9:0] RetimeWrapper_132_io_in; // @[package.scala 93:22:@41310.4]
  wire [9:0] RetimeWrapper_132_io_out; // @[package.scala 93:22:@41310.4]
  wire  RetimeWrapper_133_clock; // @[package.scala 93:22:@41322.4]
  wire  RetimeWrapper_133_reset; // @[package.scala 93:22:@41322.4]
  wire  RetimeWrapper_133_io_flow; // @[package.scala 93:22:@41322.4]
  wire [8:0] RetimeWrapper_133_io_in; // @[package.scala 93:22:@41322.4]
  wire [8:0] RetimeWrapper_133_io_out; // @[package.scala 93:22:@41322.4]
  wire  RetimeWrapper_134_clock; // @[package.scala 93:22:@41334.4]
  wire  RetimeWrapper_134_reset; // @[package.scala 93:22:@41334.4]
  wire  RetimeWrapper_134_io_flow; // @[package.scala 93:22:@41334.4]
  wire [8:0] RetimeWrapper_134_io_in; // @[package.scala 93:22:@41334.4]
  wire [8:0] RetimeWrapper_134_io_out; // @[package.scala 93:22:@41334.4]
  wire  RetimeWrapper_135_clock; // @[package.scala 93:22:@41344.4]
  wire  RetimeWrapper_135_reset; // @[package.scala 93:22:@41344.4]
  wire  RetimeWrapper_135_io_flow; // @[package.scala 93:22:@41344.4]
  wire [7:0] RetimeWrapper_135_io_in; // @[package.scala 93:22:@41344.4]
  wire [7:0] RetimeWrapper_135_io_out; // @[package.scala 93:22:@41344.4]
  wire [7:0] x516_x11_1_io_a; // @[Math.scala 150:24:@41353.4]
  wire [7:0] x516_x11_1_io_b; // @[Math.scala 150:24:@41353.4]
  wire [7:0] x516_x11_1_io_result; // @[Math.scala 150:24:@41353.4]
  wire  RetimeWrapper_136_clock; // @[package.scala 93:22:@41363.4]
  wire  RetimeWrapper_136_reset; // @[package.scala 93:22:@41363.4]
  wire  RetimeWrapper_136_io_flow; // @[package.scala 93:22:@41363.4]
  wire [7:0] RetimeWrapper_136_io_in; // @[package.scala 93:22:@41363.4]
  wire [7:0] RetimeWrapper_136_io_out; // @[package.scala 93:22:@41363.4]
  wire  RetimeWrapper_137_clock; // @[package.scala 93:22:@41372.4]
  wire  RetimeWrapper_137_reset; // @[package.scala 93:22:@41372.4]
  wire  RetimeWrapper_137_io_flow; // @[package.scala 93:22:@41372.4]
  wire [7:0] RetimeWrapper_137_io_in; // @[package.scala 93:22:@41372.4]
  wire [7:0] RetimeWrapper_137_io_out; // @[package.scala 93:22:@41372.4]
  wire [7:0] x517_x12_1_io_a; // @[Math.scala 150:24:@41381.4]
  wire [7:0] x517_x12_1_io_b; // @[Math.scala 150:24:@41381.4]
  wire [7:0] x517_x12_1_io_result; // @[Math.scala 150:24:@41381.4]
  wire [7:0] x518_x11_1_io_a; // @[Math.scala 150:24:@41391.4]
  wire [7:0] x518_x11_1_io_b; // @[Math.scala 150:24:@41391.4]
  wire [7:0] x518_x11_1_io_result; // @[Math.scala 150:24:@41391.4]
  wire  RetimeWrapper_138_clock; // @[package.scala 93:22:@41401.4]
  wire  RetimeWrapper_138_reset; // @[package.scala 93:22:@41401.4]
  wire  RetimeWrapper_138_io_flow; // @[package.scala 93:22:@41401.4]
  wire [7:0] RetimeWrapper_138_io_in; // @[package.scala 93:22:@41401.4]
  wire [7:0] RetimeWrapper_138_io_out; // @[package.scala 93:22:@41401.4]
  wire [7:0] x519_x12_1_io_a; // @[Math.scala 150:24:@41410.4]
  wire [7:0] x519_x12_1_io_b; // @[Math.scala 150:24:@41410.4]
  wire [7:0] x519_x12_1_io_result; // @[Math.scala 150:24:@41410.4]
  wire  RetimeWrapper_139_clock; // @[package.scala 93:22:@41420.4]
  wire  RetimeWrapper_139_reset; // @[package.scala 93:22:@41420.4]
  wire  RetimeWrapper_139_io_flow; // @[package.scala 93:22:@41420.4]
  wire [7:0] RetimeWrapper_139_io_in; // @[package.scala 93:22:@41420.4]
  wire [7:0] RetimeWrapper_139_io_out; // @[package.scala 93:22:@41420.4]
  wire  RetimeWrapper_140_clock; // @[package.scala 93:22:@41429.4]
  wire  RetimeWrapper_140_reset; // @[package.scala 93:22:@41429.4]
  wire  RetimeWrapper_140_io_flow; // @[package.scala 93:22:@41429.4]
  wire [7:0] RetimeWrapper_140_io_in; // @[package.scala 93:22:@41429.4]
  wire [7:0] RetimeWrapper_140_io_out; // @[package.scala 93:22:@41429.4]
  wire [7:0] x520_x11_1_io_a; // @[Math.scala 150:24:@41438.4]
  wire [7:0] x520_x11_1_io_b; // @[Math.scala 150:24:@41438.4]
  wire [7:0] x520_x11_1_io_result; // @[Math.scala 150:24:@41438.4]
  wire [7:0] x521_x12_1_io_a; // @[Math.scala 150:24:@41448.4]
  wire [7:0] x521_x12_1_io_b; // @[Math.scala 150:24:@41448.4]
  wire [7:0] x521_x12_1_io_result; // @[Math.scala 150:24:@41448.4]
  wire  RetimeWrapper_141_clock; // @[package.scala 93:22:@41458.4]
  wire  RetimeWrapper_141_reset; // @[package.scala 93:22:@41458.4]
  wire  RetimeWrapper_141_io_flow; // @[package.scala 93:22:@41458.4]
  wire [7:0] RetimeWrapper_141_io_in; // @[package.scala 93:22:@41458.4]
  wire [7:0] RetimeWrapper_141_io_out; // @[package.scala 93:22:@41458.4]
  wire [7:0] x522_x11_1_io_a; // @[Math.scala 150:24:@41467.4]
  wire [7:0] x522_x11_1_io_b; // @[Math.scala 150:24:@41467.4]
  wire [7:0] x522_x11_1_io_result; // @[Math.scala 150:24:@41467.4]
  wire  RetimeWrapper_142_clock; // @[package.scala 93:22:@41477.4]
  wire  RetimeWrapper_142_reset; // @[package.scala 93:22:@41477.4]
  wire  RetimeWrapper_142_io_flow; // @[package.scala 93:22:@41477.4]
  wire [7:0] RetimeWrapper_142_io_in; // @[package.scala 93:22:@41477.4]
  wire [7:0] RetimeWrapper_142_io_out; // @[package.scala 93:22:@41477.4]
  wire  x523_sum_1_clock; // @[Math.scala 150:24:@41486.4]
  wire  x523_sum_1_reset; // @[Math.scala 150:24:@41486.4]
  wire [7:0] x523_sum_1_io_a; // @[Math.scala 150:24:@41486.4]
  wire [7:0] x523_sum_1_io_b; // @[Math.scala 150:24:@41486.4]
  wire  x523_sum_1_io_flow; // @[Math.scala 150:24:@41486.4]
  wire [7:0] x523_sum_1_io_result; // @[Math.scala 150:24:@41486.4]
  wire  RetimeWrapper_143_clock; // @[package.scala 93:22:@41507.4]
  wire  RetimeWrapper_143_reset; // @[package.scala 93:22:@41507.4]
  wire  RetimeWrapper_143_io_flow; // @[package.scala 93:22:@41507.4]
  wire [8:0] RetimeWrapper_143_io_in; // @[package.scala 93:22:@41507.4]
  wire [8:0] RetimeWrapper_143_io_out; // @[package.scala 93:22:@41507.4]
  wire  RetimeWrapper_144_clock; // @[package.scala 93:22:@41519.4]
  wire  RetimeWrapper_144_reset; // @[package.scala 93:22:@41519.4]
  wire  RetimeWrapper_144_io_flow; // @[package.scala 93:22:@41519.4]
  wire [9:0] RetimeWrapper_144_io_in; // @[package.scala 93:22:@41519.4]
  wire [9:0] RetimeWrapper_144_io_out; // @[package.scala 93:22:@41519.4]
  wire  RetimeWrapper_145_clock; // @[package.scala 93:22:@41531.4]
  wire  RetimeWrapper_145_reset; // @[package.scala 93:22:@41531.4]
  wire  RetimeWrapper_145_io_flow; // @[package.scala 93:22:@41531.4]
  wire [8:0] RetimeWrapper_145_io_in; // @[package.scala 93:22:@41531.4]
  wire [8:0] RetimeWrapper_145_io_out; // @[package.scala 93:22:@41531.4]
  wire  RetimeWrapper_146_clock; // @[package.scala 93:22:@41543.4]
  wire  RetimeWrapper_146_reset; // @[package.scala 93:22:@41543.4]
  wire  RetimeWrapper_146_io_flow; // @[package.scala 93:22:@41543.4]
  wire [8:0] RetimeWrapper_146_io_in; // @[package.scala 93:22:@41543.4]
  wire [8:0] RetimeWrapper_146_io_out; // @[package.scala 93:22:@41543.4]
  wire  RetimeWrapper_147_clock; // @[package.scala 93:22:@41553.4]
  wire  RetimeWrapper_147_reset; // @[package.scala 93:22:@41553.4]
  wire  RetimeWrapper_147_io_flow; // @[package.scala 93:22:@41553.4]
  wire [7:0] RetimeWrapper_147_io_in; // @[package.scala 93:22:@41553.4]
  wire [7:0] RetimeWrapper_147_io_out; // @[package.scala 93:22:@41553.4]
  wire [7:0] x529_x11_1_io_a; // @[Math.scala 150:24:@41562.4]
  wire [7:0] x529_x11_1_io_b; // @[Math.scala 150:24:@41562.4]
  wire [7:0] x529_x11_1_io_result; // @[Math.scala 150:24:@41562.4]
  wire  RetimeWrapper_148_clock; // @[package.scala 93:22:@41572.4]
  wire  RetimeWrapper_148_reset; // @[package.scala 93:22:@41572.4]
  wire  RetimeWrapper_148_io_flow; // @[package.scala 93:22:@41572.4]
  wire [7:0] RetimeWrapper_148_io_in; // @[package.scala 93:22:@41572.4]
  wire [7:0] RetimeWrapper_148_io_out; // @[package.scala 93:22:@41572.4]
  wire  RetimeWrapper_149_clock; // @[package.scala 93:22:@41581.4]
  wire  RetimeWrapper_149_reset; // @[package.scala 93:22:@41581.4]
  wire  RetimeWrapper_149_io_flow; // @[package.scala 93:22:@41581.4]
  wire [7:0] RetimeWrapper_149_io_in; // @[package.scala 93:22:@41581.4]
  wire [7:0] RetimeWrapper_149_io_out; // @[package.scala 93:22:@41581.4]
  wire [7:0] x530_x12_1_io_a; // @[Math.scala 150:24:@41590.4]
  wire [7:0] x530_x12_1_io_b; // @[Math.scala 150:24:@41590.4]
  wire [7:0] x530_x12_1_io_result; // @[Math.scala 150:24:@41590.4]
  wire [7:0] x531_x11_1_io_a; // @[Math.scala 150:24:@41600.4]
  wire [7:0] x531_x11_1_io_b; // @[Math.scala 150:24:@41600.4]
  wire [7:0] x531_x11_1_io_result; // @[Math.scala 150:24:@41600.4]
  wire  RetimeWrapper_150_clock; // @[package.scala 93:22:@41610.4]
  wire  RetimeWrapper_150_reset; // @[package.scala 93:22:@41610.4]
  wire  RetimeWrapper_150_io_flow; // @[package.scala 93:22:@41610.4]
  wire [7:0] RetimeWrapper_150_io_in; // @[package.scala 93:22:@41610.4]
  wire [7:0] RetimeWrapper_150_io_out; // @[package.scala 93:22:@41610.4]
  wire [7:0] x532_x12_1_io_a; // @[Math.scala 150:24:@41619.4]
  wire [7:0] x532_x12_1_io_b; // @[Math.scala 150:24:@41619.4]
  wire [7:0] x532_x12_1_io_result; // @[Math.scala 150:24:@41619.4]
  wire  RetimeWrapper_151_clock; // @[package.scala 93:22:@41629.4]
  wire  RetimeWrapper_151_reset; // @[package.scala 93:22:@41629.4]
  wire  RetimeWrapper_151_io_flow; // @[package.scala 93:22:@41629.4]
  wire [7:0] RetimeWrapper_151_io_in; // @[package.scala 93:22:@41629.4]
  wire [7:0] RetimeWrapper_151_io_out; // @[package.scala 93:22:@41629.4]
  wire  RetimeWrapper_152_clock; // @[package.scala 93:22:@41638.4]
  wire  RetimeWrapper_152_reset; // @[package.scala 93:22:@41638.4]
  wire  RetimeWrapper_152_io_flow; // @[package.scala 93:22:@41638.4]
  wire [7:0] RetimeWrapper_152_io_in; // @[package.scala 93:22:@41638.4]
  wire [7:0] RetimeWrapper_152_io_out; // @[package.scala 93:22:@41638.4]
  wire [7:0] x533_x11_1_io_a; // @[Math.scala 150:24:@41647.4]
  wire [7:0] x533_x11_1_io_b; // @[Math.scala 150:24:@41647.4]
  wire [7:0] x533_x11_1_io_result; // @[Math.scala 150:24:@41647.4]
  wire [7:0] x534_x12_1_io_a; // @[Math.scala 150:24:@41657.4]
  wire [7:0] x534_x12_1_io_b; // @[Math.scala 150:24:@41657.4]
  wire [7:0] x534_x12_1_io_result; // @[Math.scala 150:24:@41657.4]
  wire  RetimeWrapper_153_clock; // @[package.scala 93:22:@41667.4]
  wire  RetimeWrapper_153_reset; // @[package.scala 93:22:@41667.4]
  wire  RetimeWrapper_153_io_flow; // @[package.scala 93:22:@41667.4]
  wire [7:0] RetimeWrapper_153_io_in; // @[package.scala 93:22:@41667.4]
  wire [7:0] RetimeWrapper_153_io_out; // @[package.scala 93:22:@41667.4]
  wire [7:0] x535_x11_1_io_a; // @[Math.scala 150:24:@41676.4]
  wire [7:0] x535_x11_1_io_b; // @[Math.scala 150:24:@41676.4]
  wire [7:0] x535_x11_1_io_result; // @[Math.scala 150:24:@41676.4]
  wire  RetimeWrapper_154_clock; // @[package.scala 93:22:@41686.4]
  wire  RetimeWrapper_154_reset; // @[package.scala 93:22:@41686.4]
  wire  RetimeWrapper_154_io_flow; // @[package.scala 93:22:@41686.4]
  wire [7:0] RetimeWrapper_154_io_in; // @[package.scala 93:22:@41686.4]
  wire [7:0] RetimeWrapper_154_io_out; // @[package.scala 93:22:@41686.4]
  wire  x536_sum_1_clock; // @[Math.scala 150:24:@41695.4]
  wire  x536_sum_1_reset; // @[Math.scala 150:24:@41695.4]
  wire [7:0] x536_sum_1_io_a; // @[Math.scala 150:24:@41695.4]
  wire [7:0] x536_sum_1_io_b; // @[Math.scala 150:24:@41695.4]
  wire  x536_sum_1_io_flow; // @[Math.scala 150:24:@41695.4]
  wire [7:0] x536_sum_1_io_result; // @[Math.scala 150:24:@41695.4]
  wire  RetimeWrapper_155_clock; // @[package.scala 93:22:@41712.4]
  wire  RetimeWrapper_155_reset; // @[package.scala 93:22:@41712.4]
  wire  RetimeWrapper_155_io_flow; // @[package.scala 93:22:@41712.4]
  wire [7:0] RetimeWrapper_155_io_in; // @[package.scala 93:22:@41712.4]
  wire [7:0] RetimeWrapper_155_io_out; // @[package.scala 93:22:@41712.4]
  wire  RetimeWrapper_156_clock; // @[package.scala 93:22:@41721.4]
  wire  RetimeWrapper_156_reset; // @[package.scala 93:22:@41721.4]
  wire  RetimeWrapper_156_io_flow; // @[package.scala 93:22:@41721.4]
  wire [7:0] RetimeWrapper_156_io_in; // @[package.scala 93:22:@41721.4]
  wire [7:0] RetimeWrapper_156_io_out; // @[package.scala 93:22:@41721.4]
  wire  RetimeWrapper_157_clock; // @[package.scala 93:22:@41730.4]
  wire  RetimeWrapper_157_reset; // @[package.scala 93:22:@41730.4]
  wire  RetimeWrapper_157_io_flow; // @[package.scala 93:22:@41730.4]
  wire [7:0] RetimeWrapper_157_io_in; // @[package.scala 93:22:@41730.4]
  wire [7:0] RetimeWrapper_157_io_out; // @[package.scala 93:22:@41730.4]
  wire  RetimeWrapper_158_clock; // @[package.scala 93:22:@41739.4]
  wire  RetimeWrapper_158_reset; // @[package.scala 93:22:@41739.4]
  wire  RetimeWrapper_158_io_flow; // @[package.scala 93:22:@41739.4]
  wire [7:0] RetimeWrapper_158_io_in; // @[package.scala 93:22:@41739.4]
  wire [7:0] RetimeWrapper_158_io_out; // @[package.scala 93:22:@41739.4]
  wire  RetimeWrapper_159_clock; // @[package.scala 93:22:@41758.4]
  wire  RetimeWrapper_159_reset; // @[package.scala 93:22:@41758.4]
  wire  RetimeWrapper_159_io_flow; // @[package.scala 93:22:@41758.4]
  wire [31:0] RetimeWrapper_159_io_in; // @[package.scala 93:22:@41758.4]
  wire [31:0] RetimeWrapper_159_io_out; // @[package.scala 93:22:@41758.4]
  wire  RetimeWrapper_160_clock; // @[package.scala 93:22:@41767.4]
  wire  RetimeWrapper_160_reset; // @[package.scala 93:22:@41767.4]
  wire  RetimeWrapper_160_io_flow; // @[package.scala 93:22:@41767.4]
  wire  RetimeWrapper_160_io_in; // @[package.scala 93:22:@41767.4]
  wire  RetimeWrapper_160_io_out; // @[package.scala 93:22:@41767.4]
  wire  RetimeWrapper_161_clock; // @[package.scala 93:22:@41776.4]
  wire  RetimeWrapper_161_reset; // @[package.scala 93:22:@41776.4]
  wire  RetimeWrapper_161_io_flow; // @[package.scala 93:22:@41776.4]
  wire  RetimeWrapper_161_io_in; // @[package.scala 93:22:@41776.4]
  wire  RetimeWrapper_161_io_out; // @[package.scala 93:22:@41776.4]
  wire  RetimeWrapper_162_clock; // @[package.scala 93:22:@41785.4]
  wire  RetimeWrapper_162_reset; // @[package.scala 93:22:@41785.4]
  wire  RetimeWrapper_162_io_flow; // @[package.scala 93:22:@41785.4]
  wire  RetimeWrapper_162_io_in; // @[package.scala 93:22:@41785.4]
  wire  RetimeWrapper_162_io_out; // @[package.scala 93:22:@41785.4]
  wire  b327; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 62:18:@38584.4]
  wire  b328; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 63:18:@38585.4]
  wire  _T_206; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 68:30:@38732.4]
  wire  _T_207; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 68:37:@38733.4]
  wire  _T_211; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 70:76:@38738.4]
  wire  _T_212; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 70:62:@38739.4]
  wire  _T_214; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 70:101:@38740.4]
  wire [31:0] x614_x330_D1_0_number; // @[package.scala 96:25:@38749.4 package.scala 96:25:@38750.4]
  wire [31:0] b325_number; // @[Math.scala 712:22:@38569.4 Math.scala 713:14:@38570.4]
  wire [31:0] _T_246; // @[Math.scala 499:52:@38769.4]
  wire  x334; // @[Math.scala 499:44:@38777.4]
  wire  x335; // @[Math.scala 499:44:@38784.4]
  wire  x336; // @[Math.scala 499:44:@38791.4]
  wire [31:0] _T_293; // @[Mux.scala 19:72:@38803.4]
  wire [31:0] _T_295; // @[Mux.scala 19:72:@38804.4]
  wire [31:0] _T_297; // @[Mux.scala 19:72:@38805.4]
  wire [31:0] _T_299; // @[Mux.scala 19:72:@38807.4]
  wire [31:0] x337_number; // @[Mux.scala 19:72:@38808.4]
  wire [31:0] _T_311; // @[Math.scala 406:49:@38818.4]
  wire [31:0] _T_313; // @[Math.scala 406:56:@38820.4]
  wire [31:0] _T_314; // @[Math.scala 406:56:@38821.4]
  wire  _T_326; // @[FixedPoint.scala 50:25:@38839.4]
  wire [1:0] _T_330; // @[Bitwise.scala 72:12:@38841.4]
  wire [29:0] _T_331; // @[FixedPoint.scala 18:52:@38842.4]
  wire  _T_372; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 121:101:@38943.4]
  wire  _T_376; // @[package.scala 96:25:@38951.4 package.scala 96:25:@38952.4]
  wire  _T_378; // @[implicits.scala 55:10:@38953.4]
  wire  _T_379; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 121:118:@38954.4]
  wire  _T_381; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 121:207:@38956.4]
  wire  _T_382; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 121:226:@38957.4]
  wire  x620_b327_D24; // @[package.scala 96:25:@38931.4 package.scala 96:25:@38932.4]
  wire  _T_383; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 121:252:@38958.4]
  wire  x619_b328_D24; // @[package.scala 96:25:@38922.4 package.scala 96:25:@38923.4]
  wire  _T_427; // @[package.scala 96:25:@39058.4 package.scala 96:25:@39059.4]
  wire  _T_429; // @[implicits.scala 55:10:@39060.4]
  wire  _T_430; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 144:118:@39061.4]
  wire  _T_432; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 144:207:@39063.4]
  wire  _T_433; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 144:226:@39064.4]
  wire  _T_434; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 144:252:@39065.4]
  wire  _T_475; // @[package.scala 96:25:@39156.4 package.scala 96:25:@39157.4]
  wire  _T_477; // @[implicits.scala 55:10:@39158.4]
  wire  _T_478; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 165:118:@39159.4]
  wire  _T_480; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 165:207:@39161.4]
  wire  _T_481; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 165:226:@39162.4]
  wire  _T_482; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 165:252:@39163.4]
  wire  _T_523; // @[package.scala 96:25:@39254.4 package.scala 96:25:@39255.4]
  wire  _T_525; // @[implicits.scala 55:10:@39256.4]
  wire  _T_526; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 192:166:@39257.4]
  wire  _T_528; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 192:255:@39259.4]
  wire  _T_529; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 192:274:@39260.4]
  wire  _T_530; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 192:300:@39261.4]
  wire [31:0] x632_b325_D26_number; // @[package.scala 96:25:@39275.4 package.scala 96:25:@39276.4]
  wire [31:0] _T_549; // @[Math.scala 465:37:@39295.4]
  wire [31:0] x633_x358_rdcol_D26_number; // @[package.scala 96:25:@39312.4 package.scala 96:25:@39313.4]
  wire [31:0] _T_562; // @[Math.scala 465:37:@39318.4]
  wire  x634_x366_D1; // @[package.scala 96:25:@39335.4 package.scala 96:25:@39336.4]
  wire  x367; // @[package.scala 96:25:@39326.4 package.scala 96:25:@39327.4]
  wire  x368; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 209:24:@39339.4]
  wire [31:0] x365_number; // @[Math.scala 370:22:@39289.4 Math.scala 371:14:@39290.4]
  wire [31:0] _T_581; // @[Math.scala 406:49:@39348.4]
  wire [31:0] _T_583; // @[Math.scala 406:56:@39350.4]
  wire [31:0] _T_584; // @[Math.scala 406:56:@39351.4]
  wire  _T_589; // @[FixedPoint.scala 50:25:@39357.4]
  wire [1:0] _T_593; // @[Bitwise.scala 72:12:@39359.4]
  wire [29:0] _T_594; // @[FixedPoint.scala 18:52:@39360.4]
  wire  _T_638; // @[package.scala 96:25:@39458.4 package.scala 96:25:@39459.4]
  wire  _T_640; // @[implicits.scala 55:10:@39460.4]
  wire  _T_641; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 238:194:@39461.4]
  wire  x641_x369_D22; // @[package.scala 96:25:@39446.4 package.scala 96:25:@39447.4]
  wire  _T_642; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 238:283:@39462.4]
  wire  x639_b327_D50; // @[package.scala 96:25:@39428.4 package.scala 96:25:@39429.4]
  wire  _T_643; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 238:291:@39463.4]
  wire  x636_b328_D50; // @[package.scala 96:25:@39401.4 package.scala 96:25:@39402.4]
  wire [31:0] x642_x352_rdcol_D26_number; // @[package.scala 96:25:@39479.4 package.scala 96:25:@39480.4]
  wire [31:0] _T_654; // @[Math.scala 465:37:@39485.4]
  wire  x376; // @[package.scala 96:25:@39493.4 package.scala 96:25:@39494.4]
  wire  x377; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 246:24:@39497.4]
  wire  _T_689; // @[package.scala 96:25:@39557.4 package.scala 96:25:@39558.4]
  wire  _T_691; // @[implicits.scala 55:10:@39559.4]
  wire  _T_692; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 263:194:@39560.4]
  wire  x645_x378_D22; // @[package.scala 96:25:@39536.4 package.scala 96:25:@39537.4]
  wire  _T_693; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 263:283:@39561.4]
  wire  _T_694; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 263:291:@39562.4]
  wire [31:0] x647_x346_rdcol_D26_number; // @[package.scala 96:25:@39578.4 package.scala 96:25:@39579.4]
  wire [31:0] _T_705; // @[Math.scala 465:37:@39584.4]
  wire  x382; // @[package.scala 96:25:@39592.4 package.scala 96:25:@39593.4]
  wire  x383; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 271:24:@39596.4]
  wire  _T_740; // @[package.scala 96:25:@39656.4 package.scala 96:25:@39657.4]
  wire  _T_742; // @[implicits.scala 55:10:@39658.4]
  wire  _T_743; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 288:194:@39659.4]
  wire  x650_x384_D22; // @[package.scala 96:25:@39635.4 package.scala 96:25:@39636.4]
  wire  _T_744; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 288:283:@39660.4]
  wire  _T_745; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 288:291:@39661.4]
  wire [31:0] x652_b326_D26_number; // @[package.scala 96:25:@39677.4 package.scala 96:25:@39678.4]
  wire [31:0] _T_758; // @[Math.scala 465:37:@39685.4]
  wire  x366; // @[package.scala 96:25:@39303.4 package.scala 96:25:@39304.4]
  wire  x388; // @[package.scala 96:25:@39693.4 package.scala 96:25:@39694.4]
  wire  x389; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 304:59:@39697.4]
  wire  _T_793; // @[package.scala 96:25:@39757.4 package.scala 96:25:@39758.4]
  wire  _T_795; // @[implicits.scala 55:10:@39759.4]
  wire  _T_796; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 321:194:@39760.4]
  wire  x656_x390_D23; // @[package.scala 96:25:@39745.4 package.scala 96:25:@39746.4]
  wire  _T_797; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 321:283:@39761.4]
  wire  _T_798; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 321:291:@39762.4]
  wire [31:0] x394_rdcol_number; // @[Math.scala 154:22:@39781.4 Math.scala 155:14:@39782.4]
  wire [31:0] _T_813; // @[Math.scala 465:37:@39787.4]
  wire  x395; // @[package.scala 96:25:@39795.4 package.scala 96:25:@39796.4]
  wire  x396; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 329:59:@39799.4]
  wire  _T_862; // @[package.scala 96:25:@39883.4 package.scala 96:25:@39884.4]
  wire  _T_864; // @[implicits.scala 55:10:@39885.4]
  wire  _T_865; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 350:194:@39886.4]
  wire  x658_x397_D22; // @[package.scala 96:25:@39853.4 package.scala 96:25:@39854.4]
  wire  _T_866; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 350:283:@39887.4]
  wire  _T_867; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 350:291:@39888.4]
  wire [31:0] x403_rdcol_number; // @[Math.scala 154:22:@39907.4 Math.scala 155:14:@39908.4]
  wire [31:0] _T_882; // @[Math.scala 465:37:@39913.4]
  wire  x404; // @[package.scala 96:25:@39921.4 package.scala 96:25:@39922.4]
  wire  x405; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 358:59:@39925.4]
  wire  _T_931; // @[package.scala 96:25:@40009.4 package.scala 96:25:@40010.4]
  wire  _T_933; // @[implicits.scala 55:10:@40011.4]
  wire  _T_934; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 379:194:@40012.4]
  wire  x663_x406_D22; // @[package.scala 96:25:@39988.4 package.scala 96:25:@39989.4]
  wire  _T_935; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 379:283:@40013.4]
  wire  _T_936; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 379:291:@40014.4]
  wire [31:0] x412_rdrow_number; // @[Math.scala 195:22:@40033.4 Math.scala 196:14:@40034.4]
  wire [31:0] _T_958; // @[Math.scala 465:37:@40051.4]
  wire  x414; // @[package.scala 96:25:@40059.4 package.scala 96:25:@40060.4]
  wire  x415; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 389:24:@40063.4]
  wire [31:0] x413_number; // @[Math.scala 370:22:@40045.4 Math.scala 371:14:@40046.4]
  wire [31:0] _T_974; // @[Math.scala 406:49:@40072.4]
  wire [31:0] _T_976; // @[Math.scala 406:56:@40074.4]
  wire [31:0] _T_977; // @[Math.scala 406:56:@40075.4]
  wire  _T_982; // @[FixedPoint.scala 50:25:@40081.4]
  wire [1:0] _T_986; // @[Bitwise.scala 72:12:@40083.4]
  wire [29:0] _T_987; // @[FixedPoint.scala 18:52:@40084.4]
  wire  _T_1019; // @[package.scala 96:25:@40146.4 package.scala 96:25:@40147.4]
  wire  _T_1021; // @[implicits.scala 55:10:@40148.4]
  wire  _T_1022; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 410:194:@40149.4]
  wire  x666_x416_D22; // @[package.scala 96:25:@40125.4 package.scala 96:25:@40126.4]
  wire  _T_1023; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 410:283:@40150.4]
  wire  _T_1024; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 410:291:@40151.4]
  wire  x423; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 420:59:@40162.4]
  wire  _T_1053; // @[package.scala 96:25:@40206.4 package.scala 96:25:@40207.4]
  wire  _T_1055; // @[implicits.scala 55:10:@40208.4]
  wire  _T_1056; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 435:194:@40209.4]
  wire  x669_x424_D22; // @[package.scala 96:25:@40194.4 package.scala 96:25:@40195.4]
  wire  _T_1057; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 435:283:@40210.4]
  wire  _T_1058; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 435:291:@40211.4]
  wire  x428; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 439:59:@40222.4]
  wire  _T_1085; // @[package.scala 96:25:@40264.4 package.scala 96:25:@40265.4]
  wire  _T_1087; // @[implicits.scala 55:10:@40266.4]
  wire  _T_1088; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 452:194:@40267.4]
  wire  x671_x429_D22; // @[package.scala 96:25:@40252.4 package.scala 96:25:@40253.4]
  wire  _T_1089; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 452:283:@40268.4]
  wire  _T_1090; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 452:291:@40269.4]
  wire  x672_x388_D1; // @[package.scala 96:25:@40285.4 package.scala 96:25:@40286.4]
  wire  x433; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 458:59:@40289.4]
  wire  _T_1120; // @[package.scala 96:25:@40331.4 package.scala 96:25:@40332.4]
  wire  _T_1122; // @[implicits.scala 55:10:@40333.4]
  wire  _T_1123; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 471:194:@40334.4]
  wire  x674_x434_D22; // @[package.scala 96:25:@40319.4 package.scala 96:25:@40320.4]
  wire  _T_1124; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 471:283:@40335.4]
  wire  _T_1125; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 471:291:@40336.4]
  wire  x438; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 475:59:@40347.4]
  wire  _T_1152; // @[package.scala 96:25:@40389.4 package.scala 96:25:@40390.4]
  wire  _T_1154; // @[implicits.scala 55:10:@40391.4]
  wire  _T_1155; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 488:194:@40392.4]
  wire  x676_x439_D22; // @[package.scala 96:25:@40377.4 package.scala 96:25:@40378.4]
  wire  _T_1156; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 488:283:@40393.4]
  wire  _T_1157; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 488:291:@40394.4]
  wire  x443; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 492:59:@40405.4]
  wire  _T_1184; // @[package.scala 96:25:@40447.4 package.scala 96:25:@40448.4]
  wire  _T_1186; // @[implicits.scala 55:10:@40449.4]
  wire  _T_1187; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 505:194:@40450.4]
  wire  x678_x444_D22; // @[package.scala 96:25:@40435.4 package.scala 96:25:@40436.4]
  wire  _T_1188; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 505:283:@40451.4]
  wire  _T_1189; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 505:291:@40452.4]
  wire [31:0] x448_rdrow_number; // @[Math.scala 195:22:@40471.4 Math.scala 196:14:@40472.4]
  wire [31:0] _T_1211; // @[Math.scala 465:37:@40489.4]
  wire  x450; // @[package.scala 96:25:@40497.4 package.scala 96:25:@40498.4]
  wire  x451; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 515:24:@40501.4]
  wire [31:0] x449_number; // @[Math.scala 370:22:@40483.4 Math.scala 371:14:@40484.4]
  wire [31:0] _T_1227; // @[Math.scala 406:49:@40510.4]
  wire [31:0] _T_1229; // @[Math.scala 406:56:@40512.4]
  wire [31:0] _T_1230; // @[Math.scala 406:56:@40513.4]
  wire  _T_1235; // @[FixedPoint.scala 50:25:@40519.4]
  wire [1:0] _T_1239; // @[Bitwise.scala 72:12:@40521.4]
  wire [29:0] _T_1240; // @[FixedPoint.scala 18:52:@40522.4]
  wire  _T_1269; // @[package.scala 96:25:@40575.4 package.scala 96:25:@40576.4]
  wire  _T_1271; // @[implicits.scala 55:10:@40577.4]
  wire  _T_1272; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 534:194:@40578.4]
  wire  x679_x452_D22; // @[package.scala 96:25:@40554.4 package.scala 96:25:@40555.4]
  wire  _T_1273; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 534:283:@40579.4]
  wire  _T_1274; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 534:291:@40580.4]
  wire  x459; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 544:59:@40591.4]
  wire  _T_1300; // @[package.scala 96:25:@40626.4 package.scala 96:25:@40627.4]
  wire  _T_1302; // @[implicits.scala 55:10:@40628.4]
  wire  _T_1303; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 557:194:@40629.4]
  wire  x681_x460_D22; // @[package.scala 96:25:@40614.4 package.scala 96:25:@40615.4]
  wire  _T_1304; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 557:283:@40630.4]
  wire  _T_1305; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 557:291:@40631.4]
  wire  x464; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 561:59:@40642.4]
  wire  _T_1329; // @[package.scala 96:25:@40675.4 package.scala 96:25:@40676.4]
  wire  _T_1331; // @[implicits.scala 55:10:@40677.4]
  wire  _T_1332; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 572:194:@40678.4]
  wire  x682_x465_D22; // @[package.scala 96:25:@40663.4 package.scala 96:25:@40664.4]
  wire  _T_1333; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 572:283:@40679.4]
  wire  _T_1334; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 572:291:@40680.4]
  wire  x469; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 576:59:@40691.4]
  wire  _T_1358; // @[package.scala 96:25:@40724.4 package.scala 96:25:@40725.4]
  wire  _T_1360; // @[implicits.scala 55:10:@40726.4]
  wire  _T_1361; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 587:194:@40727.4]
  wire  x683_x470_D22; // @[package.scala 96:25:@40712.4 package.scala 96:25:@40713.4]
  wire  _T_1362; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 587:283:@40728.4]
  wire  _T_1363; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 587:291:@40729.4]
  wire  x474; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 591:59:@40740.4]
  wire  _T_1387; // @[package.scala 96:25:@40773.4 package.scala 96:25:@40774.4]
  wire  _T_1389; // @[implicits.scala 55:10:@40775.4]
  wire  _T_1390; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 602:194:@40776.4]
  wire  x684_x475_D22; // @[package.scala 96:25:@40761.4 package.scala 96:25:@40762.4]
  wire  _T_1391; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 602:283:@40777.4]
  wire  _T_1392; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 602:291:@40778.4]
  wire  x479; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 606:59:@40789.4]
  wire  _T_1416; // @[package.scala 96:25:@40822.4 package.scala 96:25:@40823.4]
  wire  _T_1418; // @[implicits.scala 55:10:@40824.4]
  wire  _T_1419; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 617:194:@40825.4]
  wire  x685_x480_D22; // @[package.scala 96:25:@40810.4 package.scala 96:25:@40811.4]
  wire  _T_1420; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 617:283:@40826.4]
  wire  _T_1421; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 617:291:@40827.4]
  wire [7:0] x380_rd_0_number; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 259:29:@39548.4 sm_x542_inr_Foreach_SAMPLER_BOX.scala 263:338:@39569.4]
  wire [8:0] _GEN_0; // @[Math.scala 450:32:@40839.4]
  wire [7:0] x421_rd_0_number; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 406:29:@40137.4 sm_x542_inr_Foreach_SAMPLER_BOX.scala 410:408:@40158.4]
  wire [8:0] _GEN_1; // @[Math.scala 450:32:@40851.4]
  wire [7:0] x426_rd_0_number; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 431:29:@40197.4 sm_x542_inr_Foreach_SAMPLER_BOX.scala 435:408:@40218.4]
  wire [9:0] _GEN_2; // @[Math.scala 450:32:@40863.4]
  wire [7:0] x431_rd_0_number; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 448:29:@40255.4 sm_x542_inr_Foreach_SAMPLER_BOX.scala 452:408:@40276.4]
  wire [8:0] _GEN_3; // @[Math.scala 450:32:@40875.4]
  wire [7:0] x462_rd_0_number; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 553:29:@40617.4 sm_x542_inr_Foreach_SAMPLER_BOX.scala 557:408:@40638.4]
  wire [8:0] _GEN_4; // @[Math.scala 450:32:@40887.4]
  wire [7:0] x496_sum_number; // @[Math.scala 154:22:@41057.4 Math.scala 155:14:@41058.4]
  wire [3:0] _T_1515; // @[FixedPoint.scala 18:52:@41063.4]
  wire [7:0] x386_rd_0_number; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 284:29:@39647.4 sm_x542_inr_Foreach_SAMPLER_BOX.scala 288:338:@39668.4]
  wire [8:0] _GEN_5; // @[Math.scala 450:32:@41069.4]
  wire [8:0] _GEN_6; // @[Math.scala 450:32:@41081.4]
  wire [9:0] _GEN_7; // @[Math.scala 450:32:@41093.4]
  wire [7:0] x436_rd_0_number; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 467:29:@40322.4 sm_x542_inr_Foreach_SAMPLER_BOX.scala 471:408:@40343.4]
  wire [8:0] _GEN_8; // @[Math.scala 450:32:@41105.4]
  wire [7:0] x467_rd_0_number; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 568:29:@40666.4 sm_x542_inr_Foreach_SAMPLER_BOX.scala 572:408:@40687.4]
  wire [8:0] _GEN_9; // @[Math.scala 450:32:@41117.4]
  wire [7:0] x510_sum_number; // @[Math.scala 154:22:@41285.4 Math.scala 155:14:@41286.4]
  wire [3:0] _T_1606; // @[FixedPoint.scala 18:52:@41291.4]
  wire [7:0] x392_rd_0_number; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 317:29:@39748.4 sm_x542_inr_Foreach_SAMPLER_BOX.scala 321:408:@39769.4]
  wire [8:0] _GEN_10; // @[Math.scala 450:32:@41297.4]
  wire [9:0] _GEN_11; // @[Math.scala 450:32:@41309.4]
  wire [7:0] x441_rd_0_number; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 484:29:@40380.4 sm_x542_inr_Foreach_SAMPLER_BOX.scala 488:408:@40401.4]
  wire [8:0] _GEN_12; // @[Math.scala 450:32:@41321.4]
  wire [7:0] x472_rd_0_number; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 583:29:@40715.4 sm_x542_inr_Foreach_SAMPLER_BOX.scala 587:408:@40736.4]
  wire [8:0] _GEN_13; // @[Math.scala 450:32:@41333.4]
  wire [7:0] x523_sum_number; // @[Math.scala 154:22:@41492.4 Math.scala 155:14:@41493.4]
  wire [3:0] _T_1688; // @[FixedPoint.scala 18:52:@41498.4]
  wire [7:0] x401_rd_0_number; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 346:29:@39874.4 sm_x542_inr_Foreach_SAMPLER_BOX.scala 350:408:@39895.4]
  wire [8:0] _GEN_14; // @[Math.scala 450:32:@41506.4]
  wire [9:0] _GEN_15; // @[Math.scala 450:32:@41518.4]
  wire [7:0] x446_rd_0_number; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 501:29:@40438.4 sm_x542_inr_Foreach_SAMPLER_BOX.scala 505:408:@40459.4]
  wire [8:0] _GEN_16; // @[Math.scala 450:32:@41530.4]
  wire [7:0] x477_rd_0_number; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 598:29:@40764.4 sm_x542_inr_Foreach_SAMPLER_BOX.scala 602:408:@40785.4]
  wire [8:0] _GEN_17; // @[Math.scala 450:32:@41542.4]
  wire [7:0] x536_sum_number; // @[Math.scala 154:22:@41701.4 Math.scala 155:14:@41702.4]
  wire [3:0] _T_1772; // @[FixedPoint.scala 18:52:@41707.4]
  wire [7:0] x720_x524_D3_number; // @[package.scala 96:25:@41717.4 package.scala 96:25:@41718.4]
  wire [7:0] x722_x537_D3_number; // @[package.scala 96:25:@41735.4 package.scala 96:25:@41736.4]
  wire [15:0] _T_1797; // @[Cat.scala 30:58:@41753.4]
  wire [7:0] x721_x497_D3_number; // @[package.scala 96:25:@41726.4 package.scala 96:25:@41727.4]
  wire [7:0] x723_x511_D3_number; // @[package.scala 96:25:@41744.4 package.scala 96:25:@41745.4]
  wire [15:0] _T_1798; // @[Cat.scala 30:58:@41754.4]
  wire  _T_1811; // @[package.scala 96:25:@41790.4 package.scala 96:25:@41791.4]
  wire  _T_1813; // @[implicits.scala 55:10:@41792.4]
  wire  x724_b327_D63; // @[package.scala 96:25:@41772.4 package.scala 96:25:@41773.4]
  wire  _T_1814; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 829:117:@41793.4]
  wire  x725_b328_D63; // @[package.scala 96:25:@41781.4 package.scala 96:25:@41782.4]
  wire  _T_1815; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 829:123:@41794.4]
  wire [31:0] x616_x340_D8_number; // @[package.scala 96:25:@38895.4 package.scala 96:25:@38896.4]
  wire [31:0] x617_x344_sum_D3_number; // @[package.scala 96:25:@38904.4 package.scala 96:25:@38905.4]
  wire [31:0] x618_x610_D24_number; // @[package.scala 96:25:@38913.4 package.scala 96:25:@38914.4]
  wire [31:0] x624_x348_D7_number; // @[package.scala 96:25:@39038.4 package.scala 96:25:@39039.4]
  wire [31:0] x625_x350_sum_D2_number; // @[package.scala 96:25:@39047.4 package.scala 96:25:@39048.4]
  wire [31:0] x627_x356_sum_D2_number; // @[package.scala 96:25:@39136.4 package.scala 96:25:@39137.4]
  wire [31:0] x628_x354_D7_number; // @[package.scala 96:25:@39145.4 package.scala 96:25:@39146.4]
  wire [31:0] x629_x360_D7_number; // @[package.scala 96:25:@39225.4 package.scala 96:25:@39226.4]
  wire [31:0] x630_x362_sum_D2_number; // @[package.scala 96:25:@39234.4 package.scala 96:25:@39235.4]
  wire [31:0] x637_x360_D33_number; // @[package.scala 96:25:@39410.4 package.scala 96:25:@39411.4]
  wire [31:0] x638_x611_D8_number; // @[package.scala 96:25:@39419.4 package.scala 96:25:@39420.4]
  wire [31:0] x640_x373_sum_D1_number; // @[package.scala 96:25:@39437.4 package.scala 96:25:@39438.4]
  wire [31:0] x644_x379_sum_D1_number; // @[package.scala 96:25:@39527.4 package.scala 96:25:@39528.4]
  wire [31:0] x646_x354_D33_number; // @[package.scala 96:25:@39545.4 package.scala 96:25:@39546.4]
  wire [31:0] x649_x385_sum_D1_number; // @[package.scala 96:25:@39626.4 package.scala 96:25:@39627.4]
  wire [31:0] x651_x348_D33_number; // @[package.scala 96:25:@39644.4 package.scala 96:25:@39645.4]
  wire [31:0] x654_x340_D34_number; // @[package.scala 96:25:@39727.4 package.scala 96:25:@39728.4]
  wire [31:0] x655_x391_sum_D1_number; // @[package.scala 96:25:@39736.4 package.scala 96:25:@39737.4]
  wire [31:0] x659_x398_D7_number; // @[package.scala 96:25:@39862.4 package.scala 96:25:@39863.4]
  wire [31:0] x660_x400_sum_D1_number; // @[package.scala 96:25:@39871.4 package.scala 96:25:@39872.4]
  wire [31:0] x662_x407_D7_number; // @[package.scala 96:25:@39979.4 package.scala 96:25:@39980.4]
  wire [31:0] x664_x409_sum_D1_number; // @[package.scala 96:25:@39997.4 package.scala 96:25:@39998.4]
  wire [31:0] x420_sum_number; // @[Math.scala 154:22:@40116.4 Math.scala 155:14:@40117.4]
  wire [31:0] x667_x612_D7_number; // @[package.scala 96:25:@40134.4 package.scala 96:25:@40135.4]
  wire [31:0] x425_sum_number; // @[Math.scala 154:22:@40185.4 Math.scala 155:14:@40186.4]
  wire [31:0] x430_sum_number; // @[Math.scala 154:22:@40243.4 Math.scala 155:14:@40244.4]
  wire [31:0] x435_sum_number; // @[Math.scala 154:22:@40310.4 Math.scala 155:14:@40311.4]
  wire [31:0] x440_sum_number; // @[Math.scala 154:22:@40368.4 Math.scala 155:14:@40369.4]
  wire [31:0] x445_sum_number; // @[Math.scala 154:22:@40426.4 Math.scala 155:14:@40427.4]
  wire [31:0] x456_sum_number; // @[Math.scala 154:22:@40545.4 Math.scala 155:14:@40546.4]
  wire [31:0] x680_x613_D7_number; // @[package.scala 96:25:@40563.4 package.scala 96:25:@40564.4]
  wire [31:0] x461_sum_number; // @[Math.scala 154:22:@40605.4 Math.scala 155:14:@40606.4]
  wire [31:0] x466_sum_number; // @[Math.scala 154:22:@40654.4 Math.scala 155:14:@40655.4]
  wire [31:0] x471_sum_number; // @[Math.scala 154:22:@40703.4 Math.scala 155:14:@40704.4]
  wire [31:0] x476_sum_number; // @[Math.scala 154:22:@40752.4 Math.scala 155:14:@40753.4]
  wire [31:0] x481_sum_number; // @[Math.scala 154:22:@40801.4 Math.scala 155:14:@40802.4]
  wire [8:0] _T_1429; // @[package.scala 96:25:@40845.4 package.scala 96:25:@40846.4]
  wire [8:0] _T_1435; // @[package.scala 96:25:@40857.4 package.scala 96:25:@40858.4]
  wire [9:0] _T_1441; // @[package.scala 96:25:@40869.4 package.scala 96:25:@40870.4]
  wire [8:0] _T_1447; // @[package.scala 96:25:@40881.4 package.scala 96:25:@40882.4]
  wire [8:0] _T_1453; // @[package.scala 96:25:@40893.4 package.scala 96:25:@40894.4]
  wire [8:0] _T_1522; // @[package.scala 96:25:@41075.4 package.scala 96:25:@41076.4]
  wire [8:0] _T_1528; // @[package.scala 96:25:@41087.4 package.scala 96:25:@41088.4]
  wire [9:0] _T_1534; // @[package.scala 96:25:@41099.4 package.scala 96:25:@41100.4]
  wire [8:0] _T_1540; // @[package.scala 96:25:@41111.4 package.scala 96:25:@41112.4]
  wire [8:0] _T_1546; // @[package.scala 96:25:@41123.4 package.scala 96:25:@41124.4]
  wire [8:0] _T_1613; // @[package.scala 96:25:@41303.4 package.scala 96:25:@41304.4]
  wire [9:0] _T_1619; // @[package.scala 96:25:@41315.4 package.scala 96:25:@41316.4]
  wire [8:0] _T_1625; // @[package.scala 96:25:@41327.4 package.scala 96:25:@41328.4]
  wire [8:0] _T_1631; // @[package.scala 96:25:@41339.4 package.scala 96:25:@41340.4]
  wire [8:0] _T_1697; // @[package.scala 96:25:@41512.4 package.scala 96:25:@41513.4]
  wire [9:0] _T_1703; // @[package.scala 96:25:@41524.4 package.scala 96:25:@41525.4]
  wire [8:0] _T_1709; // @[package.scala 96:25:@41536.4 package.scala 96:25:@41537.4]
  wire [8:0] _T_1715; // @[package.scala 96:25:@41548.4 package.scala 96:25:@41549.4]
  _ _ ( // @[Math.scala 709:24:@38564.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 709:24:@38576.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  x329_lb_0 x329_lb_0 ( // @[m_x329_lb_0.scala 47:17:@38586.4]
    .clock(x329_lb_0_clock),
    .reset(x329_lb_0_reset),
    .io_rPort_17_banks_1(x329_lb_0_io_rPort_17_banks_1),
    .io_rPort_17_banks_0(x329_lb_0_io_rPort_17_banks_0),
    .io_rPort_17_ofs_0(x329_lb_0_io_rPort_17_ofs_0),
    .io_rPort_17_en_0(x329_lb_0_io_rPort_17_en_0),
    .io_rPort_17_backpressure(x329_lb_0_io_rPort_17_backpressure),
    .io_rPort_17_output_0(x329_lb_0_io_rPort_17_output_0),
    .io_rPort_16_banks_1(x329_lb_0_io_rPort_16_banks_1),
    .io_rPort_16_banks_0(x329_lb_0_io_rPort_16_banks_0),
    .io_rPort_16_ofs_0(x329_lb_0_io_rPort_16_ofs_0),
    .io_rPort_16_en_0(x329_lb_0_io_rPort_16_en_0),
    .io_rPort_16_backpressure(x329_lb_0_io_rPort_16_backpressure),
    .io_rPort_16_output_0(x329_lb_0_io_rPort_16_output_0),
    .io_rPort_15_banks_1(x329_lb_0_io_rPort_15_banks_1),
    .io_rPort_15_banks_0(x329_lb_0_io_rPort_15_banks_0),
    .io_rPort_15_ofs_0(x329_lb_0_io_rPort_15_ofs_0),
    .io_rPort_15_en_0(x329_lb_0_io_rPort_15_en_0),
    .io_rPort_15_backpressure(x329_lb_0_io_rPort_15_backpressure),
    .io_rPort_15_output_0(x329_lb_0_io_rPort_15_output_0),
    .io_rPort_14_banks_1(x329_lb_0_io_rPort_14_banks_1),
    .io_rPort_14_banks_0(x329_lb_0_io_rPort_14_banks_0),
    .io_rPort_14_ofs_0(x329_lb_0_io_rPort_14_ofs_0),
    .io_rPort_14_en_0(x329_lb_0_io_rPort_14_en_0),
    .io_rPort_14_backpressure(x329_lb_0_io_rPort_14_backpressure),
    .io_rPort_14_output_0(x329_lb_0_io_rPort_14_output_0),
    .io_rPort_13_banks_1(x329_lb_0_io_rPort_13_banks_1),
    .io_rPort_13_banks_0(x329_lb_0_io_rPort_13_banks_0),
    .io_rPort_13_ofs_0(x329_lb_0_io_rPort_13_ofs_0),
    .io_rPort_13_en_0(x329_lb_0_io_rPort_13_en_0),
    .io_rPort_13_backpressure(x329_lb_0_io_rPort_13_backpressure),
    .io_rPort_13_output_0(x329_lb_0_io_rPort_13_output_0),
    .io_rPort_12_banks_1(x329_lb_0_io_rPort_12_banks_1),
    .io_rPort_12_banks_0(x329_lb_0_io_rPort_12_banks_0),
    .io_rPort_12_ofs_0(x329_lb_0_io_rPort_12_ofs_0),
    .io_rPort_12_en_0(x329_lb_0_io_rPort_12_en_0),
    .io_rPort_12_backpressure(x329_lb_0_io_rPort_12_backpressure),
    .io_rPort_12_output_0(x329_lb_0_io_rPort_12_output_0),
    .io_rPort_11_banks_1(x329_lb_0_io_rPort_11_banks_1),
    .io_rPort_11_banks_0(x329_lb_0_io_rPort_11_banks_0),
    .io_rPort_11_ofs_0(x329_lb_0_io_rPort_11_ofs_0),
    .io_rPort_11_en_0(x329_lb_0_io_rPort_11_en_0),
    .io_rPort_11_backpressure(x329_lb_0_io_rPort_11_backpressure),
    .io_rPort_11_output_0(x329_lb_0_io_rPort_11_output_0),
    .io_rPort_10_banks_1(x329_lb_0_io_rPort_10_banks_1),
    .io_rPort_10_banks_0(x329_lb_0_io_rPort_10_banks_0),
    .io_rPort_10_ofs_0(x329_lb_0_io_rPort_10_ofs_0),
    .io_rPort_10_en_0(x329_lb_0_io_rPort_10_en_0),
    .io_rPort_10_backpressure(x329_lb_0_io_rPort_10_backpressure),
    .io_rPort_10_output_0(x329_lb_0_io_rPort_10_output_0),
    .io_rPort_9_banks_1(x329_lb_0_io_rPort_9_banks_1),
    .io_rPort_9_banks_0(x329_lb_0_io_rPort_9_banks_0),
    .io_rPort_9_ofs_0(x329_lb_0_io_rPort_9_ofs_0),
    .io_rPort_9_en_0(x329_lb_0_io_rPort_9_en_0),
    .io_rPort_9_backpressure(x329_lb_0_io_rPort_9_backpressure),
    .io_rPort_9_output_0(x329_lb_0_io_rPort_9_output_0),
    .io_rPort_8_banks_1(x329_lb_0_io_rPort_8_banks_1),
    .io_rPort_8_banks_0(x329_lb_0_io_rPort_8_banks_0),
    .io_rPort_8_ofs_0(x329_lb_0_io_rPort_8_ofs_0),
    .io_rPort_8_en_0(x329_lb_0_io_rPort_8_en_0),
    .io_rPort_8_backpressure(x329_lb_0_io_rPort_8_backpressure),
    .io_rPort_8_output_0(x329_lb_0_io_rPort_8_output_0),
    .io_rPort_7_banks_1(x329_lb_0_io_rPort_7_banks_1),
    .io_rPort_7_banks_0(x329_lb_0_io_rPort_7_banks_0),
    .io_rPort_7_ofs_0(x329_lb_0_io_rPort_7_ofs_0),
    .io_rPort_7_en_0(x329_lb_0_io_rPort_7_en_0),
    .io_rPort_7_backpressure(x329_lb_0_io_rPort_7_backpressure),
    .io_rPort_7_output_0(x329_lb_0_io_rPort_7_output_0),
    .io_rPort_6_banks_1(x329_lb_0_io_rPort_6_banks_1),
    .io_rPort_6_banks_0(x329_lb_0_io_rPort_6_banks_0),
    .io_rPort_6_ofs_0(x329_lb_0_io_rPort_6_ofs_0),
    .io_rPort_6_en_0(x329_lb_0_io_rPort_6_en_0),
    .io_rPort_6_backpressure(x329_lb_0_io_rPort_6_backpressure),
    .io_rPort_6_output_0(x329_lb_0_io_rPort_6_output_0),
    .io_rPort_5_banks_1(x329_lb_0_io_rPort_5_banks_1),
    .io_rPort_5_banks_0(x329_lb_0_io_rPort_5_banks_0),
    .io_rPort_5_ofs_0(x329_lb_0_io_rPort_5_ofs_0),
    .io_rPort_5_en_0(x329_lb_0_io_rPort_5_en_0),
    .io_rPort_5_backpressure(x329_lb_0_io_rPort_5_backpressure),
    .io_rPort_5_output_0(x329_lb_0_io_rPort_5_output_0),
    .io_rPort_4_banks_1(x329_lb_0_io_rPort_4_banks_1),
    .io_rPort_4_banks_0(x329_lb_0_io_rPort_4_banks_0),
    .io_rPort_4_ofs_0(x329_lb_0_io_rPort_4_ofs_0),
    .io_rPort_4_en_0(x329_lb_0_io_rPort_4_en_0),
    .io_rPort_4_backpressure(x329_lb_0_io_rPort_4_backpressure),
    .io_rPort_4_output_0(x329_lb_0_io_rPort_4_output_0),
    .io_rPort_3_banks_1(x329_lb_0_io_rPort_3_banks_1),
    .io_rPort_3_banks_0(x329_lb_0_io_rPort_3_banks_0),
    .io_rPort_3_ofs_0(x329_lb_0_io_rPort_3_ofs_0),
    .io_rPort_3_en_0(x329_lb_0_io_rPort_3_en_0),
    .io_rPort_3_backpressure(x329_lb_0_io_rPort_3_backpressure),
    .io_rPort_3_output_0(x329_lb_0_io_rPort_3_output_0),
    .io_rPort_2_banks_1(x329_lb_0_io_rPort_2_banks_1),
    .io_rPort_2_banks_0(x329_lb_0_io_rPort_2_banks_0),
    .io_rPort_2_ofs_0(x329_lb_0_io_rPort_2_ofs_0),
    .io_rPort_2_en_0(x329_lb_0_io_rPort_2_en_0),
    .io_rPort_2_backpressure(x329_lb_0_io_rPort_2_backpressure),
    .io_rPort_2_output_0(x329_lb_0_io_rPort_2_output_0),
    .io_rPort_1_banks_1(x329_lb_0_io_rPort_1_banks_1),
    .io_rPort_1_banks_0(x329_lb_0_io_rPort_1_banks_0),
    .io_rPort_1_ofs_0(x329_lb_0_io_rPort_1_ofs_0),
    .io_rPort_1_en_0(x329_lb_0_io_rPort_1_en_0),
    .io_rPort_1_backpressure(x329_lb_0_io_rPort_1_backpressure),
    .io_rPort_1_output_0(x329_lb_0_io_rPort_1_output_0),
    .io_rPort_0_banks_1(x329_lb_0_io_rPort_0_banks_1),
    .io_rPort_0_banks_0(x329_lb_0_io_rPort_0_banks_0),
    .io_rPort_0_ofs_0(x329_lb_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x329_lb_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x329_lb_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x329_lb_0_io_rPort_0_output_0),
    .io_wPort_3_banks_1(x329_lb_0_io_wPort_3_banks_1),
    .io_wPort_3_banks_0(x329_lb_0_io_wPort_3_banks_0),
    .io_wPort_3_ofs_0(x329_lb_0_io_wPort_3_ofs_0),
    .io_wPort_3_data_0(x329_lb_0_io_wPort_3_data_0),
    .io_wPort_3_en_0(x329_lb_0_io_wPort_3_en_0),
    .io_wPort_2_banks_1(x329_lb_0_io_wPort_2_banks_1),
    .io_wPort_2_banks_0(x329_lb_0_io_wPort_2_banks_0),
    .io_wPort_2_ofs_0(x329_lb_0_io_wPort_2_ofs_0),
    .io_wPort_2_data_0(x329_lb_0_io_wPort_2_data_0),
    .io_wPort_2_en_0(x329_lb_0_io_wPort_2_en_0),
    .io_wPort_1_banks_1(x329_lb_0_io_wPort_1_banks_1),
    .io_wPort_1_banks_0(x329_lb_0_io_wPort_1_banks_0),
    .io_wPort_1_ofs_0(x329_lb_0_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(x329_lb_0_io_wPort_1_data_0),
    .io_wPort_1_en_0(x329_lb_0_io_wPort_1_en_0),
    .io_wPort_0_banks_1(x329_lb_0_io_wPort_0_banks_1),
    .io_wPort_0_banks_0(x329_lb_0_io_wPort_0_banks_0),
    .io_wPort_0_ofs_0(x329_lb_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x329_lb_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x329_lb_0_io_wPort_0_en_0)
  );
  RetimeWrapper_260 RetimeWrapper ( // @[package.scala 93:22:@38744.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x340 x340_1 ( // @[Math.scala 366:24:@38828.4]
    .clock(x340_1_clock),
    .reset(x340_1_reset),
    .io_a(x340_1_io_a),
    .io_b(x340_1_io_b),
    .io_flow(x340_1_io_flow),
    .io_result(x340_1_io_result)
  );
  x342_mul x342_mul_1 ( // @[Math.scala 262:24:@38849.4]
    .clock(x342_mul_1_clock),
    .reset(x342_mul_1_reset),
    .io_a(x342_mul_1_io_a),
    .io_flow(x342_mul_1_io_flow),
    .io_result(x342_mul_1_io_result)
  );
  x343_div x343_div_1 ( // @[Math.scala 327:24:@38861.4]
    .clock(x343_div_1_clock),
    .reset(x343_div_1_reset),
    .io_a(x343_div_1_io_a),
    .io_flow(x343_div_1_io_flow),
    .io_result(x343_div_1_io_result)
  );
  RetimeWrapper_266 RetimeWrapper_1 ( // @[package.scala 93:22:@38871.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x344_sum x344_sum_1 ( // @[Math.scala 150:24:@38880.4]
    .clock(x344_sum_1_clock),
    .reset(x344_sum_1_reset),
    .io_a(x344_sum_1_io_a),
    .io_b(x344_sum_1_io_b),
    .io_flow(x344_sum_1_io_flow),
    .io_result(x344_sum_1_io_result)
  );
  RetimeWrapper_268 RetimeWrapper_2 ( // @[package.scala 93:22:@38890.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_269 RetimeWrapper_3 ( // @[package.scala 93:22:@38899.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_270 RetimeWrapper_4 ( // @[package.scala 93:22:@38908.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_271 RetimeWrapper_5 ( // @[package.scala 93:22:@38917.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_271 RetimeWrapper_6 ( // @[package.scala 93:22:@38926.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_273 RetimeWrapper_7 ( // @[package.scala 93:22:@38935.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_271 RetimeWrapper_8 ( // @[package.scala 93:22:@38946.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  x344_sum x346_rdcol_1 ( // @[Math.scala 150:24:@38969.4]
    .clock(x346_rdcol_1_clock),
    .reset(x346_rdcol_1_reset),
    .io_a(x346_rdcol_1_io_a),
    .io_b(x346_rdcol_1_io_b),
    .io_flow(x346_rdcol_1_io_flow),
    .io_result(x346_rdcol_1_io_result)
  );
  x340 x348_1 ( // @[Math.scala 366:24:@38983.4]
    .clock(x348_1_clock),
    .reset(x348_1_reset),
    .io_a(x348_1_io_a),
    .io_b(x348_1_io_b),
    .io_flow(x348_1_io_flow),
    .io_result(x348_1_io_result)
  );
  x343_div x349_div_1 ( // @[Math.scala 327:24:@38995.4]
    .clock(x349_div_1_clock),
    .reset(x349_div_1_reset),
    .io_a(x349_div_1_io_a),
    .io_flow(x349_div_1_io_flow),
    .io_result(x349_div_1_io_result)
  );
  RetimeWrapper_278 RetimeWrapper_9 ( // @[package.scala 93:22:@39005.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  x344_sum x350_sum_1 ( // @[Math.scala 150:24:@39014.4]
    .clock(x350_sum_1_clock),
    .reset(x350_sum_1_reset),
    .io_a(x350_sum_1_io_a),
    .io_b(x350_sum_1_io_b),
    .io_flow(x350_sum_1_io_flow),
    .io_result(x350_sum_1_io_result)
  );
  RetimeWrapper_273 RetimeWrapper_10 ( // @[package.scala 93:22:@39024.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_281 RetimeWrapper_11 ( // @[package.scala 93:22:@39033.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_282 RetimeWrapper_12 ( // @[package.scala 93:22:@39042.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_271 RetimeWrapper_13 ( // @[package.scala 93:22:@39053.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  x344_sum x352_rdcol_1 ( // @[Math.scala 150:24:@39076.4]
    .clock(x352_rdcol_1_clock),
    .reset(x352_rdcol_1_reset),
    .io_a(x352_rdcol_1_io_a),
    .io_b(x352_rdcol_1_io_b),
    .io_flow(x352_rdcol_1_io_flow),
    .io_result(x352_rdcol_1_io_result)
  );
  x340 x354_1 ( // @[Math.scala 366:24:@39090.4]
    .clock(x354_1_clock),
    .reset(x354_1_reset),
    .io_a(x354_1_io_a),
    .io_b(x354_1_io_b),
    .io_flow(x354_1_io_flow),
    .io_result(x354_1_io_result)
  );
  x343_div x355_div_1 ( // @[Math.scala 327:24:@39102.4]
    .clock(x355_div_1_clock),
    .reset(x355_div_1_reset),
    .io_a(x355_div_1_io_a),
    .io_flow(x355_div_1_io_flow),
    .io_result(x355_div_1_io_result)
  );
  x344_sum x356_sum_1 ( // @[Math.scala 150:24:@39112.4]
    .clock(x356_sum_1_clock),
    .reset(x356_sum_1_reset),
    .io_a(x356_sum_1_io_a),
    .io_b(x356_sum_1_io_b),
    .io_flow(x356_sum_1_io_flow),
    .io_result(x356_sum_1_io_result)
  );
  RetimeWrapper_273 RetimeWrapper_14 ( // @[package.scala 93:22:@39122.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_282 RetimeWrapper_15 ( // @[package.scala 93:22:@39131.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_281 RetimeWrapper_16 ( // @[package.scala 93:22:@39140.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_271 RetimeWrapper_17 ( // @[package.scala 93:22:@39151.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  x344_sum x358_rdcol_1 ( // @[Math.scala 150:24:@39174.4]
    .clock(x358_rdcol_1_clock),
    .reset(x358_rdcol_1_reset),
    .io_a(x358_rdcol_1_io_a),
    .io_b(x358_rdcol_1_io_b),
    .io_flow(x358_rdcol_1_io_flow),
    .io_result(x358_rdcol_1_io_result)
  );
  x340 x360_1 ( // @[Math.scala 366:24:@39188.4]
    .clock(x360_1_clock),
    .reset(x360_1_reset),
    .io_a(x360_1_io_a),
    .io_b(x360_1_io_b),
    .io_flow(x360_1_io_flow),
    .io_result(x360_1_io_result)
  );
  x343_div x361_div_1 ( // @[Math.scala 327:24:@39200.4]
    .clock(x361_div_1_clock),
    .reset(x361_div_1_reset),
    .io_a(x361_div_1_io_a),
    .io_flow(x361_div_1_io_flow),
    .io_result(x361_div_1_io_result)
  );
  x344_sum x362_sum_1 ( // @[Math.scala 150:24:@39210.4]
    .clock(x362_sum_1_clock),
    .reset(x362_sum_1_reset),
    .io_a(x362_sum_1_io_a),
    .io_b(x362_sum_1_io_b),
    .io_flow(x362_sum_1_io_flow),
    .io_result(x362_sum_1_io_result)
  );
  RetimeWrapper_281 RetimeWrapper_18 ( // @[package.scala 93:22:@39220.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_282 RetimeWrapper_19 ( // @[package.scala 93:22:@39229.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_273 RetimeWrapper_20 ( // @[package.scala 93:22:@39238.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_271 RetimeWrapper_21 ( // @[package.scala 93:22:@39249.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_300 RetimeWrapper_22 ( // @[package.scala 93:22:@39270.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  x340 x365_1 ( // @[Math.scala 366:24:@39283.4]
    .clock(x365_1_clock),
    .reset(x365_1_reset),
    .io_a(x365_1_io_a),
    .io_b(x365_1_io_b),
    .io_flow(x365_1_io_flow),
    .io_result(x365_1_io_result)
  );
  RetimeWrapper RetimeWrapper_23 ( // @[package.scala 93:22:@39298.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_300 RetimeWrapper_24 ( // @[package.scala 93:22:@39307.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper RetimeWrapper_25 ( // @[package.scala 93:22:@39321.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper RetimeWrapper_26 ( // @[package.scala 93:22:@39330.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  x342_mul x372_mul_1 ( // @[Math.scala 262:24:@39367.4]
    .clock(x372_mul_1_clock),
    .reset(x372_mul_1_reset),
    .io_a(x372_mul_1_io_a),
    .io_flow(x372_mul_1_io_flow),
    .io_result(x372_mul_1_io_result)
  );
  RetimeWrapper_309 RetimeWrapper_27 ( // @[package.scala 93:22:@39377.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  x344_sum x373_sum_1 ( // @[Math.scala 150:24:@39386.4]
    .clock(x373_sum_1_clock),
    .reset(x373_sum_1_reset),
    .io_a(x373_sum_1_io_a),
    .io_b(x373_sum_1_io_b),
    .io_flow(x373_sum_1_io_flow),
    .io_result(x373_sum_1_io_result)
  );
  RetimeWrapper_311 RetimeWrapper_28 ( // @[package.scala 93:22:@39396.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_312 RetimeWrapper_29 ( // @[package.scala 93:22:@39405.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_268 RetimeWrapper_30 ( // @[package.scala 93:22:@39414.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_311 RetimeWrapper_31 ( // @[package.scala 93:22:@39423.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_260 RetimeWrapper_32 ( // @[package.scala 93:22:@39432.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_316 RetimeWrapper_33 ( // @[package.scala 93:22:@39441.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_311 RetimeWrapper_34 ( // @[package.scala 93:22:@39453.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_300 RetimeWrapper_35 ( // @[package.scala 93:22:@39474.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper RetimeWrapper_36 ( // @[package.scala 93:22:@39488.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_309 RetimeWrapper_37 ( // @[package.scala 93:22:@39503.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  x344_sum x379_sum_1 ( // @[Math.scala 150:24:@39512.4]
    .clock(x379_sum_1_clock),
    .reset(x379_sum_1_reset),
    .io_a(x379_sum_1_io_a),
    .io_b(x379_sum_1_io_b),
    .io_flow(x379_sum_1_io_flow),
    .io_result(x379_sum_1_io_result)
  );
  RetimeWrapper_260 RetimeWrapper_38 ( // @[package.scala 93:22:@39522.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_316 RetimeWrapper_39 ( // @[package.scala 93:22:@39531.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_312 RetimeWrapper_40 ( // @[package.scala 93:22:@39540.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper_311 RetimeWrapper_41 ( // @[package.scala 93:22:@39552.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_300 RetimeWrapper_42 ( // @[package.scala 93:22:@39573.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper RetimeWrapper_43 ( // @[package.scala 93:22:@39587.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_309 RetimeWrapper_44 ( // @[package.scala 93:22:@39602.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  x344_sum x385_sum_1 ( // @[Math.scala 150:24:@39611.4]
    .clock(x385_sum_1_clock),
    .reset(x385_sum_1_reset),
    .io_a(x385_sum_1_io_a),
    .io_b(x385_sum_1_io_b),
    .io_flow(x385_sum_1_io_flow),
    .io_result(x385_sum_1_io_result)
  );
  RetimeWrapper_260 RetimeWrapper_45 ( // @[package.scala 93:22:@39621.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_316 RetimeWrapper_46 ( // @[package.scala 93:22:@39630.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_312 RetimeWrapper_47 ( // @[package.scala 93:22:@39639.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_311 RetimeWrapper_48 ( // @[package.scala 93:22:@39651.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_300 RetimeWrapper_49 ( // @[package.scala 93:22:@39672.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper RetimeWrapper_50 ( // @[package.scala 93:22:@39688.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_336 RetimeWrapper_51 ( // @[package.scala 93:22:@39703.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  x344_sum x391_sum_1 ( // @[Math.scala 150:24:@39712.4]
    .clock(x391_sum_1_clock),
    .reset(x391_sum_1_reset),
    .io_a(x391_sum_1_io_a),
    .io_b(x391_sum_1_io_b),
    .io_flow(x391_sum_1_io_flow),
    .io_result(x391_sum_1_io_result)
  );
  RetimeWrapper_338 RetimeWrapper_52 ( // @[package.scala 93:22:@39722.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_260 RetimeWrapper_53 ( // @[package.scala 93:22:@39731.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper_340 RetimeWrapper_54 ( // @[package.scala 93:22:@39740.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_311 RetimeWrapper_55 ( // @[package.scala 93:22:@39752.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  x344_sum x394_rdcol_1 ( // @[Math.scala 150:24:@39775.4]
    .clock(x394_rdcol_1_clock),
    .reset(x394_rdcol_1_reset),
    .io_a(x394_rdcol_1_io_a),
    .io_b(x394_rdcol_1_io_b),
    .io_flow(x394_rdcol_1_io_flow),
    .io_result(x394_rdcol_1_io_result)
  );
  RetimeWrapper RetimeWrapper_56 ( // @[package.scala 93:22:@39790.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  x340 x398_1 ( // @[Math.scala 366:24:@39807.4]
    .clock(x398_1_clock),
    .reset(x398_1_reset),
    .io_a(x398_1_io_a),
    .io_b(x398_1_io_b),
    .io_flow(x398_1_io_flow),
    .io_result(x398_1_io_result)
  );
  x343_div x399_div_1 ( // @[Math.scala 327:24:@39819.4]
    .clock(x399_div_1_clock),
    .reset(x399_div_1_reset),
    .io_a(x399_div_1_io_a),
    .io_flow(x399_div_1_io_flow),
    .io_result(x399_div_1_io_result)
  );
  RetimeWrapper_260 RetimeWrapper_57 ( // @[package.scala 93:22:@39829.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  x344_sum x400_sum_1 ( // @[Math.scala 150:24:@39838.4]
    .clock(x400_sum_1_clock),
    .reset(x400_sum_1_reset),
    .io_a(x400_sum_1_io_a),
    .io_b(x400_sum_1_io_b),
    .io_flow(x400_sum_1_io_flow),
    .io_result(x400_sum_1_io_result)
  );
  RetimeWrapper_316 RetimeWrapper_58 ( // @[package.scala 93:22:@39848.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_281 RetimeWrapper_59 ( // @[package.scala 93:22:@39857.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_260 RetimeWrapper_60 ( // @[package.scala 93:22:@39866.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_311 RetimeWrapper_61 ( // @[package.scala 93:22:@39878.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  x344_sum x403_rdcol_1 ( // @[Math.scala 150:24:@39901.4]
    .clock(x403_rdcol_1_clock),
    .reset(x403_rdcol_1_reset),
    .io_a(x403_rdcol_1_io_a),
    .io_b(x403_rdcol_1_io_b),
    .io_flow(x403_rdcol_1_io_flow),
    .io_result(x403_rdcol_1_io_result)
  );
  RetimeWrapper RetimeWrapper_62 ( // @[package.scala 93:22:@39916.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  x340 x407_1 ( // @[Math.scala 366:24:@39933.4]
    .clock(x407_1_clock),
    .reset(x407_1_reset),
    .io_a(x407_1_io_a),
    .io_b(x407_1_io_b),
    .io_flow(x407_1_io_flow),
    .io_result(x407_1_io_result)
  );
  x343_div x408_div_1 ( // @[Math.scala 327:24:@39945.4]
    .clock(x408_div_1_clock),
    .reset(x408_div_1_reset),
    .io_a(x408_div_1_io_a),
    .io_flow(x408_div_1_io_flow),
    .io_result(x408_div_1_io_result)
  );
  RetimeWrapper_260 RetimeWrapper_63 ( // @[package.scala 93:22:@39955.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  x344_sum x409_sum_1 ( // @[Math.scala 150:24:@39964.4]
    .clock(x409_sum_1_clock),
    .reset(x409_sum_1_reset),
    .io_a(x409_sum_1_io_a),
    .io_b(x409_sum_1_io_b),
    .io_flow(x409_sum_1_io_flow),
    .io_result(x409_sum_1_io_result)
  );
  RetimeWrapper_281 RetimeWrapper_64 ( // @[package.scala 93:22:@39974.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_316 RetimeWrapper_65 ( // @[package.scala 93:22:@39983.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper_260 RetimeWrapper_66 ( // @[package.scala 93:22:@39992.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper_311 RetimeWrapper_67 ( // @[package.scala 93:22:@40004.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  x412_rdrow x412_rdrow_1 ( // @[Math.scala 191:24:@40027.4]
    .clock(x412_rdrow_1_clock),
    .reset(x412_rdrow_1_reset),
    .io_a(x412_rdrow_1_io_a),
    .io_b(x412_rdrow_1_io_b),
    .io_flow(x412_rdrow_1_io_flow),
    .io_result(x412_rdrow_1_io_result)
  );
  x340 x413_1 ( // @[Math.scala 366:24:@40039.4]
    .clock(x413_1_clock),
    .reset(x413_1_reset),
    .io_a(x413_1_io_a),
    .io_b(x413_1_io_b),
    .io_flow(x413_1_io_flow),
    .io_result(x413_1_io_result)
  );
  RetimeWrapper RetimeWrapper_68 ( // @[package.scala 93:22:@40054.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  x342_mul x419_mul_1 ( // @[Math.scala 262:24:@40091.4]
    .clock(x419_mul_1_clock),
    .reset(x419_mul_1_reset),
    .io_a(x419_mul_1_io_a),
    .io_flow(x419_mul_1_io_flow),
    .io_result(x419_mul_1_io_result)
  );
  RetimeWrapper_336 RetimeWrapper_69 ( // @[package.scala 93:22:@40101.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  x344_sum x420_sum_1 ( // @[Math.scala 150:24:@40110.4]
    .clock(x420_sum_1_clock),
    .reset(x420_sum_1_reset),
    .io_a(x420_sum_1_io_a),
    .io_b(x420_sum_1_io_b),
    .io_flow(x420_sum_1_io_flow),
    .io_result(x420_sum_1_io_result)
  );
  RetimeWrapper_316 RetimeWrapper_70 ( // @[package.scala 93:22:@40120.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_281 RetimeWrapper_71 ( // @[package.scala 93:22:@40129.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  RetimeWrapper_311 RetimeWrapper_72 ( // @[package.scala 93:22:@40141.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  RetimeWrapper_336 RetimeWrapper_73 ( // @[package.scala 93:22:@40168.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  x344_sum x425_sum_1 ( // @[Math.scala 150:24:@40179.4]
    .clock(x425_sum_1_clock),
    .reset(x425_sum_1_reset),
    .io_a(x425_sum_1_io_a),
    .io_b(x425_sum_1_io_b),
    .io_flow(x425_sum_1_io_flow),
    .io_result(x425_sum_1_io_result)
  );
  RetimeWrapper_316 RetimeWrapper_74 ( // @[package.scala 93:22:@40189.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  RetimeWrapper_311 RetimeWrapper_75 ( // @[package.scala 93:22:@40201.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_336 RetimeWrapper_76 ( // @[package.scala 93:22:@40228.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  x344_sum x430_sum_1 ( // @[Math.scala 150:24:@40237.4]
    .clock(x430_sum_1_clock),
    .reset(x430_sum_1_reset),
    .io_a(x430_sum_1_io_a),
    .io_b(x430_sum_1_io_b),
    .io_flow(x430_sum_1_io_flow),
    .io_result(x430_sum_1_io_result)
  );
  RetimeWrapper_316 RetimeWrapper_77 ( // @[package.scala 93:22:@40247.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  RetimeWrapper_311 RetimeWrapper_78 ( // @[package.scala 93:22:@40259.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  RetimeWrapper RetimeWrapper_79 ( // @[package.scala 93:22:@40280.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper_382 RetimeWrapper_80 ( // @[package.scala 93:22:@40295.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  x344_sum x435_sum_1 ( // @[Math.scala 150:24:@40304.4]
    .clock(x435_sum_1_clock),
    .reset(x435_sum_1_reset),
    .io_a(x435_sum_1_io_a),
    .io_b(x435_sum_1_io_b),
    .io_flow(x435_sum_1_io_flow),
    .io_result(x435_sum_1_io_result)
  );
  RetimeWrapper_316 RetimeWrapper_81 ( // @[package.scala 93:22:@40314.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_311 RetimeWrapper_82 ( // @[package.scala 93:22:@40326.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  RetimeWrapper_282 RetimeWrapper_83 ( // @[package.scala 93:22:@40353.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  x344_sum x440_sum_1 ( // @[Math.scala 150:24:@40362.4]
    .clock(x440_sum_1_clock),
    .reset(x440_sum_1_reset),
    .io_a(x440_sum_1_io_a),
    .io_b(x440_sum_1_io_b),
    .io_flow(x440_sum_1_io_flow),
    .io_result(x440_sum_1_io_result)
  );
  RetimeWrapper_316 RetimeWrapper_84 ( // @[package.scala 93:22:@40372.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  RetimeWrapper_311 RetimeWrapper_85 ( // @[package.scala 93:22:@40384.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  RetimeWrapper_282 RetimeWrapper_86 ( // @[package.scala 93:22:@40411.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  x344_sum x445_sum_1 ( // @[Math.scala 150:24:@40420.4]
    .clock(x445_sum_1_clock),
    .reset(x445_sum_1_reset),
    .io_a(x445_sum_1_io_a),
    .io_b(x445_sum_1_io_b),
    .io_flow(x445_sum_1_io_flow),
    .io_result(x445_sum_1_io_result)
  );
  RetimeWrapper_316 RetimeWrapper_87 ( // @[package.scala 93:22:@40430.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  RetimeWrapper_311 RetimeWrapper_88 ( // @[package.scala 93:22:@40442.4]
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  x412_rdrow x448_rdrow_1 ( // @[Math.scala 191:24:@40465.4]
    .clock(x448_rdrow_1_clock),
    .reset(x448_rdrow_1_reset),
    .io_a(x448_rdrow_1_io_a),
    .io_b(x448_rdrow_1_io_b),
    .io_flow(x448_rdrow_1_io_flow),
    .io_result(x448_rdrow_1_io_result)
  );
  x340 x449_1 ( // @[Math.scala 366:24:@40477.4]
    .clock(x449_1_clock),
    .reset(x449_1_reset),
    .io_a(x449_1_io_a),
    .io_b(x449_1_io_b),
    .io_flow(x449_1_io_flow),
    .io_result(x449_1_io_result)
  );
  RetimeWrapper RetimeWrapper_89 ( // @[package.scala 93:22:@40492.4]
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  x342_mul x455_mul_1 ( // @[Math.scala 262:24:@40529.4]
    .clock(x455_mul_1_clock),
    .reset(x455_mul_1_reset),
    .io_a(x455_mul_1_io_a),
    .io_flow(x455_mul_1_io_flow),
    .io_result(x455_mul_1_io_result)
  );
  x344_sum x456_sum_1 ( // @[Math.scala 150:24:@40539.4]
    .clock(x456_sum_1_clock),
    .reset(x456_sum_1_reset),
    .io_a(x456_sum_1_io_a),
    .io_b(x456_sum_1_io_b),
    .io_flow(x456_sum_1_io_flow),
    .io_result(x456_sum_1_io_result)
  );
  RetimeWrapper_316 RetimeWrapper_90 ( // @[package.scala 93:22:@40549.4]
    .clock(RetimeWrapper_90_clock),
    .reset(RetimeWrapper_90_reset),
    .io_flow(RetimeWrapper_90_io_flow),
    .io_in(RetimeWrapper_90_io_in),
    .io_out(RetimeWrapper_90_io_out)
  );
  RetimeWrapper_281 RetimeWrapper_91 ( // @[package.scala 93:22:@40558.4]
    .clock(RetimeWrapper_91_clock),
    .reset(RetimeWrapper_91_reset),
    .io_flow(RetimeWrapper_91_io_flow),
    .io_in(RetimeWrapper_91_io_in),
    .io_out(RetimeWrapper_91_io_out)
  );
  RetimeWrapper_311 RetimeWrapper_92 ( // @[package.scala 93:22:@40570.4]
    .clock(RetimeWrapper_92_clock),
    .reset(RetimeWrapper_92_reset),
    .io_flow(RetimeWrapper_92_io_flow),
    .io_in(RetimeWrapper_92_io_in),
    .io_out(RetimeWrapper_92_io_out)
  );
  x344_sum x461_sum_1 ( // @[Math.scala 150:24:@40599.4]
    .clock(x461_sum_1_clock),
    .reset(x461_sum_1_reset),
    .io_a(x461_sum_1_io_a),
    .io_b(x461_sum_1_io_b),
    .io_flow(x461_sum_1_io_flow),
    .io_result(x461_sum_1_io_result)
  );
  RetimeWrapper_316 RetimeWrapper_93 ( // @[package.scala 93:22:@40609.4]
    .clock(RetimeWrapper_93_clock),
    .reset(RetimeWrapper_93_reset),
    .io_flow(RetimeWrapper_93_io_flow),
    .io_in(RetimeWrapper_93_io_in),
    .io_out(RetimeWrapper_93_io_out)
  );
  RetimeWrapper_311 RetimeWrapper_94 ( // @[package.scala 93:22:@40621.4]
    .clock(RetimeWrapper_94_clock),
    .reset(RetimeWrapper_94_reset),
    .io_flow(RetimeWrapper_94_io_flow),
    .io_in(RetimeWrapper_94_io_in),
    .io_out(RetimeWrapper_94_io_out)
  );
  x344_sum x466_sum_1 ( // @[Math.scala 150:24:@40648.4]
    .clock(x466_sum_1_clock),
    .reset(x466_sum_1_reset),
    .io_a(x466_sum_1_io_a),
    .io_b(x466_sum_1_io_b),
    .io_flow(x466_sum_1_io_flow),
    .io_result(x466_sum_1_io_result)
  );
  RetimeWrapper_316 RetimeWrapper_95 ( // @[package.scala 93:22:@40658.4]
    .clock(RetimeWrapper_95_clock),
    .reset(RetimeWrapper_95_reset),
    .io_flow(RetimeWrapper_95_io_flow),
    .io_in(RetimeWrapper_95_io_in),
    .io_out(RetimeWrapper_95_io_out)
  );
  RetimeWrapper_311 RetimeWrapper_96 ( // @[package.scala 93:22:@40670.4]
    .clock(RetimeWrapper_96_clock),
    .reset(RetimeWrapper_96_reset),
    .io_flow(RetimeWrapper_96_io_flow),
    .io_in(RetimeWrapper_96_io_in),
    .io_out(RetimeWrapper_96_io_out)
  );
  x344_sum x471_sum_1 ( // @[Math.scala 150:24:@40697.4]
    .clock(x471_sum_1_clock),
    .reset(x471_sum_1_reset),
    .io_a(x471_sum_1_io_a),
    .io_b(x471_sum_1_io_b),
    .io_flow(x471_sum_1_io_flow),
    .io_result(x471_sum_1_io_result)
  );
  RetimeWrapper_316 RetimeWrapper_97 ( // @[package.scala 93:22:@40707.4]
    .clock(RetimeWrapper_97_clock),
    .reset(RetimeWrapper_97_reset),
    .io_flow(RetimeWrapper_97_io_flow),
    .io_in(RetimeWrapper_97_io_in),
    .io_out(RetimeWrapper_97_io_out)
  );
  RetimeWrapper_311 RetimeWrapper_98 ( // @[package.scala 93:22:@40719.4]
    .clock(RetimeWrapper_98_clock),
    .reset(RetimeWrapper_98_reset),
    .io_flow(RetimeWrapper_98_io_flow),
    .io_in(RetimeWrapper_98_io_in),
    .io_out(RetimeWrapper_98_io_out)
  );
  x344_sum x476_sum_1 ( // @[Math.scala 150:24:@40746.4]
    .clock(x476_sum_1_clock),
    .reset(x476_sum_1_reset),
    .io_a(x476_sum_1_io_a),
    .io_b(x476_sum_1_io_b),
    .io_flow(x476_sum_1_io_flow),
    .io_result(x476_sum_1_io_result)
  );
  RetimeWrapper_316 RetimeWrapper_99 ( // @[package.scala 93:22:@40756.4]
    .clock(RetimeWrapper_99_clock),
    .reset(RetimeWrapper_99_reset),
    .io_flow(RetimeWrapper_99_io_flow),
    .io_in(RetimeWrapper_99_io_in),
    .io_out(RetimeWrapper_99_io_out)
  );
  RetimeWrapper_311 RetimeWrapper_100 ( // @[package.scala 93:22:@40768.4]
    .clock(RetimeWrapper_100_clock),
    .reset(RetimeWrapper_100_reset),
    .io_flow(RetimeWrapper_100_io_flow),
    .io_in(RetimeWrapper_100_io_in),
    .io_out(RetimeWrapper_100_io_out)
  );
  x344_sum x481_sum_1 ( // @[Math.scala 150:24:@40795.4]
    .clock(x481_sum_1_clock),
    .reset(x481_sum_1_reset),
    .io_a(x481_sum_1_io_a),
    .io_b(x481_sum_1_io_b),
    .io_flow(x481_sum_1_io_flow),
    .io_result(x481_sum_1_io_result)
  );
  RetimeWrapper_316 RetimeWrapper_101 ( // @[package.scala 93:22:@40805.4]
    .clock(RetimeWrapper_101_clock),
    .reset(RetimeWrapper_101_reset),
    .io_flow(RetimeWrapper_101_io_flow),
    .io_in(RetimeWrapper_101_io_in),
    .io_out(RetimeWrapper_101_io_out)
  );
  RetimeWrapper_311 RetimeWrapper_102 ( // @[package.scala 93:22:@40817.4]
    .clock(RetimeWrapper_102_clock),
    .reset(RetimeWrapper_102_reset),
    .io_flow(RetimeWrapper_102_io_flow),
    .io_in(RetimeWrapper_102_io_in),
    .io_out(RetimeWrapper_102_io_out)
  );
  RetimeWrapper_419 RetimeWrapper_103 ( // @[package.scala 93:22:@40840.4]
    .clock(RetimeWrapper_103_clock),
    .reset(RetimeWrapper_103_reset),
    .io_flow(RetimeWrapper_103_io_flow),
    .io_in(RetimeWrapper_103_io_in),
    .io_out(RetimeWrapper_103_io_out)
  );
  RetimeWrapper_419 RetimeWrapper_104 ( // @[package.scala 93:22:@40852.4]
    .clock(RetimeWrapper_104_clock),
    .reset(RetimeWrapper_104_reset),
    .io_flow(RetimeWrapper_104_io_flow),
    .io_in(RetimeWrapper_104_io_in),
    .io_out(RetimeWrapper_104_io_out)
  );
  RetimeWrapper_421 RetimeWrapper_105 ( // @[package.scala 93:22:@40864.4]
    .clock(RetimeWrapper_105_clock),
    .reset(RetimeWrapper_105_reset),
    .io_flow(RetimeWrapper_105_io_flow),
    .io_in(RetimeWrapper_105_io_in),
    .io_out(RetimeWrapper_105_io_out)
  );
  RetimeWrapper_419 RetimeWrapper_106 ( // @[package.scala 93:22:@40876.4]
    .clock(RetimeWrapper_106_clock),
    .reset(RetimeWrapper_106_reset),
    .io_flow(RetimeWrapper_106_io_flow),
    .io_in(RetimeWrapper_106_io_in),
    .io_out(RetimeWrapper_106_io_out)
  );
  RetimeWrapper_419 RetimeWrapper_107 ( // @[package.scala 93:22:@40888.4]
    .clock(RetimeWrapper_107_clock),
    .reset(RetimeWrapper_107_reset),
    .io_flow(RetimeWrapper_107_io_flow),
    .io_in(RetimeWrapper_107_io_in),
    .io_out(RetimeWrapper_107_io_out)
  );
  RetimeWrapper_424 RetimeWrapper_108 ( // @[package.scala 93:22:@40898.4]
    .clock(RetimeWrapper_108_clock),
    .reset(RetimeWrapper_108_reset),
    .io_flow(RetimeWrapper_108_io_flow),
    .io_in(RetimeWrapper_108_io_in),
    .io_out(RetimeWrapper_108_io_out)
  );
  RetimeWrapper_20 RetimeWrapper_109 ( // @[package.scala 93:22:@40907.4]
    .clock(RetimeWrapper_109_clock),
    .reset(RetimeWrapper_109_reset),
    .io_flow(RetimeWrapper_109_io_flow),
    .io_in(RetimeWrapper_109_io_in),
    .io_out(RetimeWrapper_109_io_out)
  );
  x489_x11 x489_x11_1 ( // @[Math.scala 150:24:@40916.4]
    .io_a(x489_x11_1_io_a),
    .io_b(x489_x11_1_io_b),
    .io_result(x489_x11_1_io_result)
  );
  RetimeWrapper_424 RetimeWrapper_110 ( // @[package.scala 93:22:@40926.4]
    .clock(RetimeWrapper_110_clock),
    .reset(RetimeWrapper_110_reset),
    .io_flow(RetimeWrapper_110_io_flow),
    .io_in(RetimeWrapper_110_io_in),
    .io_out(RetimeWrapper_110_io_out)
  );
  RetimeWrapper_20 RetimeWrapper_111 ( // @[package.scala 93:22:@40935.4]
    .clock(RetimeWrapper_111_clock),
    .reset(RetimeWrapper_111_reset),
    .io_flow(RetimeWrapper_111_io_flow),
    .io_in(RetimeWrapper_111_io_in),
    .io_out(RetimeWrapper_111_io_out)
  );
  x489_x11 x490_x12_1 ( // @[Math.scala 150:24:@40944.4]
    .io_a(x490_x12_1_io_a),
    .io_b(x490_x12_1_io_b),
    .io_result(x490_x12_1_io_result)
  );
  x489_x11 x491_x11_1 ( // @[Math.scala 150:24:@40954.4]
    .io_a(x491_x11_1_io_a),
    .io_b(x491_x11_1_io_b),
    .io_result(x491_x11_1_io_result)
  );
  RetimeWrapper_20 RetimeWrapper_112 ( // @[package.scala 93:22:@40964.4]
    .clock(RetimeWrapper_112_clock),
    .reset(RetimeWrapper_112_reset),
    .io_flow(RetimeWrapper_112_io_flow),
    .io_in(RetimeWrapper_112_io_in),
    .io_out(RetimeWrapper_112_io_out)
  );
  x489_x11 x492_x12_1 ( // @[Math.scala 150:24:@40973.4]
    .io_a(x492_x12_1_io_a),
    .io_b(x492_x12_1_io_b),
    .io_result(x492_x12_1_io_result)
  );
  RetimeWrapper_424 RetimeWrapper_113 ( // @[package.scala 93:22:@40983.4]
    .clock(RetimeWrapper_113_clock),
    .reset(RetimeWrapper_113_reset),
    .io_flow(RetimeWrapper_113_io_flow),
    .io_in(RetimeWrapper_113_io_in),
    .io_out(RetimeWrapper_113_io_out)
  );
  RetimeWrapper_424 RetimeWrapper_114 ( // @[package.scala 93:22:@40992.4]
    .clock(RetimeWrapper_114_clock),
    .reset(RetimeWrapper_114_reset),
    .io_flow(RetimeWrapper_114_io_flow),
    .io_in(RetimeWrapper_114_io_in),
    .io_out(RetimeWrapper_114_io_out)
  );
  x489_x11 x493_x11_1 ( // @[Math.scala 150:24:@41001.4]
    .io_a(x493_x11_1_io_a),
    .io_b(x493_x11_1_io_b),
    .io_result(x493_x11_1_io_result)
  );
  x489_x11 x494_x12_1 ( // @[Math.scala 150:24:@41011.4]
    .io_a(x494_x12_1_io_a),
    .io_b(x494_x12_1_io_b),
    .io_result(x494_x12_1_io_result)
  );
  RetimeWrapper_431 RetimeWrapper_115 ( // @[package.scala 93:22:@41021.4]
    .clock(RetimeWrapper_115_clock),
    .reset(RetimeWrapper_115_reset),
    .io_flow(RetimeWrapper_115_io_flow),
    .io_in(RetimeWrapper_115_io_in),
    .io_out(RetimeWrapper_115_io_out)
  );
  x489_x11 x495_x11_1 ( // @[Math.scala 150:24:@41032.4]
    .io_a(x495_x11_1_io_a),
    .io_b(x495_x11_1_io_b),
    .io_result(x495_x11_1_io_result)
  );
  RetimeWrapper_432 RetimeWrapper_116 ( // @[package.scala 93:22:@41042.4]
    .clock(RetimeWrapper_116_clock),
    .reset(RetimeWrapper_116_reset),
    .io_flow(RetimeWrapper_116_io_flow),
    .io_in(RetimeWrapper_116_io_in),
    .io_out(RetimeWrapper_116_io_out)
  );
  x496_sum x496_sum_1 ( // @[Math.scala 150:24:@41051.4]
    .clock(x496_sum_1_clock),
    .reset(x496_sum_1_reset),
    .io_a(x496_sum_1_io_a),
    .io_b(x496_sum_1_io_b),
    .io_flow(x496_sum_1_io_flow),
    .io_result(x496_sum_1_io_result)
  );
  RetimeWrapper_419 RetimeWrapper_117 ( // @[package.scala 93:22:@41070.4]
    .clock(RetimeWrapper_117_clock),
    .reset(RetimeWrapper_117_reset),
    .io_flow(RetimeWrapper_117_io_flow),
    .io_in(RetimeWrapper_117_io_in),
    .io_out(RetimeWrapper_117_io_out)
  );
  RetimeWrapper_419 RetimeWrapper_118 ( // @[package.scala 93:22:@41082.4]
    .clock(RetimeWrapper_118_clock),
    .reset(RetimeWrapper_118_reset),
    .io_flow(RetimeWrapper_118_io_flow),
    .io_in(RetimeWrapper_118_io_in),
    .io_out(RetimeWrapper_118_io_out)
  );
  RetimeWrapper_421 RetimeWrapper_119 ( // @[package.scala 93:22:@41094.4]
    .clock(RetimeWrapper_119_clock),
    .reset(RetimeWrapper_119_reset),
    .io_flow(RetimeWrapper_119_io_flow),
    .io_in(RetimeWrapper_119_io_in),
    .io_out(RetimeWrapper_119_io_out)
  );
  RetimeWrapper_419 RetimeWrapper_120 ( // @[package.scala 93:22:@41106.4]
    .clock(RetimeWrapper_120_clock),
    .reset(RetimeWrapper_120_reset),
    .io_flow(RetimeWrapper_120_io_flow),
    .io_in(RetimeWrapper_120_io_in),
    .io_out(RetimeWrapper_120_io_out)
  );
  RetimeWrapper_419 RetimeWrapper_121 ( // @[package.scala 93:22:@41118.4]
    .clock(RetimeWrapper_121_clock),
    .reset(RetimeWrapper_121_reset),
    .io_flow(RetimeWrapper_121_io_flow),
    .io_in(RetimeWrapper_121_io_in),
    .io_out(RetimeWrapper_121_io_out)
  );
  RetimeWrapper_20 RetimeWrapper_122 ( // @[package.scala 93:22:@41128.4]
    .clock(RetimeWrapper_122_clock),
    .reset(RetimeWrapper_122_reset),
    .io_flow(RetimeWrapper_122_io_flow),
    .io_in(RetimeWrapper_122_io_in),
    .io_out(RetimeWrapper_122_io_out)
  );
  RetimeWrapper_424 RetimeWrapper_123 ( // @[package.scala 93:22:@41137.4]
    .clock(RetimeWrapper_123_clock),
    .reset(RetimeWrapper_123_reset),
    .io_flow(RetimeWrapper_123_io_flow),
    .io_in(RetimeWrapper_123_io_in),
    .io_out(RetimeWrapper_123_io_out)
  );
  x489_x11 x503_x11_1 ( // @[Math.scala 150:24:@41146.4]
    .io_a(x503_x11_1_io_a),
    .io_b(x503_x11_1_io_b),
    .io_result(x503_x11_1_io_result)
  );
  RetimeWrapper_424 RetimeWrapper_124 ( // @[package.scala 93:22:@41156.4]
    .clock(RetimeWrapper_124_clock),
    .reset(RetimeWrapper_124_reset),
    .io_flow(RetimeWrapper_124_io_flow),
    .io_in(RetimeWrapper_124_io_in),
    .io_out(RetimeWrapper_124_io_out)
  );
  RetimeWrapper_20 RetimeWrapper_125 ( // @[package.scala 93:22:@41165.4]
    .clock(RetimeWrapper_125_clock),
    .reset(RetimeWrapper_125_reset),
    .io_flow(RetimeWrapper_125_io_flow),
    .io_in(RetimeWrapper_125_io_in),
    .io_out(RetimeWrapper_125_io_out)
  );
  x489_x11 x504_x12_1 ( // @[Math.scala 150:24:@41174.4]
    .io_a(x504_x12_1_io_a),
    .io_b(x504_x12_1_io_b),
    .io_result(x504_x12_1_io_result)
  );
  x489_x11 x505_x11_1 ( // @[Math.scala 150:24:@41184.4]
    .io_a(x505_x11_1_io_a),
    .io_b(x505_x11_1_io_b),
    .io_result(x505_x11_1_io_result)
  );
  RetimeWrapper_20 RetimeWrapper_126 ( // @[package.scala 93:22:@41194.4]
    .clock(RetimeWrapper_126_clock),
    .reset(RetimeWrapper_126_reset),
    .io_flow(RetimeWrapper_126_io_flow),
    .io_in(RetimeWrapper_126_io_in),
    .io_out(RetimeWrapper_126_io_out)
  );
  x489_x11 x506_x12_1 ( // @[Math.scala 150:24:@41203.4]
    .io_a(x506_x12_1_io_a),
    .io_b(x506_x12_1_io_b),
    .io_result(x506_x12_1_io_result)
  );
  RetimeWrapper_424 RetimeWrapper_127 ( // @[package.scala 93:22:@41213.4]
    .clock(RetimeWrapper_127_clock),
    .reset(RetimeWrapper_127_reset),
    .io_flow(RetimeWrapper_127_io_flow),
    .io_in(RetimeWrapper_127_io_in),
    .io_out(RetimeWrapper_127_io_out)
  );
  RetimeWrapper_424 RetimeWrapper_128 ( // @[package.scala 93:22:@41222.4]
    .clock(RetimeWrapper_128_clock),
    .reset(RetimeWrapper_128_reset),
    .io_flow(RetimeWrapper_128_io_flow),
    .io_in(RetimeWrapper_128_io_in),
    .io_out(RetimeWrapper_128_io_out)
  );
  x489_x11 x507_x11_1 ( // @[Math.scala 150:24:@41231.4]
    .io_a(x507_x11_1_io_a),
    .io_b(x507_x11_1_io_b),
    .io_result(x507_x11_1_io_result)
  );
  x489_x11 x508_x12_1 ( // @[Math.scala 150:24:@41241.4]
    .io_a(x508_x12_1_io_a),
    .io_b(x508_x12_1_io_b),
    .io_result(x508_x12_1_io_result)
  );
  RetimeWrapper_431 RetimeWrapper_129 ( // @[package.scala 93:22:@41251.4]
    .clock(RetimeWrapper_129_clock),
    .reset(RetimeWrapper_129_reset),
    .io_flow(RetimeWrapper_129_io_flow),
    .io_in(RetimeWrapper_129_io_in),
    .io_out(RetimeWrapper_129_io_out)
  );
  x489_x11 x509_x11_1 ( // @[Math.scala 150:24:@41260.4]
    .io_a(x509_x11_1_io_a),
    .io_b(x509_x11_1_io_b),
    .io_result(x509_x11_1_io_result)
  );
  RetimeWrapper_432 RetimeWrapper_130 ( // @[package.scala 93:22:@41270.4]
    .clock(RetimeWrapper_130_clock),
    .reset(RetimeWrapper_130_reset),
    .io_flow(RetimeWrapper_130_io_flow),
    .io_in(RetimeWrapper_130_io_in),
    .io_out(RetimeWrapper_130_io_out)
  );
  x496_sum x510_sum_1 ( // @[Math.scala 150:24:@41279.4]
    .clock(x510_sum_1_clock),
    .reset(x510_sum_1_reset),
    .io_a(x510_sum_1_io_a),
    .io_b(x510_sum_1_io_b),
    .io_flow(x510_sum_1_io_flow),
    .io_result(x510_sum_1_io_result)
  );
  RetimeWrapper_419 RetimeWrapper_131 ( // @[package.scala 93:22:@41298.4]
    .clock(RetimeWrapper_131_clock),
    .reset(RetimeWrapper_131_reset),
    .io_flow(RetimeWrapper_131_io_flow),
    .io_in(RetimeWrapper_131_io_in),
    .io_out(RetimeWrapper_131_io_out)
  );
  RetimeWrapper_421 RetimeWrapper_132 ( // @[package.scala 93:22:@41310.4]
    .clock(RetimeWrapper_132_clock),
    .reset(RetimeWrapper_132_reset),
    .io_flow(RetimeWrapper_132_io_flow),
    .io_in(RetimeWrapper_132_io_in),
    .io_out(RetimeWrapper_132_io_out)
  );
  RetimeWrapper_419 RetimeWrapper_133 ( // @[package.scala 93:22:@41322.4]
    .clock(RetimeWrapper_133_clock),
    .reset(RetimeWrapper_133_reset),
    .io_flow(RetimeWrapper_133_io_flow),
    .io_in(RetimeWrapper_133_io_in),
    .io_out(RetimeWrapper_133_io_out)
  );
  RetimeWrapper_419 RetimeWrapper_134 ( // @[package.scala 93:22:@41334.4]
    .clock(RetimeWrapper_134_clock),
    .reset(RetimeWrapper_134_reset),
    .io_flow(RetimeWrapper_134_io_flow),
    .io_in(RetimeWrapper_134_io_in),
    .io_out(RetimeWrapper_134_io_out)
  );
  RetimeWrapper_20 RetimeWrapper_135 ( // @[package.scala 93:22:@41344.4]
    .clock(RetimeWrapper_135_clock),
    .reset(RetimeWrapper_135_reset),
    .io_flow(RetimeWrapper_135_io_flow),
    .io_in(RetimeWrapper_135_io_in),
    .io_out(RetimeWrapper_135_io_out)
  );
  x489_x11 x516_x11_1 ( // @[Math.scala 150:24:@41353.4]
    .io_a(x516_x11_1_io_a),
    .io_b(x516_x11_1_io_b),
    .io_result(x516_x11_1_io_result)
  );
  RetimeWrapper_20 RetimeWrapper_136 ( // @[package.scala 93:22:@41363.4]
    .clock(RetimeWrapper_136_clock),
    .reset(RetimeWrapper_136_reset),
    .io_flow(RetimeWrapper_136_io_flow),
    .io_in(RetimeWrapper_136_io_in),
    .io_out(RetimeWrapper_136_io_out)
  );
  RetimeWrapper_424 RetimeWrapper_137 ( // @[package.scala 93:22:@41372.4]
    .clock(RetimeWrapper_137_clock),
    .reset(RetimeWrapper_137_reset),
    .io_flow(RetimeWrapper_137_io_flow),
    .io_in(RetimeWrapper_137_io_in),
    .io_out(RetimeWrapper_137_io_out)
  );
  x489_x11 x517_x12_1 ( // @[Math.scala 150:24:@41381.4]
    .io_a(x517_x12_1_io_a),
    .io_b(x517_x12_1_io_b),
    .io_result(x517_x12_1_io_result)
  );
  x489_x11 x518_x11_1 ( // @[Math.scala 150:24:@41391.4]
    .io_a(x518_x11_1_io_a),
    .io_b(x518_x11_1_io_b),
    .io_result(x518_x11_1_io_result)
  );
  RetimeWrapper_20 RetimeWrapper_138 ( // @[package.scala 93:22:@41401.4]
    .clock(RetimeWrapper_138_clock),
    .reset(RetimeWrapper_138_reset),
    .io_flow(RetimeWrapper_138_io_flow),
    .io_in(RetimeWrapper_138_io_in),
    .io_out(RetimeWrapper_138_io_out)
  );
  x489_x11 x519_x12_1 ( // @[Math.scala 150:24:@41410.4]
    .io_a(x519_x12_1_io_a),
    .io_b(x519_x12_1_io_b),
    .io_result(x519_x12_1_io_result)
  );
  RetimeWrapper_424 RetimeWrapper_139 ( // @[package.scala 93:22:@41420.4]
    .clock(RetimeWrapper_139_clock),
    .reset(RetimeWrapper_139_reset),
    .io_flow(RetimeWrapper_139_io_flow),
    .io_in(RetimeWrapper_139_io_in),
    .io_out(RetimeWrapper_139_io_out)
  );
  RetimeWrapper_424 RetimeWrapper_140 ( // @[package.scala 93:22:@41429.4]
    .clock(RetimeWrapper_140_clock),
    .reset(RetimeWrapper_140_reset),
    .io_flow(RetimeWrapper_140_io_flow),
    .io_in(RetimeWrapper_140_io_in),
    .io_out(RetimeWrapper_140_io_out)
  );
  x489_x11 x520_x11_1 ( // @[Math.scala 150:24:@41438.4]
    .io_a(x520_x11_1_io_a),
    .io_b(x520_x11_1_io_b),
    .io_result(x520_x11_1_io_result)
  );
  x489_x11 x521_x12_1 ( // @[Math.scala 150:24:@41448.4]
    .io_a(x521_x12_1_io_a),
    .io_b(x521_x12_1_io_b),
    .io_result(x521_x12_1_io_result)
  );
  RetimeWrapper_431 RetimeWrapper_141 ( // @[package.scala 93:22:@41458.4]
    .clock(RetimeWrapper_141_clock),
    .reset(RetimeWrapper_141_reset),
    .io_flow(RetimeWrapper_141_io_flow),
    .io_in(RetimeWrapper_141_io_in),
    .io_out(RetimeWrapper_141_io_out)
  );
  x489_x11 x522_x11_1 ( // @[Math.scala 150:24:@41467.4]
    .io_a(x522_x11_1_io_a),
    .io_b(x522_x11_1_io_b),
    .io_result(x522_x11_1_io_result)
  );
  RetimeWrapper_432 RetimeWrapper_142 ( // @[package.scala 93:22:@41477.4]
    .clock(RetimeWrapper_142_clock),
    .reset(RetimeWrapper_142_reset),
    .io_flow(RetimeWrapper_142_io_flow),
    .io_in(RetimeWrapper_142_io_in),
    .io_out(RetimeWrapper_142_io_out)
  );
  x496_sum x523_sum_1 ( // @[Math.scala 150:24:@41486.4]
    .clock(x523_sum_1_clock),
    .reset(x523_sum_1_reset),
    .io_a(x523_sum_1_io_a),
    .io_b(x523_sum_1_io_b),
    .io_flow(x523_sum_1_io_flow),
    .io_result(x523_sum_1_io_result)
  );
  RetimeWrapper_419 RetimeWrapper_143 ( // @[package.scala 93:22:@41507.4]
    .clock(RetimeWrapper_143_clock),
    .reset(RetimeWrapper_143_reset),
    .io_flow(RetimeWrapper_143_io_flow),
    .io_in(RetimeWrapper_143_io_in),
    .io_out(RetimeWrapper_143_io_out)
  );
  RetimeWrapper_421 RetimeWrapper_144 ( // @[package.scala 93:22:@41519.4]
    .clock(RetimeWrapper_144_clock),
    .reset(RetimeWrapper_144_reset),
    .io_flow(RetimeWrapper_144_io_flow),
    .io_in(RetimeWrapper_144_io_in),
    .io_out(RetimeWrapper_144_io_out)
  );
  RetimeWrapper_419 RetimeWrapper_145 ( // @[package.scala 93:22:@41531.4]
    .clock(RetimeWrapper_145_clock),
    .reset(RetimeWrapper_145_reset),
    .io_flow(RetimeWrapper_145_io_flow),
    .io_in(RetimeWrapper_145_io_in),
    .io_out(RetimeWrapper_145_io_out)
  );
  RetimeWrapper_419 RetimeWrapper_146 ( // @[package.scala 93:22:@41543.4]
    .clock(RetimeWrapper_146_clock),
    .reset(RetimeWrapper_146_reset),
    .io_flow(RetimeWrapper_146_io_flow),
    .io_in(RetimeWrapper_146_io_in),
    .io_out(RetimeWrapper_146_io_out)
  );
  RetimeWrapper_20 RetimeWrapper_147 ( // @[package.scala 93:22:@41553.4]
    .clock(RetimeWrapper_147_clock),
    .reset(RetimeWrapper_147_reset),
    .io_flow(RetimeWrapper_147_io_flow),
    .io_in(RetimeWrapper_147_io_in),
    .io_out(RetimeWrapper_147_io_out)
  );
  x489_x11 x529_x11_1 ( // @[Math.scala 150:24:@41562.4]
    .io_a(x529_x11_1_io_a),
    .io_b(x529_x11_1_io_b),
    .io_result(x529_x11_1_io_result)
  );
  RetimeWrapper_20 RetimeWrapper_148 ( // @[package.scala 93:22:@41572.4]
    .clock(RetimeWrapper_148_clock),
    .reset(RetimeWrapper_148_reset),
    .io_flow(RetimeWrapper_148_io_flow),
    .io_in(RetimeWrapper_148_io_in),
    .io_out(RetimeWrapper_148_io_out)
  );
  RetimeWrapper_424 RetimeWrapper_149 ( // @[package.scala 93:22:@41581.4]
    .clock(RetimeWrapper_149_clock),
    .reset(RetimeWrapper_149_reset),
    .io_flow(RetimeWrapper_149_io_flow),
    .io_in(RetimeWrapper_149_io_in),
    .io_out(RetimeWrapper_149_io_out)
  );
  x489_x11 x530_x12_1 ( // @[Math.scala 150:24:@41590.4]
    .io_a(x530_x12_1_io_a),
    .io_b(x530_x12_1_io_b),
    .io_result(x530_x12_1_io_result)
  );
  x489_x11 x531_x11_1 ( // @[Math.scala 150:24:@41600.4]
    .io_a(x531_x11_1_io_a),
    .io_b(x531_x11_1_io_b),
    .io_result(x531_x11_1_io_result)
  );
  RetimeWrapper_20 RetimeWrapper_150 ( // @[package.scala 93:22:@41610.4]
    .clock(RetimeWrapper_150_clock),
    .reset(RetimeWrapper_150_reset),
    .io_flow(RetimeWrapper_150_io_flow),
    .io_in(RetimeWrapper_150_io_in),
    .io_out(RetimeWrapper_150_io_out)
  );
  x489_x11 x532_x12_1 ( // @[Math.scala 150:24:@41619.4]
    .io_a(x532_x12_1_io_a),
    .io_b(x532_x12_1_io_b),
    .io_result(x532_x12_1_io_result)
  );
  RetimeWrapper_424 RetimeWrapper_151 ( // @[package.scala 93:22:@41629.4]
    .clock(RetimeWrapper_151_clock),
    .reset(RetimeWrapper_151_reset),
    .io_flow(RetimeWrapper_151_io_flow),
    .io_in(RetimeWrapper_151_io_in),
    .io_out(RetimeWrapper_151_io_out)
  );
  RetimeWrapper_424 RetimeWrapper_152 ( // @[package.scala 93:22:@41638.4]
    .clock(RetimeWrapper_152_clock),
    .reset(RetimeWrapper_152_reset),
    .io_flow(RetimeWrapper_152_io_flow),
    .io_in(RetimeWrapper_152_io_in),
    .io_out(RetimeWrapper_152_io_out)
  );
  x489_x11 x533_x11_1 ( // @[Math.scala 150:24:@41647.4]
    .io_a(x533_x11_1_io_a),
    .io_b(x533_x11_1_io_b),
    .io_result(x533_x11_1_io_result)
  );
  x489_x11 x534_x12_1 ( // @[Math.scala 150:24:@41657.4]
    .io_a(x534_x12_1_io_a),
    .io_b(x534_x12_1_io_b),
    .io_result(x534_x12_1_io_result)
  );
  RetimeWrapper_431 RetimeWrapper_153 ( // @[package.scala 93:22:@41667.4]
    .clock(RetimeWrapper_153_clock),
    .reset(RetimeWrapper_153_reset),
    .io_flow(RetimeWrapper_153_io_flow),
    .io_in(RetimeWrapper_153_io_in),
    .io_out(RetimeWrapper_153_io_out)
  );
  x489_x11 x535_x11_1 ( // @[Math.scala 150:24:@41676.4]
    .io_a(x535_x11_1_io_a),
    .io_b(x535_x11_1_io_b),
    .io_result(x535_x11_1_io_result)
  );
  RetimeWrapper_432 RetimeWrapper_154 ( // @[package.scala 93:22:@41686.4]
    .clock(RetimeWrapper_154_clock),
    .reset(RetimeWrapper_154_reset),
    .io_flow(RetimeWrapper_154_io_flow),
    .io_in(RetimeWrapper_154_io_in),
    .io_out(RetimeWrapper_154_io_out)
  );
  x496_sum x536_sum_1 ( // @[Math.scala 150:24:@41695.4]
    .clock(x536_sum_1_clock),
    .reset(x536_sum_1_reset),
    .io_a(x536_sum_1_io_a),
    .io_b(x536_sum_1_io_b),
    .io_flow(x536_sum_1_io_flow),
    .io_result(x536_sum_1_io_result)
  );
  RetimeWrapper_431 RetimeWrapper_155 ( // @[package.scala 93:22:@41712.4]
    .clock(RetimeWrapper_155_clock),
    .reset(RetimeWrapper_155_reset),
    .io_flow(RetimeWrapper_155_io_flow),
    .io_in(RetimeWrapper_155_io_in),
    .io_out(RetimeWrapper_155_io_out)
  );
  RetimeWrapper_431 RetimeWrapper_156 ( // @[package.scala 93:22:@41721.4]
    .clock(RetimeWrapper_156_clock),
    .reset(RetimeWrapper_156_reset),
    .io_flow(RetimeWrapper_156_io_flow),
    .io_in(RetimeWrapper_156_io_in),
    .io_out(RetimeWrapper_156_io_out)
  );
  RetimeWrapper_431 RetimeWrapper_157 ( // @[package.scala 93:22:@41730.4]
    .clock(RetimeWrapper_157_clock),
    .reset(RetimeWrapper_157_reset),
    .io_flow(RetimeWrapper_157_io_flow),
    .io_in(RetimeWrapper_157_io_in),
    .io_out(RetimeWrapper_157_io_out)
  );
  RetimeWrapper_431 RetimeWrapper_158 ( // @[package.scala 93:22:@41739.4]
    .clock(RetimeWrapper_158_clock),
    .reset(RetimeWrapper_158_reset),
    .io_flow(RetimeWrapper_158_io_flow),
    .io_in(RetimeWrapper_158_io_in),
    .io_out(RetimeWrapper_158_io_out)
  );
  RetimeWrapper_269 RetimeWrapper_159 ( // @[package.scala 93:22:@41758.4]
    .clock(RetimeWrapper_159_clock),
    .reset(RetimeWrapper_159_reset),
    .io_flow(RetimeWrapper_159_io_flow),
    .io_in(RetimeWrapper_159_io_in),
    .io_out(RetimeWrapper_159_io_out)
  );
  RetimeWrapper_12 RetimeWrapper_160 ( // @[package.scala 93:22:@41767.4]
    .clock(RetimeWrapper_160_clock),
    .reset(RetimeWrapper_160_reset),
    .io_flow(RetimeWrapper_160_io_flow),
    .io_in(RetimeWrapper_160_io_in),
    .io_out(RetimeWrapper_160_io_out)
  );
  RetimeWrapper_12 RetimeWrapper_161 ( // @[package.scala 93:22:@41776.4]
    .clock(RetimeWrapper_161_clock),
    .reset(RetimeWrapper_161_reset),
    .io_flow(RetimeWrapper_161_io_flow),
    .io_in(RetimeWrapper_161_io_in),
    .io_out(RetimeWrapper_161_io_out)
  );
  RetimeWrapper_12 RetimeWrapper_162 ( // @[package.scala 93:22:@41785.4]
    .clock(RetimeWrapper_162_clock),
    .reset(RetimeWrapper_162_reset),
    .io_flow(RetimeWrapper_162_io_flow),
    .io_in(RetimeWrapper_162_io_in),
    .io_out(RetimeWrapper_162_io_out)
  );
  assign b327 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 62:18:@38584.4]
  assign b328 = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 63:18:@38585.4]
  assign _T_206 = b327 & b328; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 68:30:@38732.4]
  assign _T_207 = _T_206 & io_sigsIn_datapathEn; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 68:37:@38733.4]
  assign _T_211 = io_in_x316_TID == 8'h0; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 70:76:@38738.4]
  assign _T_212 = _T_207 & _T_211; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 70:62:@38739.4]
  assign _T_214 = io_in_x316_TDEST == 8'h0; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 70:101:@38740.4]
  assign x614_x330_D1_0_number = RetimeWrapper_io_out; // @[package.scala 96:25:@38749.4 package.scala 96:25:@38750.4]
  assign b325_number = __io_result; // @[Math.scala 712:22:@38569.4 Math.scala 713:14:@38570.4]
  assign _T_246 = $signed(b325_number); // @[Math.scala 499:52:@38769.4]
  assign x334 = $signed(32'sh1) == $signed(_T_246); // @[Math.scala 499:44:@38777.4]
  assign x335 = $signed(32'sh2) == $signed(_T_246); // @[Math.scala 499:44:@38784.4]
  assign x336 = $signed(32'sh3) == $signed(_T_246); // @[Math.scala 499:44:@38791.4]
  assign _T_293 = x334 ? 32'h1 : 32'h0; // @[Mux.scala 19:72:@38803.4]
  assign _T_295 = x335 ? 32'h2 : 32'h0; // @[Mux.scala 19:72:@38804.4]
  assign _T_297 = x336 ? 32'h3 : 32'h0; // @[Mux.scala 19:72:@38805.4]
  assign _T_299 = _T_293 | _T_295; // @[Mux.scala 19:72:@38807.4]
  assign x337_number = _T_299 | _T_297; // @[Mux.scala 19:72:@38808.4]
  assign _T_311 = $signed(x337_number); // @[Math.scala 406:49:@38818.4]
  assign _T_313 = $signed(_T_311) & $signed(32'sh3); // @[Math.scala 406:56:@38820.4]
  assign _T_314 = $signed(_T_313); // @[Math.scala 406:56:@38821.4]
  assign _T_326 = x337_number[31]; // @[FixedPoint.scala 50:25:@38839.4]
  assign _T_330 = _T_326 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@38841.4]
  assign _T_331 = x337_number[31:2]; // @[FixedPoint.scala 18:52:@38842.4]
  assign _T_372 = ~ io_sigsIn_break; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 121:101:@38943.4]
  assign _T_376 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@38951.4 package.scala 96:25:@38952.4]
  assign _T_378 = io_rr ? _T_376 : 1'h0; // @[implicits.scala 55:10:@38953.4]
  assign _T_379 = _T_372 & _T_378; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 121:118:@38954.4]
  assign _T_381 = _T_379 & _T_372; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 121:207:@38956.4]
  assign _T_382 = _T_381 & io_sigsIn_backpressure; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 121:226:@38957.4]
  assign x620_b327_D24 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@38931.4 package.scala 96:25:@38932.4]
  assign _T_383 = _T_382 & x620_b327_D24; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 121:252:@38958.4]
  assign x619_b328_D24 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@38922.4 package.scala 96:25:@38923.4]
  assign _T_427 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@39058.4 package.scala 96:25:@39059.4]
  assign _T_429 = io_rr ? _T_427 : 1'h0; // @[implicits.scala 55:10:@39060.4]
  assign _T_430 = _T_372 & _T_429; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 144:118:@39061.4]
  assign _T_432 = _T_430 & _T_372; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 144:207:@39063.4]
  assign _T_433 = _T_432 & io_sigsIn_backpressure; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 144:226:@39064.4]
  assign _T_434 = _T_433 & x620_b327_D24; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 144:252:@39065.4]
  assign _T_475 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@39156.4 package.scala 96:25:@39157.4]
  assign _T_477 = io_rr ? _T_475 : 1'h0; // @[implicits.scala 55:10:@39158.4]
  assign _T_478 = _T_372 & _T_477; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 165:118:@39159.4]
  assign _T_480 = _T_478 & _T_372; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 165:207:@39161.4]
  assign _T_481 = _T_480 & io_sigsIn_backpressure; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 165:226:@39162.4]
  assign _T_482 = _T_481 & x620_b327_D24; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 165:252:@39163.4]
  assign _T_523 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@39254.4 package.scala 96:25:@39255.4]
  assign _T_525 = io_rr ? _T_523 : 1'h0; // @[implicits.scala 55:10:@39256.4]
  assign _T_526 = _T_372 & _T_525; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 192:166:@39257.4]
  assign _T_528 = _T_526 & _T_372; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 192:255:@39259.4]
  assign _T_529 = _T_528 & io_sigsIn_backpressure; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 192:274:@39260.4]
  assign _T_530 = _T_529 & x620_b327_D24; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 192:300:@39261.4]
  assign x632_b325_D26_number = RetimeWrapper_22_io_out; // @[package.scala 96:25:@39275.4 package.scala 96:25:@39276.4]
  assign _T_549 = $signed(x632_b325_D26_number); // @[Math.scala 465:37:@39295.4]
  assign x633_x358_rdcol_D26_number = RetimeWrapper_24_io_out; // @[package.scala 96:25:@39312.4 package.scala 96:25:@39313.4]
  assign _T_562 = $signed(x633_x358_rdcol_D26_number); // @[Math.scala 465:37:@39318.4]
  assign x634_x366_D1 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@39335.4 package.scala 96:25:@39336.4]
  assign x367 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@39326.4 package.scala 96:25:@39327.4]
  assign x368 = x634_x366_D1 | x367; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 209:24:@39339.4]
  assign x365_number = x365_1_io_result; // @[Math.scala 370:22:@39289.4 Math.scala 371:14:@39290.4]
  assign _T_581 = $signed(x365_number); // @[Math.scala 406:49:@39348.4]
  assign _T_583 = $signed(_T_581) & $signed(32'sh3); // @[Math.scala 406:56:@39350.4]
  assign _T_584 = $signed(_T_583); // @[Math.scala 406:56:@39351.4]
  assign _T_589 = x365_number[31]; // @[FixedPoint.scala 50:25:@39357.4]
  assign _T_593 = _T_589 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@39359.4]
  assign _T_594 = x365_number[31:2]; // @[FixedPoint.scala 18:52:@39360.4]
  assign _T_638 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@39458.4 package.scala 96:25:@39459.4]
  assign _T_640 = io_rr ? _T_638 : 1'h0; // @[implicits.scala 55:10:@39460.4]
  assign _T_641 = _T_372 & _T_640; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 238:194:@39461.4]
  assign x641_x369_D22 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@39446.4 package.scala 96:25:@39447.4]
  assign _T_642 = _T_641 & x641_x369_D22; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 238:283:@39462.4]
  assign x639_b327_D50 = RetimeWrapper_31_io_out; // @[package.scala 96:25:@39428.4 package.scala 96:25:@39429.4]
  assign _T_643 = _T_642 & x639_b327_D50; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 238:291:@39463.4]
  assign x636_b328_D50 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@39401.4 package.scala 96:25:@39402.4]
  assign x642_x352_rdcol_D26_number = RetimeWrapper_35_io_out; // @[package.scala 96:25:@39479.4 package.scala 96:25:@39480.4]
  assign _T_654 = $signed(x642_x352_rdcol_D26_number); // @[Math.scala 465:37:@39485.4]
  assign x376 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@39493.4 package.scala 96:25:@39494.4]
  assign x377 = x634_x366_D1 | x376; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 246:24:@39497.4]
  assign _T_689 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@39557.4 package.scala 96:25:@39558.4]
  assign _T_691 = io_rr ? _T_689 : 1'h0; // @[implicits.scala 55:10:@39559.4]
  assign _T_692 = _T_372 & _T_691; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 263:194:@39560.4]
  assign x645_x378_D22 = RetimeWrapper_39_io_out; // @[package.scala 96:25:@39536.4 package.scala 96:25:@39537.4]
  assign _T_693 = _T_692 & x645_x378_D22; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 263:283:@39561.4]
  assign _T_694 = _T_693 & x639_b327_D50; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 263:291:@39562.4]
  assign x647_x346_rdcol_D26_number = RetimeWrapper_42_io_out; // @[package.scala 96:25:@39578.4 package.scala 96:25:@39579.4]
  assign _T_705 = $signed(x647_x346_rdcol_D26_number); // @[Math.scala 465:37:@39584.4]
  assign x382 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@39592.4 package.scala 96:25:@39593.4]
  assign x383 = x634_x366_D1 | x382; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 271:24:@39596.4]
  assign _T_740 = RetimeWrapper_48_io_out; // @[package.scala 96:25:@39656.4 package.scala 96:25:@39657.4]
  assign _T_742 = io_rr ? _T_740 : 1'h0; // @[implicits.scala 55:10:@39658.4]
  assign _T_743 = _T_372 & _T_742; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 288:194:@39659.4]
  assign x650_x384_D22 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@39635.4 package.scala 96:25:@39636.4]
  assign _T_744 = _T_743 & x650_x384_D22; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 288:283:@39660.4]
  assign _T_745 = _T_744 & x639_b327_D50; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 288:291:@39661.4]
  assign x652_b326_D26_number = RetimeWrapper_49_io_out; // @[package.scala 96:25:@39677.4 package.scala 96:25:@39678.4]
  assign _T_758 = $signed(x652_b326_D26_number); // @[Math.scala 465:37:@39685.4]
  assign x366 = RetimeWrapper_23_io_out; // @[package.scala 96:25:@39303.4 package.scala 96:25:@39304.4]
  assign x388 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@39693.4 package.scala 96:25:@39694.4]
  assign x389 = x366 | x388; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 304:59:@39697.4]
  assign _T_793 = RetimeWrapper_55_io_out; // @[package.scala 96:25:@39757.4 package.scala 96:25:@39758.4]
  assign _T_795 = io_rr ? _T_793 : 1'h0; // @[implicits.scala 55:10:@39759.4]
  assign _T_796 = _T_372 & _T_795; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 321:194:@39760.4]
  assign x656_x390_D23 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@39745.4 package.scala 96:25:@39746.4]
  assign _T_797 = _T_796 & x656_x390_D23; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 321:283:@39761.4]
  assign _T_798 = _T_797 & x639_b327_D50; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 321:291:@39762.4]
  assign x394_rdcol_number = x394_rdcol_1_io_result; // @[Math.scala 154:22:@39781.4 Math.scala 155:14:@39782.4]
  assign _T_813 = $signed(x394_rdcol_number); // @[Math.scala 465:37:@39787.4]
  assign x395 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@39795.4 package.scala 96:25:@39796.4]
  assign x396 = x634_x366_D1 | x395; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 329:59:@39799.4]
  assign _T_862 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@39883.4 package.scala 96:25:@39884.4]
  assign _T_864 = io_rr ? _T_862 : 1'h0; // @[implicits.scala 55:10:@39885.4]
  assign _T_865 = _T_372 & _T_864; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 350:194:@39886.4]
  assign x658_x397_D22 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@39853.4 package.scala 96:25:@39854.4]
  assign _T_866 = _T_865 & x658_x397_D22; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 350:283:@39887.4]
  assign _T_867 = _T_866 & x639_b327_D50; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 350:291:@39888.4]
  assign x403_rdcol_number = x403_rdcol_1_io_result; // @[Math.scala 154:22:@39907.4 Math.scala 155:14:@39908.4]
  assign _T_882 = $signed(x403_rdcol_number); // @[Math.scala 465:37:@39913.4]
  assign x404 = RetimeWrapper_62_io_out; // @[package.scala 96:25:@39921.4 package.scala 96:25:@39922.4]
  assign x405 = x634_x366_D1 | x404; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 358:59:@39925.4]
  assign _T_931 = RetimeWrapper_67_io_out; // @[package.scala 96:25:@40009.4 package.scala 96:25:@40010.4]
  assign _T_933 = io_rr ? _T_931 : 1'h0; // @[implicits.scala 55:10:@40011.4]
  assign _T_934 = _T_372 & _T_933; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 379:194:@40012.4]
  assign x663_x406_D22 = RetimeWrapper_65_io_out; // @[package.scala 96:25:@39988.4 package.scala 96:25:@39989.4]
  assign _T_935 = _T_934 & x663_x406_D22; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 379:283:@40013.4]
  assign _T_936 = _T_935 & x639_b327_D50; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 379:291:@40014.4]
  assign x412_rdrow_number = x412_rdrow_1_io_result; // @[Math.scala 195:22:@40033.4 Math.scala 196:14:@40034.4]
  assign _T_958 = $signed(x412_rdrow_number); // @[Math.scala 465:37:@40051.4]
  assign x414 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@40059.4 package.scala 96:25:@40060.4]
  assign x415 = x414 | x367; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 389:24:@40063.4]
  assign x413_number = x413_1_io_result; // @[Math.scala 370:22:@40045.4 Math.scala 371:14:@40046.4]
  assign _T_974 = $signed(x413_number); // @[Math.scala 406:49:@40072.4]
  assign _T_976 = $signed(_T_974) & $signed(32'sh3); // @[Math.scala 406:56:@40074.4]
  assign _T_977 = $signed(_T_976); // @[Math.scala 406:56:@40075.4]
  assign _T_982 = x413_number[31]; // @[FixedPoint.scala 50:25:@40081.4]
  assign _T_986 = _T_982 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@40083.4]
  assign _T_987 = x413_number[31:2]; // @[FixedPoint.scala 18:52:@40084.4]
  assign _T_1019 = RetimeWrapper_72_io_out; // @[package.scala 96:25:@40146.4 package.scala 96:25:@40147.4]
  assign _T_1021 = io_rr ? _T_1019 : 1'h0; // @[implicits.scala 55:10:@40148.4]
  assign _T_1022 = _T_372 & _T_1021; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 410:194:@40149.4]
  assign x666_x416_D22 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@40125.4 package.scala 96:25:@40126.4]
  assign _T_1023 = _T_1022 & x666_x416_D22; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 410:283:@40150.4]
  assign _T_1024 = _T_1023 & x639_b327_D50; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 410:291:@40151.4]
  assign x423 = x414 | x376; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 420:59:@40162.4]
  assign _T_1053 = RetimeWrapper_75_io_out; // @[package.scala 96:25:@40206.4 package.scala 96:25:@40207.4]
  assign _T_1055 = io_rr ? _T_1053 : 1'h0; // @[implicits.scala 55:10:@40208.4]
  assign _T_1056 = _T_372 & _T_1055; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 435:194:@40209.4]
  assign x669_x424_D22 = RetimeWrapper_74_io_out; // @[package.scala 96:25:@40194.4 package.scala 96:25:@40195.4]
  assign _T_1057 = _T_1056 & x669_x424_D22; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 435:283:@40210.4]
  assign _T_1058 = _T_1057 & x639_b327_D50; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 435:291:@40211.4]
  assign x428 = x414 | x382; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 439:59:@40222.4]
  assign _T_1085 = RetimeWrapper_78_io_out; // @[package.scala 96:25:@40264.4 package.scala 96:25:@40265.4]
  assign _T_1087 = io_rr ? _T_1085 : 1'h0; // @[implicits.scala 55:10:@40266.4]
  assign _T_1088 = _T_372 & _T_1087; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 452:194:@40267.4]
  assign x671_x429_D22 = RetimeWrapper_77_io_out; // @[package.scala 96:25:@40252.4 package.scala 96:25:@40253.4]
  assign _T_1089 = _T_1088 & x671_x429_D22; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 452:283:@40268.4]
  assign _T_1090 = _T_1089 & x639_b327_D50; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 452:291:@40269.4]
  assign x672_x388_D1 = RetimeWrapper_79_io_out; // @[package.scala 96:25:@40285.4 package.scala 96:25:@40286.4]
  assign x433 = x414 | x672_x388_D1; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 458:59:@40289.4]
  assign _T_1120 = RetimeWrapper_82_io_out; // @[package.scala 96:25:@40331.4 package.scala 96:25:@40332.4]
  assign _T_1122 = io_rr ? _T_1120 : 1'h0; // @[implicits.scala 55:10:@40333.4]
  assign _T_1123 = _T_372 & _T_1122; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 471:194:@40334.4]
  assign x674_x434_D22 = RetimeWrapper_81_io_out; // @[package.scala 96:25:@40319.4 package.scala 96:25:@40320.4]
  assign _T_1124 = _T_1123 & x674_x434_D22; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 471:283:@40335.4]
  assign _T_1125 = _T_1124 & x639_b327_D50; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 471:291:@40336.4]
  assign x438 = x414 | x395; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 475:59:@40347.4]
  assign _T_1152 = RetimeWrapper_85_io_out; // @[package.scala 96:25:@40389.4 package.scala 96:25:@40390.4]
  assign _T_1154 = io_rr ? _T_1152 : 1'h0; // @[implicits.scala 55:10:@40391.4]
  assign _T_1155 = _T_372 & _T_1154; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 488:194:@40392.4]
  assign x676_x439_D22 = RetimeWrapper_84_io_out; // @[package.scala 96:25:@40377.4 package.scala 96:25:@40378.4]
  assign _T_1156 = _T_1155 & x676_x439_D22; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 488:283:@40393.4]
  assign _T_1157 = _T_1156 & x639_b327_D50; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 488:291:@40394.4]
  assign x443 = x414 | x404; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 492:59:@40405.4]
  assign _T_1184 = RetimeWrapper_88_io_out; // @[package.scala 96:25:@40447.4 package.scala 96:25:@40448.4]
  assign _T_1186 = io_rr ? _T_1184 : 1'h0; // @[implicits.scala 55:10:@40449.4]
  assign _T_1187 = _T_372 & _T_1186; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 505:194:@40450.4]
  assign x678_x444_D22 = RetimeWrapper_87_io_out; // @[package.scala 96:25:@40435.4 package.scala 96:25:@40436.4]
  assign _T_1188 = _T_1187 & x678_x444_D22; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 505:283:@40451.4]
  assign _T_1189 = _T_1188 & x639_b327_D50; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 505:291:@40452.4]
  assign x448_rdrow_number = x448_rdrow_1_io_result; // @[Math.scala 195:22:@40471.4 Math.scala 196:14:@40472.4]
  assign _T_1211 = $signed(x448_rdrow_number); // @[Math.scala 465:37:@40489.4]
  assign x450 = RetimeWrapper_89_io_out; // @[package.scala 96:25:@40497.4 package.scala 96:25:@40498.4]
  assign x451 = x450 | x367; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 515:24:@40501.4]
  assign x449_number = x449_1_io_result; // @[Math.scala 370:22:@40483.4 Math.scala 371:14:@40484.4]
  assign _T_1227 = $signed(x449_number); // @[Math.scala 406:49:@40510.4]
  assign _T_1229 = $signed(_T_1227) & $signed(32'sh3); // @[Math.scala 406:56:@40512.4]
  assign _T_1230 = $signed(_T_1229); // @[Math.scala 406:56:@40513.4]
  assign _T_1235 = x449_number[31]; // @[FixedPoint.scala 50:25:@40519.4]
  assign _T_1239 = _T_1235 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@40521.4]
  assign _T_1240 = x449_number[31:2]; // @[FixedPoint.scala 18:52:@40522.4]
  assign _T_1269 = RetimeWrapper_92_io_out; // @[package.scala 96:25:@40575.4 package.scala 96:25:@40576.4]
  assign _T_1271 = io_rr ? _T_1269 : 1'h0; // @[implicits.scala 55:10:@40577.4]
  assign _T_1272 = _T_372 & _T_1271; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 534:194:@40578.4]
  assign x679_x452_D22 = RetimeWrapper_90_io_out; // @[package.scala 96:25:@40554.4 package.scala 96:25:@40555.4]
  assign _T_1273 = _T_1272 & x679_x452_D22; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 534:283:@40579.4]
  assign _T_1274 = _T_1273 & x639_b327_D50; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 534:291:@40580.4]
  assign x459 = x450 | x376; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 544:59:@40591.4]
  assign _T_1300 = RetimeWrapper_94_io_out; // @[package.scala 96:25:@40626.4 package.scala 96:25:@40627.4]
  assign _T_1302 = io_rr ? _T_1300 : 1'h0; // @[implicits.scala 55:10:@40628.4]
  assign _T_1303 = _T_372 & _T_1302; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 557:194:@40629.4]
  assign x681_x460_D22 = RetimeWrapper_93_io_out; // @[package.scala 96:25:@40614.4 package.scala 96:25:@40615.4]
  assign _T_1304 = _T_1303 & x681_x460_D22; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 557:283:@40630.4]
  assign _T_1305 = _T_1304 & x639_b327_D50; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 557:291:@40631.4]
  assign x464 = x450 | x382; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 561:59:@40642.4]
  assign _T_1329 = RetimeWrapper_96_io_out; // @[package.scala 96:25:@40675.4 package.scala 96:25:@40676.4]
  assign _T_1331 = io_rr ? _T_1329 : 1'h0; // @[implicits.scala 55:10:@40677.4]
  assign _T_1332 = _T_372 & _T_1331; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 572:194:@40678.4]
  assign x682_x465_D22 = RetimeWrapper_95_io_out; // @[package.scala 96:25:@40663.4 package.scala 96:25:@40664.4]
  assign _T_1333 = _T_1332 & x682_x465_D22; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 572:283:@40679.4]
  assign _T_1334 = _T_1333 & x639_b327_D50; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 572:291:@40680.4]
  assign x469 = x450 | x672_x388_D1; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 576:59:@40691.4]
  assign _T_1358 = RetimeWrapper_98_io_out; // @[package.scala 96:25:@40724.4 package.scala 96:25:@40725.4]
  assign _T_1360 = io_rr ? _T_1358 : 1'h0; // @[implicits.scala 55:10:@40726.4]
  assign _T_1361 = _T_372 & _T_1360; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 587:194:@40727.4]
  assign x683_x470_D22 = RetimeWrapper_97_io_out; // @[package.scala 96:25:@40712.4 package.scala 96:25:@40713.4]
  assign _T_1362 = _T_1361 & x683_x470_D22; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 587:283:@40728.4]
  assign _T_1363 = _T_1362 & x639_b327_D50; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 587:291:@40729.4]
  assign x474 = x450 | x395; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 591:59:@40740.4]
  assign _T_1387 = RetimeWrapper_100_io_out; // @[package.scala 96:25:@40773.4 package.scala 96:25:@40774.4]
  assign _T_1389 = io_rr ? _T_1387 : 1'h0; // @[implicits.scala 55:10:@40775.4]
  assign _T_1390 = _T_372 & _T_1389; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 602:194:@40776.4]
  assign x684_x475_D22 = RetimeWrapper_99_io_out; // @[package.scala 96:25:@40761.4 package.scala 96:25:@40762.4]
  assign _T_1391 = _T_1390 & x684_x475_D22; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 602:283:@40777.4]
  assign _T_1392 = _T_1391 & x639_b327_D50; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 602:291:@40778.4]
  assign x479 = x450 | x404; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 606:59:@40789.4]
  assign _T_1416 = RetimeWrapper_102_io_out; // @[package.scala 96:25:@40822.4 package.scala 96:25:@40823.4]
  assign _T_1418 = io_rr ? _T_1416 : 1'h0; // @[implicits.scala 55:10:@40824.4]
  assign _T_1419 = _T_372 & _T_1418; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 617:194:@40825.4]
  assign x685_x480_D22 = RetimeWrapper_101_io_out; // @[package.scala 96:25:@40810.4 package.scala 96:25:@40811.4]
  assign _T_1420 = _T_1419 & x685_x480_D22; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 617:283:@40826.4]
  assign _T_1421 = _T_1420 & x639_b327_D50; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 617:291:@40827.4]
  assign x380_rd_0_number = x329_lb_0_io_rPort_3_output_0; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 259:29:@39548.4 sm_x542_inr_Foreach_SAMPLER_BOX.scala 263:338:@39569.4]
  assign _GEN_0 = {{1'd0}, x380_rd_0_number}; // @[Math.scala 450:32:@40839.4]
  assign x421_rd_0_number = x329_lb_0_io_rPort_2_output_0; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 406:29:@40137.4 sm_x542_inr_Foreach_SAMPLER_BOX.scala 410:408:@40158.4]
  assign _GEN_1 = {{1'd0}, x421_rd_0_number}; // @[Math.scala 450:32:@40851.4]
  assign x426_rd_0_number = x329_lb_0_io_rPort_10_output_0; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 431:29:@40197.4 sm_x542_inr_Foreach_SAMPLER_BOX.scala 435:408:@40218.4]
  assign _GEN_2 = {{2'd0}, x426_rd_0_number}; // @[Math.scala 450:32:@40863.4]
  assign x431_rd_0_number = x329_lb_0_io_rPort_9_output_0; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 448:29:@40255.4 sm_x542_inr_Foreach_SAMPLER_BOX.scala 452:408:@40276.4]
  assign _GEN_3 = {{1'd0}, x431_rd_0_number}; // @[Math.scala 450:32:@40875.4]
  assign x462_rd_0_number = x329_lb_0_io_rPort_8_output_0; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 553:29:@40617.4 sm_x542_inr_Foreach_SAMPLER_BOX.scala 557:408:@40638.4]
  assign _GEN_4 = {{1'd0}, x462_rd_0_number}; // @[Math.scala 450:32:@40887.4]
  assign x496_sum_number = x496_sum_1_io_result; // @[Math.scala 154:22:@41057.4 Math.scala 155:14:@41058.4]
  assign _T_1515 = x496_sum_number[7:4]; // @[FixedPoint.scala 18:52:@41063.4]
  assign x386_rd_0_number = x329_lb_0_io_rPort_13_output_0; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 284:29:@39647.4 sm_x542_inr_Foreach_SAMPLER_BOX.scala 288:338:@39668.4]
  assign _GEN_5 = {{1'd0}, x386_rd_0_number}; // @[Math.scala 450:32:@41069.4]
  assign _GEN_6 = {{1'd0}, x426_rd_0_number}; // @[Math.scala 450:32:@41081.4]
  assign _GEN_7 = {{2'd0}, x431_rd_0_number}; // @[Math.scala 450:32:@41093.4]
  assign x436_rd_0_number = x329_lb_0_io_rPort_1_output_0; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 467:29:@40322.4 sm_x542_inr_Foreach_SAMPLER_BOX.scala 471:408:@40343.4]
  assign _GEN_8 = {{1'd0}, x436_rd_0_number}; // @[Math.scala 450:32:@41105.4]
  assign x467_rd_0_number = x329_lb_0_io_rPort_5_output_0; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 568:29:@40666.4 sm_x542_inr_Foreach_SAMPLER_BOX.scala 572:408:@40687.4]
  assign _GEN_9 = {{1'd0}, x467_rd_0_number}; // @[Math.scala 450:32:@41117.4]
  assign x510_sum_number = x510_sum_1_io_result; // @[Math.scala 154:22:@41285.4 Math.scala 155:14:@41286.4]
  assign _T_1606 = x510_sum_number[7:4]; // @[FixedPoint.scala 18:52:@41291.4]
  assign x392_rd_0_number = x329_lb_0_io_rPort_4_output_0; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 317:29:@39748.4 sm_x542_inr_Foreach_SAMPLER_BOX.scala 321:408:@39769.4]
  assign _GEN_10 = {{1'd0}, x392_rd_0_number}; // @[Math.scala 450:32:@41297.4]
  assign _GEN_11 = {{2'd0}, x436_rd_0_number}; // @[Math.scala 450:32:@41309.4]
  assign x441_rd_0_number = x329_lb_0_io_rPort_12_output_0; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 484:29:@40380.4 sm_x542_inr_Foreach_SAMPLER_BOX.scala 488:408:@40401.4]
  assign _GEN_12 = {{1'd0}, x441_rd_0_number}; // @[Math.scala 450:32:@41321.4]
  assign x472_rd_0_number = x329_lb_0_io_rPort_0_output_0; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 583:29:@40715.4 sm_x542_inr_Foreach_SAMPLER_BOX.scala 587:408:@40736.4]
  assign _GEN_13 = {{1'd0}, x472_rd_0_number}; // @[Math.scala 450:32:@41333.4]
  assign x523_sum_number = x523_sum_1_io_result; // @[Math.scala 154:22:@41492.4 Math.scala 155:14:@41493.4]
  assign _T_1688 = x523_sum_number[7:4]; // @[FixedPoint.scala 18:52:@41498.4]
  assign x401_rd_0_number = x329_lb_0_io_rPort_16_output_0; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 346:29:@39874.4 sm_x542_inr_Foreach_SAMPLER_BOX.scala 350:408:@39895.4]
  assign _GEN_14 = {{1'd0}, x401_rd_0_number}; // @[Math.scala 450:32:@41506.4]
  assign _GEN_15 = {{2'd0}, x441_rd_0_number}; // @[Math.scala 450:32:@41518.4]
  assign x446_rd_0_number = x329_lb_0_io_rPort_14_output_0; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 501:29:@40438.4 sm_x542_inr_Foreach_SAMPLER_BOX.scala 505:408:@40459.4]
  assign _GEN_16 = {{1'd0}, x446_rd_0_number}; // @[Math.scala 450:32:@41530.4]
  assign x477_rd_0_number = x329_lb_0_io_rPort_7_output_0; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 598:29:@40764.4 sm_x542_inr_Foreach_SAMPLER_BOX.scala 602:408:@40785.4]
  assign _GEN_17 = {{1'd0}, x477_rd_0_number}; // @[Math.scala 450:32:@41542.4]
  assign x536_sum_number = x536_sum_1_io_result; // @[Math.scala 154:22:@41701.4 Math.scala 155:14:@41702.4]
  assign _T_1772 = x536_sum_number[7:4]; // @[FixedPoint.scala 18:52:@41707.4]
  assign x720_x524_D3_number = RetimeWrapper_155_io_out; // @[package.scala 96:25:@41717.4 package.scala 96:25:@41718.4]
  assign x722_x537_D3_number = RetimeWrapper_157_io_out; // @[package.scala 96:25:@41735.4 package.scala 96:25:@41736.4]
  assign _T_1797 = {x720_x524_D3_number,x722_x537_D3_number}; // @[Cat.scala 30:58:@41753.4]
  assign x721_x497_D3_number = RetimeWrapper_156_io_out; // @[package.scala 96:25:@41726.4 package.scala 96:25:@41727.4]
  assign x723_x511_D3_number = RetimeWrapper_158_io_out; // @[package.scala 96:25:@41744.4 package.scala 96:25:@41745.4]
  assign _T_1798 = {x721_x497_D3_number,x723_x511_D3_number}; // @[Cat.scala 30:58:@41754.4]
  assign _T_1811 = RetimeWrapper_162_io_out; // @[package.scala 96:25:@41790.4 package.scala 96:25:@41791.4]
  assign _T_1813 = io_rr ? _T_1811 : 1'h0; // @[implicits.scala 55:10:@41792.4]
  assign x724_b327_D63 = RetimeWrapper_160_io_out; // @[package.scala 96:25:@41772.4 package.scala 96:25:@41773.4]
  assign _T_1814 = _T_1813 & x724_b327_D63; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 829:117:@41793.4]
  assign x725_b328_D63 = RetimeWrapper_161_io_out; // @[package.scala 96:25:@41781.4 package.scala 96:25:@41782.4]
  assign _T_1815 = _T_1814 & x725_b328_D63; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 829:123:@41794.4]
  assign x616_x340_D8_number = RetimeWrapper_2_io_out; // @[package.scala 96:25:@38895.4 package.scala 96:25:@38896.4]
  assign x617_x344_sum_D3_number = RetimeWrapper_3_io_out; // @[package.scala 96:25:@38904.4 package.scala 96:25:@38905.4]
  assign x618_x610_D24_number = RetimeWrapper_4_io_out; // @[package.scala 96:25:@38913.4 package.scala 96:25:@38914.4]
  assign x624_x348_D7_number = RetimeWrapper_11_io_out; // @[package.scala 96:25:@39038.4 package.scala 96:25:@39039.4]
  assign x625_x350_sum_D2_number = RetimeWrapper_12_io_out; // @[package.scala 96:25:@39047.4 package.scala 96:25:@39048.4]
  assign x627_x356_sum_D2_number = RetimeWrapper_15_io_out; // @[package.scala 96:25:@39136.4 package.scala 96:25:@39137.4]
  assign x628_x354_D7_number = RetimeWrapper_16_io_out; // @[package.scala 96:25:@39145.4 package.scala 96:25:@39146.4]
  assign x629_x360_D7_number = RetimeWrapper_18_io_out; // @[package.scala 96:25:@39225.4 package.scala 96:25:@39226.4]
  assign x630_x362_sum_D2_number = RetimeWrapper_19_io_out; // @[package.scala 96:25:@39234.4 package.scala 96:25:@39235.4]
  assign x637_x360_D33_number = RetimeWrapper_29_io_out; // @[package.scala 96:25:@39410.4 package.scala 96:25:@39411.4]
  assign x638_x611_D8_number = RetimeWrapper_30_io_out; // @[package.scala 96:25:@39419.4 package.scala 96:25:@39420.4]
  assign x640_x373_sum_D1_number = RetimeWrapper_32_io_out; // @[package.scala 96:25:@39437.4 package.scala 96:25:@39438.4]
  assign x644_x379_sum_D1_number = RetimeWrapper_38_io_out; // @[package.scala 96:25:@39527.4 package.scala 96:25:@39528.4]
  assign x646_x354_D33_number = RetimeWrapper_40_io_out; // @[package.scala 96:25:@39545.4 package.scala 96:25:@39546.4]
  assign x649_x385_sum_D1_number = RetimeWrapper_45_io_out; // @[package.scala 96:25:@39626.4 package.scala 96:25:@39627.4]
  assign x651_x348_D33_number = RetimeWrapper_47_io_out; // @[package.scala 96:25:@39644.4 package.scala 96:25:@39645.4]
  assign x654_x340_D34_number = RetimeWrapper_52_io_out; // @[package.scala 96:25:@39727.4 package.scala 96:25:@39728.4]
  assign x655_x391_sum_D1_number = RetimeWrapper_53_io_out; // @[package.scala 96:25:@39736.4 package.scala 96:25:@39737.4]
  assign x659_x398_D7_number = RetimeWrapper_59_io_out; // @[package.scala 96:25:@39862.4 package.scala 96:25:@39863.4]
  assign x660_x400_sum_D1_number = RetimeWrapper_60_io_out; // @[package.scala 96:25:@39871.4 package.scala 96:25:@39872.4]
  assign x662_x407_D7_number = RetimeWrapper_64_io_out; // @[package.scala 96:25:@39979.4 package.scala 96:25:@39980.4]
  assign x664_x409_sum_D1_number = RetimeWrapper_66_io_out; // @[package.scala 96:25:@39997.4 package.scala 96:25:@39998.4]
  assign x420_sum_number = x420_sum_1_io_result; // @[Math.scala 154:22:@40116.4 Math.scala 155:14:@40117.4]
  assign x667_x612_D7_number = RetimeWrapper_71_io_out; // @[package.scala 96:25:@40134.4 package.scala 96:25:@40135.4]
  assign x425_sum_number = x425_sum_1_io_result; // @[Math.scala 154:22:@40185.4 Math.scala 155:14:@40186.4]
  assign x430_sum_number = x430_sum_1_io_result; // @[Math.scala 154:22:@40243.4 Math.scala 155:14:@40244.4]
  assign x435_sum_number = x435_sum_1_io_result; // @[Math.scala 154:22:@40310.4 Math.scala 155:14:@40311.4]
  assign x440_sum_number = x440_sum_1_io_result; // @[Math.scala 154:22:@40368.4 Math.scala 155:14:@40369.4]
  assign x445_sum_number = x445_sum_1_io_result; // @[Math.scala 154:22:@40426.4 Math.scala 155:14:@40427.4]
  assign x456_sum_number = x456_sum_1_io_result; // @[Math.scala 154:22:@40545.4 Math.scala 155:14:@40546.4]
  assign x680_x613_D7_number = RetimeWrapper_91_io_out; // @[package.scala 96:25:@40563.4 package.scala 96:25:@40564.4]
  assign x461_sum_number = x461_sum_1_io_result; // @[Math.scala 154:22:@40605.4 Math.scala 155:14:@40606.4]
  assign x466_sum_number = x466_sum_1_io_result; // @[Math.scala 154:22:@40654.4 Math.scala 155:14:@40655.4]
  assign x471_sum_number = x471_sum_1_io_result; // @[Math.scala 154:22:@40703.4 Math.scala 155:14:@40704.4]
  assign x476_sum_number = x476_sum_1_io_result; // @[Math.scala 154:22:@40752.4 Math.scala 155:14:@40753.4]
  assign x481_sum_number = x481_sum_1_io_result; // @[Math.scala 154:22:@40801.4 Math.scala 155:14:@40802.4]
  assign _T_1429 = RetimeWrapper_103_io_out; // @[package.scala 96:25:@40845.4 package.scala 96:25:@40846.4]
  assign _T_1435 = RetimeWrapper_104_io_out; // @[package.scala 96:25:@40857.4 package.scala 96:25:@40858.4]
  assign _T_1441 = RetimeWrapper_105_io_out; // @[package.scala 96:25:@40869.4 package.scala 96:25:@40870.4]
  assign _T_1447 = RetimeWrapper_106_io_out; // @[package.scala 96:25:@40881.4 package.scala 96:25:@40882.4]
  assign _T_1453 = RetimeWrapper_107_io_out; // @[package.scala 96:25:@40893.4 package.scala 96:25:@40894.4]
  assign _T_1522 = RetimeWrapper_117_io_out; // @[package.scala 96:25:@41075.4 package.scala 96:25:@41076.4]
  assign _T_1528 = RetimeWrapper_118_io_out; // @[package.scala 96:25:@41087.4 package.scala 96:25:@41088.4]
  assign _T_1534 = RetimeWrapper_119_io_out; // @[package.scala 96:25:@41099.4 package.scala 96:25:@41100.4]
  assign _T_1540 = RetimeWrapper_120_io_out; // @[package.scala 96:25:@41111.4 package.scala 96:25:@41112.4]
  assign _T_1546 = RetimeWrapper_121_io_out; // @[package.scala 96:25:@41123.4 package.scala 96:25:@41124.4]
  assign _T_1613 = RetimeWrapper_131_io_out; // @[package.scala 96:25:@41303.4 package.scala 96:25:@41304.4]
  assign _T_1619 = RetimeWrapper_132_io_out; // @[package.scala 96:25:@41315.4 package.scala 96:25:@41316.4]
  assign _T_1625 = RetimeWrapper_133_io_out; // @[package.scala 96:25:@41327.4 package.scala 96:25:@41328.4]
  assign _T_1631 = RetimeWrapper_134_io_out; // @[package.scala 96:25:@41339.4 package.scala 96:25:@41340.4]
  assign _T_1697 = RetimeWrapper_143_io_out; // @[package.scala 96:25:@41512.4 package.scala 96:25:@41513.4]
  assign _T_1703 = RetimeWrapper_144_io_out; // @[package.scala 96:25:@41524.4 package.scala 96:25:@41525.4]
  assign _T_1709 = RetimeWrapper_145_io_out; // @[package.scala 96:25:@41536.4 package.scala 96:25:@41537.4]
  assign _T_1715 = RetimeWrapper_146_io_out; // @[package.scala 96:25:@41548.4 package.scala 96:25:@41549.4]
  assign io_in_x316_TREADY = _T_212 & _T_214; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 68:22:@38734.4 sm_x542_inr_Foreach_SAMPLER_BOX.scala 70:22:@38742.4]
  assign io_in_x317_TVALID = _T_1815 & io_sigsIn_backpressure; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 829:22:@41796.4]
  assign io_in_x317_TDATA = {{224'd0}, RetimeWrapper_159_io_out}; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 830:24:@41797.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 710:17:@38567.4]
  assign __1_io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_1); // @[Math.scala 710:17:@38579.4]
  assign x329_lb_0_clock = clock; // @[:@38587.4]
  assign x329_lb_0_reset = reset; // @[:@38588.4]
  assign x329_lb_0_io_rPort_17_banks_1 = x662_x407_D7_number[2:0]; // @[MemInterfaceType.scala 106:58:@40017.4]
  assign x329_lb_0_io_rPort_17_banks_0 = x638_x611_D8_number[2:0]; // @[MemInterfaceType.scala 106:58:@40016.4]
  assign x329_lb_0_io_rPort_17_ofs_0 = x664_x409_sum_D1_number[7:0]; // @[MemInterfaceType.scala 107:54:@40018.4]
  assign x329_lb_0_io_rPort_17_en_0 = _T_936 & x636_b328_D50; // @[MemInterfaceType.scala 110:79:@40020.4]
  assign x329_lb_0_io_rPort_17_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@40019.4]
  assign x329_lb_0_io_rPort_16_banks_1 = x659_x398_D7_number[2:0]; // @[MemInterfaceType.scala 106:58:@39891.4]
  assign x329_lb_0_io_rPort_16_banks_0 = x638_x611_D8_number[2:0]; // @[MemInterfaceType.scala 106:58:@39890.4]
  assign x329_lb_0_io_rPort_16_ofs_0 = x660_x400_sum_D1_number[7:0]; // @[MemInterfaceType.scala 107:54:@39892.4]
  assign x329_lb_0_io_rPort_16_en_0 = _T_867 & x636_b328_D50; // @[MemInterfaceType.scala 110:79:@39894.4]
  assign x329_lb_0_io_rPort_16_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@39893.4]
  assign x329_lb_0_io_rPort_15_banks_1 = x662_x407_D7_number[2:0]; // @[MemInterfaceType.scala 106:58:@40830.4]
  assign x329_lb_0_io_rPort_15_banks_0 = x680_x613_D7_number[2:0]; // @[MemInterfaceType.scala 106:58:@40829.4]
  assign x329_lb_0_io_rPort_15_ofs_0 = x481_sum_number[7:0]; // @[MemInterfaceType.scala 107:54:@40831.4]
  assign x329_lb_0_io_rPort_15_en_0 = _T_1421 & x636_b328_D50; // @[MemInterfaceType.scala 110:79:@40833.4]
  assign x329_lb_0_io_rPort_15_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@40832.4]
  assign x329_lb_0_io_rPort_14_banks_1 = x662_x407_D7_number[2:0]; // @[MemInterfaceType.scala 106:58:@40455.4]
  assign x329_lb_0_io_rPort_14_banks_0 = x667_x612_D7_number[2:0]; // @[MemInterfaceType.scala 106:58:@40454.4]
  assign x329_lb_0_io_rPort_14_ofs_0 = x445_sum_number[7:0]; // @[MemInterfaceType.scala 107:54:@40456.4]
  assign x329_lb_0_io_rPort_14_en_0 = _T_1189 & x636_b328_D50; // @[MemInterfaceType.scala 110:79:@40458.4]
  assign x329_lb_0_io_rPort_14_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@40457.4]
  assign x329_lb_0_io_rPort_13_banks_1 = x651_x348_D33_number[2:0]; // @[MemInterfaceType.scala 106:58:@39664.4]
  assign x329_lb_0_io_rPort_13_banks_0 = x638_x611_D8_number[2:0]; // @[MemInterfaceType.scala 106:58:@39663.4]
  assign x329_lb_0_io_rPort_13_ofs_0 = x649_x385_sum_D1_number[7:0]; // @[MemInterfaceType.scala 107:54:@39665.4]
  assign x329_lb_0_io_rPort_13_en_0 = _T_745 & x636_b328_D50; // @[MemInterfaceType.scala 110:79:@39667.4]
  assign x329_lb_0_io_rPort_13_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@39666.4]
  assign x329_lb_0_io_rPort_12_banks_1 = x659_x398_D7_number[2:0]; // @[MemInterfaceType.scala 106:58:@40397.4]
  assign x329_lb_0_io_rPort_12_banks_0 = x667_x612_D7_number[2:0]; // @[MemInterfaceType.scala 106:58:@40396.4]
  assign x329_lb_0_io_rPort_12_ofs_0 = x440_sum_number[7:0]; // @[MemInterfaceType.scala 107:54:@40398.4]
  assign x329_lb_0_io_rPort_12_en_0 = _T_1157 & x636_b328_D50; // @[MemInterfaceType.scala 110:79:@40400.4]
  assign x329_lb_0_io_rPort_12_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@40399.4]
  assign x329_lb_0_io_rPort_11_banks_1 = x637_x360_D33_number[2:0]; // @[MemInterfaceType.scala 106:58:@39466.4]
  assign x329_lb_0_io_rPort_11_banks_0 = x638_x611_D8_number[2:0]; // @[MemInterfaceType.scala 106:58:@39465.4]
  assign x329_lb_0_io_rPort_11_ofs_0 = x640_x373_sum_D1_number[7:0]; // @[MemInterfaceType.scala 107:54:@39467.4]
  assign x329_lb_0_io_rPort_11_en_0 = _T_643 & x636_b328_D50; // @[MemInterfaceType.scala 110:79:@39469.4]
  assign x329_lb_0_io_rPort_11_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@39468.4]
  assign x329_lb_0_io_rPort_10_banks_1 = x646_x354_D33_number[2:0]; // @[MemInterfaceType.scala 106:58:@40214.4]
  assign x329_lb_0_io_rPort_10_banks_0 = x667_x612_D7_number[2:0]; // @[MemInterfaceType.scala 106:58:@40213.4]
  assign x329_lb_0_io_rPort_10_ofs_0 = x425_sum_number[7:0]; // @[MemInterfaceType.scala 107:54:@40215.4]
  assign x329_lb_0_io_rPort_10_en_0 = _T_1058 & x636_b328_D50; // @[MemInterfaceType.scala 110:79:@40217.4]
  assign x329_lb_0_io_rPort_10_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@40216.4]
  assign x329_lb_0_io_rPort_9_banks_1 = x651_x348_D33_number[2:0]; // @[MemInterfaceType.scala 106:58:@40272.4]
  assign x329_lb_0_io_rPort_9_banks_0 = x667_x612_D7_number[2:0]; // @[MemInterfaceType.scala 106:58:@40271.4]
  assign x329_lb_0_io_rPort_9_ofs_0 = x430_sum_number[7:0]; // @[MemInterfaceType.scala 107:54:@40273.4]
  assign x329_lb_0_io_rPort_9_en_0 = _T_1090 & x636_b328_D50; // @[MemInterfaceType.scala 110:79:@40275.4]
  assign x329_lb_0_io_rPort_9_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@40274.4]
  assign x329_lb_0_io_rPort_8_banks_1 = x646_x354_D33_number[2:0]; // @[MemInterfaceType.scala 106:58:@40634.4]
  assign x329_lb_0_io_rPort_8_banks_0 = x680_x613_D7_number[2:0]; // @[MemInterfaceType.scala 106:58:@40633.4]
  assign x329_lb_0_io_rPort_8_ofs_0 = x461_sum_number[7:0]; // @[MemInterfaceType.scala 107:54:@40635.4]
  assign x329_lb_0_io_rPort_8_en_0 = _T_1305 & x636_b328_D50; // @[MemInterfaceType.scala 110:79:@40637.4]
  assign x329_lb_0_io_rPort_8_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@40636.4]
  assign x329_lb_0_io_rPort_7_banks_1 = x659_x398_D7_number[2:0]; // @[MemInterfaceType.scala 106:58:@40781.4]
  assign x329_lb_0_io_rPort_7_banks_0 = x680_x613_D7_number[2:0]; // @[MemInterfaceType.scala 106:58:@40780.4]
  assign x329_lb_0_io_rPort_7_ofs_0 = x476_sum_number[7:0]; // @[MemInterfaceType.scala 107:54:@40782.4]
  assign x329_lb_0_io_rPort_7_en_0 = _T_1392 & x636_b328_D50; // @[MemInterfaceType.scala 110:79:@40784.4]
  assign x329_lb_0_io_rPort_7_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@40783.4]
  assign x329_lb_0_io_rPort_6_banks_1 = x637_x360_D33_number[2:0]; // @[MemInterfaceType.scala 106:58:@40583.4]
  assign x329_lb_0_io_rPort_6_banks_0 = x680_x613_D7_number[2:0]; // @[MemInterfaceType.scala 106:58:@40582.4]
  assign x329_lb_0_io_rPort_6_ofs_0 = x456_sum_number[7:0]; // @[MemInterfaceType.scala 107:54:@40584.4]
  assign x329_lb_0_io_rPort_6_en_0 = _T_1274 & x636_b328_D50; // @[MemInterfaceType.scala 110:79:@40586.4]
  assign x329_lb_0_io_rPort_6_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@40585.4]
  assign x329_lb_0_io_rPort_5_banks_1 = x651_x348_D33_number[2:0]; // @[MemInterfaceType.scala 106:58:@40683.4]
  assign x329_lb_0_io_rPort_5_banks_0 = x680_x613_D7_number[2:0]; // @[MemInterfaceType.scala 106:58:@40682.4]
  assign x329_lb_0_io_rPort_5_ofs_0 = x466_sum_number[7:0]; // @[MemInterfaceType.scala 107:54:@40684.4]
  assign x329_lb_0_io_rPort_5_en_0 = _T_1334 & x636_b328_D50; // @[MemInterfaceType.scala 110:79:@40686.4]
  assign x329_lb_0_io_rPort_5_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@40685.4]
  assign x329_lb_0_io_rPort_4_banks_1 = x654_x340_D34_number[2:0]; // @[MemInterfaceType.scala 106:58:@39765.4]
  assign x329_lb_0_io_rPort_4_banks_0 = x638_x611_D8_number[2:0]; // @[MemInterfaceType.scala 106:58:@39764.4]
  assign x329_lb_0_io_rPort_4_ofs_0 = x655_x391_sum_D1_number[7:0]; // @[MemInterfaceType.scala 107:54:@39766.4]
  assign x329_lb_0_io_rPort_4_en_0 = _T_798 & x636_b328_D50; // @[MemInterfaceType.scala 110:79:@39768.4]
  assign x329_lb_0_io_rPort_4_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@39767.4]
  assign x329_lb_0_io_rPort_3_banks_1 = x646_x354_D33_number[2:0]; // @[MemInterfaceType.scala 106:58:@39565.4]
  assign x329_lb_0_io_rPort_3_banks_0 = x638_x611_D8_number[2:0]; // @[MemInterfaceType.scala 106:58:@39564.4]
  assign x329_lb_0_io_rPort_3_ofs_0 = x644_x379_sum_D1_number[7:0]; // @[MemInterfaceType.scala 107:54:@39566.4]
  assign x329_lb_0_io_rPort_3_en_0 = _T_694 & x636_b328_D50; // @[MemInterfaceType.scala 110:79:@39568.4]
  assign x329_lb_0_io_rPort_3_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@39567.4]
  assign x329_lb_0_io_rPort_2_banks_1 = x637_x360_D33_number[2:0]; // @[MemInterfaceType.scala 106:58:@40154.4]
  assign x329_lb_0_io_rPort_2_banks_0 = x667_x612_D7_number[2:0]; // @[MemInterfaceType.scala 106:58:@40153.4]
  assign x329_lb_0_io_rPort_2_ofs_0 = x420_sum_number[7:0]; // @[MemInterfaceType.scala 107:54:@40155.4]
  assign x329_lb_0_io_rPort_2_en_0 = _T_1024 & x636_b328_D50; // @[MemInterfaceType.scala 110:79:@40157.4]
  assign x329_lb_0_io_rPort_2_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@40156.4]
  assign x329_lb_0_io_rPort_1_banks_1 = x654_x340_D34_number[2:0]; // @[MemInterfaceType.scala 106:58:@40339.4]
  assign x329_lb_0_io_rPort_1_banks_0 = x667_x612_D7_number[2:0]; // @[MemInterfaceType.scala 106:58:@40338.4]
  assign x329_lb_0_io_rPort_1_ofs_0 = x435_sum_number[7:0]; // @[MemInterfaceType.scala 107:54:@40340.4]
  assign x329_lb_0_io_rPort_1_en_0 = _T_1125 & x636_b328_D50; // @[MemInterfaceType.scala 110:79:@40342.4]
  assign x329_lb_0_io_rPort_1_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@40341.4]
  assign x329_lb_0_io_rPort_0_banks_1 = x654_x340_D34_number[2:0]; // @[MemInterfaceType.scala 106:58:@40732.4]
  assign x329_lb_0_io_rPort_0_banks_0 = x680_x613_D7_number[2:0]; // @[MemInterfaceType.scala 106:58:@40731.4]
  assign x329_lb_0_io_rPort_0_ofs_0 = x471_sum_number[7:0]; // @[MemInterfaceType.scala 107:54:@40733.4]
  assign x329_lb_0_io_rPort_0_en_0 = _T_1363 & x636_b328_D50; // @[MemInterfaceType.scala 110:79:@40735.4]
  assign x329_lb_0_io_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@40734.4]
  assign x329_lb_0_io_wPort_3_banks_1 = x629_x360_D7_number[2:0]; // @[MemInterfaceType.scala 88:58:@39264.4]
  assign x329_lb_0_io_wPort_3_banks_0 = x618_x610_D24_number[2:0]; // @[MemInterfaceType.scala 88:58:@39263.4]
  assign x329_lb_0_io_wPort_3_ofs_0 = x630_x362_sum_D2_number[7:0]; // @[MemInterfaceType.scala 89:54:@39265.4]
  assign x329_lb_0_io_wPort_3_data_0 = RetimeWrapper_20_io_out; // @[MemInterfaceType.scala 90:56:@39266.4]
  assign x329_lb_0_io_wPort_3_en_0 = _T_530 & x619_b328_D24; // @[MemInterfaceType.scala 93:57:@39268.4]
  assign x329_lb_0_io_wPort_2_banks_1 = x628_x354_D7_number[2:0]; // @[MemInterfaceType.scala 88:58:@39166.4]
  assign x329_lb_0_io_wPort_2_banks_0 = x618_x610_D24_number[2:0]; // @[MemInterfaceType.scala 88:58:@39165.4]
  assign x329_lb_0_io_wPort_2_ofs_0 = x627_x356_sum_D2_number[7:0]; // @[MemInterfaceType.scala 89:54:@39167.4]
  assign x329_lb_0_io_wPort_2_data_0 = RetimeWrapper_14_io_out; // @[MemInterfaceType.scala 90:56:@39168.4]
  assign x329_lb_0_io_wPort_2_en_0 = _T_482 & x619_b328_D24; // @[MemInterfaceType.scala 93:57:@39170.4]
  assign x329_lb_0_io_wPort_1_banks_1 = x624_x348_D7_number[2:0]; // @[MemInterfaceType.scala 88:58:@39068.4]
  assign x329_lb_0_io_wPort_1_banks_0 = x618_x610_D24_number[2:0]; // @[MemInterfaceType.scala 88:58:@39067.4]
  assign x329_lb_0_io_wPort_1_ofs_0 = x625_x350_sum_D2_number[7:0]; // @[MemInterfaceType.scala 89:54:@39069.4]
  assign x329_lb_0_io_wPort_1_data_0 = RetimeWrapper_10_io_out; // @[MemInterfaceType.scala 90:56:@39070.4]
  assign x329_lb_0_io_wPort_1_en_0 = _T_434 & x619_b328_D24; // @[MemInterfaceType.scala 93:57:@39072.4]
  assign x329_lb_0_io_wPort_0_banks_1 = x616_x340_D8_number[2:0]; // @[MemInterfaceType.scala 88:58:@38961.4]
  assign x329_lb_0_io_wPort_0_banks_0 = x618_x610_D24_number[2:0]; // @[MemInterfaceType.scala 88:58:@38960.4]
  assign x329_lb_0_io_wPort_0_ofs_0 = x617_x344_sum_D3_number[7:0]; // @[MemInterfaceType.scala 89:54:@38962.4]
  assign x329_lb_0_io_wPort_0_data_0 = RetimeWrapper_7_io_out; // @[MemInterfaceType.scala 90:56:@38963.4]
  assign x329_lb_0_io_wPort_0_en_0 = _T_383 & x619_b328_D24; // @[MemInterfaceType.scala 93:57:@38965.4]
  assign RetimeWrapper_clock = clock; // @[:@38745.4]
  assign RetimeWrapper_reset = reset; // @[:@38746.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38748.4]
  assign RetimeWrapper_io_in = io_in_x316_TDATA[31:0]; // @[package.scala 94:16:@38747.4]
  assign x340_1_clock = clock; // @[:@38829.4]
  assign x340_1_reset = reset; // @[:@38830.4]
  assign x340_1_io_a = __1_io_result; // @[Math.scala 367:17:@38831.4]
  assign x340_1_io_b = 32'h6; // @[Math.scala 368:17:@38832.4]
  assign x340_1_io_flow = io_in_x317_TREADY; // @[Math.scala 369:20:@38833.4]
  assign x342_mul_1_clock = clock; // @[:@38850.4]
  assign x342_mul_1_reset = reset; // @[:@38851.4]
  assign x342_mul_1_io_a = {_T_330,_T_331}; // @[Math.scala 263:17:@38852.4]
  assign x342_mul_1_io_flow = io_in_x317_TREADY; // @[Math.scala 265:20:@38854.4]
  assign x343_div_1_clock = clock; // @[:@38862.4]
  assign x343_div_1_reset = reset; // @[:@38863.4]
  assign x343_div_1_io_a = __1_io_result; // @[Math.scala 328:17:@38864.4]
  assign x343_div_1_io_flow = io_in_x317_TREADY; // @[Math.scala 330:20:@38866.4]
  assign RetimeWrapper_1_clock = clock; // @[:@38872.4]
  assign RetimeWrapper_1_reset = reset; // @[:@38873.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38875.4]
  assign RetimeWrapper_1_io_in = x342_mul_1_io_result; // @[package.scala 94:16:@38874.4]
  assign x344_sum_1_clock = clock; // @[:@38881.4]
  assign x344_sum_1_reset = reset; // @[:@38882.4]
  assign x344_sum_1_io_a = RetimeWrapper_1_io_out; // @[Math.scala 151:17:@38883.4]
  assign x344_sum_1_io_b = x343_div_1_io_result; // @[Math.scala 152:17:@38884.4]
  assign x344_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@38885.4]
  assign RetimeWrapper_2_clock = clock; // @[:@38891.4]
  assign RetimeWrapper_2_reset = reset; // @[:@38892.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38894.4]
  assign RetimeWrapper_2_io_in = x340_1_io_result; // @[package.scala 94:16:@38893.4]
  assign RetimeWrapper_3_clock = clock; // @[:@38900.4]
  assign RetimeWrapper_3_reset = reset; // @[:@38901.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38903.4]
  assign RetimeWrapper_3_io_in = x344_sum_1_io_result; // @[package.scala 94:16:@38902.4]
  assign RetimeWrapper_4_clock = clock; // @[:@38909.4]
  assign RetimeWrapper_4_reset = reset; // @[:@38910.4]
  assign RetimeWrapper_4_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38912.4]
  assign RetimeWrapper_4_io_in = $unsigned(_T_314); // @[package.scala 94:16:@38911.4]
  assign RetimeWrapper_5_clock = clock; // @[:@38918.4]
  assign RetimeWrapper_5_reset = reset; // @[:@38919.4]
  assign RetimeWrapper_5_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38921.4]
  assign RetimeWrapper_5_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@38920.4]
  assign RetimeWrapper_6_clock = clock; // @[:@38927.4]
  assign RetimeWrapper_6_reset = reset; // @[:@38928.4]
  assign RetimeWrapper_6_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38930.4]
  assign RetimeWrapper_6_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@38929.4]
  assign RetimeWrapper_7_clock = clock; // @[:@38936.4]
  assign RetimeWrapper_7_reset = reset; // @[:@38937.4]
  assign RetimeWrapper_7_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38939.4]
  assign RetimeWrapper_7_io_in = x614_x330_D1_0_number[7:0]; // @[package.scala 94:16:@38938.4]
  assign RetimeWrapper_8_clock = clock; // @[:@38947.4]
  assign RetimeWrapper_8_reset = reset; // @[:@38948.4]
  assign RetimeWrapper_8_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38950.4]
  assign RetimeWrapper_8_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@38949.4]
  assign x346_rdcol_1_clock = clock; // @[:@38970.4]
  assign x346_rdcol_1_reset = reset; // @[:@38971.4]
  assign x346_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@38972.4]
  assign x346_rdcol_1_io_b = 32'h1; // @[Math.scala 152:17:@38973.4]
  assign x346_rdcol_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@38974.4]
  assign x348_1_clock = clock; // @[:@38984.4]
  assign x348_1_reset = reset; // @[:@38985.4]
  assign x348_1_io_a = x346_rdcol_1_io_result; // @[Math.scala 367:17:@38986.4]
  assign x348_1_io_b = 32'h6; // @[Math.scala 368:17:@38987.4]
  assign x348_1_io_flow = io_in_x317_TREADY; // @[Math.scala 369:20:@38988.4]
  assign x349_div_1_clock = clock; // @[:@38996.4]
  assign x349_div_1_reset = reset; // @[:@38997.4]
  assign x349_div_1_io_a = x346_rdcol_1_io_result; // @[Math.scala 328:17:@38998.4]
  assign x349_div_1_io_flow = io_in_x317_TREADY; // @[Math.scala 330:20:@39000.4]
  assign RetimeWrapper_9_clock = clock; // @[:@39006.4]
  assign RetimeWrapper_9_reset = reset; // @[:@39007.4]
  assign RetimeWrapper_9_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39009.4]
  assign RetimeWrapper_9_io_in = x342_mul_1_io_result; // @[package.scala 94:16:@39008.4]
  assign x350_sum_1_clock = clock; // @[:@39015.4]
  assign x350_sum_1_reset = reset; // @[:@39016.4]
  assign x350_sum_1_io_a = RetimeWrapper_9_io_out; // @[Math.scala 151:17:@39017.4]
  assign x350_sum_1_io_b = x349_div_1_io_result; // @[Math.scala 152:17:@39018.4]
  assign x350_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@39019.4]
  assign RetimeWrapper_10_clock = clock; // @[:@39025.4]
  assign RetimeWrapper_10_reset = reset; // @[:@39026.4]
  assign RetimeWrapper_10_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39028.4]
  assign RetimeWrapper_10_io_in = x614_x330_D1_0_number[15:8]; // @[package.scala 94:16:@39027.4]
  assign RetimeWrapper_11_clock = clock; // @[:@39034.4]
  assign RetimeWrapper_11_reset = reset; // @[:@39035.4]
  assign RetimeWrapper_11_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39037.4]
  assign RetimeWrapper_11_io_in = x348_1_io_result; // @[package.scala 94:16:@39036.4]
  assign RetimeWrapper_12_clock = clock; // @[:@39043.4]
  assign RetimeWrapper_12_reset = reset; // @[:@39044.4]
  assign RetimeWrapper_12_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39046.4]
  assign RetimeWrapper_12_io_in = x350_sum_1_io_result; // @[package.scala 94:16:@39045.4]
  assign RetimeWrapper_13_clock = clock; // @[:@39054.4]
  assign RetimeWrapper_13_reset = reset; // @[:@39055.4]
  assign RetimeWrapper_13_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39057.4]
  assign RetimeWrapper_13_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@39056.4]
  assign x352_rdcol_1_clock = clock; // @[:@39077.4]
  assign x352_rdcol_1_reset = reset; // @[:@39078.4]
  assign x352_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@39079.4]
  assign x352_rdcol_1_io_b = 32'h2; // @[Math.scala 152:17:@39080.4]
  assign x352_rdcol_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@39081.4]
  assign x354_1_clock = clock; // @[:@39091.4]
  assign x354_1_reset = reset; // @[:@39092.4]
  assign x354_1_io_a = x352_rdcol_1_io_result; // @[Math.scala 367:17:@39093.4]
  assign x354_1_io_b = 32'h6; // @[Math.scala 368:17:@39094.4]
  assign x354_1_io_flow = io_in_x317_TREADY; // @[Math.scala 369:20:@39095.4]
  assign x355_div_1_clock = clock; // @[:@39103.4]
  assign x355_div_1_reset = reset; // @[:@39104.4]
  assign x355_div_1_io_a = x352_rdcol_1_io_result; // @[Math.scala 328:17:@39105.4]
  assign x355_div_1_io_flow = io_in_x317_TREADY; // @[Math.scala 330:20:@39107.4]
  assign x356_sum_1_clock = clock; // @[:@39113.4]
  assign x356_sum_1_reset = reset; // @[:@39114.4]
  assign x356_sum_1_io_a = RetimeWrapper_9_io_out; // @[Math.scala 151:17:@39115.4]
  assign x356_sum_1_io_b = x355_div_1_io_result; // @[Math.scala 152:17:@39116.4]
  assign x356_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@39117.4]
  assign RetimeWrapper_14_clock = clock; // @[:@39123.4]
  assign RetimeWrapper_14_reset = reset; // @[:@39124.4]
  assign RetimeWrapper_14_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39126.4]
  assign RetimeWrapper_14_io_in = x614_x330_D1_0_number[23:16]; // @[package.scala 94:16:@39125.4]
  assign RetimeWrapper_15_clock = clock; // @[:@39132.4]
  assign RetimeWrapper_15_reset = reset; // @[:@39133.4]
  assign RetimeWrapper_15_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39135.4]
  assign RetimeWrapper_15_io_in = x356_sum_1_io_result; // @[package.scala 94:16:@39134.4]
  assign RetimeWrapper_16_clock = clock; // @[:@39141.4]
  assign RetimeWrapper_16_reset = reset; // @[:@39142.4]
  assign RetimeWrapper_16_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39144.4]
  assign RetimeWrapper_16_io_in = x354_1_io_result; // @[package.scala 94:16:@39143.4]
  assign RetimeWrapper_17_clock = clock; // @[:@39152.4]
  assign RetimeWrapper_17_reset = reset; // @[:@39153.4]
  assign RetimeWrapper_17_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39155.4]
  assign RetimeWrapper_17_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@39154.4]
  assign x358_rdcol_1_clock = clock; // @[:@39175.4]
  assign x358_rdcol_1_reset = reset; // @[:@39176.4]
  assign x358_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@39177.4]
  assign x358_rdcol_1_io_b = 32'h3; // @[Math.scala 152:17:@39178.4]
  assign x358_rdcol_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@39179.4]
  assign x360_1_clock = clock; // @[:@39189.4]
  assign x360_1_reset = reset; // @[:@39190.4]
  assign x360_1_io_a = x358_rdcol_1_io_result; // @[Math.scala 367:17:@39191.4]
  assign x360_1_io_b = 32'h6; // @[Math.scala 368:17:@39192.4]
  assign x360_1_io_flow = io_in_x317_TREADY; // @[Math.scala 369:20:@39193.4]
  assign x361_div_1_clock = clock; // @[:@39201.4]
  assign x361_div_1_reset = reset; // @[:@39202.4]
  assign x361_div_1_io_a = x358_rdcol_1_io_result; // @[Math.scala 328:17:@39203.4]
  assign x361_div_1_io_flow = io_in_x317_TREADY; // @[Math.scala 330:20:@39205.4]
  assign x362_sum_1_clock = clock; // @[:@39211.4]
  assign x362_sum_1_reset = reset; // @[:@39212.4]
  assign x362_sum_1_io_a = RetimeWrapper_9_io_out; // @[Math.scala 151:17:@39213.4]
  assign x362_sum_1_io_b = x361_div_1_io_result; // @[Math.scala 152:17:@39214.4]
  assign x362_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@39215.4]
  assign RetimeWrapper_18_clock = clock; // @[:@39221.4]
  assign RetimeWrapper_18_reset = reset; // @[:@39222.4]
  assign RetimeWrapper_18_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39224.4]
  assign RetimeWrapper_18_io_in = x360_1_io_result; // @[package.scala 94:16:@39223.4]
  assign RetimeWrapper_19_clock = clock; // @[:@39230.4]
  assign RetimeWrapper_19_reset = reset; // @[:@39231.4]
  assign RetimeWrapper_19_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39233.4]
  assign RetimeWrapper_19_io_in = x362_sum_1_io_result; // @[package.scala 94:16:@39232.4]
  assign RetimeWrapper_20_clock = clock; // @[:@39239.4]
  assign RetimeWrapper_20_reset = reset; // @[:@39240.4]
  assign RetimeWrapper_20_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39242.4]
  assign RetimeWrapper_20_io_in = x614_x330_D1_0_number[31:24]; // @[package.scala 94:16:@39241.4]
  assign RetimeWrapper_21_clock = clock; // @[:@39250.4]
  assign RetimeWrapper_21_reset = reset; // @[:@39251.4]
  assign RetimeWrapper_21_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39253.4]
  assign RetimeWrapper_21_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@39252.4]
  assign RetimeWrapper_22_clock = clock; // @[:@39271.4]
  assign RetimeWrapper_22_reset = reset; // @[:@39272.4]
  assign RetimeWrapper_22_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39274.4]
  assign RetimeWrapper_22_io_in = __io_result; // @[package.scala 94:16:@39273.4]
  assign x365_1_clock = clock; // @[:@39284.4]
  assign x365_1_reset = reset; // @[:@39285.4]
  assign x365_1_io_a = RetimeWrapper_22_io_out; // @[Math.scala 367:17:@39286.4]
  assign x365_1_io_b = 32'h780; // @[Math.scala 368:17:@39287.4]
  assign x365_1_io_flow = io_in_x317_TREADY; // @[Math.scala 369:20:@39288.4]
  assign RetimeWrapper_23_clock = clock; // @[:@39299.4]
  assign RetimeWrapper_23_reset = reset; // @[:@39300.4]
  assign RetimeWrapper_23_io_flow = io_in_x317_TREADY; // @[package.scala 95:18:@39302.4]
  assign RetimeWrapper_23_io_in = $signed(_T_549) < $signed(32'sh0); // @[package.scala 94:16:@39301.4]
  assign RetimeWrapper_24_clock = clock; // @[:@39308.4]
  assign RetimeWrapper_24_reset = reset; // @[:@39309.4]
  assign RetimeWrapper_24_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39311.4]
  assign RetimeWrapper_24_io_in = x358_rdcol_1_io_result; // @[package.scala 94:16:@39310.4]
  assign RetimeWrapper_25_clock = clock; // @[:@39322.4]
  assign RetimeWrapper_25_reset = reset; // @[:@39323.4]
  assign RetimeWrapper_25_io_flow = io_in_x317_TREADY; // @[package.scala 95:18:@39325.4]
  assign RetimeWrapper_25_io_in = $signed(_T_562) < $signed(32'sh0); // @[package.scala 94:16:@39324.4]
  assign RetimeWrapper_26_clock = clock; // @[:@39331.4]
  assign RetimeWrapper_26_reset = reset; // @[:@39332.4]
  assign RetimeWrapper_26_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39334.4]
  assign RetimeWrapper_26_io_in = RetimeWrapper_23_io_out; // @[package.scala 94:16:@39333.4]
  assign x372_mul_1_clock = clock; // @[:@39368.4]
  assign x372_mul_1_reset = reset; // @[:@39369.4]
  assign x372_mul_1_io_a = {_T_593,_T_594}; // @[Math.scala 263:17:@39370.4]
  assign x372_mul_1_io_flow = io_in_x317_TREADY; // @[Math.scala 265:20:@39372.4]
  assign RetimeWrapper_27_clock = clock; // @[:@39378.4]
  assign RetimeWrapper_27_reset = reset; // @[:@39379.4]
  assign RetimeWrapper_27_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39381.4]
  assign RetimeWrapper_27_io_in = x361_div_1_io_result; // @[package.scala 94:16:@39380.4]
  assign x373_sum_1_clock = clock; // @[:@39387.4]
  assign x373_sum_1_reset = reset; // @[:@39388.4]
  assign x373_sum_1_io_a = x372_mul_1_io_result; // @[Math.scala 151:17:@39389.4]
  assign x373_sum_1_io_b = RetimeWrapper_27_io_out; // @[Math.scala 152:17:@39390.4]
  assign x373_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@39391.4]
  assign RetimeWrapper_28_clock = clock; // @[:@39397.4]
  assign RetimeWrapper_28_reset = reset; // @[:@39398.4]
  assign RetimeWrapper_28_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39400.4]
  assign RetimeWrapper_28_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@39399.4]
  assign RetimeWrapper_29_clock = clock; // @[:@39406.4]
  assign RetimeWrapper_29_reset = reset; // @[:@39407.4]
  assign RetimeWrapper_29_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39409.4]
  assign RetimeWrapper_29_io_in = x360_1_io_result; // @[package.scala 94:16:@39408.4]
  assign RetimeWrapper_30_clock = clock; // @[:@39415.4]
  assign RetimeWrapper_30_reset = reset; // @[:@39416.4]
  assign RetimeWrapper_30_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39418.4]
  assign RetimeWrapper_30_io_in = $unsigned(_T_584); // @[package.scala 94:16:@39417.4]
  assign RetimeWrapper_31_clock = clock; // @[:@39424.4]
  assign RetimeWrapper_31_reset = reset; // @[:@39425.4]
  assign RetimeWrapper_31_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39427.4]
  assign RetimeWrapper_31_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@39426.4]
  assign RetimeWrapper_32_clock = clock; // @[:@39433.4]
  assign RetimeWrapper_32_reset = reset; // @[:@39434.4]
  assign RetimeWrapper_32_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39436.4]
  assign RetimeWrapper_32_io_in = x373_sum_1_io_result; // @[package.scala 94:16:@39435.4]
  assign RetimeWrapper_33_clock = clock; // @[:@39442.4]
  assign RetimeWrapper_33_reset = reset; // @[:@39443.4]
  assign RetimeWrapper_33_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39445.4]
  assign RetimeWrapper_33_io_in = ~ x368; // @[package.scala 94:16:@39444.4]
  assign RetimeWrapper_34_clock = clock; // @[:@39454.4]
  assign RetimeWrapper_34_reset = reset; // @[:@39455.4]
  assign RetimeWrapper_34_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39457.4]
  assign RetimeWrapper_34_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@39456.4]
  assign RetimeWrapper_35_clock = clock; // @[:@39475.4]
  assign RetimeWrapper_35_reset = reset; // @[:@39476.4]
  assign RetimeWrapper_35_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39478.4]
  assign RetimeWrapper_35_io_in = x352_rdcol_1_io_result; // @[package.scala 94:16:@39477.4]
  assign RetimeWrapper_36_clock = clock; // @[:@39489.4]
  assign RetimeWrapper_36_reset = reset; // @[:@39490.4]
  assign RetimeWrapper_36_io_flow = io_in_x317_TREADY; // @[package.scala 95:18:@39492.4]
  assign RetimeWrapper_36_io_in = $signed(_T_654) < $signed(32'sh0); // @[package.scala 94:16:@39491.4]
  assign RetimeWrapper_37_clock = clock; // @[:@39504.4]
  assign RetimeWrapper_37_reset = reset; // @[:@39505.4]
  assign RetimeWrapper_37_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39507.4]
  assign RetimeWrapper_37_io_in = x355_div_1_io_result; // @[package.scala 94:16:@39506.4]
  assign x379_sum_1_clock = clock; // @[:@39513.4]
  assign x379_sum_1_reset = reset; // @[:@39514.4]
  assign x379_sum_1_io_a = x372_mul_1_io_result; // @[Math.scala 151:17:@39515.4]
  assign x379_sum_1_io_b = RetimeWrapper_37_io_out; // @[Math.scala 152:17:@39516.4]
  assign x379_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@39517.4]
  assign RetimeWrapper_38_clock = clock; // @[:@39523.4]
  assign RetimeWrapper_38_reset = reset; // @[:@39524.4]
  assign RetimeWrapper_38_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39526.4]
  assign RetimeWrapper_38_io_in = x379_sum_1_io_result; // @[package.scala 94:16:@39525.4]
  assign RetimeWrapper_39_clock = clock; // @[:@39532.4]
  assign RetimeWrapper_39_reset = reset; // @[:@39533.4]
  assign RetimeWrapper_39_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39535.4]
  assign RetimeWrapper_39_io_in = ~ x377; // @[package.scala 94:16:@39534.4]
  assign RetimeWrapper_40_clock = clock; // @[:@39541.4]
  assign RetimeWrapper_40_reset = reset; // @[:@39542.4]
  assign RetimeWrapper_40_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39544.4]
  assign RetimeWrapper_40_io_in = x354_1_io_result; // @[package.scala 94:16:@39543.4]
  assign RetimeWrapper_41_clock = clock; // @[:@39553.4]
  assign RetimeWrapper_41_reset = reset; // @[:@39554.4]
  assign RetimeWrapper_41_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39556.4]
  assign RetimeWrapper_41_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@39555.4]
  assign RetimeWrapper_42_clock = clock; // @[:@39574.4]
  assign RetimeWrapper_42_reset = reset; // @[:@39575.4]
  assign RetimeWrapper_42_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39577.4]
  assign RetimeWrapper_42_io_in = x346_rdcol_1_io_result; // @[package.scala 94:16:@39576.4]
  assign RetimeWrapper_43_clock = clock; // @[:@39588.4]
  assign RetimeWrapper_43_reset = reset; // @[:@39589.4]
  assign RetimeWrapper_43_io_flow = io_in_x317_TREADY; // @[package.scala 95:18:@39591.4]
  assign RetimeWrapper_43_io_in = $signed(_T_705) < $signed(32'sh0); // @[package.scala 94:16:@39590.4]
  assign RetimeWrapper_44_clock = clock; // @[:@39603.4]
  assign RetimeWrapper_44_reset = reset; // @[:@39604.4]
  assign RetimeWrapper_44_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39606.4]
  assign RetimeWrapper_44_io_in = x349_div_1_io_result; // @[package.scala 94:16:@39605.4]
  assign x385_sum_1_clock = clock; // @[:@39612.4]
  assign x385_sum_1_reset = reset; // @[:@39613.4]
  assign x385_sum_1_io_a = x372_mul_1_io_result; // @[Math.scala 151:17:@39614.4]
  assign x385_sum_1_io_b = RetimeWrapper_44_io_out; // @[Math.scala 152:17:@39615.4]
  assign x385_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@39616.4]
  assign RetimeWrapper_45_clock = clock; // @[:@39622.4]
  assign RetimeWrapper_45_reset = reset; // @[:@39623.4]
  assign RetimeWrapper_45_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39625.4]
  assign RetimeWrapper_45_io_in = x385_sum_1_io_result; // @[package.scala 94:16:@39624.4]
  assign RetimeWrapper_46_clock = clock; // @[:@39631.4]
  assign RetimeWrapper_46_reset = reset; // @[:@39632.4]
  assign RetimeWrapper_46_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39634.4]
  assign RetimeWrapper_46_io_in = ~ x383; // @[package.scala 94:16:@39633.4]
  assign RetimeWrapper_47_clock = clock; // @[:@39640.4]
  assign RetimeWrapper_47_reset = reset; // @[:@39641.4]
  assign RetimeWrapper_47_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39643.4]
  assign RetimeWrapper_47_io_in = x348_1_io_result; // @[package.scala 94:16:@39642.4]
  assign RetimeWrapper_48_clock = clock; // @[:@39652.4]
  assign RetimeWrapper_48_reset = reset; // @[:@39653.4]
  assign RetimeWrapper_48_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39655.4]
  assign RetimeWrapper_48_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@39654.4]
  assign RetimeWrapper_49_clock = clock; // @[:@39673.4]
  assign RetimeWrapper_49_reset = reset; // @[:@39674.4]
  assign RetimeWrapper_49_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39676.4]
  assign RetimeWrapper_49_io_in = __1_io_result; // @[package.scala 94:16:@39675.4]
  assign RetimeWrapper_50_clock = clock; // @[:@39689.4]
  assign RetimeWrapper_50_reset = reset; // @[:@39690.4]
  assign RetimeWrapper_50_io_flow = io_in_x317_TREADY; // @[package.scala 95:18:@39692.4]
  assign RetimeWrapper_50_io_in = $signed(_T_758) < $signed(32'sh0); // @[package.scala 94:16:@39691.4]
  assign RetimeWrapper_51_clock = clock; // @[:@39704.4]
  assign RetimeWrapper_51_reset = reset; // @[:@39705.4]
  assign RetimeWrapper_51_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39707.4]
  assign RetimeWrapper_51_io_in = x343_div_1_io_result; // @[package.scala 94:16:@39706.4]
  assign x391_sum_1_clock = clock; // @[:@39713.4]
  assign x391_sum_1_reset = reset; // @[:@39714.4]
  assign x391_sum_1_io_a = x372_mul_1_io_result; // @[Math.scala 151:17:@39715.4]
  assign x391_sum_1_io_b = RetimeWrapper_51_io_out; // @[Math.scala 152:17:@39716.4]
  assign x391_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@39717.4]
  assign RetimeWrapper_52_clock = clock; // @[:@39723.4]
  assign RetimeWrapper_52_reset = reset; // @[:@39724.4]
  assign RetimeWrapper_52_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39726.4]
  assign RetimeWrapper_52_io_in = x340_1_io_result; // @[package.scala 94:16:@39725.4]
  assign RetimeWrapper_53_clock = clock; // @[:@39732.4]
  assign RetimeWrapper_53_reset = reset; // @[:@39733.4]
  assign RetimeWrapper_53_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39735.4]
  assign RetimeWrapper_53_io_in = x391_sum_1_io_result; // @[package.scala 94:16:@39734.4]
  assign RetimeWrapper_54_clock = clock; // @[:@39741.4]
  assign RetimeWrapper_54_reset = reset; // @[:@39742.4]
  assign RetimeWrapper_54_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39744.4]
  assign RetimeWrapper_54_io_in = ~ x389; // @[package.scala 94:16:@39743.4]
  assign RetimeWrapper_55_clock = clock; // @[:@39753.4]
  assign RetimeWrapper_55_reset = reset; // @[:@39754.4]
  assign RetimeWrapper_55_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39756.4]
  assign RetimeWrapper_55_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@39755.4]
  assign x394_rdcol_1_clock = clock; // @[:@39776.4]
  assign x394_rdcol_1_reset = reset; // @[:@39777.4]
  assign x394_rdcol_1_io_a = RetimeWrapper_49_io_out; // @[Math.scala 151:17:@39778.4]
  assign x394_rdcol_1_io_b = 32'hffffffff; // @[Math.scala 152:17:@39779.4]
  assign x394_rdcol_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@39780.4]
  assign RetimeWrapper_56_clock = clock; // @[:@39791.4]
  assign RetimeWrapper_56_reset = reset; // @[:@39792.4]
  assign RetimeWrapper_56_io_flow = io_in_x317_TREADY; // @[package.scala 95:18:@39794.4]
  assign RetimeWrapper_56_io_in = $signed(_T_813) < $signed(32'sh0); // @[package.scala 94:16:@39793.4]
  assign x398_1_clock = clock; // @[:@39808.4]
  assign x398_1_reset = reset; // @[:@39809.4]
  assign x398_1_io_a = x394_rdcol_1_io_result; // @[Math.scala 367:17:@39810.4]
  assign x398_1_io_b = 32'h6; // @[Math.scala 368:17:@39811.4]
  assign x398_1_io_flow = io_in_x317_TREADY; // @[Math.scala 369:20:@39812.4]
  assign x399_div_1_clock = clock; // @[:@39820.4]
  assign x399_div_1_reset = reset; // @[:@39821.4]
  assign x399_div_1_io_a = x394_rdcol_1_io_result; // @[Math.scala 328:17:@39822.4]
  assign x399_div_1_io_flow = io_in_x317_TREADY; // @[Math.scala 330:20:@39824.4]
  assign RetimeWrapper_57_clock = clock; // @[:@39830.4]
  assign RetimeWrapper_57_reset = reset; // @[:@39831.4]
  assign RetimeWrapper_57_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39833.4]
  assign RetimeWrapper_57_io_in = x399_div_1_io_result; // @[package.scala 94:16:@39832.4]
  assign x400_sum_1_clock = clock; // @[:@39839.4]
  assign x400_sum_1_reset = reset; // @[:@39840.4]
  assign x400_sum_1_io_a = x372_mul_1_io_result; // @[Math.scala 151:17:@39841.4]
  assign x400_sum_1_io_b = RetimeWrapper_57_io_out; // @[Math.scala 152:17:@39842.4]
  assign x400_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@39843.4]
  assign RetimeWrapper_58_clock = clock; // @[:@39849.4]
  assign RetimeWrapper_58_reset = reset; // @[:@39850.4]
  assign RetimeWrapper_58_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39852.4]
  assign RetimeWrapper_58_io_in = ~ x396; // @[package.scala 94:16:@39851.4]
  assign RetimeWrapper_59_clock = clock; // @[:@39858.4]
  assign RetimeWrapper_59_reset = reset; // @[:@39859.4]
  assign RetimeWrapper_59_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39861.4]
  assign RetimeWrapper_59_io_in = x398_1_io_result; // @[package.scala 94:16:@39860.4]
  assign RetimeWrapper_60_clock = clock; // @[:@39867.4]
  assign RetimeWrapper_60_reset = reset; // @[:@39868.4]
  assign RetimeWrapper_60_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39870.4]
  assign RetimeWrapper_60_io_in = x400_sum_1_io_result; // @[package.scala 94:16:@39869.4]
  assign RetimeWrapper_61_clock = clock; // @[:@39879.4]
  assign RetimeWrapper_61_reset = reset; // @[:@39880.4]
  assign RetimeWrapper_61_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39882.4]
  assign RetimeWrapper_61_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@39881.4]
  assign x403_rdcol_1_clock = clock; // @[:@39902.4]
  assign x403_rdcol_1_reset = reset; // @[:@39903.4]
  assign x403_rdcol_1_io_a = RetimeWrapper_49_io_out; // @[Math.scala 151:17:@39904.4]
  assign x403_rdcol_1_io_b = 32'hfffffffe; // @[Math.scala 152:17:@39905.4]
  assign x403_rdcol_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@39906.4]
  assign RetimeWrapper_62_clock = clock; // @[:@39917.4]
  assign RetimeWrapper_62_reset = reset; // @[:@39918.4]
  assign RetimeWrapper_62_io_flow = io_in_x317_TREADY; // @[package.scala 95:18:@39920.4]
  assign RetimeWrapper_62_io_in = $signed(_T_882) < $signed(32'sh0); // @[package.scala 94:16:@39919.4]
  assign x407_1_clock = clock; // @[:@39934.4]
  assign x407_1_reset = reset; // @[:@39935.4]
  assign x407_1_io_a = x403_rdcol_1_io_result; // @[Math.scala 367:17:@39936.4]
  assign x407_1_io_b = 32'h6; // @[Math.scala 368:17:@39937.4]
  assign x407_1_io_flow = io_in_x317_TREADY; // @[Math.scala 369:20:@39938.4]
  assign x408_div_1_clock = clock; // @[:@39946.4]
  assign x408_div_1_reset = reset; // @[:@39947.4]
  assign x408_div_1_io_a = x403_rdcol_1_io_result; // @[Math.scala 328:17:@39948.4]
  assign x408_div_1_io_flow = io_in_x317_TREADY; // @[Math.scala 330:20:@39950.4]
  assign RetimeWrapper_63_clock = clock; // @[:@39956.4]
  assign RetimeWrapper_63_reset = reset; // @[:@39957.4]
  assign RetimeWrapper_63_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39959.4]
  assign RetimeWrapper_63_io_in = x408_div_1_io_result; // @[package.scala 94:16:@39958.4]
  assign x409_sum_1_clock = clock; // @[:@39965.4]
  assign x409_sum_1_reset = reset; // @[:@39966.4]
  assign x409_sum_1_io_a = x372_mul_1_io_result; // @[Math.scala 151:17:@39967.4]
  assign x409_sum_1_io_b = RetimeWrapper_63_io_out; // @[Math.scala 152:17:@39968.4]
  assign x409_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@39969.4]
  assign RetimeWrapper_64_clock = clock; // @[:@39975.4]
  assign RetimeWrapper_64_reset = reset; // @[:@39976.4]
  assign RetimeWrapper_64_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39978.4]
  assign RetimeWrapper_64_io_in = x407_1_io_result; // @[package.scala 94:16:@39977.4]
  assign RetimeWrapper_65_clock = clock; // @[:@39984.4]
  assign RetimeWrapper_65_reset = reset; // @[:@39985.4]
  assign RetimeWrapper_65_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39987.4]
  assign RetimeWrapper_65_io_in = ~ x405; // @[package.scala 94:16:@39986.4]
  assign RetimeWrapper_66_clock = clock; // @[:@39993.4]
  assign RetimeWrapper_66_reset = reset; // @[:@39994.4]
  assign RetimeWrapper_66_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39996.4]
  assign RetimeWrapper_66_io_in = x409_sum_1_io_result; // @[package.scala 94:16:@39995.4]
  assign RetimeWrapper_67_clock = clock; // @[:@40005.4]
  assign RetimeWrapper_67_reset = reset; // @[:@40006.4]
  assign RetimeWrapper_67_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40008.4]
  assign RetimeWrapper_67_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@40007.4]
  assign x412_rdrow_1_clock = clock; // @[:@40028.4]
  assign x412_rdrow_1_reset = reset; // @[:@40029.4]
  assign x412_rdrow_1_io_a = RetimeWrapper_22_io_out; // @[Math.scala 192:17:@40030.4]
  assign x412_rdrow_1_io_b = 32'h1; // @[Math.scala 193:17:@40031.4]
  assign x412_rdrow_1_io_flow = io_in_x317_TREADY; // @[Math.scala 194:20:@40032.4]
  assign x413_1_clock = clock; // @[:@40040.4]
  assign x413_1_reset = reset; // @[:@40041.4]
  assign x413_1_io_a = x412_rdrow_1_io_result; // @[Math.scala 367:17:@40042.4]
  assign x413_1_io_b = 32'h780; // @[Math.scala 368:17:@40043.4]
  assign x413_1_io_flow = io_in_x317_TREADY; // @[Math.scala 369:20:@40044.4]
  assign RetimeWrapper_68_clock = clock; // @[:@40055.4]
  assign RetimeWrapper_68_reset = reset; // @[:@40056.4]
  assign RetimeWrapper_68_io_flow = io_in_x317_TREADY; // @[package.scala 95:18:@40058.4]
  assign RetimeWrapper_68_io_in = $signed(_T_958) < $signed(32'sh0); // @[package.scala 94:16:@40057.4]
  assign x419_mul_1_clock = clock; // @[:@40092.4]
  assign x419_mul_1_reset = reset; // @[:@40093.4]
  assign x419_mul_1_io_a = {_T_986,_T_987}; // @[Math.scala 263:17:@40094.4]
  assign x419_mul_1_io_flow = io_in_x317_TREADY; // @[Math.scala 265:20:@40096.4]
  assign RetimeWrapper_69_clock = clock; // @[:@40102.4]
  assign RetimeWrapper_69_reset = reset; // @[:@40103.4]
  assign RetimeWrapper_69_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40105.4]
  assign RetimeWrapper_69_io_in = x361_div_1_io_result; // @[package.scala 94:16:@40104.4]
  assign x420_sum_1_clock = clock; // @[:@40111.4]
  assign x420_sum_1_reset = reset; // @[:@40112.4]
  assign x420_sum_1_io_a = x419_mul_1_io_result; // @[Math.scala 151:17:@40113.4]
  assign x420_sum_1_io_b = RetimeWrapper_69_io_out; // @[Math.scala 152:17:@40114.4]
  assign x420_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@40115.4]
  assign RetimeWrapper_70_clock = clock; // @[:@40121.4]
  assign RetimeWrapper_70_reset = reset; // @[:@40122.4]
  assign RetimeWrapper_70_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40124.4]
  assign RetimeWrapper_70_io_in = ~ x415; // @[package.scala 94:16:@40123.4]
  assign RetimeWrapper_71_clock = clock; // @[:@40130.4]
  assign RetimeWrapper_71_reset = reset; // @[:@40131.4]
  assign RetimeWrapper_71_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40133.4]
  assign RetimeWrapper_71_io_in = $unsigned(_T_977); // @[package.scala 94:16:@40132.4]
  assign RetimeWrapper_72_clock = clock; // @[:@40142.4]
  assign RetimeWrapper_72_reset = reset; // @[:@40143.4]
  assign RetimeWrapper_72_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40145.4]
  assign RetimeWrapper_72_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@40144.4]
  assign RetimeWrapper_73_clock = clock; // @[:@40169.4]
  assign RetimeWrapper_73_reset = reset; // @[:@40170.4]
  assign RetimeWrapper_73_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40172.4]
  assign RetimeWrapper_73_io_in = x355_div_1_io_result; // @[package.scala 94:16:@40171.4]
  assign x425_sum_1_clock = clock; // @[:@40180.4]
  assign x425_sum_1_reset = reset; // @[:@40181.4]
  assign x425_sum_1_io_a = x419_mul_1_io_result; // @[Math.scala 151:17:@40182.4]
  assign x425_sum_1_io_b = RetimeWrapper_73_io_out; // @[Math.scala 152:17:@40183.4]
  assign x425_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@40184.4]
  assign RetimeWrapper_74_clock = clock; // @[:@40190.4]
  assign RetimeWrapper_74_reset = reset; // @[:@40191.4]
  assign RetimeWrapper_74_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40193.4]
  assign RetimeWrapper_74_io_in = ~ x423; // @[package.scala 94:16:@40192.4]
  assign RetimeWrapper_75_clock = clock; // @[:@40202.4]
  assign RetimeWrapper_75_reset = reset; // @[:@40203.4]
  assign RetimeWrapper_75_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40205.4]
  assign RetimeWrapper_75_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@40204.4]
  assign RetimeWrapper_76_clock = clock; // @[:@40229.4]
  assign RetimeWrapper_76_reset = reset; // @[:@40230.4]
  assign RetimeWrapper_76_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40232.4]
  assign RetimeWrapper_76_io_in = x349_div_1_io_result; // @[package.scala 94:16:@40231.4]
  assign x430_sum_1_clock = clock; // @[:@40238.4]
  assign x430_sum_1_reset = reset; // @[:@40239.4]
  assign x430_sum_1_io_a = x419_mul_1_io_result; // @[Math.scala 151:17:@40240.4]
  assign x430_sum_1_io_b = RetimeWrapper_76_io_out; // @[Math.scala 152:17:@40241.4]
  assign x430_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@40242.4]
  assign RetimeWrapper_77_clock = clock; // @[:@40248.4]
  assign RetimeWrapper_77_reset = reset; // @[:@40249.4]
  assign RetimeWrapper_77_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40251.4]
  assign RetimeWrapper_77_io_in = ~ x428; // @[package.scala 94:16:@40250.4]
  assign RetimeWrapper_78_clock = clock; // @[:@40260.4]
  assign RetimeWrapper_78_reset = reset; // @[:@40261.4]
  assign RetimeWrapper_78_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40263.4]
  assign RetimeWrapper_78_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@40262.4]
  assign RetimeWrapper_79_clock = clock; // @[:@40281.4]
  assign RetimeWrapper_79_reset = reset; // @[:@40282.4]
  assign RetimeWrapper_79_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40284.4]
  assign RetimeWrapper_79_io_in = RetimeWrapper_50_io_out; // @[package.scala 94:16:@40283.4]
  assign RetimeWrapper_80_clock = clock; // @[:@40296.4]
  assign RetimeWrapper_80_reset = reset; // @[:@40297.4]
  assign RetimeWrapper_80_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40299.4]
  assign RetimeWrapper_80_io_in = x343_div_1_io_result; // @[package.scala 94:16:@40298.4]
  assign x435_sum_1_clock = clock; // @[:@40305.4]
  assign x435_sum_1_reset = reset; // @[:@40306.4]
  assign x435_sum_1_io_a = x419_mul_1_io_result; // @[Math.scala 151:17:@40307.4]
  assign x435_sum_1_io_b = RetimeWrapper_80_io_out; // @[Math.scala 152:17:@40308.4]
  assign x435_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@40309.4]
  assign RetimeWrapper_81_clock = clock; // @[:@40315.4]
  assign RetimeWrapper_81_reset = reset; // @[:@40316.4]
  assign RetimeWrapper_81_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40318.4]
  assign RetimeWrapper_81_io_in = ~ x433; // @[package.scala 94:16:@40317.4]
  assign RetimeWrapper_82_clock = clock; // @[:@40327.4]
  assign RetimeWrapper_82_reset = reset; // @[:@40328.4]
  assign RetimeWrapper_82_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40330.4]
  assign RetimeWrapper_82_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@40329.4]
  assign RetimeWrapper_83_clock = clock; // @[:@40354.4]
  assign RetimeWrapper_83_reset = reset; // @[:@40355.4]
  assign RetimeWrapper_83_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40357.4]
  assign RetimeWrapper_83_io_in = x399_div_1_io_result; // @[package.scala 94:16:@40356.4]
  assign x440_sum_1_clock = clock; // @[:@40363.4]
  assign x440_sum_1_reset = reset; // @[:@40364.4]
  assign x440_sum_1_io_a = x419_mul_1_io_result; // @[Math.scala 151:17:@40365.4]
  assign x440_sum_1_io_b = RetimeWrapper_83_io_out; // @[Math.scala 152:17:@40366.4]
  assign x440_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@40367.4]
  assign RetimeWrapper_84_clock = clock; // @[:@40373.4]
  assign RetimeWrapper_84_reset = reset; // @[:@40374.4]
  assign RetimeWrapper_84_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40376.4]
  assign RetimeWrapper_84_io_in = ~ x438; // @[package.scala 94:16:@40375.4]
  assign RetimeWrapper_85_clock = clock; // @[:@40385.4]
  assign RetimeWrapper_85_reset = reset; // @[:@40386.4]
  assign RetimeWrapper_85_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40388.4]
  assign RetimeWrapper_85_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@40387.4]
  assign RetimeWrapper_86_clock = clock; // @[:@40412.4]
  assign RetimeWrapper_86_reset = reset; // @[:@40413.4]
  assign RetimeWrapper_86_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40415.4]
  assign RetimeWrapper_86_io_in = x408_div_1_io_result; // @[package.scala 94:16:@40414.4]
  assign x445_sum_1_clock = clock; // @[:@40421.4]
  assign x445_sum_1_reset = reset; // @[:@40422.4]
  assign x445_sum_1_io_a = x419_mul_1_io_result; // @[Math.scala 151:17:@40423.4]
  assign x445_sum_1_io_b = RetimeWrapper_86_io_out; // @[Math.scala 152:17:@40424.4]
  assign x445_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@40425.4]
  assign RetimeWrapper_87_clock = clock; // @[:@40431.4]
  assign RetimeWrapper_87_reset = reset; // @[:@40432.4]
  assign RetimeWrapper_87_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40434.4]
  assign RetimeWrapper_87_io_in = ~ x443; // @[package.scala 94:16:@40433.4]
  assign RetimeWrapper_88_clock = clock; // @[:@40443.4]
  assign RetimeWrapper_88_reset = reset; // @[:@40444.4]
  assign RetimeWrapper_88_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40446.4]
  assign RetimeWrapper_88_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@40445.4]
  assign x448_rdrow_1_clock = clock; // @[:@40466.4]
  assign x448_rdrow_1_reset = reset; // @[:@40467.4]
  assign x448_rdrow_1_io_a = RetimeWrapper_22_io_out; // @[Math.scala 192:17:@40468.4]
  assign x448_rdrow_1_io_b = 32'h2; // @[Math.scala 193:17:@40469.4]
  assign x448_rdrow_1_io_flow = io_in_x317_TREADY; // @[Math.scala 194:20:@40470.4]
  assign x449_1_clock = clock; // @[:@40478.4]
  assign x449_1_reset = reset; // @[:@40479.4]
  assign x449_1_io_a = x448_rdrow_1_io_result; // @[Math.scala 367:17:@40480.4]
  assign x449_1_io_b = 32'h780; // @[Math.scala 368:17:@40481.4]
  assign x449_1_io_flow = io_in_x317_TREADY; // @[Math.scala 369:20:@40482.4]
  assign RetimeWrapper_89_clock = clock; // @[:@40493.4]
  assign RetimeWrapper_89_reset = reset; // @[:@40494.4]
  assign RetimeWrapper_89_io_flow = io_in_x317_TREADY; // @[package.scala 95:18:@40496.4]
  assign RetimeWrapper_89_io_in = $signed(_T_1211) < $signed(32'sh0); // @[package.scala 94:16:@40495.4]
  assign x455_mul_1_clock = clock; // @[:@40530.4]
  assign x455_mul_1_reset = reset; // @[:@40531.4]
  assign x455_mul_1_io_a = {_T_1239,_T_1240}; // @[Math.scala 263:17:@40532.4]
  assign x455_mul_1_io_flow = io_in_x317_TREADY; // @[Math.scala 265:20:@40534.4]
  assign x456_sum_1_clock = clock; // @[:@40540.4]
  assign x456_sum_1_reset = reset; // @[:@40541.4]
  assign x456_sum_1_io_a = x455_mul_1_io_result; // @[Math.scala 151:17:@40542.4]
  assign x456_sum_1_io_b = RetimeWrapper_69_io_out; // @[Math.scala 152:17:@40543.4]
  assign x456_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@40544.4]
  assign RetimeWrapper_90_clock = clock; // @[:@40550.4]
  assign RetimeWrapper_90_reset = reset; // @[:@40551.4]
  assign RetimeWrapper_90_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40553.4]
  assign RetimeWrapper_90_io_in = ~ x451; // @[package.scala 94:16:@40552.4]
  assign RetimeWrapper_91_clock = clock; // @[:@40559.4]
  assign RetimeWrapper_91_reset = reset; // @[:@40560.4]
  assign RetimeWrapper_91_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40562.4]
  assign RetimeWrapper_91_io_in = $unsigned(_T_1230); // @[package.scala 94:16:@40561.4]
  assign RetimeWrapper_92_clock = clock; // @[:@40571.4]
  assign RetimeWrapper_92_reset = reset; // @[:@40572.4]
  assign RetimeWrapper_92_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40574.4]
  assign RetimeWrapper_92_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@40573.4]
  assign x461_sum_1_clock = clock; // @[:@40600.4]
  assign x461_sum_1_reset = reset; // @[:@40601.4]
  assign x461_sum_1_io_a = x455_mul_1_io_result; // @[Math.scala 151:17:@40602.4]
  assign x461_sum_1_io_b = RetimeWrapper_73_io_out; // @[Math.scala 152:17:@40603.4]
  assign x461_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@40604.4]
  assign RetimeWrapper_93_clock = clock; // @[:@40610.4]
  assign RetimeWrapper_93_reset = reset; // @[:@40611.4]
  assign RetimeWrapper_93_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40613.4]
  assign RetimeWrapper_93_io_in = ~ x459; // @[package.scala 94:16:@40612.4]
  assign RetimeWrapper_94_clock = clock; // @[:@40622.4]
  assign RetimeWrapper_94_reset = reset; // @[:@40623.4]
  assign RetimeWrapper_94_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40625.4]
  assign RetimeWrapper_94_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@40624.4]
  assign x466_sum_1_clock = clock; // @[:@40649.4]
  assign x466_sum_1_reset = reset; // @[:@40650.4]
  assign x466_sum_1_io_a = x455_mul_1_io_result; // @[Math.scala 151:17:@40651.4]
  assign x466_sum_1_io_b = RetimeWrapper_76_io_out; // @[Math.scala 152:17:@40652.4]
  assign x466_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@40653.4]
  assign RetimeWrapper_95_clock = clock; // @[:@40659.4]
  assign RetimeWrapper_95_reset = reset; // @[:@40660.4]
  assign RetimeWrapper_95_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40662.4]
  assign RetimeWrapper_95_io_in = ~ x464; // @[package.scala 94:16:@40661.4]
  assign RetimeWrapper_96_clock = clock; // @[:@40671.4]
  assign RetimeWrapper_96_reset = reset; // @[:@40672.4]
  assign RetimeWrapper_96_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40674.4]
  assign RetimeWrapper_96_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@40673.4]
  assign x471_sum_1_clock = clock; // @[:@40698.4]
  assign x471_sum_1_reset = reset; // @[:@40699.4]
  assign x471_sum_1_io_a = x455_mul_1_io_result; // @[Math.scala 151:17:@40700.4]
  assign x471_sum_1_io_b = RetimeWrapper_80_io_out; // @[Math.scala 152:17:@40701.4]
  assign x471_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@40702.4]
  assign RetimeWrapper_97_clock = clock; // @[:@40708.4]
  assign RetimeWrapper_97_reset = reset; // @[:@40709.4]
  assign RetimeWrapper_97_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40711.4]
  assign RetimeWrapper_97_io_in = ~ x469; // @[package.scala 94:16:@40710.4]
  assign RetimeWrapper_98_clock = clock; // @[:@40720.4]
  assign RetimeWrapper_98_reset = reset; // @[:@40721.4]
  assign RetimeWrapper_98_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40723.4]
  assign RetimeWrapper_98_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@40722.4]
  assign x476_sum_1_clock = clock; // @[:@40747.4]
  assign x476_sum_1_reset = reset; // @[:@40748.4]
  assign x476_sum_1_io_a = x455_mul_1_io_result; // @[Math.scala 151:17:@40749.4]
  assign x476_sum_1_io_b = RetimeWrapper_83_io_out; // @[Math.scala 152:17:@40750.4]
  assign x476_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@40751.4]
  assign RetimeWrapper_99_clock = clock; // @[:@40757.4]
  assign RetimeWrapper_99_reset = reset; // @[:@40758.4]
  assign RetimeWrapper_99_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40760.4]
  assign RetimeWrapper_99_io_in = ~ x474; // @[package.scala 94:16:@40759.4]
  assign RetimeWrapper_100_clock = clock; // @[:@40769.4]
  assign RetimeWrapper_100_reset = reset; // @[:@40770.4]
  assign RetimeWrapper_100_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40772.4]
  assign RetimeWrapper_100_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@40771.4]
  assign x481_sum_1_clock = clock; // @[:@40796.4]
  assign x481_sum_1_reset = reset; // @[:@40797.4]
  assign x481_sum_1_io_a = x455_mul_1_io_result; // @[Math.scala 151:17:@40798.4]
  assign x481_sum_1_io_b = RetimeWrapper_86_io_out; // @[Math.scala 152:17:@40799.4]
  assign x481_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@40800.4]
  assign RetimeWrapper_101_clock = clock; // @[:@40806.4]
  assign RetimeWrapper_101_reset = reset; // @[:@40807.4]
  assign RetimeWrapper_101_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40809.4]
  assign RetimeWrapper_101_io_in = ~ x479; // @[package.scala 94:16:@40808.4]
  assign RetimeWrapper_102_clock = clock; // @[:@40818.4]
  assign RetimeWrapper_102_reset = reset; // @[:@40819.4]
  assign RetimeWrapper_102_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40821.4]
  assign RetimeWrapper_102_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@40820.4]
  assign RetimeWrapper_103_clock = clock; // @[:@40841.4]
  assign RetimeWrapper_103_reset = reset; // @[:@40842.4]
  assign RetimeWrapper_103_io_flow = io_in_x317_TREADY; // @[package.scala 95:18:@40844.4]
  assign RetimeWrapper_103_io_in = _GEN_0 << 1; // @[package.scala 94:16:@40843.4]
  assign RetimeWrapper_104_clock = clock; // @[:@40853.4]
  assign RetimeWrapper_104_reset = reset; // @[:@40854.4]
  assign RetimeWrapper_104_io_flow = io_in_x317_TREADY; // @[package.scala 95:18:@40856.4]
  assign RetimeWrapper_104_io_in = _GEN_1 << 1; // @[package.scala 94:16:@40855.4]
  assign RetimeWrapper_105_clock = clock; // @[:@40865.4]
  assign RetimeWrapper_105_reset = reset; // @[:@40866.4]
  assign RetimeWrapper_105_io_flow = io_in_x317_TREADY; // @[package.scala 95:18:@40868.4]
  assign RetimeWrapper_105_io_in = _GEN_2 << 2; // @[package.scala 94:16:@40867.4]
  assign RetimeWrapper_106_clock = clock; // @[:@40877.4]
  assign RetimeWrapper_106_reset = reset; // @[:@40878.4]
  assign RetimeWrapper_106_io_flow = io_in_x317_TREADY; // @[package.scala 95:18:@40880.4]
  assign RetimeWrapper_106_io_in = _GEN_3 << 1; // @[package.scala 94:16:@40879.4]
  assign RetimeWrapper_107_clock = clock; // @[:@40889.4]
  assign RetimeWrapper_107_reset = reset; // @[:@40890.4]
  assign RetimeWrapper_107_io_flow = io_in_x317_TREADY; // @[package.scala 95:18:@40892.4]
  assign RetimeWrapper_107_io_in = _GEN_4 << 1; // @[package.scala 94:16:@40891.4]
  assign RetimeWrapper_108_clock = clock; // @[:@40899.4]
  assign RetimeWrapper_108_reset = reset; // @[:@40900.4]
  assign RetimeWrapper_108_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40902.4]
  assign RetimeWrapper_108_io_in = x329_lb_0_io_rPort_11_output_0; // @[package.scala 94:16:@40901.4]
  assign RetimeWrapper_109_clock = clock; // @[:@40908.4]
  assign RetimeWrapper_109_reset = reset; // @[:@40909.4]
  assign RetimeWrapper_109_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40911.4]
  assign RetimeWrapper_109_io_in = _T_1429[7:0]; // @[package.scala 94:16:@40910.4]
  assign x489_x11_1_io_a = RetimeWrapper_108_io_out; // @[Math.scala 151:17:@40919.4]
  assign x489_x11_1_io_b = RetimeWrapper_109_io_out; // @[Math.scala 152:17:@40920.4]
  assign RetimeWrapper_110_clock = clock; // @[:@40927.4]
  assign RetimeWrapper_110_reset = reset; // @[:@40928.4]
  assign RetimeWrapper_110_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40930.4]
  assign RetimeWrapper_110_io_in = x329_lb_0_io_rPort_13_output_0; // @[package.scala 94:16:@40929.4]
  assign RetimeWrapper_111_clock = clock; // @[:@40936.4]
  assign RetimeWrapper_111_reset = reset; // @[:@40937.4]
  assign RetimeWrapper_111_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40939.4]
  assign RetimeWrapper_111_io_in = _T_1435[7:0]; // @[package.scala 94:16:@40938.4]
  assign x490_x12_1_io_a = RetimeWrapper_110_io_out; // @[Math.scala 151:17:@40947.4]
  assign x490_x12_1_io_b = RetimeWrapper_111_io_out; // @[Math.scala 152:17:@40948.4]
  assign x491_x11_1_io_a = _T_1441[7:0]; // @[Math.scala 151:17:@40957.4]
  assign x491_x11_1_io_b = _T_1447[7:0]; // @[Math.scala 152:17:@40958.4]
  assign RetimeWrapper_112_clock = clock; // @[:@40965.4]
  assign RetimeWrapper_112_reset = reset; // @[:@40966.4]
  assign RetimeWrapper_112_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40968.4]
  assign RetimeWrapper_112_io_in = x329_lb_0_io_rPort_6_output_0; // @[package.scala 94:16:@40967.4]
  assign x492_x12_1_io_a = RetimeWrapper_112_io_out; // @[Math.scala 151:17:@40976.4]
  assign x492_x12_1_io_b = _T_1453[7:0]; // @[Math.scala 152:17:@40977.4]
  assign RetimeWrapper_113_clock = clock; // @[:@40984.4]
  assign RetimeWrapper_113_reset = reset; // @[:@40985.4]
  assign RetimeWrapper_113_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40987.4]
  assign RetimeWrapper_113_io_in = x490_x12_1_io_result; // @[package.scala 94:16:@40986.4]
  assign RetimeWrapper_114_clock = clock; // @[:@40993.4]
  assign RetimeWrapper_114_reset = reset; // @[:@40994.4]
  assign RetimeWrapper_114_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40996.4]
  assign RetimeWrapper_114_io_in = x489_x11_1_io_result; // @[package.scala 94:16:@40995.4]
  assign x493_x11_1_io_a = RetimeWrapper_114_io_out; // @[Math.scala 151:17:@41004.4]
  assign x493_x11_1_io_b = RetimeWrapper_113_io_out; // @[Math.scala 152:17:@41005.4]
  assign x494_x12_1_io_a = x491_x11_1_io_result; // @[Math.scala 151:17:@41014.4]
  assign x494_x12_1_io_b = x492_x12_1_io_result; // @[Math.scala 152:17:@41015.4]
  assign RetimeWrapper_115_clock = clock; // @[:@41022.4]
  assign RetimeWrapper_115_reset = reset; // @[:@41023.4]
  assign RetimeWrapper_115_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41025.4]
  assign RetimeWrapper_115_io_in = x494_x12_1_io_result; // @[package.scala 94:16:@41024.4]
  assign x495_x11_1_io_a = x493_x11_1_io_result; // @[Math.scala 151:17:@41035.4]
  assign x495_x11_1_io_b = RetimeWrapper_115_io_out; // @[Math.scala 152:17:@41036.4]
  assign RetimeWrapper_116_clock = clock; // @[:@41043.4]
  assign RetimeWrapper_116_reset = reset; // @[:@41044.4]
  assign RetimeWrapper_116_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41046.4]
  assign RetimeWrapper_116_io_in = x329_lb_0_io_rPort_5_output_0; // @[package.scala 94:16:@41045.4]
  assign x496_sum_1_clock = clock; // @[:@41052.4]
  assign x496_sum_1_reset = reset; // @[:@41053.4]
  assign x496_sum_1_io_a = x495_x11_1_io_result; // @[Math.scala 151:17:@41054.4]
  assign x496_sum_1_io_b = RetimeWrapper_116_io_out; // @[Math.scala 152:17:@41055.4]
  assign x496_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@41056.4]
  assign RetimeWrapper_117_clock = clock; // @[:@41071.4]
  assign RetimeWrapper_117_reset = reset; // @[:@41072.4]
  assign RetimeWrapper_117_io_flow = io_in_x317_TREADY; // @[package.scala 95:18:@41074.4]
  assign RetimeWrapper_117_io_in = _GEN_5 << 1; // @[package.scala 94:16:@41073.4]
  assign RetimeWrapper_118_clock = clock; // @[:@41083.4]
  assign RetimeWrapper_118_reset = reset; // @[:@41084.4]
  assign RetimeWrapper_118_io_flow = io_in_x317_TREADY; // @[package.scala 95:18:@41086.4]
  assign RetimeWrapper_118_io_in = _GEN_6 << 1; // @[package.scala 94:16:@41085.4]
  assign RetimeWrapper_119_clock = clock; // @[:@41095.4]
  assign RetimeWrapper_119_reset = reset; // @[:@41096.4]
  assign RetimeWrapper_119_io_flow = io_in_x317_TREADY; // @[package.scala 95:18:@41098.4]
  assign RetimeWrapper_119_io_in = _GEN_7 << 2; // @[package.scala 94:16:@41097.4]
  assign RetimeWrapper_120_clock = clock; // @[:@41107.4]
  assign RetimeWrapper_120_reset = reset; // @[:@41108.4]
  assign RetimeWrapper_120_io_flow = io_in_x317_TREADY; // @[package.scala 95:18:@41110.4]
  assign RetimeWrapper_120_io_in = _GEN_8 << 1; // @[package.scala 94:16:@41109.4]
  assign RetimeWrapper_121_clock = clock; // @[:@41119.4]
  assign RetimeWrapper_121_reset = reset; // @[:@41120.4]
  assign RetimeWrapper_121_io_flow = io_in_x317_TREADY; // @[package.scala 95:18:@41122.4]
  assign RetimeWrapper_121_io_in = _GEN_9 << 1; // @[package.scala 94:16:@41121.4]
  assign RetimeWrapper_122_clock = clock; // @[:@41129.4]
  assign RetimeWrapper_122_reset = reset; // @[:@41130.4]
  assign RetimeWrapper_122_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41132.4]
  assign RetimeWrapper_122_io_in = _T_1522[7:0]; // @[package.scala 94:16:@41131.4]
  assign RetimeWrapper_123_clock = clock; // @[:@41138.4]
  assign RetimeWrapper_123_reset = reset; // @[:@41139.4]
  assign RetimeWrapper_123_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41141.4]
  assign RetimeWrapper_123_io_in = x329_lb_0_io_rPort_3_output_0; // @[package.scala 94:16:@41140.4]
  assign x503_x11_1_io_a = RetimeWrapper_123_io_out; // @[Math.scala 151:17:@41149.4]
  assign x503_x11_1_io_b = RetimeWrapper_122_io_out; // @[Math.scala 152:17:@41150.4]
  assign RetimeWrapper_124_clock = clock; // @[:@41157.4]
  assign RetimeWrapper_124_reset = reset; // @[:@41158.4]
  assign RetimeWrapper_124_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41160.4]
  assign RetimeWrapper_124_io_in = x329_lb_0_io_rPort_4_output_0; // @[package.scala 94:16:@41159.4]
  assign RetimeWrapper_125_clock = clock; // @[:@41166.4]
  assign RetimeWrapper_125_reset = reset; // @[:@41167.4]
  assign RetimeWrapper_125_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41169.4]
  assign RetimeWrapper_125_io_in = _T_1528[7:0]; // @[package.scala 94:16:@41168.4]
  assign x504_x12_1_io_a = RetimeWrapper_124_io_out; // @[Math.scala 151:17:@41177.4]
  assign x504_x12_1_io_b = RetimeWrapper_125_io_out; // @[Math.scala 152:17:@41178.4]
  assign x505_x11_1_io_a = _T_1534[7:0]; // @[Math.scala 151:17:@41187.4]
  assign x505_x11_1_io_b = _T_1540[7:0]; // @[Math.scala 152:17:@41188.4]
  assign RetimeWrapper_126_clock = clock; // @[:@41195.4]
  assign RetimeWrapper_126_reset = reset; // @[:@41196.4]
  assign RetimeWrapper_126_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41198.4]
  assign RetimeWrapper_126_io_in = x329_lb_0_io_rPort_8_output_0; // @[package.scala 94:16:@41197.4]
  assign x506_x12_1_io_a = RetimeWrapper_126_io_out; // @[Math.scala 151:17:@41206.4]
  assign x506_x12_1_io_b = _T_1546[7:0]; // @[Math.scala 152:17:@41207.4]
  assign RetimeWrapper_127_clock = clock; // @[:@41214.4]
  assign RetimeWrapper_127_reset = reset; // @[:@41215.4]
  assign RetimeWrapper_127_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41217.4]
  assign RetimeWrapper_127_io_in = x503_x11_1_io_result; // @[package.scala 94:16:@41216.4]
  assign RetimeWrapper_128_clock = clock; // @[:@41223.4]
  assign RetimeWrapper_128_reset = reset; // @[:@41224.4]
  assign RetimeWrapper_128_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41226.4]
  assign RetimeWrapper_128_io_in = x504_x12_1_io_result; // @[package.scala 94:16:@41225.4]
  assign x507_x11_1_io_a = RetimeWrapper_127_io_out; // @[Math.scala 151:17:@41234.4]
  assign x507_x11_1_io_b = RetimeWrapper_128_io_out; // @[Math.scala 152:17:@41235.4]
  assign x508_x12_1_io_a = x505_x11_1_io_result; // @[Math.scala 151:17:@41244.4]
  assign x508_x12_1_io_b = x506_x12_1_io_result; // @[Math.scala 152:17:@41245.4]
  assign RetimeWrapper_129_clock = clock; // @[:@41252.4]
  assign RetimeWrapper_129_reset = reset; // @[:@41253.4]
  assign RetimeWrapper_129_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41255.4]
  assign RetimeWrapper_129_io_in = x508_x12_1_io_result; // @[package.scala 94:16:@41254.4]
  assign x509_x11_1_io_a = x507_x11_1_io_result; // @[Math.scala 151:17:@41263.4]
  assign x509_x11_1_io_b = RetimeWrapper_129_io_out; // @[Math.scala 152:17:@41264.4]
  assign RetimeWrapper_130_clock = clock; // @[:@41271.4]
  assign RetimeWrapper_130_reset = reset; // @[:@41272.4]
  assign RetimeWrapper_130_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41274.4]
  assign RetimeWrapper_130_io_in = x329_lb_0_io_rPort_0_output_0; // @[package.scala 94:16:@41273.4]
  assign x510_sum_1_clock = clock; // @[:@41280.4]
  assign x510_sum_1_reset = reset; // @[:@41281.4]
  assign x510_sum_1_io_a = x509_x11_1_io_result; // @[Math.scala 151:17:@41282.4]
  assign x510_sum_1_io_b = RetimeWrapper_130_io_out; // @[Math.scala 152:17:@41283.4]
  assign x510_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@41284.4]
  assign RetimeWrapper_131_clock = clock; // @[:@41299.4]
  assign RetimeWrapper_131_reset = reset; // @[:@41300.4]
  assign RetimeWrapper_131_io_flow = io_in_x317_TREADY; // @[package.scala 95:18:@41302.4]
  assign RetimeWrapper_131_io_in = _GEN_10 << 1; // @[package.scala 94:16:@41301.4]
  assign RetimeWrapper_132_clock = clock; // @[:@41311.4]
  assign RetimeWrapper_132_reset = reset; // @[:@41312.4]
  assign RetimeWrapper_132_io_flow = io_in_x317_TREADY; // @[package.scala 95:18:@41314.4]
  assign RetimeWrapper_132_io_in = _GEN_11 << 2; // @[package.scala 94:16:@41313.4]
  assign RetimeWrapper_133_clock = clock; // @[:@41323.4]
  assign RetimeWrapper_133_reset = reset; // @[:@41324.4]
  assign RetimeWrapper_133_io_flow = io_in_x317_TREADY; // @[package.scala 95:18:@41326.4]
  assign RetimeWrapper_133_io_in = _GEN_12 << 1; // @[package.scala 94:16:@41325.4]
  assign RetimeWrapper_134_clock = clock; // @[:@41335.4]
  assign RetimeWrapper_134_reset = reset; // @[:@41336.4]
  assign RetimeWrapper_134_io_flow = io_in_x317_TREADY; // @[package.scala 95:18:@41338.4]
  assign RetimeWrapper_134_io_in = _GEN_13 << 1; // @[package.scala 94:16:@41337.4]
  assign RetimeWrapper_135_clock = clock; // @[:@41345.4]
  assign RetimeWrapper_135_reset = reset; // @[:@41346.4]
  assign RetimeWrapper_135_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41348.4]
  assign RetimeWrapper_135_io_in = _T_1613[7:0]; // @[package.scala 94:16:@41347.4]
  assign x516_x11_1_io_a = RetimeWrapper_110_io_out; // @[Math.scala 151:17:@41356.4]
  assign x516_x11_1_io_b = RetimeWrapper_135_io_out; // @[Math.scala 152:17:@41357.4]
  assign RetimeWrapper_136_clock = clock; // @[:@41364.4]
  assign RetimeWrapper_136_reset = reset; // @[:@41365.4]
  assign RetimeWrapper_136_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41367.4]
  assign RetimeWrapper_136_io_in = _T_1447[7:0]; // @[package.scala 94:16:@41366.4]
  assign RetimeWrapper_137_clock = clock; // @[:@41373.4]
  assign RetimeWrapper_137_reset = reset; // @[:@41374.4]
  assign RetimeWrapper_137_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41376.4]
  assign RetimeWrapper_137_io_in = x329_lb_0_io_rPort_16_output_0; // @[package.scala 94:16:@41375.4]
  assign x517_x12_1_io_a = RetimeWrapper_137_io_out; // @[Math.scala 151:17:@41384.4]
  assign x517_x12_1_io_b = RetimeWrapper_136_io_out; // @[Math.scala 152:17:@41385.4]
  assign x518_x11_1_io_a = _T_1619[7:0]; // @[Math.scala 151:17:@41394.4]
  assign x518_x11_1_io_b = _T_1625[7:0]; // @[Math.scala 152:17:@41395.4]
  assign RetimeWrapper_138_clock = clock; // @[:@41402.4]
  assign RetimeWrapper_138_reset = reset; // @[:@41403.4]
  assign RetimeWrapper_138_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41405.4]
  assign RetimeWrapper_138_io_in = x329_lb_0_io_rPort_5_output_0; // @[package.scala 94:16:@41404.4]
  assign x519_x12_1_io_a = RetimeWrapper_138_io_out; // @[Math.scala 151:17:@41413.4]
  assign x519_x12_1_io_b = _T_1631[7:0]; // @[Math.scala 152:17:@41414.4]
  assign RetimeWrapper_139_clock = clock; // @[:@41421.4]
  assign RetimeWrapper_139_reset = reset; // @[:@41422.4]
  assign RetimeWrapper_139_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41424.4]
  assign RetimeWrapper_139_io_in = x517_x12_1_io_result; // @[package.scala 94:16:@41423.4]
  assign RetimeWrapper_140_clock = clock; // @[:@41430.4]
  assign RetimeWrapper_140_reset = reset; // @[:@41431.4]
  assign RetimeWrapper_140_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41433.4]
  assign RetimeWrapper_140_io_in = x516_x11_1_io_result; // @[package.scala 94:16:@41432.4]
  assign x520_x11_1_io_a = RetimeWrapper_140_io_out; // @[Math.scala 151:17:@41441.4]
  assign x520_x11_1_io_b = RetimeWrapper_139_io_out; // @[Math.scala 152:17:@41442.4]
  assign x521_x12_1_io_a = x518_x11_1_io_result; // @[Math.scala 151:17:@41451.4]
  assign x521_x12_1_io_b = x519_x12_1_io_result; // @[Math.scala 152:17:@41452.4]
  assign RetimeWrapper_141_clock = clock; // @[:@41459.4]
  assign RetimeWrapper_141_reset = reset; // @[:@41460.4]
  assign RetimeWrapper_141_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41462.4]
  assign RetimeWrapper_141_io_in = x521_x12_1_io_result; // @[package.scala 94:16:@41461.4]
  assign x522_x11_1_io_a = x520_x11_1_io_result; // @[Math.scala 151:17:@41470.4]
  assign x522_x11_1_io_b = RetimeWrapper_141_io_out; // @[Math.scala 152:17:@41471.4]
  assign RetimeWrapper_142_clock = clock; // @[:@41478.4]
  assign RetimeWrapper_142_reset = reset; // @[:@41479.4]
  assign RetimeWrapper_142_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41481.4]
  assign RetimeWrapper_142_io_in = x329_lb_0_io_rPort_7_output_0; // @[package.scala 94:16:@41480.4]
  assign x523_sum_1_clock = clock; // @[:@41487.4]
  assign x523_sum_1_reset = reset; // @[:@41488.4]
  assign x523_sum_1_io_a = x522_x11_1_io_result; // @[Math.scala 151:17:@41489.4]
  assign x523_sum_1_io_b = RetimeWrapper_142_io_out; // @[Math.scala 152:17:@41490.4]
  assign x523_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@41491.4]
  assign RetimeWrapper_143_clock = clock; // @[:@41508.4]
  assign RetimeWrapper_143_reset = reset; // @[:@41509.4]
  assign RetimeWrapper_143_io_flow = io_in_x317_TREADY; // @[package.scala 95:18:@41511.4]
  assign RetimeWrapper_143_io_in = _GEN_14 << 1; // @[package.scala 94:16:@41510.4]
  assign RetimeWrapper_144_clock = clock; // @[:@41520.4]
  assign RetimeWrapper_144_reset = reset; // @[:@41521.4]
  assign RetimeWrapper_144_io_flow = io_in_x317_TREADY; // @[package.scala 95:18:@41523.4]
  assign RetimeWrapper_144_io_in = _GEN_15 << 2; // @[package.scala 94:16:@41522.4]
  assign RetimeWrapper_145_clock = clock; // @[:@41532.4]
  assign RetimeWrapper_145_reset = reset; // @[:@41533.4]
  assign RetimeWrapper_145_io_flow = io_in_x317_TREADY; // @[package.scala 95:18:@41535.4]
  assign RetimeWrapper_145_io_in = _GEN_16 << 1; // @[package.scala 94:16:@41534.4]
  assign RetimeWrapper_146_clock = clock; // @[:@41544.4]
  assign RetimeWrapper_146_reset = reset; // @[:@41545.4]
  assign RetimeWrapper_146_io_flow = io_in_x317_TREADY; // @[package.scala 95:18:@41547.4]
  assign RetimeWrapper_146_io_in = _GEN_17 << 1; // @[package.scala 94:16:@41546.4]
  assign RetimeWrapper_147_clock = clock; // @[:@41554.4]
  assign RetimeWrapper_147_reset = reset; // @[:@41555.4]
  assign RetimeWrapper_147_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41557.4]
  assign RetimeWrapper_147_io_in = _T_1697[7:0]; // @[package.scala 94:16:@41556.4]
  assign x529_x11_1_io_a = RetimeWrapper_124_io_out; // @[Math.scala 151:17:@41565.4]
  assign x529_x11_1_io_b = RetimeWrapper_147_io_out; // @[Math.scala 152:17:@41566.4]
  assign RetimeWrapper_148_clock = clock; // @[:@41573.4]
  assign RetimeWrapper_148_reset = reset; // @[:@41574.4]
  assign RetimeWrapper_148_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41576.4]
  assign RetimeWrapper_148_io_in = _T_1540[7:0]; // @[package.scala 94:16:@41575.4]
  assign RetimeWrapper_149_clock = clock; // @[:@41582.4]
  assign RetimeWrapper_149_reset = reset; // @[:@41583.4]
  assign RetimeWrapper_149_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41585.4]
  assign RetimeWrapper_149_io_in = x329_lb_0_io_rPort_17_output_0; // @[package.scala 94:16:@41584.4]
  assign x530_x12_1_io_a = RetimeWrapper_149_io_out; // @[Math.scala 151:17:@41593.4]
  assign x530_x12_1_io_b = RetimeWrapper_148_io_out; // @[Math.scala 152:17:@41594.4]
  assign x531_x11_1_io_a = _T_1703[7:0]; // @[Math.scala 151:17:@41603.4]
  assign x531_x11_1_io_b = _T_1709[7:0]; // @[Math.scala 152:17:@41604.4]
  assign RetimeWrapper_150_clock = clock; // @[:@41611.4]
  assign RetimeWrapper_150_reset = reset; // @[:@41612.4]
  assign RetimeWrapper_150_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41614.4]
  assign RetimeWrapper_150_io_in = x329_lb_0_io_rPort_0_output_0; // @[package.scala 94:16:@41613.4]
  assign x532_x12_1_io_a = RetimeWrapper_150_io_out; // @[Math.scala 151:17:@41622.4]
  assign x532_x12_1_io_b = _T_1715[7:0]; // @[Math.scala 152:17:@41623.4]
  assign RetimeWrapper_151_clock = clock; // @[:@41630.4]
  assign RetimeWrapper_151_reset = reset; // @[:@41631.4]
  assign RetimeWrapper_151_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41633.4]
  assign RetimeWrapper_151_io_in = x530_x12_1_io_result; // @[package.scala 94:16:@41632.4]
  assign RetimeWrapper_152_clock = clock; // @[:@41639.4]
  assign RetimeWrapper_152_reset = reset; // @[:@41640.4]
  assign RetimeWrapper_152_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41642.4]
  assign RetimeWrapper_152_io_in = x529_x11_1_io_result; // @[package.scala 94:16:@41641.4]
  assign x533_x11_1_io_a = RetimeWrapper_152_io_out; // @[Math.scala 151:17:@41650.4]
  assign x533_x11_1_io_b = RetimeWrapper_151_io_out; // @[Math.scala 152:17:@41651.4]
  assign x534_x12_1_io_a = x531_x11_1_io_result; // @[Math.scala 151:17:@41660.4]
  assign x534_x12_1_io_b = x532_x12_1_io_result; // @[Math.scala 152:17:@41661.4]
  assign RetimeWrapper_153_clock = clock; // @[:@41668.4]
  assign RetimeWrapper_153_reset = reset; // @[:@41669.4]
  assign RetimeWrapper_153_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41671.4]
  assign RetimeWrapper_153_io_in = x534_x12_1_io_result; // @[package.scala 94:16:@41670.4]
  assign x535_x11_1_io_a = x533_x11_1_io_result; // @[Math.scala 151:17:@41679.4]
  assign x535_x11_1_io_b = RetimeWrapper_153_io_out; // @[Math.scala 152:17:@41680.4]
  assign RetimeWrapper_154_clock = clock; // @[:@41687.4]
  assign RetimeWrapper_154_reset = reset; // @[:@41688.4]
  assign RetimeWrapper_154_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41690.4]
  assign RetimeWrapper_154_io_in = x329_lb_0_io_rPort_15_output_0; // @[package.scala 94:16:@41689.4]
  assign x536_sum_1_clock = clock; // @[:@41696.4]
  assign x536_sum_1_reset = reset; // @[:@41697.4]
  assign x536_sum_1_io_a = x535_x11_1_io_result; // @[Math.scala 151:17:@41698.4]
  assign x536_sum_1_io_b = RetimeWrapper_154_io_out; // @[Math.scala 152:17:@41699.4]
  assign x536_sum_1_io_flow = io_in_x317_TREADY; // @[Math.scala 153:20:@41700.4]
  assign RetimeWrapper_155_clock = clock; // @[:@41713.4]
  assign RetimeWrapper_155_reset = reset; // @[:@41714.4]
  assign RetimeWrapper_155_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41716.4]
  assign RetimeWrapper_155_io_in = {4'h0,_T_1688}; // @[package.scala 94:16:@41715.4]
  assign RetimeWrapper_156_clock = clock; // @[:@41722.4]
  assign RetimeWrapper_156_reset = reset; // @[:@41723.4]
  assign RetimeWrapper_156_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41725.4]
  assign RetimeWrapper_156_io_in = {4'h0,_T_1515}; // @[package.scala 94:16:@41724.4]
  assign RetimeWrapper_157_clock = clock; // @[:@41731.4]
  assign RetimeWrapper_157_reset = reset; // @[:@41732.4]
  assign RetimeWrapper_157_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41734.4]
  assign RetimeWrapper_157_io_in = {4'h0,_T_1772}; // @[package.scala 94:16:@41733.4]
  assign RetimeWrapper_158_clock = clock; // @[:@41740.4]
  assign RetimeWrapper_158_reset = reset; // @[:@41741.4]
  assign RetimeWrapper_158_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41743.4]
  assign RetimeWrapper_158_io_in = {4'h0,_T_1606}; // @[package.scala 94:16:@41742.4]
  assign RetimeWrapper_159_clock = clock; // @[:@41759.4]
  assign RetimeWrapper_159_reset = reset; // @[:@41760.4]
  assign RetimeWrapper_159_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41762.4]
  assign RetimeWrapper_159_io_in = {_T_1798,_T_1797}; // @[package.scala 94:16:@41761.4]
  assign RetimeWrapper_160_clock = clock; // @[:@41768.4]
  assign RetimeWrapper_160_reset = reset; // @[:@41769.4]
  assign RetimeWrapper_160_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41771.4]
  assign RetimeWrapper_160_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@41770.4]
  assign RetimeWrapper_161_clock = clock; // @[:@41777.4]
  assign RetimeWrapper_161_reset = reset; // @[:@41778.4]
  assign RetimeWrapper_161_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41780.4]
  assign RetimeWrapper_161_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@41779.4]
  assign RetimeWrapper_162_clock = clock; // @[:@41786.4]
  assign RetimeWrapper_162_reset = reset; // @[:@41787.4]
  assign RetimeWrapper_162_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41789.4]
  assign RetimeWrapper_162_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@41788.4]
endmodule
module x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1( // @[:@41807.2]
  input          clock, // @[:@41808.4]
  input          reset, // @[:@41809.4]
  input          io_in_x316_TVALID, // @[:@41810.4]
  output         io_in_x316_TREADY, // @[:@41810.4]
  input  [255:0] io_in_x316_TDATA, // @[:@41810.4]
  input  [7:0]   io_in_x316_TID, // @[:@41810.4]
  input  [7:0]   io_in_x316_TDEST, // @[:@41810.4]
  output         io_in_x317_TVALID, // @[:@41810.4]
  input          io_in_x317_TREADY, // @[:@41810.4]
  output [255:0] io_in_x317_TDATA, // @[:@41810.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@41810.4]
  input          io_sigsIn_smChildAcks_0, // @[:@41810.4]
  output         io_sigsOut_smDoneIn_0, // @[:@41810.4]
  output         io_sigsOut_smCtrCopyDone_0, // @[:@41810.4]
  input          io_rr // @[:@41810.4]
);
  wire  x324_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@41820.4]
  wire  x324_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@41820.4]
  wire  x324_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@41820.4]
  wire  x324_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@41820.4]
  wire [31:0] x324_ctrchain_io_output_counts_1; // @[SpatialBlocks.scala 37:22:@41820.4]
  wire [31:0] x324_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@41820.4]
  wire  x324_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@41820.4]
  wire  x324_ctrchain_io_output_oobs_1; // @[SpatialBlocks.scala 37:22:@41820.4]
  wire  x324_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@41820.4]
  wire  x542_inr_Foreach_SAMPLER_BOX_sm_clock; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 32:18:@41880.4]
  wire  x542_inr_Foreach_SAMPLER_BOX_sm_reset; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 32:18:@41880.4]
  wire  x542_inr_Foreach_SAMPLER_BOX_sm_io_enable; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 32:18:@41880.4]
  wire  x542_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 32:18:@41880.4]
  wire  x542_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 32:18:@41880.4]
  wire  x542_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 32:18:@41880.4]
  wire  x542_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 32:18:@41880.4]
  wire  x542_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 32:18:@41880.4]
  wire  x542_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 32:18:@41880.4]
  wire  x542_inr_Foreach_SAMPLER_BOX_sm_io_parentAck; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 32:18:@41880.4]
  wire  x542_inr_Foreach_SAMPLER_BOX_sm_io_backpressure; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 32:18:@41880.4]
  wire  x542_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 32:18:@41880.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@41908.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@41908.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@41908.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@41908.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@41908.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@41950.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@41950.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@41950.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@41950.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@41950.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@41958.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@41958.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@41958.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@41958.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@41958.4]
  wire  x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_clock; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 842:24:@41993.4]
  wire  x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_reset; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 842:24:@41993.4]
  wire  x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x316_TREADY; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 842:24:@41993.4]
  wire [255:0] x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x316_TDATA; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 842:24:@41993.4]
  wire [7:0] x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x316_TID; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 842:24:@41993.4]
  wire [7:0] x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x316_TDEST; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 842:24:@41993.4]
  wire  x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x317_TVALID; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 842:24:@41993.4]
  wire  x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x317_TREADY; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 842:24:@41993.4]
  wire [255:0] x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x317_TDATA; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 842:24:@41993.4]
  wire  x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 842:24:@41993.4]
  wire  x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 842:24:@41993.4]
  wire  x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 842:24:@41993.4]
  wire [31:0] x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 842:24:@41993.4]
  wire [31:0] x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 842:24:@41993.4]
  wire  x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 842:24:@41993.4]
  wire  x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 842:24:@41993.4]
  wire  x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_rr; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 842:24:@41993.4]
  wire  _T_239; // @[package.scala 96:25:@41913.4 package.scala 96:25:@41914.4]
  wire  x542_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[sm_x543_outr_UnitPipe.scala 68:66:@41919.4]
  wire  _T_252; // @[package.scala 96:25:@41955.4 package.scala 96:25:@41956.4]
  wire  _T_258; // @[package.scala 96:25:@41963.4 package.scala 96:25:@41964.4]
  wire  _T_261; // @[SpatialBlocks.scala 138:93:@41966.4]
  wire  x542_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn; // @[SpatialBlocks.scala 138:90:@41967.4]
  wire  _T_263; // @[SpatialBlocks.scala 157:36:@41975.4]
  wire  _T_264; // @[SpatialBlocks.scala 157:78:@41976.4]
  wire  _T_271; // @[SpatialBlocks.scala 159:58:@41988.4]
  x324_ctrchain x324_ctrchain ( // @[SpatialBlocks.scala 37:22:@41820.4]
    .clock(x324_ctrchain_clock),
    .reset(x324_ctrchain_reset),
    .io_input_reset(x324_ctrchain_io_input_reset),
    .io_input_enable(x324_ctrchain_io_input_enable),
    .io_output_counts_1(x324_ctrchain_io_output_counts_1),
    .io_output_counts_0(x324_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x324_ctrchain_io_output_oobs_0),
    .io_output_oobs_1(x324_ctrchain_io_output_oobs_1),
    .io_output_done(x324_ctrchain_io_output_done)
  );
  x542_inr_Foreach_SAMPLER_BOX_sm x542_inr_Foreach_SAMPLER_BOX_sm ( // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 32:18:@41880.4]
    .clock(x542_inr_Foreach_SAMPLER_BOX_sm_clock),
    .reset(x542_inr_Foreach_SAMPLER_BOX_sm_reset),
    .io_enable(x542_inr_Foreach_SAMPLER_BOX_sm_io_enable),
    .io_done(x542_inr_Foreach_SAMPLER_BOX_sm_io_done),
    .io_doneLatch(x542_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch),
    .io_ctrDone(x542_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone),
    .io_datapathEn(x542_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn),
    .io_ctrInc(x542_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc),
    .io_ctrRst(x542_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst),
    .io_parentAck(x542_inr_Foreach_SAMPLER_BOX_sm_io_parentAck),
    .io_backpressure(x542_inr_Foreach_SAMPLER_BOX_sm_io_backpressure),
    .io_break(x542_inr_Foreach_SAMPLER_BOX_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@41908.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@41950.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@41958.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1 x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1 ( // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 842:24:@41993.4]
    .clock(x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_clock),
    .reset(x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_reset),
    .io_in_x316_TREADY(x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x316_TREADY),
    .io_in_x316_TDATA(x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x316_TDATA),
    .io_in_x316_TID(x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x316_TID),
    .io_in_x316_TDEST(x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x316_TDEST),
    .io_in_x317_TVALID(x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x317_TVALID),
    .io_in_x317_TREADY(x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x317_TREADY),
    .io_in_x317_TDATA(x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x317_TDATA),
    .io_sigsIn_backpressure(x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_1(x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsIn_cchainOutputs_0_oobs_1(x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1),
    .io_rr(x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_rr)
  );
  assign _T_239 = RetimeWrapper_io_out; // @[package.scala 96:25:@41913.4 package.scala 96:25:@41914.4]
  assign x542_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure = io_in_x316_TVALID | x542_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x543_outr_UnitPipe.scala 68:66:@41919.4]
  assign _T_252 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@41955.4 package.scala 96:25:@41956.4]
  assign _T_258 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@41963.4 package.scala 96:25:@41964.4]
  assign _T_261 = ~ _T_258; // @[SpatialBlocks.scala 138:93:@41966.4]
  assign x542_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn = _T_252 & _T_261; // @[SpatialBlocks.scala 138:90:@41967.4]
  assign _T_263 = x542_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@41975.4]
  assign _T_264 = ~ x542_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@41976.4]
  assign _T_271 = x542_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[SpatialBlocks.scala 159:58:@41988.4]
  assign io_in_x316_TREADY = x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x316_TREADY; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 48:23:@42051.4]
  assign io_in_x317_TVALID = x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x317_TVALID; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 49:23:@42061.4]
  assign io_in_x317_TDATA = x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x317_TDATA; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 49:23:@42059.4]
  assign io_sigsOut_smDoneIn_0 = x542_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[SpatialBlocks.scala 156:53:@41973.4]
  assign io_sigsOut_smCtrCopyDone_0 = x542_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[SpatialBlocks.scala 168:125:@41992.4]
  assign x324_ctrchain_clock = clock; // @[:@41821.4]
  assign x324_ctrchain_reset = reset; // @[:@41822.4]
  assign x324_ctrchain_io_input_reset = x542_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@41991.4]
  assign x324_ctrchain_io_input_enable = _T_271 & x542_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 132:75:@41943.4 SpatialBlocks.scala 159:42:@41990.4]
  assign x542_inr_Foreach_SAMPLER_BOX_sm_clock = clock; // @[:@41881.4]
  assign x542_inr_Foreach_SAMPLER_BOX_sm_reset = reset; // @[:@41882.4]
  assign x542_inr_Foreach_SAMPLER_BOX_sm_io_enable = x542_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn & x542_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 140:18:@41970.4]
  assign x542_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone = io_rr ? _T_239 : 1'h0; // @[sm_x543_outr_UnitPipe.scala 66:50:@41916.4]
  assign x542_inr_Foreach_SAMPLER_BOX_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@41972.4]
  assign x542_inr_Foreach_SAMPLER_BOX_sm_io_backpressure = io_in_x317_TREADY | x542_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@41944.4]
  assign x542_inr_Foreach_SAMPLER_BOX_sm_io_break = 1'h0; // @[sm_x543_outr_UnitPipe.scala 70:48:@41922.4]
  assign RetimeWrapper_clock = clock; // @[:@41909.4]
  assign RetimeWrapper_reset = reset; // @[:@41910.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@41912.4]
  assign RetimeWrapper_io_in = x324_ctrchain_io_output_done; // @[package.scala 94:16:@41911.4]
  assign RetimeWrapper_1_clock = clock; // @[:@41951.4]
  assign RetimeWrapper_1_reset = reset; // @[:@41952.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@41954.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@41953.4]
  assign RetimeWrapper_2_clock = clock; // @[:@41959.4]
  assign RetimeWrapper_2_reset = reset; // @[:@41960.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@41962.4]
  assign RetimeWrapper_2_io_in = x542_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[package.scala 94:16:@41961.4]
  assign x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_clock = clock; // @[:@41994.4]
  assign x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_reset = reset; // @[:@41995.4]
  assign x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x316_TDATA = io_in_x316_TDATA; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 48:23:@42050.4]
  assign x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x316_TID = io_in_x316_TID; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 48:23:@42046.4]
  assign x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x316_TDEST = io_in_x316_TDEST; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 48:23:@42045.4]
  assign x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x317_TREADY = io_in_x317_TREADY; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 49:23:@42060.4]
  assign x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure = io_in_x317_TREADY | x542_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 847:22:@42078.4]
  assign x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn = _T_263 & _T_264; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 847:22:@42076.4]
  assign x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break = x542_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 847:22:@42074.4]
  assign x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1 = x324_ctrchain_io_output_counts_1; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 847:22:@42069.4]
  assign x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = x324_ctrchain_io_output_counts_0; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 847:22:@42068.4]
  assign x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x324_ctrchain_io_output_oobs_0; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 847:22:@42066.4]
  assign x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1 = x324_ctrchain_io_output_oobs_1; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 847:22:@42067.4]
  assign x542_inr_Foreach_SAMPLER_BOX_kernelx542_inr_Foreach_SAMPLER_BOX_concrete1_io_rr = io_rr; // @[sm_x542_inr_Foreach_SAMPLER_BOX.scala 846:18:@42062.4]
endmodule
module RootController_kernelRootController_concrete1( // @[:@42092.2]
  input          clock, // @[:@42093.4]
  input          reset, // @[:@42094.4]
  input          io_in_x316_TVALID, // @[:@42095.4]
  output         io_in_x316_TREADY, // @[:@42095.4]
  input  [255:0] io_in_x316_TDATA, // @[:@42095.4]
  input  [7:0]   io_in_x316_TID, // @[:@42095.4]
  input  [7:0]   io_in_x316_TDEST, // @[:@42095.4]
  output         io_in_x317_TVALID, // @[:@42095.4]
  input          io_in_x317_TREADY, // @[:@42095.4]
  output [255:0] io_in_x317_TDATA, // @[:@42095.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@42095.4]
  input          io_sigsIn_smChildAcks_0, // @[:@42095.4]
  output         io_sigsOut_smDoneIn_0, // @[:@42095.4]
  input          io_rr // @[:@42095.4]
);
  wire  x543_outr_UnitPipe_sm_clock; // @[sm_x543_outr_UnitPipe.scala 32:18:@42237.4]
  wire  x543_outr_UnitPipe_sm_reset; // @[sm_x543_outr_UnitPipe.scala 32:18:@42237.4]
  wire  x543_outr_UnitPipe_sm_io_enable; // @[sm_x543_outr_UnitPipe.scala 32:18:@42237.4]
  wire  x543_outr_UnitPipe_sm_io_done; // @[sm_x543_outr_UnitPipe.scala 32:18:@42237.4]
  wire  x543_outr_UnitPipe_sm_io_parentAck; // @[sm_x543_outr_UnitPipe.scala 32:18:@42237.4]
  wire  x543_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x543_outr_UnitPipe.scala 32:18:@42237.4]
  wire  x543_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x543_outr_UnitPipe.scala 32:18:@42237.4]
  wire  x543_outr_UnitPipe_sm_io_childAck_0; // @[sm_x543_outr_UnitPipe.scala 32:18:@42237.4]
  wire  x543_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x543_outr_UnitPipe.scala 32:18:@42237.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@42289.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@42289.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@42289.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@42289.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@42289.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@42297.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@42297.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@42297.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@42297.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@42297.4]
  wire  x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_clock; // @[sm_x543_outr_UnitPipe.scala 75:24:@42327.4]
  wire  x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_reset; // @[sm_x543_outr_UnitPipe.scala 75:24:@42327.4]
  wire  x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_io_in_x316_TVALID; // @[sm_x543_outr_UnitPipe.scala 75:24:@42327.4]
  wire  x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_io_in_x316_TREADY; // @[sm_x543_outr_UnitPipe.scala 75:24:@42327.4]
  wire [255:0] x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_io_in_x316_TDATA; // @[sm_x543_outr_UnitPipe.scala 75:24:@42327.4]
  wire [7:0] x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_io_in_x316_TID; // @[sm_x543_outr_UnitPipe.scala 75:24:@42327.4]
  wire [7:0] x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_io_in_x316_TDEST; // @[sm_x543_outr_UnitPipe.scala 75:24:@42327.4]
  wire  x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_io_in_x317_TVALID; // @[sm_x543_outr_UnitPipe.scala 75:24:@42327.4]
  wire  x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_io_in_x317_TREADY; // @[sm_x543_outr_UnitPipe.scala 75:24:@42327.4]
  wire [255:0] x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_io_in_x317_TDATA; // @[sm_x543_outr_UnitPipe.scala 75:24:@42327.4]
  wire  x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x543_outr_UnitPipe.scala 75:24:@42327.4]
  wire  x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x543_outr_UnitPipe.scala 75:24:@42327.4]
  wire  x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x543_outr_UnitPipe.scala 75:24:@42327.4]
  wire  x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x543_outr_UnitPipe.scala 75:24:@42327.4]
  wire  x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_io_rr; // @[sm_x543_outr_UnitPipe.scala 75:24:@42327.4]
  wire  _T_246; // @[package.scala 96:25:@42294.4 package.scala 96:25:@42295.4]
  wire  _T_252; // @[package.scala 96:25:@42302.4 package.scala 96:25:@42303.4]
  wire  _T_255; // @[SpatialBlocks.scala 138:93:@42305.4]
  x543_outr_UnitPipe_sm x543_outr_UnitPipe_sm ( // @[sm_x543_outr_UnitPipe.scala 32:18:@42237.4]
    .clock(x543_outr_UnitPipe_sm_clock),
    .reset(x543_outr_UnitPipe_sm_reset),
    .io_enable(x543_outr_UnitPipe_sm_io_enable),
    .io_done(x543_outr_UnitPipe_sm_io_done),
    .io_parentAck(x543_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x543_outr_UnitPipe_sm_io_doneIn_0),
    .io_enableOut_0(x543_outr_UnitPipe_sm_io_enableOut_0),
    .io_childAck_0(x543_outr_UnitPipe_sm_io_childAck_0),
    .io_ctrCopyDone_0(x543_outr_UnitPipe_sm_io_ctrCopyDone_0)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@42289.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@42297.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1 x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1 ( // @[sm_x543_outr_UnitPipe.scala 75:24:@42327.4]
    .clock(x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_clock),
    .reset(x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_reset),
    .io_in_x316_TVALID(x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_io_in_x316_TVALID),
    .io_in_x316_TREADY(x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_io_in_x316_TREADY),
    .io_in_x316_TDATA(x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_io_in_x316_TDATA),
    .io_in_x316_TID(x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_io_in_x316_TID),
    .io_in_x316_TDEST(x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_io_in_x316_TDEST),
    .io_in_x317_TVALID(x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_io_in_x317_TVALID),
    .io_in_x317_TREADY(x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_io_in_x317_TREADY),
    .io_in_x317_TDATA(x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_io_in_x317_TDATA),
    .io_sigsIn_smEnableOuts_0(x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smCtrCopyDone_0(x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_rr(x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_246 = RetimeWrapper_io_out; // @[package.scala 96:25:@42294.4 package.scala 96:25:@42295.4]
  assign _T_252 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@42302.4 package.scala 96:25:@42303.4]
  assign _T_255 = ~ _T_252; // @[SpatialBlocks.scala 138:93:@42305.4]
  assign io_in_x316_TREADY = x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_io_in_x316_TREADY; // @[sm_x543_outr_UnitPipe.scala 48:23:@42383.4]
  assign io_in_x317_TVALID = x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_io_in_x317_TVALID; // @[sm_x543_outr_UnitPipe.scala 49:23:@42393.4]
  assign io_in_x317_TDATA = x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_io_in_x317_TDATA; // @[sm_x543_outr_UnitPipe.scala 49:23:@42391.4]
  assign io_sigsOut_smDoneIn_0 = x543_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@42312.4]
  assign x543_outr_UnitPipe_sm_clock = clock; // @[:@42238.4]
  assign x543_outr_UnitPipe_sm_reset = reset; // @[:@42239.4]
  assign x543_outr_UnitPipe_sm_io_enable = _T_246 & _T_255; // @[SpatialBlocks.scala 140:18:@42309.4]
  assign x543_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@42311.4]
  assign x543_outr_UnitPipe_sm_io_doneIn_0 = x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@42281.4]
  assign x543_outr_UnitPipe_sm_io_ctrCopyDone_0 = x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 161:90:@42326.4]
  assign RetimeWrapper_clock = clock; // @[:@42290.4]
  assign RetimeWrapper_reset = reset; // @[:@42291.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@42293.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@42292.4]
  assign RetimeWrapper_1_clock = clock; // @[:@42298.4]
  assign RetimeWrapper_1_reset = reset; // @[:@42299.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@42301.4]
  assign RetimeWrapper_1_io_in = x543_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@42300.4]
  assign x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_clock = clock; // @[:@42328.4]
  assign x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_reset = reset; // @[:@42329.4]
  assign x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_io_in_x316_TVALID = io_in_x316_TVALID; // @[sm_x543_outr_UnitPipe.scala 48:23:@42384.4]
  assign x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_io_in_x316_TDATA = io_in_x316_TDATA; // @[sm_x543_outr_UnitPipe.scala 48:23:@42382.4]
  assign x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_io_in_x316_TID = io_in_x316_TID; // @[sm_x543_outr_UnitPipe.scala 48:23:@42378.4]
  assign x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_io_in_x316_TDEST = io_in_x316_TDEST; // @[sm_x543_outr_UnitPipe.scala 48:23:@42377.4]
  assign x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_io_in_x317_TREADY = io_in_x317_TREADY; // @[sm_x543_outr_UnitPipe.scala 49:23:@42392.4]
  assign x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x543_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x543_outr_UnitPipe.scala 80:22:@42402.4]
  assign x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x543_outr_UnitPipe_sm_io_childAck_0; // @[sm_x543_outr_UnitPipe.scala 80:22:@42400.4]
  assign x543_outr_UnitPipe_kernelx543_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x543_outr_UnitPipe.scala 79:18:@42394.4]
endmodule
module AccelUnit( // @[:@42422.2]
  input          clock, // @[:@42423.4]
  input          reset, // @[:@42424.4]
  input          io_enable, // @[:@42425.4]
  output         io_done, // @[:@42425.4]
  input          io_reset, // @[:@42425.4]
  input          io_memStreams_loads_0_cmd_ready, // @[:@42425.4]
  output         io_memStreams_loads_0_cmd_valid, // @[:@42425.4]
  output [63:0]  io_memStreams_loads_0_cmd_bits_addr, // @[:@42425.4]
  output [31:0]  io_memStreams_loads_0_cmd_bits_size, // @[:@42425.4]
  output         io_memStreams_loads_0_data_ready, // @[:@42425.4]
  input          io_memStreams_loads_0_data_valid, // @[:@42425.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_0, // @[:@42425.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_1, // @[:@42425.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_2, // @[:@42425.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_3, // @[:@42425.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_4, // @[:@42425.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_5, // @[:@42425.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_6, // @[:@42425.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_7, // @[:@42425.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_8, // @[:@42425.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_9, // @[:@42425.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_10, // @[:@42425.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_11, // @[:@42425.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_12, // @[:@42425.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_13, // @[:@42425.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_14, // @[:@42425.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_15, // @[:@42425.4]
  input          io_memStreams_stores_0_cmd_ready, // @[:@42425.4]
  output         io_memStreams_stores_0_cmd_valid, // @[:@42425.4]
  output [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@42425.4]
  output [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@42425.4]
  input          io_memStreams_stores_0_data_ready, // @[:@42425.4]
  output         io_memStreams_stores_0_data_valid, // @[:@42425.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_0, // @[:@42425.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_1, // @[:@42425.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_2, // @[:@42425.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_3, // @[:@42425.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_4, // @[:@42425.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_5, // @[:@42425.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_6, // @[:@42425.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_7, // @[:@42425.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_8, // @[:@42425.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_9, // @[:@42425.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_10, // @[:@42425.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_11, // @[:@42425.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_12, // @[:@42425.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_13, // @[:@42425.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_14, // @[:@42425.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_15, // @[:@42425.4]
  output [15:0]  io_memStreams_stores_0_data_bits_wstrb, // @[:@42425.4]
  output         io_memStreams_stores_0_wresp_ready, // @[:@42425.4]
  input          io_memStreams_stores_0_wresp_valid, // @[:@42425.4]
  input          io_memStreams_stores_0_wresp_bits, // @[:@42425.4]
  input          io_memStreams_gathers_0_cmd_ready, // @[:@42425.4]
  output         io_memStreams_gathers_0_cmd_valid, // @[:@42425.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_0, // @[:@42425.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_1, // @[:@42425.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_2, // @[:@42425.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_3, // @[:@42425.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_4, // @[:@42425.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_5, // @[:@42425.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_6, // @[:@42425.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_7, // @[:@42425.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_8, // @[:@42425.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_9, // @[:@42425.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_10, // @[:@42425.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_11, // @[:@42425.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_12, // @[:@42425.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_13, // @[:@42425.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_14, // @[:@42425.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_15, // @[:@42425.4]
  output         io_memStreams_gathers_0_data_ready, // @[:@42425.4]
  input          io_memStreams_gathers_0_data_valid, // @[:@42425.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_0, // @[:@42425.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_1, // @[:@42425.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_2, // @[:@42425.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_3, // @[:@42425.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_4, // @[:@42425.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_5, // @[:@42425.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_6, // @[:@42425.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_7, // @[:@42425.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_8, // @[:@42425.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_9, // @[:@42425.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_10, // @[:@42425.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_11, // @[:@42425.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_12, // @[:@42425.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_13, // @[:@42425.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_14, // @[:@42425.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_15, // @[:@42425.4]
  input          io_memStreams_scatters_0_cmd_ready, // @[:@42425.4]
  output         io_memStreams_scatters_0_cmd_valid, // @[:@42425.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_0, // @[:@42425.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_1, // @[:@42425.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_2, // @[:@42425.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_3, // @[:@42425.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_4, // @[:@42425.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_5, // @[:@42425.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_6, // @[:@42425.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_7, // @[:@42425.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_8, // @[:@42425.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_9, // @[:@42425.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_10, // @[:@42425.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_11, // @[:@42425.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_12, // @[:@42425.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_13, // @[:@42425.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_14, // @[:@42425.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_15, // @[:@42425.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_0, // @[:@42425.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_1, // @[:@42425.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_2, // @[:@42425.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_3, // @[:@42425.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_4, // @[:@42425.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_5, // @[:@42425.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_6, // @[:@42425.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_7, // @[:@42425.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_8, // @[:@42425.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_9, // @[:@42425.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_10, // @[:@42425.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_11, // @[:@42425.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_12, // @[:@42425.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_13, // @[:@42425.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_14, // @[:@42425.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_15, // @[:@42425.4]
  output         io_memStreams_scatters_0_wresp_ready, // @[:@42425.4]
  input          io_memStreams_scatters_0_wresp_valid, // @[:@42425.4]
  input          io_memStreams_scatters_0_wresp_bits, // @[:@42425.4]
  input          io_axiStreamsIn_0_TVALID, // @[:@42425.4]
  output         io_axiStreamsIn_0_TREADY, // @[:@42425.4]
  input  [255:0] io_axiStreamsIn_0_TDATA, // @[:@42425.4]
  input  [31:0]  io_axiStreamsIn_0_TSTRB, // @[:@42425.4]
  input  [31:0]  io_axiStreamsIn_0_TKEEP, // @[:@42425.4]
  input          io_axiStreamsIn_0_TLAST, // @[:@42425.4]
  input  [7:0]   io_axiStreamsIn_0_TID, // @[:@42425.4]
  input  [7:0]   io_axiStreamsIn_0_TDEST, // @[:@42425.4]
  input  [31:0]  io_axiStreamsIn_0_TUSER, // @[:@42425.4]
  output         io_axiStreamsOut_0_TVALID, // @[:@42425.4]
  input          io_axiStreamsOut_0_TREADY, // @[:@42425.4]
  output [255:0] io_axiStreamsOut_0_TDATA, // @[:@42425.4]
  output [31:0]  io_axiStreamsOut_0_TSTRB, // @[:@42425.4]
  output [31:0]  io_axiStreamsOut_0_TKEEP, // @[:@42425.4]
  output         io_axiStreamsOut_0_TLAST, // @[:@42425.4]
  output [7:0]   io_axiStreamsOut_0_TID, // @[:@42425.4]
  output [7:0]   io_axiStreamsOut_0_TDEST, // @[:@42425.4]
  output [31:0]  io_axiStreamsOut_0_TUSER, // @[:@42425.4]
  output         io_heap_0_req_valid, // @[:@42425.4]
  output         io_heap_0_req_bits_allocDealloc, // @[:@42425.4]
  output [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@42425.4]
  input          io_heap_0_resp_valid, // @[:@42425.4]
  input          io_heap_0_resp_bits_allocDealloc, // @[:@42425.4]
  input  [63:0]  io_heap_0_resp_bits_sizeAddr, // @[:@42425.4]
  input  [63:0]  io_argIns_0, // @[:@42425.4]
  input  [63:0]  io_argIns_1, // @[:@42425.4]
  input          io_argOuts_0_port_ready, // @[:@42425.4]
  output         io_argOuts_0_port_valid, // @[:@42425.4]
  output [63:0]  io_argOuts_0_port_bits, // @[:@42425.4]
  input  [63:0]  io_argOuts_0_echo // @[:@42425.4]
);
  wire  SingleCounter_clock; // @[Main.scala 35:32:@42588.4]
  wire  SingleCounter_reset; // @[Main.scala 35:32:@42588.4]
  wire  SingleCounter_io_input_reset; // @[Main.scala 35:32:@42588.4]
  wire  SingleCounter_io_output_done; // @[Main.scala 35:32:@42588.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@42606.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@42606.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@42606.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@42606.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@42606.4]
  wire  SRFF_clock; // @[Main.scala 39:28:@42615.4]
  wire  SRFF_reset; // @[Main.scala 39:28:@42615.4]
  wire  SRFF_io_input_set; // @[Main.scala 39:28:@42615.4]
  wire  SRFF_io_input_reset; // @[Main.scala 39:28:@42615.4]
  wire  SRFF_io_input_asyn_reset; // @[Main.scala 39:28:@42615.4]
  wire  SRFF_io_output; // @[Main.scala 39:28:@42615.4]
  wire  RootController_sm_clock; // @[sm_RootController.scala 32:18:@42654.4]
  wire  RootController_sm_reset; // @[sm_RootController.scala 32:18:@42654.4]
  wire  RootController_sm_io_enable; // @[sm_RootController.scala 32:18:@42654.4]
  wire  RootController_sm_io_done; // @[sm_RootController.scala 32:18:@42654.4]
  wire  RootController_sm_io_rst; // @[sm_RootController.scala 32:18:@42654.4]
  wire  RootController_sm_io_ctrDone; // @[sm_RootController.scala 32:18:@42654.4]
  wire  RootController_sm_io_ctrInc; // @[sm_RootController.scala 32:18:@42654.4]
  wire  RootController_sm_io_doneIn_0; // @[sm_RootController.scala 32:18:@42654.4]
  wire  RootController_sm_io_enableOut_0; // @[sm_RootController.scala 32:18:@42654.4]
  wire  RootController_sm_io_childAck_0; // @[sm_RootController.scala 32:18:@42654.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@42686.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@42686.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@42686.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@42686.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@42686.4]
  wire  RootController_kernelRootController_concrete1_clock; // @[sm_RootController.scala 73:24:@42748.4]
  wire  RootController_kernelRootController_concrete1_reset; // @[sm_RootController.scala 73:24:@42748.4]
  wire  RootController_kernelRootController_concrete1_io_in_x316_TVALID; // @[sm_RootController.scala 73:24:@42748.4]
  wire  RootController_kernelRootController_concrete1_io_in_x316_TREADY; // @[sm_RootController.scala 73:24:@42748.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x316_TDATA; // @[sm_RootController.scala 73:24:@42748.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x316_TID; // @[sm_RootController.scala 73:24:@42748.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x316_TDEST; // @[sm_RootController.scala 73:24:@42748.4]
  wire  RootController_kernelRootController_concrete1_io_in_x317_TVALID; // @[sm_RootController.scala 73:24:@42748.4]
  wire  RootController_kernelRootController_concrete1_io_in_x317_TREADY; // @[sm_RootController.scala 73:24:@42748.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x317_TDATA; // @[sm_RootController.scala 73:24:@42748.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_RootController.scala 73:24:@42748.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0; // @[sm_RootController.scala 73:24:@42748.4]
  wire  RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[sm_RootController.scala 73:24:@42748.4]
  wire  RootController_kernelRootController_concrete1_io_rr; // @[sm_RootController.scala 73:24:@42748.4]
  wire  _T_599; // @[package.scala 96:25:@42611.4 package.scala 96:25:@42612.4]
  wire  _T_664; // @[Main.scala 41:50:@42682.4]
  wire  _T_665; // @[Main.scala 41:59:@42683.4]
  wire  _T_677; // @[package.scala 100:49:@42703.4]
  reg  _T_680; // @[package.scala 48:56:@42704.4]
  reg [31:0] _RAND_0;
  SingleCounter SingleCounter ( // @[Main.scala 35:32:@42588.4]
    .clock(SingleCounter_clock),
    .reset(SingleCounter_reset),
    .io_input_reset(SingleCounter_io_input_reset),
    .io_output_done(SingleCounter_io_output_done)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@42606.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  SRFF SRFF ( // @[Main.scala 39:28:@42615.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  RootController_sm RootController_sm ( // @[sm_RootController.scala 32:18:@42654.4]
    .clock(RootController_sm_clock),
    .reset(RootController_sm_reset),
    .io_enable(RootController_sm_io_enable),
    .io_done(RootController_sm_io_done),
    .io_rst(RootController_sm_io_rst),
    .io_ctrDone(RootController_sm_io_ctrDone),
    .io_ctrInc(RootController_sm_io_ctrInc),
    .io_doneIn_0(RootController_sm_io_doneIn_0),
    .io_enableOut_0(RootController_sm_io_enableOut_0),
    .io_childAck_0(RootController_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@42686.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RootController_kernelRootController_concrete1 RootController_kernelRootController_concrete1 ( // @[sm_RootController.scala 73:24:@42748.4]
    .clock(RootController_kernelRootController_concrete1_clock),
    .reset(RootController_kernelRootController_concrete1_reset),
    .io_in_x316_TVALID(RootController_kernelRootController_concrete1_io_in_x316_TVALID),
    .io_in_x316_TREADY(RootController_kernelRootController_concrete1_io_in_x316_TREADY),
    .io_in_x316_TDATA(RootController_kernelRootController_concrete1_io_in_x316_TDATA),
    .io_in_x316_TID(RootController_kernelRootController_concrete1_io_in_x316_TID),
    .io_in_x316_TDEST(RootController_kernelRootController_concrete1_io_in_x316_TDEST),
    .io_in_x317_TVALID(RootController_kernelRootController_concrete1_io_in_x317_TVALID),
    .io_in_x317_TREADY(RootController_kernelRootController_concrete1_io_in_x317_TREADY),
    .io_in_x317_TDATA(RootController_kernelRootController_concrete1_io_in_x317_TDATA),
    .io_sigsIn_smEnableOuts_0(RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(RootController_kernelRootController_concrete1_io_rr)
  );
  assign _T_599 = RetimeWrapper_io_out; // @[package.scala 96:25:@42611.4 package.scala 96:25:@42612.4]
  assign _T_664 = io_enable & _T_599; // @[Main.scala 41:50:@42682.4]
  assign _T_665 = ~ SRFF_io_output; // @[Main.scala 41:59:@42683.4]
  assign _T_677 = RootController_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@42703.4]
  assign io_done = SRFF_io_output; // @[Main.scala 48:23:@42702.4]
  assign io_memStreams_loads_0_cmd_valid = 1'h0;
  assign io_memStreams_loads_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_loads_0_cmd_bits_size = 32'h0;
  assign io_memStreams_loads_0_data_ready = 1'h0;
  assign io_memStreams_stores_0_cmd_valid = 1'h0;
  assign io_memStreams_stores_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_stores_0_cmd_bits_size = 32'h0;
  assign io_memStreams_stores_0_data_valid = 1'h0;
  assign io_memStreams_stores_0_data_bits_wdata_0 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_1 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_2 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_3 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_4 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_5 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_6 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_7 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_8 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_9 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_10 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_11 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_12 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_13 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_14 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_15 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wstrb = 16'h0;
  assign io_memStreams_stores_0_wresp_ready = 1'h0;
  assign io_memStreams_gathers_0_cmd_valid = 1'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_0 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_1 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_2 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_3 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_4 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_5 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_6 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_7 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_8 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_9 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_10 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_11 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_12 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_13 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_14 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_15 = 64'h0;
  assign io_memStreams_gathers_0_data_ready = 1'h0;
  assign io_memStreams_scatters_0_cmd_valid = 1'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_0 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_1 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_2 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_3 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_4 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_5 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_6 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_7 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_8 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_9 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_10 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_11 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_12 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_13 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_14 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_15 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_0 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_1 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_2 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_3 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_4 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_5 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_6 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_7 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_8 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_9 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_10 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_11 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_12 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_13 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_14 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_15 = 32'h0;
  assign io_memStreams_scatters_0_wresp_ready = 1'h0;
  assign io_axiStreamsIn_0_TREADY = RootController_kernelRootController_concrete1_io_in_x316_TREADY; // @[sm_RootController.scala 48:23:@42804.4]
  assign io_axiStreamsOut_0_TVALID = RootController_kernelRootController_concrete1_io_in_x317_TVALID; // @[sm_RootController.scala 49:23:@42814.4]
  assign io_axiStreamsOut_0_TDATA = RootController_kernelRootController_concrete1_io_in_x317_TDATA; // @[sm_RootController.scala 49:23:@42812.4]
  assign io_axiStreamsOut_0_TSTRB = 32'hffffffff; // @[sm_RootController.scala 49:23:@42811.4]
  assign io_axiStreamsOut_0_TKEEP = 32'hffffffff; // @[sm_RootController.scala 49:23:@42810.4]
  assign io_axiStreamsOut_0_TLAST = 1'h0; // @[sm_RootController.scala 49:23:@42809.4]
  assign io_axiStreamsOut_0_TID = 8'h0; // @[sm_RootController.scala 49:23:@42808.4]
  assign io_axiStreamsOut_0_TDEST = 8'h0; // @[sm_RootController.scala 49:23:@42807.4]
  assign io_axiStreamsOut_0_TUSER = 32'h4; // @[sm_RootController.scala 49:23:@42806.4]
  assign io_heap_0_req_valid = 1'h0;
  assign io_heap_0_req_bits_allocDealloc = 1'h0;
  assign io_heap_0_req_bits_sizeAddr = 64'h0;
  assign io_argOuts_0_port_valid = 1'h0;
  assign io_argOuts_0_port_bits = 64'h0;
  assign SingleCounter_clock = clock; // @[:@42589.4]
  assign SingleCounter_reset = reset; // @[:@42590.4]
  assign SingleCounter_io_input_reset = reset; // @[Main.scala 36:79:@42604.4]
  assign RetimeWrapper_clock = clock; // @[:@42607.4]
  assign RetimeWrapper_reset = reset; // @[:@42608.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@42610.4]
  assign RetimeWrapper_io_in = SingleCounter_io_output_done; // @[package.scala 94:16:@42609.4]
  assign SRFF_clock = clock; // @[:@42616.4]
  assign SRFF_reset = reset; // @[:@42617.4]
  assign SRFF_io_input_set = RootController_sm_io_done; // @[Main.scala 57:29:@42842.4]
  assign SRFF_io_input_reset = RetimeWrapper_1_io_out; // @[Main.scala 46:31:@42700.4]
  assign SRFF_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[Main.scala 47:36:@42701.4]
  assign RootController_sm_clock = clock; // @[:@42655.4]
  assign RootController_sm_reset = reset; // @[:@42656.4]
  assign RootController_sm_io_enable = _T_664 & _T_665; // @[Main.scala 45:33:@42699.4 SpatialBlocks.scala 140:18:@42733.4]
  assign RootController_sm_io_rst = RetimeWrapper_1_io_out; // @[SpatialBlocks.scala 134:15:@42727.4]
  assign RootController_sm_io_ctrDone = RootController_sm_io_ctrInc & _T_680; // @[Main.scala 49:34:@42707.4]
  assign RootController_sm_io_doneIn_0 = RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@42724.4]
  assign RetimeWrapper_1_clock = clock; // @[:@42687.4]
  assign RetimeWrapper_1_reset = reset; // @[:@42688.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@42690.4]
  assign RetimeWrapper_1_io_in = reset | io_reset; // @[package.scala 94:16:@42689.4]
  assign RootController_kernelRootController_concrete1_clock = clock; // @[:@42749.4]
  assign RootController_kernelRootController_concrete1_reset = reset; // @[:@42750.4]
  assign RootController_kernelRootController_concrete1_io_in_x316_TVALID = io_axiStreamsIn_0_TVALID; // @[sm_RootController.scala 48:23:@42805.4]
  assign RootController_kernelRootController_concrete1_io_in_x316_TDATA = io_axiStreamsIn_0_TDATA; // @[sm_RootController.scala 48:23:@42803.4]
  assign RootController_kernelRootController_concrete1_io_in_x316_TID = io_axiStreamsIn_0_TID; // @[sm_RootController.scala 48:23:@42799.4]
  assign RootController_kernelRootController_concrete1_io_in_x316_TDEST = io_axiStreamsIn_0_TDEST; // @[sm_RootController.scala 48:23:@42798.4]
  assign RootController_kernelRootController_concrete1_io_in_x317_TREADY = io_axiStreamsOut_0_TREADY; // @[sm_RootController.scala 49:23:@42813.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0 = RootController_sm_io_enableOut_0; // @[sm_RootController.scala 78:22:@42823.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0 = RootController_sm_io_childAck_0; // @[sm_RootController.scala 78:22:@42821.4]
  assign RootController_kernelRootController_concrete1_io_rr = RetimeWrapper_io_out; // @[sm_RootController.scala 77:18:@42815.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_680 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_680 <= 1'h0;
    end else begin
      _T_680 <= _T_677;
    end
  end
endmodule
module SpatialIP( // @[:@42844.2]
  input         clock, // @[:@42845.4]
  input         reset, // @[:@42846.4]
  input  [31:0] io_raddr, // @[:@42847.4]
  input         io_wen, // @[:@42847.4]
  input  [31:0] io_waddr, // @[:@42847.4]
  input  [63:0] io_wdata, // @[:@42847.4]
  output [63:0] io_rdata // @[:@42847.4]
);
  wire  accel_clock; // @[Instantiator.scala 53:44:@42849.4]
  wire  accel_reset; // @[Instantiator.scala 53:44:@42849.4]
  wire  accel_io_enable; // @[Instantiator.scala 53:44:@42849.4]
  wire  accel_io_done; // @[Instantiator.scala 53:44:@42849.4]
  wire  accel_io_reset; // @[Instantiator.scala 53:44:@42849.4]
  wire  accel_io_memStreams_loads_0_cmd_ready; // @[Instantiator.scala 53:44:@42849.4]
  wire  accel_io_memStreams_loads_0_cmd_valid; // @[Instantiator.scala 53:44:@42849.4]
  wire [63:0] accel_io_memStreams_loads_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_loads_0_cmd_bits_size; // @[Instantiator.scala 53:44:@42849.4]
  wire  accel_io_memStreams_loads_0_data_ready; // @[Instantiator.scala 53:44:@42849.4]
  wire  accel_io_memStreams_loads_0_data_valid; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_0; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_1; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_2; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_3; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_4; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_5; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_6; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_7; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_8; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_9; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_10; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_11; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_12; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_13; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_14; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_15; // @[Instantiator.scala 53:44:@42849.4]
  wire  accel_io_memStreams_stores_0_cmd_ready; // @[Instantiator.scala 53:44:@42849.4]
  wire  accel_io_memStreams_stores_0_cmd_valid; // @[Instantiator.scala 53:44:@42849.4]
  wire [63:0] accel_io_memStreams_stores_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_stores_0_cmd_bits_size; // @[Instantiator.scala 53:44:@42849.4]
  wire  accel_io_memStreams_stores_0_data_ready; // @[Instantiator.scala 53:44:@42849.4]
  wire  accel_io_memStreams_stores_0_data_valid; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_1; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_2; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_3; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_4; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_5; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_6; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_7; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_8; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_9; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_10; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_11; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_12; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_13; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_14; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_15; // @[Instantiator.scala 53:44:@42849.4]
  wire [15:0] accel_io_memStreams_stores_0_data_bits_wstrb; // @[Instantiator.scala 53:44:@42849.4]
  wire  accel_io_memStreams_stores_0_wresp_ready; // @[Instantiator.scala 53:44:@42849.4]
  wire  accel_io_memStreams_stores_0_wresp_valid; // @[Instantiator.scala 53:44:@42849.4]
  wire  accel_io_memStreams_stores_0_wresp_bits; // @[Instantiator.scala 53:44:@42849.4]
  wire  accel_io_memStreams_gathers_0_cmd_ready; // @[Instantiator.scala 53:44:@42849.4]
  wire  accel_io_memStreams_gathers_0_cmd_valid; // @[Instantiator.scala 53:44:@42849.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_0; // @[Instantiator.scala 53:44:@42849.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_1; // @[Instantiator.scala 53:44:@42849.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_2; // @[Instantiator.scala 53:44:@42849.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_3; // @[Instantiator.scala 53:44:@42849.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_4; // @[Instantiator.scala 53:44:@42849.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_5; // @[Instantiator.scala 53:44:@42849.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_6; // @[Instantiator.scala 53:44:@42849.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_7; // @[Instantiator.scala 53:44:@42849.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_8; // @[Instantiator.scala 53:44:@42849.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_9; // @[Instantiator.scala 53:44:@42849.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_10; // @[Instantiator.scala 53:44:@42849.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_11; // @[Instantiator.scala 53:44:@42849.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_12; // @[Instantiator.scala 53:44:@42849.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_13; // @[Instantiator.scala 53:44:@42849.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_14; // @[Instantiator.scala 53:44:@42849.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_15; // @[Instantiator.scala 53:44:@42849.4]
  wire  accel_io_memStreams_gathers_0_data_ready; // @[Instantiator.scala 53:44:@42849.4]
  wire  accel_io_memStreams_gathers_0_data_valid; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_0; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_1; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_2; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_3; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_4; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_5; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_6; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_7; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_8; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_9; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_10; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_11; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_12; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_13; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_14; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_15; // @[Instantiator.scala 53:44:@42849.4]
  wire  accel_io_memStreams_scatters_0_cmd_ready; // @[Instantiator.scala 53:44:@42849.4]
  wire  accel_io_memStreams_scatters_0_cmd_valid; // @[Instantiator.scala 53:44:@42849.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0; // @[Instantiator.scala 53:44:@42849.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1; // @[Instantiator.scala 53:44:@42849.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2; // @[Instantiator.scala 53:44:@42849.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3; // @[Instantiator.scala 53:44:@42849.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4; // @[Instantiator.scala 53:44:@42849.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5; // @[Instantiator.scala 53:44:@42849.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6; // @[Instantiator.scala 53:44:@42849.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7; // @[Instantiator.scala 53:44:@42849.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8; // @[Instantiator.scala 53:44:@42849.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9; // @[Instantiator.scala 53:44:@42849.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10; // @[Instantiator.scala 53:44:@42849.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11; // @[Instantiator.scala 53:44:@42849.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12; // @[Instantiator.scala 53:44:@42849.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13; // @[Instantiator.scala 53:44:@42849.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14; // @[Instantiator.scala 53:44:@42849.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_0; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_1; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_2; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_3; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_4; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_5; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_6; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_7; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_8; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_9; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_10; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_11; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_12; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_13; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_14; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_15; // @[Instantiator.scala 53:44:@42849.4]
  wire  accel_io_memStreams_scatters_0_wresp_ready; // @[Instantiator.scala 53:44:@42849.4]
  wire  accel_io_memStreams_scatters_0_wresp_valid; // @[Instantiator.scala 53:44:@42849.4]
  wire  accel_io_memStreams_scatters_0_wresp_bits; // @[Instantiator.scala 53:44:@42849.4]
  wire  accel_io_axiStreamsIn_0_TVALID; // @[Instantiator.scala 53:44:@42849.4]
  wire  accel_io_axiStreamsIn_0_TREADY; // @[Instantiator.scala 53:44:@42849.4]
  wire [255:0] accel_io_axiStreamsIn_0_TDATA; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_axiStreamsIn_0_TSTRB; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_axiStreamsIn_0_TKEEP; // @[Instantiator.scala 53:44:@42849.4]
  wire  accel_io_axiStreamsIn_0_TLAST; // @[Instantiator.scala 53:44:@42849.4]
  wire [7:0] accel_io_axiStreamsIn_0_TID; // @[Instantiator.scala 53:44:@42849.4]
  wire [7:0] accel_io_axiStreamsIn_0_TDEST; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_axiStreamsIn_0_TUSER; // @[Instantiator.scala 53:44:@42849.4]
  wire  accel_io_axiStreamsOut_0_TVALID; // @[Instantiator.scala 53:44:@42849.4]
  wire  accel_io_axiStreamsOut_0_TREADY; // @[Instantiator.scala 53:44:@42849.4]
  wire [255:0] accel_io_axiStreamsOut_0_TDATA; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_axiStreamsOut_0_TSTRB; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_axiStreamsOut_0_TKEEP; // @[Instantiator.scala 53:44:@42849.4]
  wire  accel_io_axiStreamsOut_0_TLAST; // @[Instantiator.scala 53:44:@42849.4]
  wire [7:0] accel_io_axiStreamsOut_0_TID; // @[Instantiator.scala 53:44:@42849.4]
  wire [7:0] accel_io_axiStreamsOut_0_TDEST; // @[Instantiator.scala 53:44:@42849.4]
  wire [31:0] accel_io_axiStreamsOut_0_TUSER; // @[Instantiator.scala 53:44:@42849.4]
  wire  accel_io_heap_0_req_valid; // @[Instantiator.scala 53:44:@42849.4]
  wire  accel_io_heap_0_req_bits_allocDealloc; // @[Instantiator.scala 53:44:@42849.4]
  wire [63:0] accel_io_heap_0_req_bits_sizeAddr; // @[Instantiator.scala 53:44:@42849.4]
  wire  accel_io_heap_0_resp_valid; // @[Instantiator.scala 53:44:@42849.4]
  wire  accel_io_heap_0_resp_bits_allocDealloc; // @[Instantiator.scala 53:44:@42849.4]
  wire [63:0] accel_io_heap_0_resp_bits_sizeAddr; // @[Instantiator.scala 53:44:@42849.4]
  wire [63:0] accel_io_argIns_0; // @[Instantiator.scala 53:44:@42849.4]
  wire [63:0] accel_io_argIns_1; // @[Instantiator.scala 53:44:@42849.4]
  wire  accel_io_argOuts_0_port_ready; // @[Instantiator.scala 53:44:@42849.4]
  wire  accel_io_argOuts_0_port_valid; // @[Instantiator.scala 53:44:@42849.4]
  wire [63:0] accel_io_argOuts_0_port_bits; // @[Instantiator.scala 53:44:@42849.4]
  wire [63:0] accel_io_argOuts_0_echo; // @[Instantiator.scala 53:44:@42849.4]
  AccelUnit accel ( // @[Instantiator.scala 53:44:@42849.4]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_enable(accel_io_enable),
    .io_done(accel_io_done),
    .io_reset(accel_io_reset),
    .io_memStreams_loads_0_cmd_ready(accel_io_memStreams_loads_0_cmd_ready),
    .io_memStreams_loads_0_cmd_valid(accel_io_memStreams_loads_0_cmd_valid),
    .io_memStreams_loads_0_cmd_bits_addr(accel_io_memStreams_loads_0_cmd_bits_addr),
    .io_memStreams_loads_0_cmd_bits_size(accel_io_memStreams_loads_0_cmd_bits_size),
    .io_memStreams_loads_0_data_ready(accel_io_memStreams_loads_0_data_ready),
    .io_memStreams_loads_0_data_valid(accel_io_memStreams_loads_0_data_valid),
    .io_memStreams_loads_0_data_bits_rdata_0(accel_io_memStreams_loads_0_data_bits_rdata_0),
    .io_memStreams_loads_0_data_bits_rdata_1(accel_io_memStreams_loads_0_data_bits_rdata_1),
    .io_memStreams_loads_0_data_bits_rdata_2(accel_io_memStreams_loads_0_data_bits_rdata_2),
    .io_memStreams_loads_0_data_bits_rdata_3(accel_io_memStreams_loads_0_data_bits_rdata_3),
    .io_memStreams_loads_0_data_bits_rdata_4(accel_io_memStreams_loads_0_data_bits_rdata_4),
    .io_memStreams_loads_0_data_bits_rdata_5(accel_io_memStreams_loads_0_data_bits_rdata_5),
    .io_memStreams_loads_0_data_bits_rdata_6(accel_io_memStreams_loads_0_data_bits_rdata_6),
    .io_memStreams_loads_0_data_bits_rdata_7(accel_io_memStreams_loads_0_data_bits_rdata_7),
    .io_memStreams_loads_0_data_bits_rdata_8(accel_io_memStreams_loads_0_data_bits_rdata_8),
    .io_memStreams_loads_0_data_bits_rdata_9(accel_io_memStreams_loads_0_data_bits_rdata_9),
    .io_memStreams_loads_0_data_bits_rdata_10(accel_io_memStreams_loads_0_data_bits_rdata_10),
    .io_memStreams_loads_0_data_bits_rdata_11(accel_io_memStreams_loads_0_data_bits_rdata_11),
    .io_memStreams_loads_0_data_bits_rdata_12(accel_io_memStreams_loads_0_data_bits_rdata_12),
    .io_memStreams_loads_0_data_bits_rdata_13(accel_io_memStreams_loads_0_data_bits_rdata_13),
    .io_memStreams_loads_0_data_bits_rdata_14(accel_io_memStreams_loads_0_data_bits_rdata_14),
    .io_memStreams_loads_0_data_bits_rdata_15(accel_io_memStreams_loads_0_data_bits_rdata_15),
    .io_memStreams_stores_0_cmd_ready(accel_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(accel_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(accel_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(accel_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(accel_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(accel_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(accel_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wdata_1(accel_io_memStreams_stores_0_data_bits_wdata_1),
    .io_memStreams_stores_0_data_bits_wdata_2(accel_io_memStreams_stores_0_data_bits_wdata_2),
    .io_memStreams_stores_0_data_bits_wdata_3(accel_io_memStreams_stores_0_data_bits_wdata_3),
    .io_memStreams_stores_0_data_bits_wdata_4(accel_io_memStreams_stores_0_data_bits_wdata_4),
    .io_memStreams_stores_0_data_bits_wdata_5(accel_io_memStreams_stores_0_data_bits_wdata_5),
    .io_memStreams_stores_0_data_bits_wdata_6(accel_io_memStreams_stores_0_data_bits_wdata_6),
    .io_memStreams_stores_0_data_bits_wdata_7(accel_io_memStreams_stores_0_data_bits_wdata_7),
    .io_memStreams_stores_0_data_bits_wdata_8(accel_io_memStreams_stores_0_data_bits_wdata_8),
    .io_memStreams_stores_0_data_bits_wdata_9(accel_io_memStreams_stores_0_data_bits_wdata_9),
    .io_memStreams_stores_0_data_bits_wdata_10(accel_io_memStreams_stores_0_data_bits_wdata_10),
    .io_memStreams_stores_0_data_bits_wdata_11(accel_io_memStreams_stores_0_data_bits_wdata_11),
    .io_memStreams_stores_0_data_bits_wdata_12(accel_io_memStreams_stores_0_data_bits_wdata_12),
    .io_memStreams_stores_0_data_bits_wdata_13(accel_io_memStreams_stores_0_data_bits_wdata_13),
    .io_memStreams_stores_0_data_bits_wdata_14(accel_io_memStreams_stores_0_data_bits_wdata_14),
    .io_memStreams_stores_0_data_bits_wdata_15(accel_io_memStreams_stores_0_data_bits_wdata_15),
    .io_memStreams_stores_0_data_bits_wstrb(accel_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(accel_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(accel_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(accel_io_memStreams_stores_0_wresp_bits),
    .io_memStreams_gathers_0_cmd_ready(accel_io_memStreams_gathers_0_cmd_ready),
    .io_memStreams_gathers_0_cmd_valid(accel_io_memStreams_gathers_0_cmd_valid),
    .io_memStreams_gathers_0_cmd_bits_addr_0(accel_io_memStreams_gathers_0_cmd_bits_addr_0),
    .io_memStreams_gathers_0_cmd_bits_addr_1(accel_io_memStreams_gathers_0_cmd_bits_addr_1),
    .io_memStreams_gathers_0_cmd_bits_addr_2(accel_io_memStreams_gathers_0_cmd_bits_addr_2),
    .io_memStreams_gathers_0_cmd_bits_addr_3(accel_io_memStreams_gathers_0_cmd_bits_addr_3),
    .io_memStreams_gathers_0_cmd_bits_addr_4(accel_io_memStreams_gathers_0_cmd_bits_addr_4),
    .io_memStreams_gathers_0_cmd_bits_addr_5(accel_io_memStreams_gathers_0_cmd_bits_addr_5),
    .io_memStreams_gathers_0_cmd_bits_addr_6(accel_io_memStreams_gathers_0_cmd_bits_addr_6),
    .io_memStreams_gathers_0_cmd_bits_addr_7(accel_io_memStreams_gathers_0_cmd_bits_addr_7),
    .io_memStreams_gathers_0_cmd_bits_addr_8(accel_io_memStreams_gathers_0_cmd_bits_addr_8),
    .io_memStreams_gathers_0_cmd_bits_addr_9(accel_io_memStreams_gathers_0_cmd_bits_addr_9),
    .io_memStreams_gathers_0_cmd_bits_addr_10(accel_io_memStreams_gathers_0_cmd_bits_addr_10),
    .io_memStreams_gathers_0_cmd_bits_addr_11(accel_io_memStreams_gathers_0_cmd_bits_addr_11),
    .io_memStreams_gathers_0_cmd_bits_addr_12(accel_io_memStreams_gathers_0_cmd_bits_addr_12),
    .io_memStreams_gathers_0_cmd_bits_addr_13(accel_io_memStreams_gathers_0_cmd_bits_addr_13),
    .io_memStreams_gathers_0_cmd_bits_addr_14(accel_io_memStreams_gathers_0_cmd_bits_addr_14),
    .io_memStreams_gathers_0_cmd_bits_addr_15(accel_io_memStreams_gathers_0_cmd_bits_addr_15),
    .io_memStreams_gathers_0_data_ready(accel_io_memStreams_gathers_0_data_ready),
    .io_memStreams_gathers_0_data_valid(accel_io_memStreams_gathers_0_data_valid),
    .io_memStreams_gathers_0_data_bits_0(accel_io_memStreams_gathers_0_data_bits_0),
    .io_memStreams_gathers_0_data_bits_1(accel_io_memStreams_gathers_0_data_bits_1),
    .io_memStreams_gathers_0_data_bits_2(accel_io_memStreams_gathers_0_data_bits_2),
    .io_memStreams_gathers_0_data_bits_3(accel_io_memStreams_gathers_0_data_bits_3),
    .io_memStreams_gathers_0_data_bits_4(accel_io_memStreams_gathers_0_data_bits_4),
    .io_memStreams_gathers_0_data_bits_5(accel_io_memStreams_gathers_0_data_bits_5),
    .io_memStreams_gathers_0_data_bits_6(accel_io_memStreams_gathers_0_data_bits_6),
    .io_memStreams_gathers_0_data_bits_7(accel_io_memStreams_gathers_0_data_bits_7),
    .io_memStreams_gathers_0_data_bits_8(accel_io_memStreams_gathers_0_data_bits_8),
    .io_memStreams_gathers_0_data_bits_9(accel_io_memStreams_gathers_0_data_bits_9),
    .io_memStreams_gathers_0_data_bits_10(accel_io_memStreams_gathers_0_data_bits_10),
    .io_memStreams_gathers_0_data_bits_11(accel_io_memStreams_gathers_0_data_bits_11),
    .io_memStreams_gathers_0_data_bits_12(accel_io_memStreams_gathers_0_data_bits_12),
    .io_memStreams_gathers_0_data_bits_13(accel_io_memStreams_gathers_0_data_bits_13),
    .io_memStreams_gathers_0_data_bits_14(accel_io_memStreams_gathers_0_data_bits_14),
    .io_memStreams_gathers_0_data_bits_15(accel_io_memStreams_gathers_0_data_bits_15),
    .io_memStreams_scatters_0_cmd_ready(accel_io_memStreams_scatters_0_cmd_ready),
    .io_memStreams_scatters_0_cmd_valid(accel_io_memStreams_scatters_0_cmd_valid),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_0(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_1(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_2(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_3(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_4(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_5(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_6(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_7(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_8(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_9(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_10(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_11(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_12(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_13(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_14(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_15(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15),
    .io_memStreams_scatters_0_cmd_bits_wdata_0(accel_io_memStreams_scatters_0_cmd_bits_wdata_0),
    .io_memStreams_scatters_0_cmd_bits_wdata_1(accel_io_memStreams_scatters_0_cmd_bits_wdata_1),
    .io_memStreams_scatters_0_cmd_bits_wdata_2(accel_io_memStreams_scatters_0_cmd_bits_wdata_2),
    .io_memStreams_scatters_0_cmd_bits_wdata_3(accel_io_memStreams_scatters_0_cmd_bits_wdata_3),
    .io_memStreams_scatters_0_cmd_bits_wdata_4(accel_io_memStreams_scatters_0_cmd_bits_wdata_4),
    .io_memStreams_scatters_0_cmd_bits_wdata_5(accel_io_memStreams_scatters_0_cmd_bits_wdata_5),
    .io_memStreams_scatters_0_cmd_bits_wdata_6(accel_io_memStreams_scatters_0_cmd_bits_wdata_6),
    .io_memStreams_scatters_0_cmd_bits_wdata_7(accel_io_memStreams_scatters_0_cmd_bits_wdata_7),
    .io_memStreams_scatters_0_cmd_bits_wdata_8(accel_io_memStreams_scatters_0_cmd_bits_wdata_8),
    .io_memStreams_scatters_0_cmd_bits_wdata_9(accel_io_memStreams_scatters_0_cmd_bits_wdata_9),
    .io_memStreams_scatters_0_cmd_bits_wdata_10(accel_io_memStreams_scatters_0_cmd_bits_wdata_10),
    .io_memStreams_scatters_0_cmd_bits_wdata_11(accel_io_memStreams_scatters_0_cmd_bits_wdata_11),
    .io_memStreams_scatters_0_cmd_bits_wdata_12(accel_io_memStreams_scatters_0_cmd_bits_wdata_12),
    .io_memStreams_scatters_0_cmd_bits_wdata_13(accel_io_memStreams_scatters_0_cmd_bits_wdata_13),
    .io_memStreams_scatters_0_cmd_bits_wdata_14(accel_io_memStreams_scatters_0_cmd_bits_wdata_14),
    .io_memStreams_scatters_0_cmd_bits_wdata_15(accel_io_memStreams_scatters_0_cmd_bits_wdata_15),
    .io_memStreams_scatters_0_wresp_ready(accel_io_memStreams_scatters_0_wresp_ready),
    .io_memStreams_scatters_0_wresp_valid(accel_io_memStreams_scatters_0_wresp_valid),
    .io_memStreams_scatters_0_wresp_bits(accel_io_memStreams_scatters_0_wresp_bits),
    .io_axiStreamsIn_0_TVALID(accel_io_axiStreamsIn_0_TVALID),
    .io_axiStreamsIn_0_TREADY(accel_io_axiStreamsIn_0_TREADY),
    .io_axiStreamsIn_0_TDATA(accel_io_axiStreamsIn_0_TDATA),
    .io_axiStreamsIn_0_TSTRB(accel_io_axiStreamsIn_0_TSTRB),
    .io_axiStreamsIn_0_TKEEP(accel_io_axiStreamsIn_0_TKEEP),
    .io_axiStreamsIn_0_TLAST(accel_io_axiStreamsIn_0_TLAST),
    .io_axiStreamsIn_0_TID(accel_io_axiStreamsIn_0_TID),
    .io_axiStreamsIn_0_TDEST(accel_io_axiStreamsIn_0_TDEST),
    .io_axiStreamsIn_0_TUSER(accel_io_axiStreamsIn_0_TUSER),
    .io_axiStreamsOut_0_TVALID(accel_io_axiStreamsOut_0_TVALID),
    .io_axiStreamsOut_0_TREADY(accel_io_axiStreamsOut_0_TREADY),
    .io_axiStreamsOut_0_TDATA(accel_io_axiStreamsOut_0_TDATA),
    .io_axiStreamsOut_0_TSTRB(accel_io_axiStreamsOut_0_TSTRB),
    .io_axiStreamsOut_0_TKEEP(accel_io_axiStreamsOut_0_TKEEP),
    .io_axiStreamsOut_0_TLAST(accel_io_axiStreamsOut_0_TLAST),
    .io_axiStreamsOut_0_TID(accel_io_axiStreamsOut_0_TID),
    .io_axiStreamsOut_0_TDEST(accel_io_axiStreamsOut_0_TDEST),
    .io_axiStreamsOut_0_TUSER(accel_io_axiStreamsOut_0_TUSER),
    .io_heap_0_req_valid(accel_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(accel_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(accel_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(accel_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(accel_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(accel_io_heap_0_resp_bits_sizeAddr),
    .io_argIns_0(accel_io_argIns_0),
    .io_argIns_1(accel_io_argIns_1),
    .io_argOuts_0_port_ready(accel_io_argOuts_0_port_ready),
    .io_argOuts_0_port_valid(accel_io_argOuts_0_port_valid),
    .io_argOuts_0_port_bits(accel_io_argOuts_0_port_bits),
    .io_argOuts_0_echo(accel_io_argOuts_0_echo)
  );
  assign io_rdata = 64'h0;
  assign accel_clock = clock; // @[:@42850.4]
  assign accel_reset = reset; // @[:@42851.4]
  assign accel_io_enable = 1'h0;
  assign accel_io_reset = 1'h0;
  assign accel_io_memStreams_loads_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_loads_0_data_valid = 1'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_0 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_1 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_2 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_3 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_4 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_5 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_6 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_7 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_8 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_9 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_10 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_11 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_12 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_13 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_14 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_15 = 32'h0;
  assign accel_io_memStreams_stores_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_stores_0_data_ready = 1'h0;
  assign accel_io_memStreams_stores_0_wresp_valid = 1'h0;
  assign accel_io_memStreams_stores_0_wresp_bits = 1'h0;
  assign accel_io_memStreams_gathers_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_gathers_0_data_valid = 1'h0;
  assign accel_io_memStreams_gathers_0_data_bits_0 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_1 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_2 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_3 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_4 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_5 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_6 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_7 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_8 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_9 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_10 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_11 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_12 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_13 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_14 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_15 = 32'h0;
  assign accel_io_memStreams_scatters_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_scatters_0_wresp_valid = 1'h0;
  assign accel_io_memStreams_scatters_0_wresp_bits = 1'h0;
  assign accel_io_axiStreamsIn_0_TVALID = 1'h0;
  assign accel_io_axiStreamsIn_0_TDATA = 256'h0;
  assign accel_io_axiStreamsIn_0_TSTRB = 32'h0;
  assign accel_io_axiStreamsIn_0_TKEEP = 32'h0;
  assign accel_io_axiStreamsIn_0_TLAST = 1'h0;
  assign accel_io_axiStreamsIn_0_TID = 8'h0;
  assign accel_io_axiStreamsIn_0_TDEST = 8'h0;
  assign accel_io_axiStreamsIn_0_TUSER = 32'h0;
  assign accel_io_axiStreamsOut_0_TREADY = 1'h0;
  assign accel_io_heap_0_resp_valid = 1'h0;
  assign accel_io_heap_0_resp_bits_allocDealloc = 1'h0;
  assign accel_io_heap_0_resp_bits_sizeAddr = 64'h0;
  assign accel_io_argIns_0 = 64'h0;
  assign accel_io_argIns_1 = 64'h0;
  assign accel_io_argOuts_0_port_ready = 1'h0;
  assign accel_io_argOuts_0_echo = 64'h0;
endmodule
