// Latency = 4
module top(
  input CLK/*verilator public*/, 
  input [7:0] I_0_0_0/*verilator public*/, 
  output [7:0] O_0_0_0/*verilator public*/, 
  input [7:0] I_1_0_0/*verilator public*/, 
  output [7:0] O_1_0_0/*verilator public*/, 
  output valid_down/*verilator public*/, 
  input valid_up/*verilator public*/
);
  wire dontcare;
  wire [31:0] io_output_counts_1;
  wire [31:0] io_output_counts_0;

  x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1 sampler_box ( // @[m_x55_ctr_0.scala 26:17:@1721.4]
    .clock(CLK), // @[:@1296.4]
    .reset('b0), // @[:@1297.4]
    .io_in_x275_TREADY(dontcare), // @[:@1298.4]
    .io_in_x275_TDATA({I_0_0_0,I_1_0_0}), // @[:@1298.4]
    .io_in_x275_TID(8'h0),
    .io_in_x275_TDEST(8'h0),
    .io_in_x276_TVALID(valid_down), // @[:@1298.4]
    .io_in_x276_TDATA({O_0_0_0,O_1_0_0}), // @[:@1298.4]
    .io_in_x276_TREADY(1'b1), // @[:@1298.4]
    .io_sigsIn_datapathEn(valid_up), // @[:@1298.4]
    .io_sigsIn_backpressure(1'b1), // @[:@20563.4]
    .io_sigsIn_break(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_1(io_output_counts_1), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_0(io_output_counts_0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_0(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_1(1'b0), // @[:@20563.4]
    .io_rr('b1) // @[:@1298.4]
  );

  wire dontcare2;

  wire io_output_oobs_0;
  wire io_output_oobs_1;
  x283_ctrchain cchain ( // @[:@2879.2]
    .clock(CLK), // @[:@2880.4]
    .reset(1'b0), // @[:@2881.4]
    .io_input_reset(1'b0), // @[:@2882.4]
    .io_input_enable(valid_up), // @[:@2882.4]
    .io_output_counts_1(io_output_counts_1), // @[:@2882.4]
    .io_output_counts_0(io_output_counts_0), // @[:@2882.4]
    .io_output_oobs_0(io_output_oobs_0), // @[:@2882.4]
    .io_output_oobs_1(io_output_oobs_1), // @[:@2882.4]
    .io_output_done(dontcare2) // @[:@2882.4]
  );

endmodule

module RetimeShiftRegister
#(
    parameter WIDTH = 1,
    parameter STAGES = 1)
(
    input clock,
    input reset,
    input flow,
    input [WIDTH-1:0] init,
    input [WIDTH-1:0] in,
    output reg [WIDTH-1:0] out
);
  integer i;
  reg [WIDTH-1:0] sr[STAGES:0]; // Create 'STAGES' number of register, each 'WIDTH' bits wide

   /* synopsys dc_tcl_script_begin
    set_ungroup [current_design] true
    set_flatten true -effort high -phase true -design [current_design]
    set_dont_retime [current_design] false
    set_optimize_registers true -design [current_design]
    */
  always @(posedge clock) begin
    if (reset) begin
      for(i=0; i<STAGES; i=i+1) begin
        sr[i] <= init;
      end
    end else begin
      if (flow) begin 
        sr[0] <= in;
        for(i=1; i<STAGES; i=i+1) begin
          sr[i] <= sr[i-1];
        end
      end
    end
  end

  always @(*) begin
    out = sr[STAGES-1];
  end
endmodule

module FF( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  output [31:0] io_rPort_0_output_0, // @[:@6.4]
  input  [31:0] io_wPort_0_data_0, // @[:@6.4]
  input         io_wPort_0_reset, // @[:@6.4]
  input         io_wPort_0_en_0 // @[:@6.4]
);
  reg [31:0] ff; // @[MemPrimitives.scala 173:19:@21.4]
  reg [31:0] _RAND_0;
  wire [31:0] _T_68; // @[MemPrimitives.scala 177:32:@23.4]
  wire [31:0] _T_69; // @[MemPrimitives.scala 177:12:@24.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 177:32:@23.4]
  assign _T_69 = io_wPort_0_reset ? 32'h0 : _T_68; // @[MemPrimitives.scala 177:12:@24.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 178:34:@26.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 32'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 32'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SRFF( // @[:@28.2]
  input   clock, // @[:@29.4]
  input   reset, // @[:@30.4]
  input   io_input_set, // @[:@31.4]
  input   io_input_reset, // @[:@31.4]
  input   io_input_asyn_reset, // @[:@31.4]
  output  io_output // @[:@31.4]
);
  reg  _T_15; // @[SRFF.scala 20:21:@33.4]
  reg [31:0] _RAND_0;
  wire  _T_19; // @[SRFF.scala 21:74:@34.4]
  wire  _T_20; // @[SRFF.scala 21:48:@35.4]
  wire  _T_21; // @[SRFF.scala 21:14:@36.4]
  assign _T_19 = io_input_reset ? 1'h0 : _T_15; // @[SRFF.scala 21:74:@34.4]
  assign _T_20 = io_input_set ? 1'h1 : _T_19; // @[SRFF.scala 21:48:@35.4]
  assign _T_21 = io_input_asyn_reset ? 1'h0 : _T_20; // @[SRFF.scala 21:14:@36.4]
  assign io_output = io_input_asyn_reset ? 1'h0 : _T_15; // @[SRFF.scala 22:15:@39.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_15 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_15 <= 1'h0;
    end else begin
      if (io_input_asyn_reset) begin
        _T_15 <= 1'h0;
      end else begin
        if (io_input_set) begin
          _T_15 <= 1'h1;
        end else begin
          if (io_input_reset) begin
            _T_15 <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module SingleCounter( // @[:@41.2]
  input   clock, // @[:@42.4]
  input   reset, // @[:@43.4]
  input   io_input_reset, // @[:@44.4]
  output  io_output_done // @[:@44.4]
);
  wire  bases_0_clock; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_reset; // @[Counter.scala 253:53:@57.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 253:53:@57.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 253:53:@57.4]
  wire  SRFF_clock; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_set; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_output; // @[Counter.scala 255:22:@73.4]
  wire [31:0] _T_48; // @[Counter.scala 279:52:@101.4]
  wire [32:0] _T_50; // @[Counter.scala 283:33:@102.4]
  wire [31:0] _T_51; // @[Counter.scala 283:33:@103.4]
  wire [31:0] _T_52; // @[Counter.scala 283:33:@104.4]
  wire  _T_57; // @[Counter.scala 285:18:@106.4]
  wire [31:0] _T_68; // @[Counter.scala 291:115:@114.4]
  wire [31:0] _T_71; // @[Counter.scala 291:152:@117.4]
  wire [31:0] _T_72; // @[Counter.scala 291:74:@118.4]
  FF bases_0 ( // @[Counter.scala 253:53:@57.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 255:22:@73.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 279:52:@101.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@102.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@103.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 283:33:@104.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh14); // @[Counter.scala 285:18:@106.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 291:115:@114.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 291:152:@117.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 291:74:@118.4]
  assign io_output_done = $signed(_T_52) >= $signed(32'sh14); // @[Counter.scala 325:20:@127.4]
  assign bases_0_clock = clock; // @[:@58.4]
  assign bases_0_reset = reset; // @[:@59.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 291:31:@120.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 273:27:@99.4]
  assign bases_0_io_wPort_0_en_0 = 1'h1; // @[Counter.scala 276:29:@100.4]
  assign SRFF_clock = clock; // @[:@74.4]
  assign SRFF_reset = reset; // @[:@75.4]
  assign SRFF_io_input_set = io_input_reset == 1'h0; // @[Counter.scala 256:23:@78.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 257:25:@80.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 258:30:@81.4]
endmodule
module RetimeWrapper( // @[:@144.2]
  input   clock, // @[:@145.4]
  input   reset, // @[:@146.4]
  input   io_flow, // @[:@147.4]
  input   io_in, // @[:@147.4]
  output  io_out // @[:@147.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@149.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@149.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@162.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@161.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@160.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@159.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@158.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@156.4]
endmodule
module RootController_sm( // @[:@312.2]
  input   clock, // @[:@313.4]
  input   reset, // @[:@314.4]
  input   io_enable, // @[:@315.4]
  output  io_done, // @[:@315.4]
  input   io_rst, // @[:@315.4]
  input   io_ctrDone, // @[:@315.4]
  output  io_ctrInc, // @[:@315.4]
  input   io_doneIn_0, // @[:@315.4]
  output  io_enableOut_0, // @[:@315.4]
  output  io_childAck_0 // @[:@315.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@318.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@321.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@338.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@433.4]
  wire  finished; // @[Controllers.scala 81:26:@324.4]
  wire  synchronize; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  wire  _T_122; // @[Controllers.scala 128:33:@371.4]
  wire  _T_124; // @[Controllers.scala 128:54:@372.4]
  wire  _T_125; // @[Controllers.scala 128:52:@373.4]
  wire  _T_126; // @[Controllers.scala 128:66:@374.4]
  wire  _T_128; // @[Controllers.scala 128:98:@376.4]
  wire  _T_129; // @[Controllers.scala 128:96:@377.4]
  wire  _T_131; // @[Controllers.scala 128:123:@378.4]
  wire  _T_133; // @[Controllers.scala 129:48:@381.4]
  wire  _T_138; // @[Controllers.scala 130:52:@386.4]
  wire  _T_139; // @[Controllers.scala 130:50:@387.4]
  wire  _T_147; // @[Controllers.scala 130:129:@393.4]
  wire  _T_150; // @[Controllers.scala 131:45:@396.4]
  wire  _T_154; // @[Controllers.scala 213:68:@402.4]
  wire  _T_156; // @[Controllers.scala 213:90:@404.4]
  wire  _T_158; // @[Controllers.scala 213:132:@406.4]
  wire  _T_159; // @[Controllers.scala 213:130:@407.4]
  wire  _T_160; // @[Controllers.scala 213:156:@408.4]
  reg  _T_166; // @[package.scala 48:56:@412.4]
  reg [31:0] _RAND_0;
  reg  _T_180; // @[package.scala 48:56:@430.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@318.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@321.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@338.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@357.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@416.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@433.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  assign finished = done_0_io_output | io_done; // @[Controllers.scala 81:26:@324.4]
  assign synchronize = RetimeWrapper_io_out; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  assign _T_122 = done_0_io_output == 1'h0; // @[Controllers.scala 128:33:@371.4]
  assign _T_124 = io_ctrDone == 1'h0; // @[Controllers.scala 128:54:@372.4]
  assign _T_125 = _T_122 & _T_124; // @[Controllers.scala 128:52:@373.4]
  assign _T_126 = _T_125 & io_enable; // @[Controllers.scala 128:66:@374.4]
  assign _T_128 = ~ iterDone_0_io_output; // @[Controllers.scala 128:98:@376.4]
  assign _T_129 = _T_126 & _T_128; // @[Controllers.scala 128:96:@377.4]
  assign _T_131 = io_doneIn_0 == 1'h0; // @[Controllers.scala 128:123:@378.4]
  assign _T_133 = io_doneIn_0 | io_rst; // @[Controllers.scala 129:48:@381.4]
  assign _T_138 = synchronize == 1'h0; // @[Controllers.scala 130:52:@386.4]
  assign _T_139 = io_doneIn_0 & _T_138; // @[Controllers.scala 130:50:@387.4]
  assign _T_147 = finished == 1'h0; // @[Controllers.scala 130:129:@393.4]
  assign _T_150 = io_rst == 1'h0; // @[Controllers.scala 131:45:@396.4]
  assign _T_154 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@402.4]
  assign _T_156 = _T_154 & _T_128; // @[Controllers.scala 213:90:@404.4]
  assign _T_158 = ~ done_0_io_output; // @[Controllers.scala 213:132:@406.4]
  assign _T_159 = _T_156 & _T_158; // @[Controllers.scala 213:130:@407.4]
  assign _T_160 = ~ io_ctrDone; // @[Controllers.scala 213:156:@408.4]
  assign io_done = RetimeWrapper_2_io_out; // @[Controllers.scala 245:13:@440.4]
  assign io_ctrInc = io_doneIn_0; // @[Controllers.scala 122:17:@356.4]
  assign io_enableOut_0 = _T_159 & _T_160; // @[Controllers.scala 213:55:@410.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@401.4]
  assign active_0_clock = clock; // @[:@319.4]
  assign active_0_reset = reset; // @[:@320.4]
  assign active_0_io_input_set = _T_129 & _T_131; // @[Controllers.scala 128:30:@380.4]
  assign active_0_io_input_reset = _T_133 | done_0_io_output; // @[Controllers.scala 129:32:@385.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@326.4]
  assign done_0_clock = clock; // @[:@322.4]
  assign done_0_reset = reset; // @[:@323.4]
  assign done_0_io_input_set = io_ctrDone & _T_150; // @[Controllers.scala 131:28:@399.4]
  assign done_0_io_input_reset = io_rst | done_0_io_output; // @[Controllers.scala 86:33:@336.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@327.4]
  assign iterDone_0_clock = clock; // @[:@339.4]
  assign iterDone_0_reset = reset; // @[:@340.4]
  assign iterDone_0_io_input_set = _T_139 & _T_147; // @[Controllers.scala 130:32:@395.4]
  assign iterDone_0_io_input_reset = synchronize | io_rst; // @[Controllers.scala 92:37:@350.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@341.4]
  assign RetimeWrapper_clock = clock; // @[:@358.4]
  assign RetimeWrapper_reset = reset; // @[:@359.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@361.4]
  assign RetimeWrapper_io_in = io_doneIn_0; // @[package.scala 94:16:@360.4]
  assign RetimeWrapper_1_clock = clock; // @[:@417.4]
  assign RetimeWrapper_1_reset = reset; // @[:@418.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@420.4]
  assign RetimeWrapper_1_io_in = done_0_io_output & _T_166; // @[package.scala 94:16:@419.4]
  assign RetimeWrapper_2_clock = clock; // @[:@434.4]
  assign RetimeWrapper_2_reset = reset; // @[:@435.4]
  assign RetimeWrapper_2_io_flow = io_enable; // @[package.scala 95:18:@437.4]
  assign RetimeWrapper_2_io_in = done_0_io_output & _T_180; // @[package.scala 94:16:@436.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_166 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_180 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_166 <= 1'h0;
    end else begin
      _T_166 <= _T_122;
    end
    if (reset) begin
      _T_180 <= 1'h0;
    end else begin
      _T_180 <= _T_122;
    end
  end
endmodule
module x493_outr_UnitPipe_sm( // @[:@2389.2]
  input   clock, // @[:@2390.4]
  input   reset, // @[:@2391.4]
  input   io_enable, // @[:@2392.4]
  output  io_done, // @[:@2392.4]
  input   io_parentAck, // @[:@2392.4]
  input   io_doneIn_0, // @[:@2392.4]
  output  io_enableOut_0, // @[:@2392.4]
  output  io_childAck_0, // @[:@2392.4]
  input   io_ctrCopyDone_0 // @[:@2392.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@2395.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@2395.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@2395.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@2395.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@2395.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@2395.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@2398.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@2398.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@2398.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@2398.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@2398.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@2398.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@2415.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@2415.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@2415.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@2415.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@2415.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@2415.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@2446.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@2446.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@2446.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@2446.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@2446.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@2460.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@2460.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@2460.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@2460.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@2460.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@2478.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@2478.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@2478.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@2478.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@2478.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@2515.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@2515.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@2515.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@2515.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@2515.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@2532.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@2532.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@2532.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@2532.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@2532.4]
  wire  _T_105; // @[Controllers.scala 165:35:@2430.4]
  wire  _T_107; // @[Controllers.scala 165:60:@2431.4]
  wire  _T_108; // @[Controllers.scala 165:58:@2432.4]
  wire  _T_110; // @[Controllers.scala 165:76:@2433.4]
  wire  _T_111; // @[Controllers.scala 165:74:@2434.4]
  wire  _T_115; // @[Controllers.scala 165:109:@2437.4]
  wire  _T_118; // @[Controllers.scala 165:141:@2439.4]
  wire  _T_126; // @[package.scala 96:25:@2451.4 package.scala 96:25:@2452.4]
  wire  _T_130; // @[Controllers.scala 167:54:@2454.4]
  wire  _T_131; // @[Controllers.scala 167:52:@2455.4]
  wire  _T_138; // @[package.scala 96:25:@2465.4 package.scala 96:25:@2466.4]
  wire  _T_156; // @[package.scala 96:25:@2483.4 package.scala 96:25:@2484.4]
  wire  _T_160; // @[Controllers.scala 169:67:@2486.4]
  wire  _T_161; // @[Controllers.scala 169:86:@2487.4]
  wire  _T_174; // @[Controllers.scala 213:68:@2501.4]
  wire  _T_176; // @[Controllers.scala 213:90:@2503.4]
  wire  _T_178; // @[Controllers.scala 213:132:@2505.4]
  reg  _T_186; // @[package.scala 48:56:@2511.4]
  reg [31:0] _RAND_0;
  wire  _T_187; // @[package.scala 100:41:@2513.4]
  reg  _T_200; // @[package.scala 48:56:@2529.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@2395.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@2398.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@2415.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@2446.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@2460.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@2478.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@2515.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@2532.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_105 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@2430.4]
  assign _T_107 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@2431.4]
  assign _T_108 = _T_105 & _T_107; // @[Controllers.scala 165:58:@2432.4]
  assign _T_110 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@2433.4]
  assign _T_111 = _T_108 & _T_110; // @[Controllers.scala 165:74:@2434.4]
  assign _T_115 = _T_111 & io_enable; // @[Controllers.scala 165:109:@2437.4]
  assign _T_118 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@2439.4]
  assign _T_126 = RetimeWrapper_io_out; // @[package.scala 96:25:@2451.4 package.scala 96:25:@2452.4]
  assign _T_130 = _T_126 == 1'h0; // @[Controllers.scala 167:54:@2454.4]
  assign _T_131 = io_doneIn_0 | _T_130; // @[Controllers.scala 167:52:@2455.4]
  assign _T_138 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@2465.4 package.scala 96:25:@2466.4]
  assign _T_156 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@2483.4 package.scala 96:25:@2484.4]
  assign _T_160 = _T_156 == 1'h0; // @[Controllers.scala 169:67:@2486.4]
  assign _T_161 = _T_160 & io_enable; // @[Controllers.scala 169:86:@2487.4]
  assign _T_174 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@2501.4]
  assign _T_176 = _T_174 & _T_105; // @[Controllers.scala 213:90:@2503.4]
  assign _T_178 = ~ done_0_io_output; // @[Controllers.scala 213:132:@2505.4]
  assign _T_187 = done_0_io_output & _T_186; // @[package.scala 100:41:@2513.4]
  assign io_done = RetimeWrapper_4_io_out; // @[Controllers.scala 245:13:@2539.4]
  assign io_enableOut_0 = _T_176 & _T_178; // @[Controllers.scala 213:55:@2509.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@2500.4]
  assign active_0_clock = clock; // @[:@2396.4]
  assign active_0_reset = reset; // @[:@2397.4]
  assign active_0_io_input_set = _T_115 & _T_118; // @[Controllers.scala 165:32:@2441.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@2445.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@2403.4]
  assign done_0_clock = clock; // @[:@2399.4]
  assign done_0_reset = reset; // @[:@2400.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_161; // @[Controllers.scala 169:30:@2491.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@2413.4 Controllers.scala 170:32:@2498.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@2404.4]
  assign iterDone_0_clock = clock; // @[:@2416.4]
  assign iterDone_0_reset = reset; // @[:@2417.4]
  assign iterDone_0_io_input_set = _T_131 & io_enable; // @[Controllers.scala 167:34:@2459.4]
  assign iterDone_0_io_input_reset = _T_138 | io_parentAck; // @[Controllers.scala 92:37:@2427.4 Controllers.scala 168:36:@2475.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@2418.4]
  assign RetimeWrapper_clock = clock; // @[:@2447.4]
  assign RetimeWrapper_reset = reset; // @[:@2448.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@2450.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@2449.4]
  assign RetimeWrapper_1_clock = clock; // @[:@2461.4]
  assign RetimeWrapper_1_reset = reset; // @[:@2462.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@2464.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@2463.4]
  assign RetimeWrapper_2_clock = clock; // @[:@2479.4]
  assign RetimeWrapper_2_reset = reset; // @[:@2480.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@2482.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@2481.4]
  assign RetimeWrapper_3_clock = clock; // @[:@2516.4]
  assign RetimeWrapper_3_reset = reset; // @[:@2517.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@2519.4]
  assign RetimeWrapper_3_io_in = _T_187 | io_parentAck; // @[package.scala 94:16:@2518.4]
  assign RetimeWrapper_4_clock = clock; // @[:@2533.4]
  assign RetimeWrapper_4_reset = reset; // @[:@2534.4]
  assign RetimeWrapper_4_io_flow = io_enable; // @[package.scala 95:18:@2536.4]
  assign RetimeWrapper_4_io_in = done_0_io_output & _T_200; // @[package.scala 94:16:@2535.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_186 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_200 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_186 <= 1'h0;
    end else begin
      _T_186 <= _T_110;
    end
    if (reset) begin
      _T_200 <= 1'h0;
    end else begin
      _T_200 <= _T_110;
    end
  end
endmodule
module SingleCounter_1( // @[:@2659.2]
  input         clock, // @[:@2660.4]
  input         reset, // @[:@2661.4]
  input         io_input_reset, // @[:@2662.4]
  input         io_input_enable, // @[:@2662.4]
  output [31:0] io_output_count_0, // @[:@2662.4]
  output        io_output_oobs_0, // @[:@2662.4]
  output        io_output_done, // @[:@2662.4]
  output        io_output_saturated // @[:@2662.4]
);
  wire  bases_0_clock; // @[Counter.scala 253:53:@2675.4]
  wire  bases_0_reset; // @[Counter.scala 253:53:@2675.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 253:53:@2675.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 253:53:@2675.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 253:53:@2675.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 253:53:@2675.4]
  wire  SRFF_clock; // @[Counter.scala 255:22:@2691.4]
  wire  SRFF_reset; // @[Counter.scala 255:22:@2691.4]
  wire  SRFF_io_input_set; // @[Counter.scala 255:22:@2691.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 255:22:@2691.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 255:22:@2691.4]
  wire  SRFF_io_output; // @[Counter.scala 255:22:@2691.4]
  wire  _T_36; // @[Counter.scala 256:45:@2694.4]
  wire [31:0] _T_48; // @[Counter.scala 279:52:@2719.4]
  wire [32:0] _T_50; // @[Counter.scala 283:33:@2720.4]
  wire [31:0] _T_51; // @[Counter.scala 283:33:@2721.4]
  wire [31:0] _T_52; // @[Counter.scala 283:33:@2722.4]
  wire  _T_57; // @[Counter.scala 285:18:@2724.4]
  wire [31:0] _T_68; // @[Counter.scala 291:115:@2732.4]
  wire [31:0] _T_71; // @[Counter.scala 291:152:@2735.4]
  wire [31:0] _T_72; // @[Counter.scala 291:74:@2736.4]
  wire  _T_75; // @[Counter.scala 314:102:@2740.4]
  wire  _T_77; // @[Counter.scala 314:130:@2741.4]
  FF bases_0 ( // @[Counter.scala 253:53:@2675.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 255:22:@2691.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 256:45:@2694.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 279:52:@2719.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@2720.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@2721.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 283:33:@2722.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh4); // @[Counter.scala 285:18:@2724.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 291:115:@2732.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 291:152:@2735.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 291:74:@2736.4]
  assign _T_75 = $signed(_T_48) < $signed(32'sh0); // @[Counter.scala 314:102:@2740.4]
  assign _T_77 = $signed(_T_48) >= $signed(32'sh4); // @[Counter.scala 314:130:@2741.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 296:28:@2739.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 314:60:@2743.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 325:20:@2745.4]
  assign io_output_saturated = $signed(_T_52) >= $signed(32'sh4); // @[Counter.scala 332:25:@2748.4]
  assign bases_0_clock = clock; // @[:@2676.4]
  assign bases_0_reset = reset; // @[:@2677.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 291:31:@2738.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 273:27:@2717.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 276:29:@2718.4]
  assign SRFF_clock = clock; // @[:@2692.4]
  assign SRFF_reset = reset; // @[:@2693.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 256:23:@2696.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 257:25:@2698.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 258:30:@2699.4]
endmodule
module SingleCounter_2( // @[:@2788.2]
  input         clock, // @[:@2789.4]
  input         reset, // @[:@2790.4]
  input         io_setup_saturate, // @[:@2791.4]
  input         io_input_reset, // @[:@2791.4]
  input         io_input_enable, // @[:@2791.4]
  output [31:0] io_output_count_0, // @[:@2791.4]
  output        io_output_oobs_0, // @[:@2791.4]
  output        io_output_done // @[:@2791.4]
);
  wire  bases_0_clock; // @[Counter.scala 253:53:@2804.4]
  wire  bases_0_reset; // @[Counter.scala 253:53:@2804.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 253:53:@2804.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 253:53:@2804.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 253:53:@2804.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 253:53:@2804.4]
  wire  SRFF_clock; // @[Counter.scala 255:22:@2820.4]
  wire  SRFF_reset; // @[Counter.scala 255:22:@2820.4]
  wire  SRFF_io_input_set; // @[Counter.scala 255:22:@2820.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 255:22:@2820.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 255:22:@2820.4]
  wire  SRFF_io_output; // @[Counter.scala 255:22:@2820.4]
  wire  _T_36; // @[Counter.scala 256:45:@2823.4]
  wire [31:0] _T_48; // @[Counter.scala 279:52:@2848.4]
  wire [32:0] _T_50; // @[Counter.scala 283:33:@2849.4]
  wire [31:0] _T_51; // @[Counter.scala 283:33:@2850.4]
  wire [31:0] _T_52; // @[Counter.scala 283:33:@2851.4]
  wire  _T_57; // @[Counter.scala 285:18:@2853.4]
  wire [31:0] _T_68; // @[Counter.scala 291:115:@2861.4]
  wire [31:0] _T_70; // @[Counter.scala 291:85:@2863.4]
  wire [31:0] _T_71; // @[Counter.scala 291:152:@2864.4]
  wire [31:0] _T_72; // @[Counter.scala 291:74:@2865.4]
  wire  _T_75; // @[Counter.scala 314:102:@2869.4]
  wire  _T_77; // @[Counter.scala 314:130:@2870.4]
  FF bases_0 ( // @[Counter.scala 253:53:@2804.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 255:22:@2820.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 256:45:@2823.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 279:52:@2848.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh2); // @[Counter.scala 283:33:@2849.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh2); // @[Counter.scala 283:33:@2850.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 283:33:@2851.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh4); // @[Counter.scala 285:18:@2853.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 291:115:@2861.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 32'h0; // @[Counter.scala 291:85:@2863.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 291:152:@2864.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 291:74:@2865.4]
  assign _T_75 = $signed(_T_48) < $signed(32'sh0); // @[Counter.scala 314:102:@2869.4]
  assign _T_77 = $signed(_T_48) >= $signed(32'sh4); // @[Counter.scala 314:130:@2870.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 296:28:@2868.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 314:60:@2872.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 325:20:@2874.4]
  assign bases_0_clock = clock; // @[:@2805.4]
  assign bases_0_reset = reset; // @[:@2806.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 291:31:@2867.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 273:27:@2846.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 276:29:@2847.4]
  assign SRFF_clock = clock; // @[:@2821.4]
  assign SRFF_reset = reset; // @[:@2822.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 256:23:@2825.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 257:25:@2827.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 258:30:@2828.4]
endmodule
module x283_ctrchain( // @[:@2879.2]
  input         clock, // @[:@2880.4]
  input         reset, // @[:@2881.4]
  input         io_input_reset, // @[:@2882.4]
  input         io_input_enable, // @[:@2882.4]
  output [31:0] io_output_counts_1, // @[:@2882.4]
  output [31:0] io_output_counts_0, // @[:@2882.4]
  output        io_output_oobs_0, // @[:@2882.4]
  output        io_output_oobs_1, // @[:@2882.4]
  output        io_output_done // @[:@2882.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_reset; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 505:46:@2884.4]
  wire [31:0] ctrs_0_io_output_count_0; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_io_output_saturated; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_1_clock; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_reset; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_io_setup_saturate; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_io_input_reset; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_io_input_enable; // @[Counter.scala 505:46:@2887.4]
  wire [31:0] ctrs_1_io_output_count_0; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_io_output_oobs_0; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_io_output_done; // @[Counter.scala 505:46:@2887.4]
  wire  isDone; // @[Counter.scala 533:51:@2904.4]
  reg  wasDone; // @[Counter.scala 534:24:@2905.4]
  reg [31:0] _RAND_0;
  wire  _T_64; // @[Counter.scala 538:69:@2913.4]
  wire  _T_66; // @[Counter.scala 538:80:@2914.4]
  reg  doneLatch; // @[Counter.scala 542:26:@2919.4]
  reg [31:0] _RAND_1;
  wire  _T_73; // @[Counter.scala 543:48:@2920.4]
  wire  _T_74; // @[Counter.scala 543:19:@2921.4]
  SingleCounter_1 ctrs_0 ( // @[Counter.scala 505:46:@2884.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done),
    .io_output_saturated(ctrs_0_io_output_saturated)
  );
  SingleCounter_2 ctrs_1 ( // @[Counter.scala 505:46:@2887.4]
    .clock(ctrs_1_clock),
    .reset(ctrs_1_reset),
    .io_setup_saturate(ctrs_1_io_setup_saturate),
    .io_input_reset(ctrs_1_io_input_reset),
    .io_input_enable(ctrs_1_io_input_enable),
    .io_output_count_0(ctrs_1_io_output_count_0),
    .io_output_oobs_0(ctrs_1_io_output_oobs_0),
    .io_output_done(ctrs_1_io_output_done)
  );
  assign isDone = ctrs_0_io_output_done & ctrs_1_io_output_done; // @[Counter.scala 533:51:@2904.4]
  assign _T_64 = io_input_enable & isDone; // @[Counter.scala 538:69:@2913.4]
  assign _T_66 = wasDone == 1'h0; // @[Counter.scala 538:80:@2914.4]
  assign _T_73 = isDone ? 1'h1 : doneLatch; // @[Counter.scala 543:48:@2920.4]
  assign _T_74 = io_input_reset ? 1'h0 : _T_73; // @[Counter.scala 543:19:@2921.4]
  assign io_output_counts_1 = ctrs_1_io_output_count_0; // @[Counter.scala 549:32:@2926.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 549:32:@2923.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 550:30:@2925.4]
  assign io_output_oobs_1 = ctrs_1_io_output_oobs_0 | doneLatch; // @[Counter.scala 550:30:@2928.4]
  assign io_output_done = _T_64 & _T_66; // @[Counter.scala 538:18:@2916.4]
  assign ctrs_0_clock = clock; // @[:@2885.4]
  assign ctrs_0_reset = reset; // @[:@2886.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 512:24:@2893.4]
  assign ctrs_0_io_input_enable = ctrs_1_io_output_done & io_input_enable; // @[Counter.scala 518:29:@2900.4]
  assign ctrs_1_clock = clock; // @[:@2888.4]
  assign ctrs_1_reset = reset; // @[:@2889.4]
  assign ctrs_1_io_setup_saturate = ctrs_0_io_output_saturated; // @[Counter.scala 524:31:@2903.4]
  assign ctrs_1_io_input_reset = io_input_reset; // @[Counter.scala 512:24:@2897.4]
  assign ctrs_1_io_input_enable = io_input_enable; // @[Counter.scala 516:33:@2898.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= isDone;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (isDone) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module RetimeWrapper_12( // @[:@2968.2]
  input   clock, // @[:@2969.4]
  input   reset, // @[:@2970.4]
  input   io_flow, // @[:@2971.4]
  input   io_in, // @[:@2971.4]
  output  io_out // @[:@2971.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(37)) sr ( // @[RetimeShiftRegister.scala 15:20:@2973.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@2986.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@2985.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@2984.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@2983.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@2982.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@2980.4]
endmodule
module RetimeWrapper_16( // @[:@3096.2]
  input   clock, // @[:@3097.4]
  input   reset, // @[:@3098.4]
  input   io_flow, // @[:@3099.4]
  input   io_in, // @[:@3099.4]
  output  io_out // @[:@3099.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(36)) sr ( // @[RetimeShiftRegister.scala 15:20:@3101.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3114.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3113.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3112.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3111.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3110.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3108.4]
endmodule
module x492_inr_Foreach_SAMPLER_BOX_sm( // @[:@3116.2]
  input   clock, // @[:@3117.4]
  input   reset, // @[:@3118.4]
  input   io_enable, // @[:@3119.4]
  output  io_done, // @[:@3119.4]
  output  io_doneLatch, // @[:@3119.4]
  input   io_ctrDone, // @[:@3119.4]
  output  io_datapathEn, // @[:@3119.4]
  output  io_ctrInc, // @[:@3119.4]
  output  io_ctrRst, // @[:@3119.4]
  input   io_parentAck, // @[:@3119.4]
  input   io_backpressure, // @[:@3119.4]
  input   io_break // @[:@3119.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@3121.4]
  wire  active_reset; // @[Controllers.scala 261:22:@3121.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@3121.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@3121.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@3121.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@3121.4]
  wire  done_clock; // @[Controllers.scala 262:20:@3124.4]
  wire  done_reset; // @[Controllers.scala 262:20:@3124.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@3124.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@3124.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@3124.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@3124.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3158.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3158.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3158.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@3158.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@3158.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@3180.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@3180.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@3180.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@3180.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@3180.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@3192.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@3192.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@3192.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@3192.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@3192.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@3200.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@3200.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@3200.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@3200.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@3200.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@3216.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@3216.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@3216.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@3216.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@3216.4]
  wire  _T_80; // @[Controllers.scala 264:48:@3129.4]
  wire  _T_81; // @[Controllers.scala 264:46:@3130.4]
  wire  _T_82; // @[Controllers.scala 264:62:@3131.4]
  wire  _T_83; // @[Controllers.scala 264:60:@3132.4]
  wire  _T_100; // @[package.scala 100:49:@3149.4]
  reg  _T_103; // @[package.scala 48:56:@3150.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@3163.4 package.scala 96:25:@3164.4]
  wire  _T_110; // @[package.scala 100:49:@3165.4]
  reg  _T_113; // @[package.scala 48:56:@3166.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@3168.4]
  wire  _T_118; // @[Controllers.scala 283:41:@3173.4]
  wire  _T_119; // @[Controllers.scala 283:59:@3174.4]
  wire  _T_121; // @[Controllers.scala 284:37:@3177.4]
  wire  _T_124; // @[package.scala 96:25:@3185.4 package.scala 96:25:@3186.4]
  wire  _T_126; // @[package.scala 100:49:@3187.4]
  reg  _T_129; // @[package.scala 48:56:@3188.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@3210.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@3212.4]
  reg  _T_153; // @[package.scala 48:56:@3213.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@3221.4 package.scala 96:25:@3222.4]
  wire  _T_158; // @[Controllers.scala 292:61:@3223.4]
  wire  _T_159; // @[Controllers.scala 292:24:@3224.4]
  SRFF active ( // @[Controllers.scala 261:22:@3121.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@3124.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_12 RetimeWrapper ( // @[package.scala 93:22:@3158.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_12 RetimeWrapper_1 ( // @[package.scala 93:22:@3180.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@3192.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@3200.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_16 RetimeWrapper_4 ( // @[package.scala 93:22:@3216.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@3129.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@3130.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@3131.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@3132.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@3149.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@3163.4 package.scala 96:25:@3164.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@3165.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@3168.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@3173.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@3174.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@3177.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@3185.4 package.scala 96:25:@3186.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@3187.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@3212.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@3221.4 package.scala 96:25:@3222.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@3223.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@3224.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@3191.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@3226.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@3176.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@3179.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@3171.4]
  assign active_clock = clock; // @[:@3122.4]
  assign active_reset = reset; // @[:@3123.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@3134.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@3138.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@3139.4]
  assign done_clock = clock; // @[:@3125.4]
  assign done_reset = reset; // @[:@3126.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@3154.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@3147.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@3148.4]
  assign RetimeWrapper_clock = clock; // @[:@3159.4]
  assign RetimeWrapper_reset = reset; // @[:@3160.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@3162.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@3161.4]
  assign RetimeWrapper_1_clock = clock; // @[:@3181.4]
  assign RetimeWrapper_1_reset = reset; // @[:@3182.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@3184.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@3183.4]
  assign RetimeWrapper_2_clock = clock; // @[:@3193.4]
  assign RetimeWrapper_2_reset = reset; // @[:@3194.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@3196.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@3195.4]
  assign RetimeWrapper_3_clock = clock; // @[:@3201.4]
  assign RetimeWrapper_3_reset = reset; // @[:@3202.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@3204.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@3203.4]
  assign RetimeWrapper_4_clock = clock; // @[:@3217.4]
  assign RetimeWrapper_4_reset = reset; // @[:@3218.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@3220.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@3219.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module SimBlackBoxesfix2fixBox( // @[:@3332.2]
  input  [31:0] io_a, // @[:@3335.4]
  output [31:0] io_b // @[:@3335.4]
);
  assign io_b = io_a; // @[SimBlackBoxes.scala 99:40:@3345.4]
endmodule
module _( // @[:@3347.2]
  input  [31:0] io_b, // @[:@3350.4]
  output [31:0] io_result // @[:@3350.4]
);
  wire [31:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@3355.4]
  wire [31:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@3355.4]
  SimBlackBoxesfix2fixBox SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@3355.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@3368.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@3363.4]
endmodule
module RetimeWrapper_21( // @[:@3452.2]
  input        clock, // @[:@3453.4]
  input        reset, // @[:@3454.4]
  input        io_flow, // @[:@3455.4]
  input  [7:0] io_in, // @[:@3455.4]
  output [7:0] io_out // @[:@3455.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@3457.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3470.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3469.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@3468.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3467.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3466.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3464.4]
endmodule
module Mem1D_4( // @[:@3472.2]
  input        clock, // @[:@3473.4]
  input        reset, // @[:@3474.4]
  input        io_r_ofs_0, // @[:@3475.4]
  input        io_r_backpressure, // @[:@3475.4]
  input        io_w_ofs_0, // @[:@3475.4]
  input  [7:0] io_w_data_0, // @[:@3475.4]
  input        io_w_en_0, // @[:@3475.4]
  output [7:0] io_output // @[:@3475.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3485.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3485.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3485.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@3485.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@3485.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@3494.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@3494.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@3494.4]
  wire [7:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@3494.4]
  wire [7:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@3494.4]
  reg [7:0] _T_127; // @[MemPrimitives.scala 560:26:@3479.4]
  reg [31:0] _RAND_0;
  wire  _T_130; // @[MemPrimitives.scala 561:61:@3481.4]
  wire  _T_131; // @[MemPrimitives.scala 561:44:@3482.4]
  wire [7:0] _T_132; // @[MemPrimitives.scala 561:19:@3483.4]
  wire  _T_135; // @[package.scala 96:25:@3490.4 package.scala 96:25:@3491.4]
  wire  _T_137; // @[Mux.scala 46:19:@3492.4]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@3485.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_1 ( // @[package.scala 93:22:@3494.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign _T_130 = io_w_ofs_0 == 1'h0; // @[MemPrimitives.scala 561:61:@3481.4]
  assign _T_131 = io_w_en_0 & _T_130; // @[MemPrimitives.scala 561:44:@3482.4]
  assign _T_132 = _T_131 ? io_w_data_0 : _T_127; // @[MemPrimitives.scala 561:19:@3483.4]
  assign _T_135 = RetimeWrapper_io_out; // @[package.scala 96:25:@3490.4 package.scala 96:25:@3491.4]
  assign _T_137 = 1'h0 == _T_135; // @[Mux.scala 46:19:@3492.4]
  assign io_output = RetimeWrapper_1_io_out; // @[MemPrimitives.scala 565:17:@3501.4]
  assign RetimeWrapper_clock = clock; // @[:@3486.4]
  assign RetimeWrapper_reset = reset; // @[:@3487.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@3489.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@3488.4]
  assign RetimeWrapper_1_clock = clock; // @[:@3495.4]
  assign RetimeWrapper_1_reset = reset; // @[:@3496.4]
  assign RetimeWrapper_1_io_flow = io_r_backpressure; // @[package.scala 95:18:@3498.4]
  assign RetimeWrapper_1_io_in = _T_137 ? _T_127 : 8'h0; // @[package.scala 94:16:@3497.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_127 = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_127 <= 8'h0;
    end else begin
      if (_T_131) begin
        _T_127 <= io_w_data_0;
      end
    end
  end
endmodule
module StickySelects( // @[:@4928.2]
  input   clock, // @[:@4929.4]
  input   reset, // @[:@4930.4]
  input   io_ins_0, // @[:@4931.4]
  input   io_ins_1, // @[:@4931.4]
  input   io_ins_2, // @[:@4931.4]
  input   io_ins_3, // @[:@4931.4]
  input   io_ins_4, // @[:@4931.4]
  input   io_ins_5, // @[:@4931.4]
  output  io_outs_0, // @[:@4931.4]
  output  io_outs_1, // @[:@4931.4]
  output  io_outs_2, // @[:@4931.4]
  output  io_outs_3, // @[:@4931.4]
  output  io_outs_4, // @[:@4931.4]
  output  io_outs_5 // @[:@4931.4]
);
  reg  _T_19; // @[StickySelects.scala 21:22:@4933.4]
  reg [31:0] _RAND_0;
  wire  _T_20; // @[StickySelects.scala 22:54:@4934.4]
  wire  _T_21; // @[StickySelects.scala 22:54:@4935.4]
  wire  _T_22; // @[StickySelects.scala 22:54:@4936.4]
  wire  _T_23; // @[StickySelects.scala 22:54:@4937.4]
  wire  _T_25; // @[StickySelects.scala 24:52:@4938.4]
  wire  _T_26; // @[StickySelects.scala 24:21:@4939.4]
  reg  _T_29; // @[StickySelects.scala 21:22:@4941.4]
  reg [31:0] _RAND_1;
  wire  _T_30; // @[StickySelects.scala 22:54:@4942.4]
  wire  _T_31; // @[StickySelects.scala 22:54:@4943.4]
  wire  _T_32; // @[StickySelects.scala 22:54:@4944.4]
  wire  _T_33; // @[StickySelects.scala 22:54:@4945.4]
  wire  _T_35; // @[StickySelects.scala 24:52:@4946.4]
  wire  _T_36; // @[StickySelects.scala 24:21:@4947.4]
  reg  _T_39; // @[StickySelects.scala 21:22:@4949.4]
  reg [31:0] _RAND_2;
  wire  _T_40; // @[StickySelects.scala 22:54:@4950.4]
  wire  _T_41; // @[StickySelects.scala 22:54:@4951.4]
  wire  _T_42; // @[StickySelects.scala 22:54:@4952.4]
  wire  _T_43; // @[StickySelects.scala 22:54:@4953.4]
  wire  _T_45; // @[StickySelects.scala 24:52:@4954.4]
  wire  _T_46; // @[StickySelects.scala 24:21:@4955.4]
  reg  _T_49; // @[StickySelects.scala 21:22:@4957.4]
  reg [31:0] _RAND_3;
  wire  _T_51; // @[StickySelects.scala 22:54:@4959.4]
  wire  _T_52; // @[StickySelects.scala 22:54:@4960.4]
  wire  _T_53; // @[StickySelects.scala 22:54:@4961.4]
  wire  _T_55; // @[StickySelects.scala 24:52:@4962.4]
  wire  _T_56; // @[StickySelects.scala 24:21:@4963.4]
  reg  _T_59; // @[StickySelects.scala 21:22:@4965.4]
  reg [31:0] _RAND_4;
  wire  _T_62; // @[StickySelects.scala 22:54:@4968.4]
  wire  _T_63; // @[StickySelects.scala 22:54:@4969.4]
  wire  _T_65; // @[StickySelects.scala 24:52:@4970.4]
  wire  _T_66; // @[StickySelects.scala 24:21:@4971.4]
  reg  _T_69; // @[StickySelects.scala 21:22:@4973.4]
  reg [31:0] _RAND_5;
  wire  _T_73; // @[StickySelects.scala 22:54:@4977.4]
  wire  _T_75; // @[StickySelects.scala 24:52:@4978.4]
  wire  _T_76; // @[StickySelects.scala 24:21:@4979.4]
  assign _T_20 = io_ins_1 | io_ins_2; // @[StickySelects.scala 22:54:@4934.4]
  assign _T_21 = _T_20 | io_ins_3; // @[StickySelects.scala 22:54:@4935.4]
  assign _T_22 = _T_21 | io_ins_4; // @[StickySelects.scala 22:54:@4936.4]
  assign _T_23 = _T_22 | io_ins_5; // @[StickySelects.scala 22:54:@4937.4]
  assign _T_25 = io_ins_0 | _T_19; // @[StickySelects.scala 24:52:@4938.4]
  assign _T_26 = _T_23 ? 1'h0 : _T_25; // @[StickySelects.scala 24:21:@4939.4]
  assign _T_30 = io_ins_0 | io_ins_2; // @[StickySelects.scala 22:54:@4942.4]
  assign _T_31 = _T_30 | io_ins_3; // @[StickySelects.scala 22:54:@4943.4]
  assign _T_32 = _T_31 | io_ins_4; // @[StickySelects.scala 22:54:@4944.4]
  assign _T_33 = _T_32 | io_ins_5; // @[StickySelects.scala 22:54:@4945.4]
  assign _T_35 = io_ins_1 | _T_29; // @[StickySelects.scala 24:52:@4946.4]
  assign _T_36 = _T_33 ? 1'h0 : _T_35; // @[StickySelects.scala 24:21:@4947.4]
  assign _T_40 = io_ins_0 | io_ins_1; // @[StickySelects.scala 22:54:@4950.4]
  assign _T_41 = _T_40 | io_ins_3; // @[StickySelects.scala 22:54:@4951.4]
  assign _T_42 = _T_41 | io_ins_4; // @[StickySelects.scala 22:54:@4952.4]
  assign _T_43 = _T_42 | io_ins_5; // @[StickySelects.scala 22:54:@4953.4]
  assign _T_45 = io_ins_2 | _T_39; // @[StickySelects.scala 24:52:@4954.4]
  assign _T_46 = _T_43 ? 1'h0 : _T_45; // @[StickySelects.scala 24:21:@4955.4]
  assign _T_51 = _T_40 | io_ins_2; // @[StickySelects.scala 22:54:@4959.4]
  assign _T_52 = _T_51 | io_ins_4; // @[StickySelects.scala 22:54:@4960.4]
  assign _T_53 = _T_52 | io_ins_5; // @[StickySelects.scala 22:54:@4961.4]
  assign _T_55 = io_ins_3 | _T_49; // @[StickySelects.scala 24:52:@4962.4]
  assign _T_56 = _T_53 ? 1'h0 : _T_55; // @[StickySelects.scala 24:21:@4963.4]
  assign _T_62 = _T_51 | io_ins_3; // @[StickySelects.scala 22:54:@4968.4]
  assign _T_63 = _T_62 | io_ins_5; // @[StickySelects.scala 22:54:@4969.4]
  assign _T_65 = io_ins_4 | _T_59; // @[StickySelects.scala 24:52:@4970.4]
  assign _T_66 = _T_63 ? 1'h0 : _T_65; // @[StickySelects.scala 24:21:@4971.4]
  assign _T_73 = _T_62 | io_ins_4; // @[StickySelects.scala 22:54:@4977.4]
  assign _T_75 = io_ins_5 | _T_69; // @[StickySelects.scala 24:52:@4978.4]
  assign _T_76 = _T_73 ? 1'h0 : _T_75; // @[StickySelects.scala 24:21:@4979.4]
  assign io_outs_0 = _T_23 ? 1'h0 : _T_25; // @[StickySelects.scala 28:52:@4981.4]
  assign io_outs_1 = _T_33 ? 1'h0 : _T_35; // @[StickySelects.scala 28:52:@4982.4]
  assign io_outs_2 = _T_43 ? 1'h0 : _T_45; // @[StickySelects.scala 28:52:@4983.4]
  assign io_outs_3 = _T_53 ? 1'h0 : _T_55; // @[StickySelects.scala 28:52:@4984.4]
  assign io_outs_4 = _T_63 ? 1'h0 : _T_65; // @[StickySelects.scala 28:52:@4985.4]
  assign io_outs_5 = _T_73 ? 1'h0 : _T_75; // @[StickySelects.scala 28:52:@4986.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_29 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_39 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_49 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_59 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_69 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (_T_23) begin
        _T_19 <= 1'h0;
      end else begin
        _T_19 <= _T_25;
      end
    end
    if (reset) begin
      _T_29 <= 1'h0;
    end else begin
      if (_T_33) begin
        _T_29 <= 1'h0;
      end else begin
        _T_29 <= _T_35;
      end
    end
    if (reset) begin
      _T_39 <= 1'h0;
    end else begin
      if (_T_43) begin
        _T_39 <= 1'h0;
      end else begin
        _T_39 <= _T_45;
      end
    end
    if (reset) begin
      _T_49 <= 1'h0;
    end else begin
      if (_T_53) begin
        _T_49 <= 1'h0;
      end else begin
        _T_49 <= _T_55;
      end
    end
    if (reset) begin
      _T_59 <= 1'h0;
    end else begin
      if (_T_63) begin
        _T_59 <= 1'h0;
      end else begin
        _T_59 <= _T_65;
      end
    end
    if (reset) begin
      _T_69 <= 1'h0;
    end else begin
      if (_T_73) begin
        _T_69 <= 1'h0;
      end else begin
        _T_69 <= _T_75;
      end
    end
  end
endmodule
module RetimeWrapper_52( // @[:@5900.2]
  input   clock, // @[:@5901.4]
  input   reset, // @[:@5902.4]
  input   io_flow, // @[:@5903.4]
  input   io_in, // @[:@5903.4]
  output  io_out // @[:@5903.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@5905.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@5905.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@5905.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@5905.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@5905.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@5905.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@5905.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@5918.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@5917.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@5916.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@5915.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@5914.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@5912.4]
endmodule
module x288_lb_0( // @[:@8960.2]
  input        clock, // @[:@8961.4]
  input        reset, // @[:@8962.4]
  input  [2:0] io_rPort_11_banks_1, // @[:@8963.4]
  input  [2:0] io_rPort_11_banks_0, // @[:@8963.4]
  input        io_rPort_11_ofs_0, // @[:@8963.4]
  input        io_rPort_11_en_0, // @[:@8963.4]
  input        io_rPort_11_backpressure, // @[:@8963.4]
  output [7:0] io_rPort_11_output_0, // @[:@8963.4]
  input  [2:0] io_rPort_10_banks_1, // @[:@8963.4]
  input  [2:0] io_rPort_10_banks_0, // @[:@8963.4]
  input        io_rPort_10_ofs_0, // @[:@8963.4]
  input        io_rPort_10_en_0, // @[:@8963.4]
  input        io_rPort_10_backpressure, // @[:@8963.4]
  output [7:0] io_rPort_10_output_0, // @[:@8963.4]
  input  [2:0] io_rPort_9_banks_1, // @[:@8963.4]
  input  [2:0] io_rPort_9_banks_0, // @[:@8963.4]
  input        io_rPort_9_ofs_0, // @[:@8963.4]
  input        io_rPort_9_en_0, // @[:@8963.4]
  input        io_rPort_9_backpressure, // @[:@8963.4]
  output [7:0] io_rPort_9_output_0, // @[:@8963.4]
  input  [2:0] io_rPort_8_banks_1, // @[:@8963.4]
  input  [2:0] io_rPort_8_banks_0, // @[:@8963.4]
  input        io_rPort_8_ofs_0, // @[:@8963.4]
  input        io_rPort_8_en_0, // @[:@8963.4]
  input        io_rPort_8_backpressure, // @[:@8963.4]
  output [7:0] io_rPort_8_output_0, // @[:@8963.4]
  input  [2:0] io_rPort_7_banks_1, // @[:@8963.4]
  input  [2:0] io_rPort_7_banks_0, // @[:@8963.4]
  input        io_rPort_7_ofs_0, // @[:@8963.4]
  input        io_rPort_7_en_0, // @[:@8963.4]
  input        io_rPort_7_backpressure, // @[:@8963.4]
  output [7:0] io_rPort_7_output_0, // @[:@8963.4]
  input  [2:0] io_rPort_6_banks_1, // @[:@8963.4]
  input  [2:0] io_rPort_6_banks_0, // @[:@8963.4]
  input        io_rPort_6_ofs_0, // @[:@8963.4]
  input        io_rPort_6_en_0, // @[:@8963.4]
  input        io_rPort_6_backpressure, // @[:@8963.4]
  output [7:0] io_rPort_6_output_0, // @[:@8963.4]
  input  [2:0] io_rPort_5_banks_1, // @[:@8963.4]
  input  [2:0] io_rPort_5_banks_0, // @[:@8963.4]
  input        io_rPort_5_ofs_0, // @[:@8963.4]
  input        io_rPort_5_en_0, // @[:@8963.4]
  input        io_rPort_5_backpressure, // @[:@8963.4]
  output [7:0] io_rPort_5_output_0, // @[:@8963.4]
  input  [2:0] io_rPort_4_banks_1, // @[:@8963.4]
  input  [2:0] io_rPort_4_banks_0, // @[:@8963.4]
  input        io_rPort_4_ofs_0, // @[:@8963.4]
  input        io_rPort_4_en_0, // @[:@8963.4]
  input        io_rPort_4_backpressure, // @[:@8963.4]
  output [7:0] io_rPort_4_output_0, // @[:@8963.4]
  input  [2:0] io_rPort_3_banks_1, // @[:@8963.4]
  input  [2:0] io_rPort_3_banks_0, // @[:@8963.4]
  input        io_rPort_3_ofs_0, // @[:@8963.4]
  input        io_rPort_3_en_0, // @[:@8963.4]
  input        io_rPort_3_backpressure, // @[:@8963.4]
  output [7:0] io_rPort_3_output_0, // @[:@8963.4]
  input  [2:0] io_rPort_2_banks_1, // @[:@8963.4]
  input  [2:0] io_rPort_2_banks_0, // @[:@8963.4]
  input        io_rPort_2_ofs_0, // @[:@8963.4]
  input        io_rPort_2_en_0, // @[:@8963.4]
  input        io_rPort_2_backpressure, // @[:@8963.4]
  output [7:0] io_rPort_2_output_0, // @[:@8963.4]
  input  [2:0] io_rPort_1_banks_1, // @[:@8963.4]
  input  [2:0] io_rPort_1_banks_0, // @[:@8963.4]
  input        io_rPort_1_ofs_0, // @[:@8963.4]
  input        io_rPort_1_en_0, // @[:@8963.4]
  input        io_rPort_1_backpressure, // @[:@8963.4]
  output [7:0] io_rPort_1_output_0, // @[:@8963.4]
  input  [2:0] io_rPort_0_banks_1, // @[:@8963.4]
  input  [2:0] io_rPort_0_banks_0, // @[:@8963.4]
  input        io_rPort_0_ofs_0, // @[:@8963.4]
  input        io_rPort_0_en_0, // @[:@8963.4]
  input        io_rPort_0_backpressure, // @[:@8963.4]
  output [7:0] io_rPort_0_output_0, // @[:@8963.4]
  input  [2:0] io_wPort_1_banks_1, // @[:@8963.4]
  input  [2:0] io_wPort_1_banks_0, // @[:@8963.4]
  input        io_wPort_1_ofs_0, // @[:@8963.4]
  input  [7:0] io_wPort_1_data_0, // @[:@8963.4]
  input        io_wPort_1_en_0, // @[:@8963.4]
  input  [2:0] io_wPort_0_banks_1, // @[:@8963.4]
  input  [2:0] io_wPort_0_banks_0, // @[:@8963.4]
  input        io_wPort_0_ofs_0, // @[:@8963.4]
  input  [7:0] io_wPort_0_data_0, // @[:@8963.4]
  input        io_wPort_0_en_0 // @[:@8963.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@9054.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@9054.4]
  wire  Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9054.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9054.4]
  wire  Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9054.4]
  wire [7:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@9054.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@9054.4]
  wire [7:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@9054.4]
  wire  Mem1D_1_clock; // @[MemPrimitives.scala 64:21:@9070.4]
  wire  Mem1D_1_reset; // @[MemPrimitives.scala 64:21:@9070.4]
  wire  Mem1D_1_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9070.4]
  wire  Mem1D_1_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9070.4]
  wire  Mem1D_1_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9070.4]
  wire [7:0] Mem1D_1_io_w_data_0; // @[MemPrimitives.scala 64:21:@9070.4]
  wire  Mem1D_1_io_w_en_0; // @[MemPrimitives.scala 64:21:@9070.4]
  wire [7:0] Mem1D_1_io_output; // @[MemPrimitives.scala 64:21:@9070.4]
  wire  Mem1D_2_clock; // @[MemPrimitives.scala 64:21:@9086.4]
  wire  Mem1D_2_reset; // @[MemPrimitives.scala 64:21:@9086.4]
  wire  Mem1D_2_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9086.4]
  wire  Mem1D_2_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9086.4]
  wire  Mem1D_2_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9086.4]
  wire [7:0] Mem1D_2_io_w_data_0; // @[MemPrimitives.scala 64:21:@9086.4]
  wire  Mem1D_2_io_w_en_0; // @[MemPrimitives.scala 64:21:@9086.4]
  wire [7:0] Mem1D_2_io_output; // @[MemPrimitives.scala 64:21:@9086.4]
  wire  Mem1D_3_clock; // @[MemPrimitives.scala 64:21:@9102.4]
  wire  Mem1D_3_reset; // @[MemPrimitives.scala 64:21:@9102.4]
  wire  Mem1D_3_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9102.4]
  wire  Mem1D_3_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9102.4]
  wire  Mem1D_3_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9102.4]
  wire [7:0] Mem1D_3_io_w_data_0; // @[MemPrimitives.scala 64:21:@9102.4]
  wire  Mem1D_3_io_w_en_0; // @[MemPrimitives.scala 64:21:@9102.4]
  wire [7:0] Mem1D_3_io_output; // @[MemPrimitives.scala 64:21:@9102.4]
  wire  Mem1D_4_clock; // @[MemPrimitives.scala 64:21:@9118.4]
  wire  Mem1D_4_reset; // @[MemPrimitives.scala 64:21:@9118.4]
  wire  Mem1D_4_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9118.4]
  wire  Mem1D_4_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9118.4]
  wire  Mem1D_4_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9118.4]
  wire [7:0] Mem1D_4_io_w_data_0; // @[MemPrimitives.scala 64:21:@9118.4]
  wire  Mem1D_4_io_w_en_0; // @[MemPrimitives.scala 64:21:@9118.4]
  wire [7:0] Mem1D_4_io_output; // @[MemPrimitives.scala 64:21:@9118.4]
  wire  Mem1D_5_clock; // @[MemPrimitives.scala 64:21:@9134.4]
  wire  Mem1D_5_reset; // @[MemPrimitives.scala 64:21:@9134.4]
  wire  Mem1D_5_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9134.4]
  wire  Mem1D_5_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9134.4]
  wire  Mem1D_5_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9134.4]
  wire [7:0] Mem1D_5_io_w_data_0; // @[MemPrimitives.scala 64:21:@9134.4]
  wire  Mem1D_5_io_w_en_0; // @[MemPrimitives.scala 64:21:@9134.4]
  wire [7:0] Mem1D_5_io_output; // @[MemPrimitives.scala 64:21:@9134.4]
  wire  Mem1D_6_clock; // @[MemPrimitives.scala 64:21:@9150.4]
  wire  Mem1D_6_reset; // @[MemPrimitives.scala 64:21:@9150.4]
  wire  Mem1D_6_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9150.4]
  wire  Mem1D_6_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9150.4]
  wire  Mem1D_6_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9150.4]
  wire [7:0] Mem1D_6_io_w_data_0; // @[MemPrimitives.scala 64:21:@9150.4]
  wire  Mem1D_6_io_w_en_0; // @[MemPrimitives.scala 64:21:@9150.4]
  wire [7:0] Mem1D_6_io_output; // @[MemPrimitives.scala 64:21:@9150.4]
  wire  Mem1D_7_clock; // @[MemPrimitives.scala 64:21:@9166.4]
  wire  Mem1D_7_reset; // @[MemPrimitives.scala 64:21:@9166.4]
  wire  Mem1D_7_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9166.4]
  wire  Mem1D_7_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9166.4]
  wire  Mem1D_7_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9166.4]
  wire [7:0] Mem1D_7_io_w_data_0; // @[MemPrimitives.scala 64:21:@9166.4]
  wire  Mem1D_7_io_w_en_0; // @[MemPrimitives.scala 64:21:@9166.4]
  wire [7:0] Mem1D_7_io_output; // @[MemPrimitives.scala 64:21:@9166.4]
  wire  Mem1D_8_clock; // @[MemPrimitives.scala 64:21:@9182.4]
  wire  Mem1D_8_reset; // @[MemPrimitives.scala 64:21:@9182.4]
  wire  Mem1D_8_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9182.4]
  wire  Mem1D_8_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9182.4]
  wire  Mem1D_8_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9182.4]
  wire [7:0] Mem1D_8_io_w_data_0; // @[MemPrimitives.scala 64:21:@9182.4]
  wire  Mem1D_8_io_w_en_0; // @[MemPrimitives.scala 64:21:@9182.4]
  wire [7:0] Mem1D_8_io_output; // @[MemPrimitives.scala 64:21:@9182.4]
  wire  Mem1D_9_clock; // @[MemPrimitives.scala 64:21:@9198.4]
  wire  Mem1D_9_reset; // @[MemPrimitives.scala 64:21:@9198.4]
  wire  Mem1D_9_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9198.4]
  wire  Mem1D_9_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9198.4]
  wire  Mem1D_9_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9198.4]
  wire [7:0] Mem1D_9_io_w_data_0; // @[MemPrimitives.scala 64:21:@9198.4]
  wire  Mem1D_9_io_w_en_0; // @[MemPrimitives.scala 64:21:@9198.4]
  wire [7:0] Mem1D_9_io_output; // @[MemPrimitives.scala 64:21:@9198.4]
  wire  Mem1D_10_clock; // @[MemPrimitives.scala 64:21:@9214.4]
  wire  Mem1D_10_reset; // @[MemPrimitives.scala 64:21:@9214.4]
  wire  Mem1D_10_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9214.4]
  wire  Mem1D_10_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9214.4]
  wire  Mem1D_10_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9214.4]
  wire [7:0] Mem1D_10_io_w_data_0; // @[MemPrimitives.scala 64:21:@9214.4]
  wire  Mem1D_10_io_w_en_0; // @[MemPrimitives.scala 64:21:@9214.4]
  wire [7:0] Mem1D_10_io_output; // @[MemPrimitives.scala 64:21:@9214.4]
  wire  Mem1D_11_clock; // @[MemPrimitives.scala 64:21:@9230.4]
  wire  Mem1D_11_reset; // @[MemPrimitives.scala 64:21:@9230.4]
  wire  Mem1D_11_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9230.4]
  wire  Mem1D_11_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9230.4]
  wire  Mem1D_11_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9230.4]
  wire [7:0] Mem1D_11_io_w_data_0; // @[MemPrimitives.scala 64:21:@9230.4]
  wire  Mem1D_11_io_w_en_0; // @[MemPrimitives.scala 64:21:@9230.4]
  wire [7:0] Mem1D_11_io_output; // @[MemPrimitives.scala 64:21:@9230.4]
  wire  Mem1D_12_clock; // @[MemPrimitives.scala 64:21:@9246.4]
  wire  Mem1D_12_reset; // @[MemPrimitives.scala 64:21:@9246.4]
  wire  Mem1D_12_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9246.4]
  wire  Mem1D_12_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9246.4]
  wire  Mem1D_12_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9246.4]
  wire [7:0] Mem1D_12_io_w_data_0; // @[MemPrimitives.scala 64:21:@9246.4]
  wire  Mem1D_12_io_w_en_0; // @[MemPrimitives.scala 64:21:@9246.4]
  wire [7:0] Mem1D_12_io_output; // @[MemPrimitives.scala 64:21:@9246.4]
  wire  Mem1D_13_clock; // @[MemPrimitives.scala 64:21:@9262.4]
  wire  Mem1D_13_reset; // @[MemPrimitives.scala 64:21:@9262.4]
  wire  Mem1D_13_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9262.4]
  wire  Mem1D_13_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9262.4]
  wire  Mem1D_13_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9262.4]
  wire [7:0] Mem1D_13_io_w_data_0; // @[MemPrimitives.scala 64:21:@9262.4]
  wire  Mem1D_13_io_w_en_0; // @[MemPrimitives.scala 64:21:@9262.4]
  wire [7:0] Mem1D_13_io_output; // @[MemPrimitives.scala 64:21:@9262.4]
  wire  Mem1D_14_clock; // @[MemPrimitives.scala 64:21:@9278.4]
  wire  Mem1D_14_reset; // @[MemPrimitives.scala 64:21:@9278.4]
  wire  Mem1D_14_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9278.4]
  wire  Mem1D_14_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9278.4]
  wire  Mem1D_14_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9278.4]
  wire [7:0] Mem1D_14_io_w_data_0; // @[MemPrimitives.scala 64:21:@9278.4]
  wire  Mem1D_14_io_w_en_0; // @[MemPrimitives.scala 64:21:@9278.4]
  wire [7:0] Mem1D_14_io_output; // @[MemPrimitives.scala 64:21:@9278.4]
  wire  Mem1D_15_clock; // @[MemPrimitives.scala 64:21:@9294.4]
  wire  Mem1D_15_reset; // @[MemPrimitives.scala 64:21:@9294.4]
  wire  Mem1D_15_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9294.4]
  wire  Mem1D_15_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9294.4]
  wire  Mem1D_15_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9294.4]
  wire [7:0] Mem1D_15_io_w_data_0; // @[MemPrimitives.scala 64:21:@9294.4]
  wire  Mem1D_15_io_w_en_0; // @[MemPrimitives.scala 64:21:@9294.4]
  wire [7:0] Mem1D_15_io_output; // @[MemPrimitives.scala 64:21:@9294.4]
  wire  StickySelects_clock; // @[MemPrimitives.scala 121:29:@9526.4]
  wire  StickySelects_reset; // @[MemPrimitives.scala 121:29:@9526.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 121:29:@9526.4]
  wire  StickySelects_io_ins_1; // @[MemPrimitives.scala 121:29:@9526.4]
  wire  StickySelects_io_ins_2; // @[MemPrimitives.scala 121:29:@9526.4]
  wire  StickySelects_io_ins_3; // @[MemPrimitives.scala 121:29:@9526.4]
  wire  StickySelects_io_ins_4; // @[MemPrimitives.scala 121:29:@9526.4]
  wire  StickySelects_io_ins_5; // @[MemPrimitives.scala 121:29:@9526.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 121:29:@9526.4]
  wire  StickySelects_io_outs_1; // @[MemPrimitives.scala 121:29:@9526.4]
  wire  StickySelects_io_outs_2; // @[MemPrimitives.scala 121:29:@9526.4]
  wire  StickySelects_io_outs_3; // @[MemPrimitives.scala 121:29:@9526.4]
  wire  StickySelects_io_outs_4; // @[MemPrimitives.scala 121:29:@9526.4]
  wire  StickySelects_io_outs_5; // @[MemPrimitives.scala 121:29:@9526.4]
  wire  StickySelects_1_clock; // @[MemPrimitives.scala 121:29:@9588.4]
  wire  StickySelects_1_reset; // @[MemPrimitives.scala 121:29:@9588.4]
  wire  StickySelects_1_io_ins_0; // @[MemPrimitives.scala 121:29:@9588.4]
  wire  StickySelects_1_io_ins_1; // @[MemPrimitives.scala 121:29:@9588.4]
  wire  StickySelects_1_io_ins_2; // @[MemPrimitives.scala 121:29:@9588.4]
  wire  StickySelects_1_io_ins_3; // @[MemPrimitives.scala 121:29:@9588.4]
  wire  StickySelects_1_io_ins_4; // @[MemPrimitives.scala 121:29:@9588.4]
  wire  StickySelects_1_io_ins_5; // @[MemPrimitives.scala 121:29:@9588.4]
  wire  StickySelects_1_io_outs_0; // @[MemPrimitives.scala 121:29:@9588.4]
  wire  StickySelects_1_io_outs_1; // @[MemPrimitives.scala 121:29:@9588.4]
  wire  StickySelects_1_io_outs_2; // @[MemPrimitives.scala 121:29:@9588.4]
  wire  StickySelects_1_io_outs_3; // @[MemPrimitives.scala 121:29:@9588.4]
  wire  StickySelects_1_io_outs_4; // @[MemPrimitives.scala 121:29:@9588.4]
  wire  StickySelects_1_io_outs_5; // @[MemPrimitives.scala 121:29:@9588.4]
  wire  StickySelects_2_clock; // @[MemPrimitives.scala 121:29:@9650.4]
  wire  StickySelects_2_reset; // @[MemPrimitives.scala 121:29:@9650.4]
  wire  StickySelects_2_io_ins_0; // @[MemPrimitives.scala 121:29:@9650.4]
  wire  StickySelects_2_io_ins_1; // @[MemPrimitives.scala 121:29:@9650.4]
  wire  StickySelects_2_io_ins_2; // @[MemPrimitives.scala 121:29:@9650.4]
  wire  StickySelects_2_io_ins_3; // @[MemPrimitives.scala 121:29:@9650.4]
  wire  StickySelects_2_io_ins_4; // @[MemPrimitives.scala 121:29:@9650.4]
  wire  StickySelects_2_io_ins_5; // @[MemPrimitives.scala 121:29:@9650.4]
  wire  StickySelects_2_io_outs_0; // @[MemPrimitives.scala 121:29:@9650.4]
  wire  StickySelects_2_io_outs_1; // @[MemPrimitives.scala 121:29:@9650.4]
  wire  StickySelects_2_io_outs_2; // @[MemPrimitives.scala 121:29:@9650.4]
  wire  StickySelects_2_io_outs_3; // @[MemPrimitives.scala 121:29:@9650.4]
  wire  StickySelects_2_io_outs_4; // @[MemPrimitives.scala 121:29:@9650.4]
  wire  StickySelects_2_io_outs_5; // @[MemPrimitives.scala 121:29:@9650.4]
  wire  StickySelects_3_clock; // @[MemPrimitives.scala 121:29:@9712.4]
  wire  StickySelects_3_reset; // @[MemPrimitives.scala 121:29:@9712.4]
  wire  StickySelects_3_io_ins_0; // @[MemPrimitives.scala 121:29:@9712.4]
  wire  StickySelects_3_io_ins_1; // @[MemPrimitives.scala 121:29:@9712.4]
  wire  StickySelects_3_io_ins_2; // @[MemPrimitives.scala 121:29:@9712.4]
  wire  StickySelects_3_io_ins_3; // @[MemPrimitives.scala 121:29:@9712.4]
  wire  StickySelects_3_io_ins_4; // @[MemPrimitives.scala 121:29:@9712.4]
  wire  StickySelects_3_io_ins_5; // @[MemPrimitives.scala 121:29:@9712.4]
  wire  StickySelects_3_io_outs_0; // @[MemPrimitives.scala 121:29:@9712.4]
  wire  StickySelects_3_io_outs_1; // @[MemPrimitives.scala 121:29:@9712.4]
  wire  StickySelects_3_io_outs_2; // @[MemPrimitives.scala 121:29:@9712.4]
  wire  StickySelects_3_io_outs_3; // @[MemPrimitives.scala 121:29:@9712.4]
  wire  StickySelects_3_io_outs_4; // @[MemPrimitives.scala 121:29:@9712.4]
  wire  StickySelects_3_io_outs_5; // @[MemPrimitives.scala 121:29:@9712.4]
  wire  StickySelects_4_clock; // @[MemPrimitives.scala 121:29:@9774.4]
  wire  StickySelects_4_reset; // @[MemPrimitives.scala 121:29:@9774.4]
  wire  StickySelects_4_io_ins_0; // @[MemPrimitives.scala 121:29:@9774.4]
  wire  StickySelects_4_io_ins_1; // @[MemPrimitives.scala 121:29:@9774.4]
  wire  StickySelects_4_io_ins_2; // @[MemPrimitives.scala 121:29:@9774.4]
  wire  StickySelects_4_io_ins_3; // @[MemPrimitives.scala 121:29:@9774.4]
  wire  StickySelects_4_io_ins_4; // @[MemPrimitives.scala 121:29:@9774.4]
  wire  StickySelects_4_io_ins_5; // @[MemPrimitives.scala 121:29:@9774.4]
  wire  StickySelects_4_io_outs_0; // @[MemPrimitives.scala 121:29:@9774.4]
  wire  StickySelects_4_io_outs_1; // @[MemPrimitives.scala 121:29:@9774.4]
  wire  StickySelects_4_io_outs_2; // @[MemPrimitives.scala 121:29:@9774.4]
  wire  StickySelects_4_io_outs_3; // @[MemPrimitives.scala 121:29:@9774.4]
  wire  StickySelects_4_io_outs_4; // @[MemPrimitives.scala 121:29:@9774.4]
  wire  StickySelects_4_io_outs_5; // @[MemPrimitives.scala 121:29:@9774.4]
  wire  StickySelects_5_clock; // @[MemPrimitives.scala 121:29:@9836.4]
  wire  StickySelects_5_reset; // @[MemPrimitives.scala 121:29:@9836.4]
  wire  StickySelects_5_io_ins_0; // @[MemPrimitives.scala 121:29:@9836.4]
  wire  StickySelects_5_io_ins_1; // @[MemPrimitives.scala 121:29:@9836.4]
  wire  StickySelects_5_io_ins_2; // @[MemPrimitives.scala 121:29:@9836.4]
  wire  StickySelects_5_io_ins_3; // @[MemPrimitives.scala 121:29:@9836.4]
  wire  StickySelects_5_io_ins_4; // @[MemPrimitives.scala 121:29:@9836.4]
  wire  StickySelects_5_io_ins_5; // @[MemPrimitives.scala 121:29:@9836.4]
  wire  StickySelects_5_io_outs_0; // @[MemPrimitives.scala 121:29:@9836.4]
  wire  StickySelects_5_io_outs_1; // @[MemPrimitives.scala 121:29:@9836.4]
  wire  StickySelects_5_io_outs_2; // @[MemPrimitives.scala 121:29:@9836.4]
  wire  StickySelects_5_io_outs_3; // @[MemPrimitives.scala 121:29:@9836.4]
  wire  StickySelects_5_io_outs_4; // @[MemPrimitives.scala 121:29:@9836.4]
  wire  StickySelects_5_io_outs_5; // @[MemPrimitives.scala 121:29:@9836.4]
  wire  StickySelects_6_clock; // @[MemPrimitives.scala 121:29:@9898.4]
  wire  StickySelects_6_reset; // @[MemPrimitives.scala 121:29:@9898.4]
  wire  StickySelects_6_io_ins_0; // @[MemPrimitives.scala 121:29:@9898.4]
  wire  StickySelects_6_io_ins_1; // @[MemPrimitives.scala 121:29:@9898.4]
  wire  StickySelects_6_io_ins_2; // @[MemPrimitives.scala 121:29:@9898.4]
  wire  StickySelects_6_io_ins_3; // @[MemPrimitives.scala 121:29:@9898.4]
  wire  StickySelects_6_io_ins_4; // @[MemPrimitives.scala 121:29:@9898.4]
  wire  StickySelects_6_io_ins_5; // @[MemPrimitives.scala 121:29:@9898.4]
  wire  StickySelects_6_io_outs_0; // @[MemPrimitives.scala 121:29:@9898.4]
  wire  StickySelects_6_io_outs_1; // @[MemPrimitives.scala 121:29:@9898.4]
  wire  StickySelects_6_io_outs_2; // @[MemPrimitives.scala 121:29:@9898.4]
  wire  StickySelects_6_io_outs_3; // @[MemPrimitives.scala 121:29:@9898.4]
  wire  StickySelects_6_io_outs_4; // @[MemPrimitives.scala 121:29:@9898.4]
  wire  StickySelects_6_io_outs_5; // @[MemPrimitives.scala 121:29:@9898.4]
  wire  StickySelects_7_clock; // @[MemPrimitives.scala 121:29:@9960.4]
  wire  StickySelects_7_reset; // @[MemPrimitives.scala 121:29:@9960.4]
  wire  StickySelects_7_io_ins_0; // @[MemPrimitives.scala 121:29:@9960.4]
  wire  StickySelects_7_io_ins_1; // @[MemPrimitives.scala 121:29:@9960.4]
  wire  StickySelects_7_io_ins_2; // @[MemPrimitives.scala 121:29:@9960.4]
  wire  StickySelects_7_io_ins_3; // @[MemPrimitives.scala 121:29:@9960.4]
  wire  StickySelects_7_io_ins_4; // @[MemPrimitives.scala 121:29:@9960.4]
  wire  StickySelects_7_io_ins_5; // @[MemPrimitives.scala 121:29:@9960.4]
  wire  StickySelects_7_io_outs_0; // @[MemPrimitives.scala 121:29:@9960.4]
  wire  StickySelects_7_io_outs_1; // @[MemPrimitives.scala 121:29:@9960.4]
  wire  StickySelects_7_io_outs_2; // @[MemPrimitives.scala 121:29:@9960.4]
  wire  StickySelects_7_io_outs_3; // @[MemPrimitives.scala 121:29:@9960.4]
  wire  StickySelects_7_io_outs_4; // @[MemPrimitives.scala 121:29:@9960.4]
  wire  StickySelects_7_io_outs_5; // @[MemPrimitives.scala 121:29:@9960.4]
  wire  StickySelects_8_clock; // @[MemPrimitives.scala 121:29:@10022.4]
  wire  StickySelects_8_reset; // @[MemPrimitives.scala 121:29:@10022.4]
  wire  StickySelects_8_io_ins_0; // @[MemPrimitives.scala 121:29:@10022.4]
  wire  StickySelects_8_io_ins_1; // @[MemPrimitives.scala 121:29:@10022.4]
  wire  StickySelects_8_io_ins_2; // @[MemPrimitives.scala 121:29:@10022.4]
  wire  StickySelects_8_io_ins_3; // @[MemPrimitives.scala 121:29:@10022.4]
  wire  StickySelects_8_io_ins_4; // @[MemPrimitives.scala 121:29:@10022.4]
  wire  StickySelects_8_io_ins_5; // @[MemPrimitives.scala 121:29:@10022.4]
  wire  StickySelects_8_io_outs_0; // @[MemPrimitives.scala 121:29:@10022.4]
  wire  StickySelects_8_io_outs_1; // @[MemPrimitives.scala 121:29:@10022.4]
  wire  StickySelects_8_io_outs_2; // @[MemPrimitives.scala 121:29:@10022.4]
  wire  StickySelects_8_io_outs_3; // @[MemPrimitives.scala 121:29:@10022.4]
  wire  StickySelects_8_io_outs_4; // @[MemPrimitives.scala 121:29:@10022.4]
  wire  StickySelects_8_io_outs_5; // @[MemPrimitives.scala 121:29:@10022.4]
  wire  StickySelects_9_clock; // @[MemPrimitives.scala 121:29:@10084.4]
  wire  StickySelects_9_reset; // @[MemPrimitives.scala 121:29:@10084.4]
  wire  StickySelects_9_io_ins_0; // @[MemPrimitives.scala 121:29:@10084.4]
  wire  StickySelects_9_io_ins_1; // @[MemPrimitives.scala 121:29:@10084.4]
  wire  StickySelects_9_io_ins_2; // @[MemPrimitives.scala 121:29:@10084.4]
  wire  StickySelects_9_io_ins_3; // @[MemPrimitives.scala 121:29:@10084.4]
  wire  StickySelects_9_io_ins_4; // @[MemPrimitives.scala 121:29:@10084.4]
  wire  StickySelects_9_io_ins_5; // @[MemPrimitives.scala 121:29:@10084.4]
  wire  StickySelects_9_io_outs_0; // @[MemPrimitives.scala 121:29:@10084.4]
  wire  StickySelects_9_io_outs_1; // @[MemPrimitives.scala 121:29:@10084.4]
  wire  StickySelects_9_io_outs_2; // @[MemPrimitives.scala 121:29:@10084.4]
  wire  StickySelects_9_io_outs_3; // @[MemPrimitives.scala 121:29:@10084.4]
  wire  StickySelects_9_io_outs_4; // @[MemPrimitives.scala 121:29:@10084.4]
  wire  StickySelects_9_io_outs_5; // @[MemPrimitives.scala 121:29:@10084.4]
  wire  StickySelects_10_clock; // @[MemPrimitives.scala 121:29:@10146.4]
  wire  StickySelects_10_reset; // @[MemPrimitives.scala 121:29:@10146.4]
  wire  StickySelects_10_io_ins_0; // @[MemPrimitives.scala 121:29:@10146.4]
  wire  StickySelects_10_io_ins_1; // @[MemPrimitives.scala 121:29:@10146.4]
  wire  StickySelects_10_io_ins_2; // @[MemPrimitives.scala 121:29:@10146.4]
  wire  StickySelects_10_io_ins_3; // @[MemPrimitives.scala 121:29:@10146.4]
  wire  StickySelects_10_io_ins_4; // @[MemPrimitives.scala 121:29:@10146.4]
  wire  StickySelects_10_io_ins_5; // @[MemPrimitives.scala 121:29:@10146.4]
  wire  StickySelects_10_io_outs_0; // @[MemPrimitives.scala 121:29:@10146.4]
  wire  StickySelects_10_io_outs_1; // @[MemPrimitives.scala 121:29:@10146.4]
  wire  StickySelects_10_io_outs_2; // @[MemPrimitives.scala 121:29:@10146.4]
  wire  StickySelects_10_io_outs_3; // @[MemPrimitives.scala 121:29:@10146.4]
  wire  StickySelects_10_io_outs_4; // @[MemPrimitives.scala 121:29:@10146.4]
  wire  StickySelects_10_io_outs_5; // @[MemPrimitives.scala 121:29:@10146.4]
  wire  StickySelects_11_clock; // @[MemPrimitives.scala 121:29:@10208.4]
  wire  StickySelects_11_reset; // @[MemPrimitives.scala 121:29:@10208.4]
  wire  StickySelects_11_io_ins_0; // @[MemPrimitives.scala 121:29:@10208.4]
  wire  StickySelects_11_io_ins_1; // @[MemPrimitives.scala 121:29:@10208.4]
  wire  StickySelects_11_io_ins_2; // @[MemPrimitives.scala 121:29:@10208.4]
  wire  StickySelects_11_io_ins_3; // @[MemPrimitives.scala 121:29:@10208.4]
  wire  StickySelects_11_io_ins_4; // @[MemPrimitives.scala 121:29:@10208.4]
  wire  StickySelects_11_io_ins_5; // @[MemPrimitives.scala 121:29:@10208.4]
  wire  StickySelects_11_io_outs_0; // @[MemPrimitives.scala 121:29:@10208.4]
  wire  StickySelects_11_io_outs_1; // @[MemPrimitives.scala 121:29:@10208.4]
  wire  StickySelects_11_io_outs_2; // @[MemPrimitives.scala 121:29:@10208.4]
  wire  StickySelects_11_io_outs_3; // @[MemPrimitives.scala 121:29:@10208.4]
  wire  StickySelects_11_io_outs_4; // @[MemPrimitives.scala 121:29:@10208.4]
  wire  StickySelects_11_io_outs_5; // @[MemPrimitives.scala 121:29:@10208.4]
  wire  StickySelects_12_clock; // @[MemPrimitives.scala 121:29:@10270.4]
  wire  StickySelects_12_reset; // @[MemPrimitives.scala 121:29:@10270.4]
  wire  StickySelects_12_io_ins_0; // @[MemPrimitives.scala 121:29:@10270.4]
  wire  StickySelects_12_io_ins_1; // @[MemPrimitives.scala 121:29:@10270.4]
  wire  StickySelects_12_io_ins_2; // @[MemPrimitives.scala 121:29:@10270.4]
  wire  StickySelects_12_io_ins_3; // @[MemPrimitives.scala 121:29:@10270.4]
  wire  StickySelects_12_io_ins_4; // @[MemPrimitives.scala 121:29:@10270.4]
  wire  StickySelects_12_io_ins_5; // @[MemPrimitives.scala 121:29:@10270.4]
  wire  StickySelects_12_io_outs_0; // @[MemPrimitives.scala 121:29:@10270.4]
  wire  StickySelects_12_io_outs_1; // @[MemPrimitives.scala 121:29:@10270.4]
  wire  StickySelects_12_io_outs_2; // @[MemPrimitives.scala 121:29:@10270.4]
  wire  StickySelects_12_io_outs_3; // @[MemPrimitives.scala 121:29:@10270.4]
  wire  StickySelects_12_io_outs_4; // @[MemPrimitives.scala 121:29:@10270.4]
  wire  StickySelects_12_io_outs_5; // @[MemPrimitives.scala 121:29:@10270.4]
  wire  StickySelects_13_clock; // @[MemPrimitives.scala 121:29:@10332.4]
  wire  StickySelects_13_reset; // @[MemPrimitives.scala 121:29:@10332.4]
  wire  StickySelects_13_io_ins_0; // @[MemPrimitives.scala 121:29:@10332.4]
  wire  StickySelects_13_io_ins_1; // @[MemPrimitives.scala 121:29:@10332.4]
  wire  StickySelects_13_io_ins_2; // @[MemPrimitives.scala 121:29:@10332.4]
  wire  StickySelects_13_io_ins_3; // @[MemPrimitives.scala 121:29:@10332.4]
  wire  StickySelects_13_io_ins_4; // @[MemPrimitives.scala 121:29:@10332.4]
  wire  StickySelects_13_io_ins_5; // @[MemPrimitives.scala 121:29:@10332.4]
  wire  StickySelects_13_io_outs_0; // @[MemPrimitives.scala 121:29:@10332.4]
  wire  StickySelects_13_io_outs_1; // @[MemPrimitives.scala 121:29:@10332.4]
  wire  StickySelects_13_io_outs_2; // @[MemPrimitives.scala 121:29:@10332.4]
  wire  StickySelects_13_io_outs_3; // @[MemPrimitives.scala 121:29:@10332.4]
  wire  StickySelects_13_io_outs_4; // @[MemPrimitives.scala 121:29:@10332.4]
  wire  StickySelects_13_io_outs_5; // @[MemPrimitives.scala 121:29:@10332.4]
  wire  StickySelects_14_clock; // @[MemPrimitives.scala 121:29:@10394.4]
  wire  StickySelects_14_reset; // @[MemPrimitives.scala 121:29:@10394.4]
  wire  StickySelects_14_io_ins_0; // @[MemPrimitives.scala 121:29:@10394.4]
  wire  StickySelects_14_io_ins_1; // @[MemPrimitives.scala 121:29:@10394.4]
  wire  StickySelects_14_io_ins_2; // @[MemPrimitives.scala 121:29:@10394.4]
  wire  StickySelects_14_io_ins_3; // @[MemPrimitives.scala 121:29:@10394.4]
  wire  StickySelects_14_io_ins_4; // @[MemPrimitives.scala 121:29:@10394.4]
  wire  StickySelects_14_io_ins_5; // @[MemPrimitives.scala 121:29:@10394.4]
  wire  StickySelects_14_io_outs_0; // @[MemPrimitives.scala 121:29:@10394.4]
  wire  StickySelects_14_io_outs_1; // @[MemPrimitives.scala 121:29:@10394.4]
  wire  StickySelects_14_io_outs_2; // @[MemPrimitives.scala 121:29:@10394.4]
  wire  StickySelects_14_io_outs_3; // @[MemPrimitives.scala 121:29:@10394.4]
  wire  StickySelects_14_io_outs_4; // @[MemPrimitives.scala 121:29:@10394.4]
  wire  StickySelects_14_io_outs_5; // @[MemPrimitives.scala 121:29:@10394.4]
  wire  StickySelects_15_clock; // @[MemPrimitives.scala 121:29:@10456.4]
  wire  StickySelects_15_reset; // @[MemPrimitives.scala 121:29:@10456.4]
  wire  StickySelects_15_io_ins_0; // @[MemPrimitives.scala 121:29:@10456.4]
  wire  StickySelects_15_io_ins_1; // @[MemPrimitives.scala 121:29:@10456.4]
  wire  StickySelects_15_io_ins_2; // @[MemPrimitives.scala 121:29:@10456.4]
  wire  StickySelects_15_io_ins_3; // @[MemPrimitives.scala 121:29:@10456.4]
  wire  StickySelects_15_io_ins_4; // @[MemPrimitives.scala 121:29:@10456.4]
  wire  StickySelects_15_io_ins_5; // @[MemPrimitives.scala 121:29:@10456.4]
  wire  StickySelects_15_io_outs_0; // @[MemPrimitives.scala 121:29:@10456.4]
  wire  StickySelects_15_io_outs_1; // @[MemPrimitives.scala 121:29:@10456.4]
  wire  StickySelects_15_io_outs_2; // @[MemPrimitives.scala 121:29:@10456.4]
  wire  StickySelects_15_io_outs_3; // @[MemPrimitives.scala 121:29:@10456.4]
  wire  StickySelects_15_io_outs_4; // @[MemPrimitives.scala 121:29:@10456.4]
  wire  StickySelects_15_io_outs_5; // @[MemPrimitives.scala 121:29:@10456.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@10519.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@10519.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@10519.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@10519.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@10519.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@10527.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@10527.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@10527.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@10527.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@10527.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@10535.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@10535.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@10535.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@10535.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@10535.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@10543.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@10543.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@10543.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@10543.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@10543.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@10551.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@10551.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@10551.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@10551.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@10551.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@10559.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@10559.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@10559.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@10559.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@10559.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@10567.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@10567.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@10567.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@10567.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@10567.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@10575.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@10575.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@10575.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@10575.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@10575.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@10615.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@10615.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@10615.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@10615.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@10615.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@10623.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@10623.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@10623.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@10623.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@10623.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@10631.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@10631.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@10631.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@10631.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@10631.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@10639.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@10639.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@10639.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@10639.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@10639.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@10647.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@10647.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@10647.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@10647.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@10647.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@10655.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@10655.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@10655.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@10655.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@10655.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@10663.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@10663.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@10663.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@10663.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@10663.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@10671.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@10671.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@10671.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@10671.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@10671.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@10711.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@10711.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@10711.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@10711.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@10711.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@10719.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@10719.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@10719.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@10719.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@10719.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@10727.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@10727.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@10727.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@10727.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@10727.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@10735.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@10735.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@10735.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@10735.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@10735.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@10743.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@10743.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@10743.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@10743.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@10743.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@10751.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@10751.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@10751.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@10751.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@10751.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@10759.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@10759.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@10759.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@10759.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@10759.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@10767.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@10767.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@10767.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@10767.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@10767.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@10807.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@10807.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@10807.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@10807.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@10807.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@10815.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@10815.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@10815.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@10815.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@10815.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@10823.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@10823.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@10823.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@10823.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@10823.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@10831.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@10831.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@10831.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@10831.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@10831.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@10839.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@10839.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@10839.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@10839.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@10839.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@10847.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@10847.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@10847.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@10847.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@10847.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@10855.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@10855.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@10855.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@10855.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@10855.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@10863.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@10863.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@10863.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@10863.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@10863.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@10903.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@10903.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@10903.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@10903.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@10903.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@10911.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@10911.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@10911.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@10911.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@10911.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@10919.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@10919.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@10919.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@10919.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@10919.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@10927.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@10927.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@10927.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@10927.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@10927.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@10935.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@10935.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@10935.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@10935.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@10935.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@10943.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@10943.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@10943.4]
  wire  RetimeWrapper_37_io_in; // @[package.scala 93:22:@10943.4]
  wire  RetimeWrapper_37_io_out; // @[package.scala 93:22:@10943.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@10951.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@10951.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@10951.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@10951.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@10951.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@10959.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@10959.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@10959.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@10959.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@10959.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@10999.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@10999.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@10999.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@10999.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@10999.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@11007.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@11007.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@11007.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@11007.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@11007.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@11015.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@11015.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@11015.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@11015.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@11015.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@11023.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@11023.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@11023.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@11023.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@11023.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@11031.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@11031.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@11031.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@11031.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@11031.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@11039.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@11039.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@11039.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@11039.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@11039.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@11047.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@11047.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@11047.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@11047.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@11047.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@11055.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@11055.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@11055.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@11055.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@11055.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@11095.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@11095.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@11095.4]
  wire  RetimeWrapper_48_io_in; // @[package.scala 93:22:@11095.4]
  wire  RetimeWrapper_48_io_out; // @[package.scala 93:22:@11095.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@11103.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@11103.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@11103.4]
  wire  RetimeWrapper_49_io_in; // @[package.scala 93:22:@11103.4]
  wire  RetimeWrapper_49_io_out; // @[package.scala 93:22:@11103.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@11111.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@11111.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@11111.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@11111.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@11111.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@11119.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@11119.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@11119.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@11119.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@11119.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@11127.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@11127.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@11127.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@11127.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@11127.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@11135.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@11135.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@11135.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@11135.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@11135.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@11143.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@11143.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@11143.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@11143.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@11143.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@11151.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@11151.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@11151.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@11151.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@11151.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@11191.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@11191.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@11191.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@11191.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@11191.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@11199.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@11199.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@11199.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@11199.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@11199.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@11207.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@11207.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@11207.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@11207.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@11207.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@11215.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@11215.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@11215.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@11215.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@11215.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@11223.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@11223.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@11223.4]
  wire  RetimeWrapper_60_io_in; // @[package.scala 93:22:@11223.4]
  wire  RetimeWrapper_60_io_out; // @[package.scala 93:22:@11223.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@11231.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@11231.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@11231.4]
  wire  RetimeWrapper_61_io_in; // @[package.scala 93:22:@11231.4]
  wire  RetimeWrapper_61_io_out; // @[package.scala 93:22:@11231.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@11239.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@11239.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@11239.4]
  wire  RetimeWrapper_62_io_in; // @[package.scala 93:22:@11239.4]
  wire  RetimeWrapper_62_io_out; // @[package.scala 93:22:@11239.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@11247.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@11247.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@11247.4]
  wire  RetimeWrapper_63_io_in; // @[package.scala 93:22:@11247.4]
  wire  RetimeWrapper_63_io_out; // @[package.scala 93:22:@11247.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@11287.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@11287.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@11287.4]
  wire  RetimeWrapper_64_io_in; // @[package.scala 93:22:@11287.4]
  wire  RetimeWrapper_64_io_out; // @[package.scala 93:22:@11287.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@11295.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@11295.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@11295.4]
  wire  RetimeWrapper_65_io_in; // @[package.scala 93:22:@11295.4]
  wire  RetimeWrapper_65_io_out; // @[package.scala 93:22:@11295.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@11303.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@11303.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@11303.4]
  wire  RetimeWrapper_66_io_in; // @[package.scala 93:22:@11303.4]
  wire  RetimeWrapper_66_io_out; // @[package.scala 93:22:@11303.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@11311.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@11311.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@11311.4]
  wire  RetimeWrapper_67_io_in; // @[package.scala 93:22:@11311.4]
  wire  RetimeWrapper_67_io_out; // @[package.scala 93:22:@11311.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@11319.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@11319.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@11319.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@11319.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@11319.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@11327.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@11327.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@11327.4]
  wire  RetimeWrapper_69_io_in; // @[package.scala 93:22:@11327.4]
  wire  RetimeWrapper_69_io_out; // @[package.scala 93:22:@11327.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@11335.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@11335.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@11335.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@11335.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@11335.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@11343.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@11343.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@11343.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@11343.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@11343.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@11383.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@11383.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@11383.4]
  wire  RetimeWrapper_72_io_in; // @[package.scala 93:22:@11383.4]
  wire  RetimeWrapper_72_io_out; // @[package.scala 93:22:@11383.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@11391.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@11391.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@11391.4]
  wire  RetimeWrapper_73_io_in; // @[package.scala 93:22:@11391.4]
  wire  RetimeWrapper_73_io_out; // @[package.scala 93:22:@11391.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@11399.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@11399.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@11399.4]
  wire  RetimeWrapper_74_io_in; // @[package.scala 93:22:@11399.4]
  wire  RetimeWrapper_74_io_out; // @[package.scala 93:22:@11399.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@11407.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@11407.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@11407.4]
  wire  RetimeWrapper_75_io_in; // @[package.scala 93:22:@11407.4]
  wire  RetimeWrapper_75_io_out; // @[package.scala 93:22:@11407.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@11415.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@11415.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@11415.4]
  wire  RetimeWrapper_76_io_in; // @[package.scala 93:22:@11415.4]
  wire  RetimeWrapper_76_io_out; // @[package.scala 93:22:@11415.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@11423.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@11423.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@11423.4]
  wire  RetimeWrapper_77_io_in; // @[package.scala 93:22:@11423.4]
  wire  RetimeWrapper_77_io_out; // @[package.scala 93:22:@11423.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@11431.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@11431.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@11431.4]
  wire  RetimeWrapper_78_io_in; // @[package.scala 93:22:@11431.4]
  wire  RetimeWrapper_78_io_out; // @[package.scala 93:22:@11431.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@11439.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@11439.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@11439.4]
  wire  RetimeWrapper_79_io_in; // @[package.scala 93:22:@11439.4]
  wire  RetimeWrapper_79_io_out; // @[package.scala 93:22:@11439.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@11479.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@11479.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@11479.4]
  wire  RetimeWrapper_80_io_in; // @[package.scala 93:22:@11479.4]
  wire  RetimeWrapper_80_io_out; // @[package.scala 93:22:@11479.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@11487.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@11487.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@11487.4]
  wire  RetimeWrapper_81_io_in; // @[package.scala 93:22:@11487.4]
  wire  RetimeWrapper_81_io_out; // @[package.scala 93:22:@11487.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@11495.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@11495.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@11495.4]
  wire  RetimeWrapper_82_io_in; // @[package.scala 93:22:@11495.4]
  wire  RetimeWrapper_82_io_out; // @[package.scala 93:22:@11495.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@11503.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@11503.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@11503.4]
  wire  RetimeWrapper_83_io_in; // @[package.scala 93:22:@11503.4]
  wire  RetimeWrapper_83_io_out; // @[package.scala 93:22:@11503.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@11511.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@11511.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@11511.4]
  wire  RetimeWrapper_84_io_in; // @[package.scala 93:22:@11511.4]
  wire  RetimeWrapper_84_io_out; // @[package.scala 93:22:@11511.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@11519.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@11519.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@11519.4]
  wire  RetimeWrapper_85_io_in; // @[package.scala 93:22:@11519.4]
  wire  RetimeWrapper_85_io_out; // @[package.scala 93:22:@11519.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@11527.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@11527.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@11527.4]
  wire  RetimeWrapper_86_io_in; // @[package.scala 93:22:@11527.4]
  wire  RetimeWrapper_86_io_out; // @[package.scala 93:22:@11527.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@11535.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@11535.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@11535.4]
  wire  RetimeWrapper_87_io_in; // @[package.scala 93:22:@11535.4]
  wire  RetimeWrapper_87_io_out; // @[package.scala 93:22:@11535.4]
  wire  RetimeWrapper_88_clock; // @[package.scala 93:22:@11575.4]
  wire  RetimeWrapper_88_reset; // @[package.scala 93:22:@11575.4]
  wire  RetimeWrapper_88_io_flow; // @[package.scala 93:22:@11575.4]
  wire  RetimeWrapper_88_io_in; // @[package.scala 93:22:@11575.4]
  wire  RetimeWrapper_88_io_out; // @[package.scala 93:22:@11575.4]
  wire  RetimeWrapper_89_clock; // @[package.scala 93:22:@11583.4]
  wire  RetimeWrapper_89_reset; // @[package.scala 93:22:@11583.4]
  wire  RetimeWrapper_89_io_flow; // @[package.scala 93:22:@11583.4]
  wire  RetimeWrapper_89_io_in; // @[package.scala 93:22:@11583.4]
  wire  RetimeWrapper_89_io_out; // @[package.scala 93:22:@11583.4]
  wire  RetimeWrapper_90_clock; // @[package.scala 93:22:@11591.4]
  wire  RetimeWrapper_90_reset; // @[package.scala 93:22:@11591.4]
  wire  RetimeWrapper_90_io_flow; // @[package.scala 93:22:@11591.4]
  wire  RetimeWrapper_90_io_in; // @[package.scala 93:22:@11591.4]
  wire  RetimeWrapper_90_io_out; // @[package.scala 93:22:@11591.4]
  wire  RetimeWrapper_91_clock; // @[package.scala 93:22:@11599.4]
  wire  RetimeWrapper_91_reset; // @[package.scala 93:22:@11599.4]
  wire  RetimeWrapper_91_io_flow; // @[package.scala 93:22:@11599.4]
  wire  RetimeWrapper_91_io_in; // @[package.scala 93:22:@11599.4]
  wire  RetimeWrapper_91_io_out; // @[package.scala 93:22:@11599.4]
  wire  RetimeWrapper_92_clock; // @[package.scala 93:22:@11607.4]
  wire  RetimeWrapper_92_reset; // @[package.scala 93:22:@11607.4]
  wire  RetimeWrapper_92_io_flow; // @[package.scala 93:22:@11607.4]
  wire  RetimeWrapper_92_io_in; // @[package.scala 93:22:@11607.4]
  wire  RetimeWrapper_92_io_out; // @[package.scala 93:22:@11607.4]
  wire  RetimeWrapper_93_clock; // @[package.scala 93:22:@11615.4]
  wire  RetimeWrapper_93_reset; // @[package.scala 93:22:@11615.4]
  wire  RetimeWrapper_93_io_flow; // @[package.scala 93:22:@11615.4]
  wire  RetimeWrapper_93_io_in; // @[package.scala 93:22:@11615.4]
  wire  RetimeWrapper_93_io_out; // @[package.scala 93:22:@11615.4]
  wire  RetimeWrapper_94_clock; // @[package.scala 93:22:@11623.4]
  wire  RetimeWrapper_94_reset; // @[package.scala 93:22:@11623.4]
  wire  RetimeWrapper_94_io_flow; // @[package.scala 93:22:@11623.4]
  wire  RetimeWrapper_94_io_in; // @[package.scala 93:22:@11623.4]
  wire  RetimeWrapper_94_io_out; // @[package.scala 93:22:@11623.4]
  wire  RetimeWrapper_95_clock; // @[package.scala 93:22:@11631.4]
  wire  RetimeWrapper_95_reset; // @[package.scala 93:22:@11631.4]
  wire  RetimeWrapper_95_io_flow; // @[package.scala 93:22:@11631.4]
  wire  RetimeWrapper_95_io_in; // @[package.scala 93:22:@11631.4]
  wire  RetimeWrapper_95_io_out; // @[package.scala 93:22:@11631.4]
  wire  _T_444; // @[MemPrimitives.scala 82:210:@9310.4]
  wire  _T_446; // @[MemPrimitives.scala 82:210:@9311.4]
  wire  _T_447; // @[MemPrimitives.scala 82:228:@9312.4]
  wire  _T_448; // @[MemPrimitives.scala 83:102:@9313.4]
  wire [9:0] _T_450; // @[Cat.scala 30:58:@9315.4]
  wire  _T_455; // @[MemPrimitives.scala 82:210:@9322.4]
  wire  _T_457; // @[MemPrimitives.scala 82:210:@9323.4]
  wire  _T_458; // @[MemPrimitives.scala 82:228:@9324.4]
  wire  _T_459; // @[MemPrimitives.scala 83:102:@9325.4]
  wire [9:0] _T_461; // @[Cat.scala 30:58:@9327.4]
  wire  _T_468; // @[MemPrimitives.scala 82:210:@9335.4]
  wire  _T_469; // @[MemPrimitives.scala 82:228:@9336.4]
  wire  _T_470; // @[MemPrimitives.scala 83:102:@9337.4]
  wire [9:0] _T_472; // @[Cat.scala 30:58:@9339.4]
  wire  _T_479; // @[MemPrimitives.scala 82:210:@9347.4]
  wire  _T_480; // @[MemPrimitives.scala 82:228:@9348.4]
  wire  _T_481; // @[MemPrimitives.scala 83:102:@9349.4]
  wire [9:0] _T_483; // @[Cat.scala 30:58:@9351.4]
  wire  _T_488; // @[MemPrimitives.scala 82:210:@9358.4]
  wire  _T_491; // @[MemPrimitives.scala 82:228:@9360.4]
  wire  _T_492; // @[MemPrimitives.scala 83:102:@9361.4]
  wire [9:0] _T_494; // @[Cat.scala 30:58:@9363.4]
  wire  _T_499; // @[MemPrimitives.scala 82:210:@9370.4]
  wire  _T_502; // @[MemPrimitives.scala 82:228:@9372.4]
  wire  _T_503; // @[MemPrimitives.scala 83:102:@9373.4]
  wire [9:0] _T_505; // @[Cat.scala 30:58:@9375.4]
  wire  _T_513; // @[MemPrimitives.scala 82:228:@9384.4]
  wire  _T_514; // @[MemPrimitives.scala 83:102:@9385.4]
  wire [9:0] _T_516; // @[Cat.scala 30:58:@9387.4]
  wire  _T_524; // @[MemPrimitives.scala 82:228:@9396.4]
  wire  _T_525; // @[MemPrimitives.scala 83:102:@9397.4]
  wire [9:0] _T_527; // @[Cat.scala 30:58:@9399.4]
  wire  _T_532; // @[MemPrimitives.scala 82:210:@9406.4]
  wire  _T_535; // @[MemPrimitives.scala 82:228:@9408.4]
  wire  _T_536; // @[MemPrimitives.scala 83:102:@9409.4]
  wire [9:0] _T_538; // @[Cat.scala 30:58:@9411.4]
  wire  _T_543; // @[MemPrimitives.scala 82:210:@9418.4]
  wire  _T_546; // @[MemPrimitives.scala 82:228:@9420.4]
  wire  _T_547; // @[MemPrimitives.scala 83:102:@9421.4]
  wire [9:0] _T_549; // @[Cat.scala 30:58:@9423.4]
  wire  _T_557; // @[MemPrimitives.scala 82:228:@9432.4]
  wire  _T_558; // @[MemPrimitives.scala 83:102:@9433.4]
  wire [9:0] _T_560; // @[Cat.scala 30:58:@9435.4]
  wire  _T_568; // @[MemPrimitives.scala 82:228:@9444.4]
  wire  _T_569; // @[MemPrimitives.scala 83:102:@9445.4]
  wire [9:0] _T_571; // @[Cat.scala 30:58:@9447.4]
  wire  _T_576; // @[MemPrimitives.scala 82:210:@9454.4]
  wire  _T_579; // @[MemPrimitives.scala 82:228:@9456.4]
  wire  _T_580; // @[MemPrimitives.scala 83:102:@9457.4]
  wire [9:0] _T_582; // @[Cat.scala 30:58:@9459.4]
  wire  _T_587; // @[MemPrimitives.scala 82:210:@9466.4]
  wire  _T_590; // @[MemPrimitives.scala 82:228:@9468.4]
  wire  _T_591; // @[MemPrimitives.scala 83:102:@9469.4]
  wire [9:0] _T_593; // @[Cat.scala 30:58:@9471.4]
  wire  _T_601; // @[MemPrimitives.scala 82:228:@9480.4]
  wire  _T_602; // @[MemPrimitives.scala 83:102:@9481.4]
  wire [9:0] _T_604; // @[Cat.scala 30:58:@9483.4]
  wire  _T_612; // @[MemPrimitives.scala 82:228:@9492.4]
  wire  _T_613; // @[MemPrimitives.scala 83:102:@9493.4]
  wire [9:0] _T_615; // @[Cat.scala 30:58:@9495.4]
  wire  _T_620; // @[MemPrimitives.scala 110:210:@9502.4]
  wire  _T_622; // @[MemPrimitives.scala 110:210:@9503.4]
  wire  _T_623; // @[MemPrimitives.scala 110:228:@9504.4]
  wire  _T_626; // @[MemPrimitives.scala 110:210:@9506.4]
  wire  _T_628; // @[MemPrimitives.scala 110:210:@9507.4]
  wire  _T_629; // @[MemPrimitives.scala 110:228:@9508.4]
  wire  _T_632; // @[MemPrimitives.scala 110:210:@9510.4]
  wire  _T_634; // @[MemPrimitives.scala 110:210:@9511.4]
  wire  _T_635; // @[MemPrimitives.scala 110:228:@9512.4]
  wire  _T_638; // @[MemPrimitives.scala 110:210:@9514.4]
  wire  _T_640; // @[MemPrimitives.scala 110:210:@9515.4]
  wire  _T_641; // @[MemPrimitives.scala 110:228:@9516.4]
  wire  _T_644; // @[MemPrimitives.scala 110:210:@9518.4]
  wire  _T_646; // @[MemPrimitives.scala 110:210:@9519.4]
  wire  _T_647; // @[MemPrimitives.scala 110:228:@9520.4]
  wire  _T_650; // @[MemPrimitives.scala 110:210:@9522.4]
  wire  _T_652; // @[MemPrimitives.scala 110:210:@9523.4]
  wire  _T_653; // @[MemPrimitives.scala 110:228:@9524.4]
  wire  _T_655; // @[MemPrimitives.scala 123:41:@9535.4]
  wire  _T_656; // @[MemPrimitives.scala 123:41:@9536.4]
  wire  _T_657; // @[MemPrimitives.scala 123:41:@9537.4]
  wire  _T_658; // @[MemPrimitives.scala 123:41:@9538.4]
  wire  _T_659; // @[MemPrimitives.scala 123:41:@9539.4]
  wire  _T_660; // @[MemPrimitives.scala 123:41:@9540.4]
  wire [2:0] _T_662; // @[Cat.scala 30:58:@9542.4]
  wire [2:0] _T_664; // @[Cat.scala 30:58:@9544.4]
  wire [2:0] _T_666; // @[Cat.scala 30:58:@9546.4]
  wire [2:0] _T_668; // @[Cat.scala 30:58:@9548.4]
  wire [2:0] _T_670; // @[Cat.scala 30:58:@9550.4]
  wire [2:0] _T_672; // @[Cat.scala 30:58:@9552.4]
  wire [2:0] _T_673; // @[Mux.scala 31:69:@9553.4]
  wire [2:0] _T_674; // @[Mux.scala 31:69:@9554.4]
  wire [2:0] _T_675; // @[Mux.scala 31:69:@9555.4]
  wire [2:0] _T_676; // @[Mux.scala 31:69:@9556.4]
  wire [2:0] _T_677; // @[Mux.scala 31:69:@9557.4]
  wire  _T_682; // @[MemPrimitives.scala 110:210:@9564.4]
  wire  _T_684; // @[MemPrimitives.scala 110:210:@9565.4]
  wire  _T_685; // @[MemPrimitives.scala 110:228:@9566.4]
  wire  _T_688; // @[MemPrimitives.scala 110:210:@9568.4]
  wire  _T_690; // @[MemPrimitives.scala 110:210:@9569.4]
  wire  _T_691; // @[MemPrimitives.scala 110:228:@9570.4]
  wire  _T_694; // @[MemPrimitives.scala 110:210:@9572.4]
  wire  _T_696; // @[MemPrimitives.scala 110:210:@9573.4]
  wire  _T_697; // @[MemPrimitives.scala 110:228:@9574.4]
  wire  _T_700; // @[MemPrimitives.scala 110:210:@9576.4]
  wire  _T_702; // @[MemPrimitives.scala 110:210:@9577.4]
  wire  _T_703; // @[MemPrimitives.scala 110:228:@9578.4]
  wire  _T_706; // @[MemPrimitives.scala 110:210:@9580.4]
  wire  _T_708; // @[MemPrimitives.scala 110:210:@9581.4]
  wire  _T_709; // @[MemPrimitives.scala 110:228:@9582.4]
  wire  _T_712; // @[MemPrimitives.scala 110:210:@9584.4]
  wire  _T_714; // @[MemPrimitives.scala 110:210:@9585.4]
  wire  _T_715; // @[MemPrimitives.scala 110:228:@9586.4]
  wire  _T_717; // @[MemPrimitives.scala 123:41:@9597.4]
  wire  _T_718; // @[MemPrimitives.scala 123:41:@9598.4]
  wire  _T_719; // @[MemPrimitives.scala 123:41:@9599.4]
  wire  _T_720; // @[MemPrimitives.scala 123:41:@9600.4]
  wire  _T_721; // @[MemPrimitives.scala 123:41:@9601.4]
  wire  _T_722; // @[MemPrimitives.scala 123:41:@9602.4]
  wire [2:0] _T_724; // @[Cat.scala 30:58:@9604.4]
  wire [2:0] _T_726; // @[Cat.scala 30:58:@9606.4]
  wire [2:0] _T_728; // @[Cat.scala 30:58:@9608.4]
  wire [2:0] _T_730; // @[Cat.scala 30:58:@9610.4]
  wire [2:0] _T_732; // @[Cat.scala 30:58:@9612.4]
  wire [2:0] _T_734; // @[Cat.scala 30:58:@9614.4]
  wire [2:0] _T_735; // @[Mux.scala 31:69:@9615.4]
  wire [2:0] _T_736; // @[Mux.scala 31:69:@9616.4]
  wire [2:0] _T_737; // @[Mux.scala 31:69:@9617.4]
  wire [2:0] _T_738; // @[Mux.scala 31:69:@9618.4]
  wire [2:0] _T_739; // @[Mux.scala 31:69:@9619.4]
  wire  _T_746; // @[MemPrimitives.scala 110:210:@9627.4]
  wire  _T_747; // @[MemPrimitives.scala 110:228:@9628.4]
  wire  _T_752; // @[MemPrimitives.scala 110:210:@9631.4]
  wire  _T_753; // @[MemPrimitives.scala 110:228:@9632.4]
  wire  _T_758; // @[MemPrimitives.scala 110:210:@9635.4]
  wire  _T_759; // @[MemPrimitives.scala 110:228:@9636.4]
  wire  _T_764; // @[MemPrimitives.scala 110:210:@9639.4]
  wire  _T_765; // @[MemPrimitives.scala 110:228:@9640.4]
  wire  _T_770; // @[MemPrimitives.scala 110:210:@9643.4]
  wire  _T_771; // @[MemPrimitives.scala 110:228:@9644.4]
  wire  _T_776; // @[MemPrimitives.scala 110:210:@9647.4]
  wire  _T_777; // @[MemPrimitives.scala 110:228:@9648.4]
  wire  _T_779; // @[MemPrimitives.scala 123:41:@9659.4]
  wire  _T_780; // @[MemPrimitives.scala 123:41:@9660.4]
  wire  _T_781; // @[MemPrimitives.scala 123:41:@9661.4]
  wire  _T_782; // @[MemPrimitives.scala 123:41:@9662.4]
  wire  _T_783; // @[MemPrimitives.scala 123:41:@9663.4]
  wire  _T_784; // @[MemPrimitives.scala 123:41:@9664.4]
  wire [2:0] _T_786; // @[Cat.scala 30:58:@9666.4]
  wire [2:0] _T_788; // @[Cat.scala 30:58:@9668.4]
  wire [2:0] _T_790; // @[Cat.scala 30:58:@9670.4]
  wire [2:0] _T_792; // @[Cat.scala 30:58:@9672.4]
  wire [2:0] _T_794; // @[Cat.scala 30:58:@9674.4]
  wire [2:0] _T_796; // @[Cat.scala 30:58:@9676.4]
  wire [2:0] _T_797; // @[Mux.scala 31:69:@9677.4]
  wire [2:0] _T_798; // @[Mux.scala 31:69:@9678.4]
  wire [2:0] _T_799; // @[Mux.scala 31:69:@9679.4]
  wire [2:0] _T_800; // @[Mux.scala 31:69:@9680.4]
  wire [2:0] _T_801; // @[Mux.scala 31:69:@9681.4]
  wire  _T_808; // @[MemPrimitives.scala 110:210:@9689.4]
  wire  _T_809; // @[MemPrimitives.scala 110:228:@9690.4]
  wire  _T_814; // @[MemPrimitives.scala 110:210:@9693.4]
  wire  _T_815; // @[MemPrimitives.scala 110:228:@9694.4]
  wire  _T_820; // @[MemPrimitives.scala 110:210:@9697.4]
  wire  _T_821; // @[MemPrimitives.scala 110:228:@9698.4]
  wire  _T_826; // @[MemPrimitives.scala 110:210:@9701.4]
  wire  _T_827; // @[MemPrimitives.scala 110:228:@9702.4]
  wire  _T_832; // @[MemPrimitives.scala 110:210:@9705.4]
  wire  _T_833; // @[MemPrimitives.scala 110:228:@9706.4]
  wire  _T_838; // @[MemPrimitives.scala 110:210:@9709.4]
  wire  _T_839; // @[MemPrimitives.scala 110:228:@9710.4]
  wire  _T_841; // @[MemPrimitives.scala 123:41:@9721.4]
  wire  _T_842; // @[MemPrimitives.scala 123:41:@9722.4]
  wire  _T_843; // @[MemPrimitives.scala 123:41:@9723.4]
  wire  _T_844; // @[MemPrimitives.scala 123:41:@9724.4]
  wire  _T_845; // @[MemPrimitives.scala 123:41:@9725.4]
  wire  _T_846; // @[MemPrimitives.scala 123:41:@9726.4]
  wire [2:0] _T_848; // @[Cat.scala 30:58:@9728.4]
  wire [2:0] _T_850; // @[Cat.scala 30:58:@9730.4]
  wire [2:0] _T_852; // @[Cat.scala 30:58:@9732.4]
  wire [2:0] _T_854; // @[Cat.scala 30:58:@9734.4]
  wire [2:0] _T_856; // @[Cat.scala 30:58:@9736.4]
  wire [2:0] _T_858; // @[Cat.scala 30:58:@9738.4]
  wire [2:0] _T_859; // @[Mux.scala 31:69:@9739.4]
  wire [2:0] _T_860; // @[Mux.scala 31:69:@9740.4]
  wire [2:0] _T_861; // @[Mux.scala 31:69:@9741.4]
  wire [2:0] _T_862; // @[Mux.scala 31:69:@9742.4]
  wire [2:0] _T_863; // @[Mux.scala 31:69:@9743.4]
  wire  _T_868; // @[MemPrimitives.scala 110:210:@9750.4]
  wire  _T_871; // @[MemPrimitives.scala 110:228:@9752.4]
  wire  _T_874; // @[MemPrimitives.scala 110:210:@9754.4]
  wire  _T_877; // @[MemPrimitives.scala 110:228:@9756.4]
  wire  _T_880; // @[MemPrimitives.scala 110:210:@9758.4]
  wire  _T_883; // @[MemPrimitives.scala 110:228:@9760.4]
  wire  _T_886; // @[MemPrimitives.scala 110:210:@9762.4]
  wire  _T_889; // @[MemPrimitives.scala 110:228:@9764.4]
  wire  _T_892; // @[MemPrimitives.scala 110:210:@9766.4]
  wire  _T_895; // @[MemPrimitives.scala 110:228:@9768.4]
  wire  _T_898; // @[MemPrimitives.scala 110:210:@9770.4]
  wire  _T_901; // @[MemPrimitives.scala 110:228:@9772.4]
  wire  _T_903; // @[MemPrimitives.scala 123:41:@9783.4]
  wire  _T_904; // @[MemPrimitives.scala 123:41:@9784.4]
  wire  _T_905; // @[MemPrimitives.scala 123:41:@9785.4]
  wire  _T_906; // @[MemPrimitives.scala 123:41:@9786.4]
  wire  _T_907; // @[MemPrimitives.scala 123:41:@9787.4]
  wire  _T_908; // @[MemPrimitives.scala 123:41:@9788.4]
  wire [2:0] _T_910; // @[Cat.scala 30:58:@9790.4]
  wire [2:0] _T_912; // @[Cat.scala 30:58:@9792.4]
  wire [2:0] _T_914; // @[Cat.scala 30:58:@9794.4]
  wire [2:0] _T_916; // @[Cat.scala 30:58:@9796.4]
  wire [2:0] _T_918; // @[Cat.scala 30:58:@9798.4]
  wire [2:0] _T_920; // @[Cat.scala 30:58:@9800.4]
  wire [2:0] _T_921; // @[Mux.scala 31:69:@9801.4]
  wire [2:0] _T_922; // @[Mux.scala 31:69:@9802.4]
  wire [2:0] _T_923; // @[Mux.scala 31:69:@9803.4]
  wire [2:0] _T_924; // @[Mux.scala 31:69:@9804.4]
  wire [2:0] _T_925; // @[Mux.scala 31:69:@9805.4]
  wire  _T_930; // @[MemPrimitives.scala 110:210:@9812.4]
  wire  _T_933; // @[MemPrimitives.scala 110:228:@9814.4]
  wire  _T_936; // @[MemPrimitives.scala 110:210:@9816.4]
  wire  _T_939; // @[MemPrimitives.scala 110:228:@9818.4]
  wire  _T_942; // @[MemPrimitives.scala 110:210:@9820.4]
  wire  _T_945; // @[MemPrimitives.scala 110:228:@9822.4]
  wire  _T_948; // @[MemPrimitives.scala 110:210:@9824.4]
  wire  _T_951; // @[MemPrimitives.scala 110:228:@9826.4]
  wire  _T_954; // @[MemPrimitives.scala 110:210:@9828.4]
  wire  _T_957; // @[MemPrimitives.scala 110:228:@9830.4]
  wire  _T_960; // @[MemPrimitives.scala 110:210:@9832.4]
  wire  _T_963; // @[MemPrimitives.scala 110:228:@9834.4]
  wire  _T_965; // @[MemPrimitives.scala 123:41:@9845.4]
  wire  _T_966; // @[MemPrimitives.scala 123:41:@9846.4]
  wire  _T_967; // @[MemPrimitives.scala 123:41:@9847.4]
  wire  _T_968; // @[MemPrimitives.scala 123:41:@9848.4]
  wire  _T_969; // @[MemPrimitives.scala 123:41:@9849.4]
  wire  _T_970; // @[MemPrimitives.scala 123:41:@9850.4]
  wire [2:0] _T_972; // @[Cat.scala 30:58:@9852.4]
  wire [2:0] _T_974; // @[Cat.scala 30:58:@9854.4]
  wire [2:0] _T_976; // @[Cat.scala 30:58:@9856.4]
  wire [2:0] _T_978; // @[Cat.scala 30:58:@9858.4]
  wire [2:0] _T_980; // @[Cat.scala 30:58:@9860.4]
  wire [2:0] _T_982; // @[Cat.scala 30:58:@9862.4]
  wire [2:0] _T_983; // @[Mux.scala 31:69:@9863.4]
  wire [2:0] _T_984; // @[Mux.scala 31:69:@9864.4]
  wire [2:0] _T_985; // @[Mux.scala 31:69:@9865.4]
  wire [2:0] _T_986; // @[Mux.scala 31:69:@9866.4]
  wire [2:0] _T_987; // @[Mux.scala 31:69:@9867.4]
  wire  _T_995; // @[MemPrimitives.scala 110:228:@9876.4]
  wire  _T_1001; // @[MemPrimitives.scala 110:228:@9880.4]
  wire  _T_1007; // @[MemPrimitives.scala 110:228:@9884.4]
  wire  _T_1013; // @[MemPrimitives.scala 110:228:@9888.4]
  wire  _T_1019; // @[MemPrimitives.scala 110:228:@9892.4]
  wire  _T_1025; // @[MemPrimitives.scala 110:228:@9896.4]
  wire  _T_1027; // @[MemPrimitives.scala 123:41:@9907.4]
  wire  _T_1028; // @[MemPrimitives.scala 123:41:@9908.4]
  wire  _T_1029; // @[MemPrimitives.scala 123:41:@9909.4]
  wire  _T_1030; // @[MemPrimitives.scala 123:41:@9910.4]
  wire  _T_1031; // @[MemPrimitives.scala 123:41:@9911.4]
  wire  _T_1032; // @[MemPrimitives.scala 123:41:@9912.4]
  wire [2:0] _T_1034; // @[Cat.scala 30:58:@9914.4]
  wire [2:0] _T_1036; // @[Cat.scala 30:58:@9916.4]
  wire [2:0] _T_1038; // @[Cat.scala 30:58:@9918.4]
  wire [2:0] _T_1040; // @[Cat.scala 30:58:@9920.4]
  wire [2:0] _T_1042; // @[Cat.scala 30:58:@9922.4]
  wire [2:0] _T_1044; // @[Cat.scala 30:58:@9924.4]
  wire [2:0] _T_1045; // @[Mux.scala 31:69:@9925.4]
  wire [2:0] _T_1046; // @[Mux.scala 31:69:@9926.4]
  wire [2:0] _T_1047; // @[Mux.scala 31:69:@9927.4]
  wire [2:0] _T_1048; // @[Mux.scala 31:69:@9928.4]
  wire [2:0] _T_1049; // @[Mux.scala 31:69:@9929.4]
  wire  _T_1057; // @[MemPrimitives.scala 110:228:@9938.4]
  wire  _T_1063; // @[MemPrimitives.scala 110:228:@9942.4]
  wire  _T_1069; // @[MemPrimitives.scala 110:228:@9946.4]
  wire  _T_1075; // @[MemPrimitives.scala 110:228:@9950.4]
  wire  _T_1081; // @[MemPrimitives.scala 110:228:@9954.4]
  wire  _T_1087; // @[MemPrimitives.scala 110:228:@9958.4]
  wire  _T_1089; // @[MemPrimitives.scala 123:41:@9969.4]
  wire  _T_1090; // @[MemPrimitives.scala 123:41:@9970.4]
  wire  _T_1091; // @[MemPrimitives.scala 123:41:@9971.4]
  wire  _T_1092; // @[MemPrimitives.scala 123:41:@9972.4]
  wire  _T_1093; // @[MemPrimitives.scala 123:41:@9973.4]
  wire  _T_1094; // @[MemPrimitives.scala 123:41:@9974.4]
  wire [2:0] _T_1096; // @[Cat.scala 30:58:@9976.4]
  wire [2:0] _T_1098; // @[Cat.scala 30:58:@9978.4]
  wire [2:0] _T_1100; // @[Cat.scala 30:58:@9980.4]
  wire [2:0] _T_1102; // @[Cat.scala 30:58:@9982.4]
  wire [2:0] _T_1104; // @[Cat.scala 30:58:@9984.4]
  wire [2:0] _T_1106; // @[Cat.scala 30:58:@9986.4]
  wire [2:0] _T_1107; // @[Mux.scala 31:69:@9987.4]
  wire [2:0] _T_1108; // @[Mux.scala 31:69:@9988.4]
  wire [2:0] _T_1109; // @[Mux.scala 31:69:@9989.4]
  wire [2:0] _T_1110; // @[Mux.scala 31:69:@9990.4]
  wire [2:0] _T_1111; // @[Mux.scala 31:69:@9991.4]
  wire  _T_1116; // @[MemPrimitives.scala 110:210:@9998.4]
  wire  _T_1119; // @[MemPrimitives.scala 110:228:@10000.4]
  wire  _T_1122; // @[MemPrimitives.scala 110:210:@10002.4]
  wire  _T_1125; // @[MemPrimitives.scala 110:228:@10004.4]
  wire  _T_1128; // @[MemPrimitives.scala 110:210:@10006.4]
  wire  _T_1131; // @[MemPrimitives.scala 110:228:@10008.4]
  wire  _T_1134; // @[MemPrimitives.scala 110:210:@10010.4]
  wire  _T_1137; // @[MemPrimitives.scala 110:228:@10012.4]
  wire  _T_1140; // @[MemPrimitives.scala 110:210:@10014.4]
  wire  _T_1143; // @[MemPrimitives.scala 110:228:@10016.4]
  wire  _T_1146; // @[MemPrimitives.scala 110:210:@10018.4]
  wire  _T_1149; // @[MemPrimitives.scala 110:228:@10020.4]
  wire  _T_1151; // @[MemPrimitives.scala 123:41:@10031.4]
  wire  _T_1152; // @[MemPrimitives.scala 123:41:@10032.4]
  wire  _T_1153; // @[MemPrimitives.scala 123:41:@10033.4]
  wire  _T_1154; // @[MemPrimitives.scala 123:41:@10034.4]
  wire  _T_1155; // @[MemPrimitives.scala 123:41:@10035.4]
  wire  _T_1156; // @[MemPrimitives.scala 123:41:@10036.4]
  wire [2:0] _T_1158; // @[Cat.scala 30:58:@10038.4]
  wire [2:0] _T_1160; // @[Cat.scala 30:58:@10040.4]
  wire [2:0] _T_1162; // @[Cat.scala 30:58:@10042.4]
  wire [2:0] _T_1164; // @[Cat.scala 30:58:@10044.4]
  wire [2:0] _T_1166; // @[Cat.scala 30:58:@10046.4]
  wire [2:0] _T_1168; // @[Cat.scala 30:58:@10048.4]
  wire [2:0] _T_1169; // @[Mux.scala 31:69:@10049.4]
  wire [2:0] _T_1170; // @[Mux.scala 31:69:@10050.4]
  wire [2:0] _T_1171; // @[Mux.scala 31:69:@10051.4]
  wire [2:0] _T_1172; // @[Mux.scala 31:69:@10052.4]
  wire [2:0] _T_1173; // @[Mux.scala 31:69:@10053.4]
  wire  _T_1178; // @[MemPrimitives.scala 110:210:@10060.4]
  wire  _T_1181; // @[MemPrimitives.scala 110:228:@10062.4]
  wire  _T_1184; // @[MemPrimitives.scala 110:210:@10064.4]
  wire  _T_1187; // @[MemPrimitives.scala 110:228:@10066.4]
  wire  _T_1190; // @[MemPrimitives.scala 110:210:@10068.4]
  wire  _T_1193; // @[MemPrimitives.scala 110:228:@10070.4]
  wire  _T_1196; // @[MemPrimitives.scala 110:210:@10072.4]
  wire  _T_1199; // @[MemPrimitives.scala 110:228:@10074.4]
  wire  _T_1202; // @[MemPrimitives.scala 110:210:@10076.4]
  wire  _T_1205; // @[MemPrimitives.scala 110:228:@10078.4]
  wire  _T_1208; // @[MemPrimitives.scala 110:210:@10080.4]
  wire  _T_1211; // @[MemPrimitives.scala 110:228:@10082.4]
  wire  _T_1213; // @[MemPrimitives.scala 123:41:@10093.4]
  wire  _T_1214; // @[MemPrimitives.scala 123:41:@10094.4]
  wire  _T_1215; // @[MemPrimitives.scala 123:41:@10095.4]
  wire  _T_1216; // @[MemPrimitives.scala 123:41:@10096.4]
  wire  _T_1217; // @[MemPrimitives.scala 123:41:@10097.4]
  wire  _T_1218; // @[MemPrimitives.scala 123:41:@10098.4]
  wire [2:0] _T_1220; // @[Cat.scala 30:58:@10100.4]
  wire [2:0] _T_1222; // @[Cat.scala 30:58:@10102.4]
  wire [2:0] _T_1224; // @[Cat.scala 30:58:@10104.4]
  wire [2:0] _T_1226; // @[Cat.scala 30:58:@10106.4]
  wire [2:0] _T_1228; // @[Cat.scala 30:58:@10108.4]
  wire [2:0] _T_1230; // @[Cat.scala 30:58:@10110.4]
  wire [2:0] _T_1231; // @[Mux.scala 31:69:@10111.4]
  wire [2:0] _T_1232; // @[Mux.scala 31:69:@10112.4]
  wire [2:0] _T_1233; // @[Mux.scala 31:69:@10113.4]
  wire [2:0] _T_1234; // @[Mux.scala 31:69:@10114.4]
  wire [2:0] _T_1235; // @[Mux.scala 31:69:@10115.4]
  wire  _T_1243; // @[MemPrimitives.scala 110:228:@10124.4]
  wire  _T_1249; // @[MemPrimitives.scala 110:228:@10128.4]
  wire  _T_1255; // @[MemPrimitives.scala 110:228:@10132.4]
  wire  _T_1261; // @[MemPrimitives.scala 110:228:@10136.4]
  wire  _T_1267; // @[MemPrimitives.scala 110:228:@10140.4]
  wire  _T_1273; // @[MemPrimitives.scala 110:228:@10144.4]
  wire  _T_1275; // @[MemPrimitives.scala 123:41:@10155.4]
  wire  _T_1276; // @[MemPrimitives.scala 123:41:@10156.4]
  wire  _T_1277; // @[MemPrimitives.scala 123:41:@10157.4]
  wire  _T_1278; // @[MemPrimitives.scala 123:41:@10158.4]
  wire  _T_1279; // @[MemPrimitives.scala 123:41:@10159.4]
  wire  _T_1280; // @[MemPrimitives.scala 123:41:@10160.4]
  wire [2:0] _T_1282; // @[Cat.scala 30:58:@10162.4]
  wire [2:0] _T_1284; // @[Cat.scala 30:58:@10164.4]
  wire [2:0] _T_1286; // @[Cat.scala 30:58:@10166.4]
  wire [2:0] _T_1288; // @[Cat.scala 30:58:@10168.4]
  wire [2:0] _T_1290; // @[Cat.scala 30:58:@10170.4]
  wire [2:0] _T_1292; // @[Cat.scala 30:58:@10172.4]
  wire [2:0] _T_1293; // @[Mux.scala 31:69:@10173.4]
  wire [2:0] _T_1294; // @[Mux.scala 31:69:@10174.4]
  wire [2:0] _T_1295; // @[Mux.scala 31:69:@10175.4]
  wire [2:0] _T_1296; // @[Mux.scala 31:69:@10176.4]
  wire [2:0] _T_1297; // @[Mux.scala 31:69:@10177.4]
  wire  _T_1305; // @[MemPrimitives.scala 110:228:@10186.4]
  wire  _T_1311; // @[MemPrimitives.scala 110:228:@10190.4]
  wire  _T_1317; // @[MemPrimitives.scala 110:228:@10194.4]
  wire  _T_1323; // @[MemPrimitives.scala 110:228:@10198.4]
  wire  _T_1329; // @[MemPrimitives.scala 110:228:@10202.4]
  wire  _T_1335; // @[MemPrimitives.scala 110:228:@10206.4]
  wire  _T_1337; // @[MemPrimitives.scala 123:41:@10217.4]
  wire  _T_1338; // @[MemPrimitives.scala 123:41:@10218.4]
  wire  _T_1339; // @[MemPrimitives.scala 123:41:@10219.4]
  wire  _T_1340; // @[MemPrimitives.scala 123:41:@10220.4]
  wire  _T_1341; // @[MemPrimitives.scala 123:41:@10221.4]
  wire  _T_1342; // @[MemPrimitives.scala 123:41:@10222.4]
  wire [2:0] _T_1344; // @[Cat.scala 30:58:@10224.4]
  wire [2:0] _T_1346; // @[Cat.scala 30:58:@10226.4]
  wire [2:0] _T_1348; // @[Cat.scala 30:58:@10228.4]
  wire [2:0] _T_1350; // @[Cat.scala 30:58:@10230.4]
  wire [2:0] _T_1352; // @[Cat.scala 30:58:@10232.4]
  wire [2:0] _T_1354; // @[Cat.scala 30:58:@10234.4]
  wire [2:0] _T_1355; // @[Mux.scala 31:69:@10235.4]
  wire [2:0] _T_1356; // @[Mux.scala 31:69:@10236.4]
  wire [2:0] _T_1357; // @[Mux.scala 31:69:@10237.4]
  wire [2:0] _T_1358; // @[Mux.scala 31:69:@10238.4]
  wire [2:0] _T_1359; // @[Mux.scala 31:69:@10239.4]
  wire  _T_1364; // @[MemPrimitives.scala 110:210:@10246.4]
  wire  _T_1367; // @[MemPrimitives.scala 110:228:@10248.4]
  wire  _T_1370; // @[MemPrimitives.scala 110:210:@10250.4]
  wire  _T_1373; // @[MemPrimitives.scala 110:228:@10252.4]
  wire  _T_1376; // @[MemPrimitives.scala 110:210:@10254.4]
  wire  _T_1379; // @[MemPrimitives.scala 110:228:@10256.4]
  wire  _T_1382; // @[MemPrimitives.scala 110:210:@10258.4]
  wire  _T_1385; // @[MemPrimitives.scala 110:228:@10260.4]
  wire  _T_1388; // @[MemPrimitives.scala 110:210:@10262.4]
  wire  _T_1391; // @[MemPrimitives.scala 110:228:@10264.4]
  wire  _T_1394; // @[MemPrimitives.scala 110:210:@10266.4]
  wire  _T_1397; // @[MemPrimitives.scala 110:228:@10268.4]
  wire  _T_1399; // @[MemPrimitives.scala 123:41:@10279.4]
  wire  _T_1400; // @[MemPrimitives.scala 123:41:@10280.4]
  wire  _T_1401; // @[MemPrimitives.scala 123:41:@10281.4]
  wire  _T_1402; // @[MemPrimitives.scala 123:41:@10282.4]
  wire  _T_1403; // @[MemPrimitives.scala 123:41:@10283.4]
  wire  _T_1404; // @[MemPrimitives.scala 123:41:@10284.4]
  wire [2:0] _T_1406; // @[Cat.scala 30:58:@10286.4]
  wire [2:0] _T_1408; // @[Cat.scala 30:58:@10288.4]
  wire [2:0] _T_1410; // @[Cat.scala 30:58:@10290.4]
  wire [2:0] _T_1412; // @[Cat.scala 30:58:@10292.4]
  wire [2:0] _T_1414; // @[Cat.scala 30:58:@10294.4]
  wire [2:0] _T_1416; // @[Cat.scala 30:58:@10296.4]
  wire [2:0] _T_1417; // @[Mux.scala 31:69:@10297.4]
  wire [2:0] _T_1418; // @[Mux.scala 31:69:@10298.4]
  wire [2:0] _T_1419; // @[Mux.scala 31:69:@10299.4]
  wire [2:0] _T_1420; // @[Mux.scala 31:69:@10300.4]
  wire [2:0] _T_1421; // @[Mux.scala 31:69:@10301.4]
  wire  _T_1426; // @[MemPrimitives.scala 110:210:@10308.4]
  wire  _T_1429; // @[MemPrimitives.scala 110:228:@10310.4]
  wire  _T_1432; // @[MemPrimitives.scala 110:210:@10312.4]
  wire  _T_1435; // @[MemPrimitives.scala 110:228:@10314.4]
  wire  _T_1438; // @[MemPrimitives.scala 110:210:@10316.4]
  wire  _T_1441; // @[MemPrimitives.scala 110:228:@10318.4]
  wire  _T_1444; // @[MemPrimitives.scala 110:210:@10320.4]
  wire  _T_1447; // @[MemPrimitives.scala 110:228:@10322.4]
  wire  _T_1450; // @[MemPrimitives.scala 110:210:@10324.4]
  wire  _T_1453; // @[MemPrimitives.scala 110:228:@10326.4]
  wire  _T_1456; // @[MemPrimitives.scala 110:210:@10328.4]
  wire  _T_1459; // @[MemPrimitives.scala 110:228:@10330.4]
  wire  _T_1461; // @[MemPrimitives.scala 123:41:@10341.4]
  wire  _T_1462; // @[MemPrimitives.scala 123:41:@10342.4]
  wire  _T_1463; // @[MemPrimitives.scala 123:41:@10343.4]
  wire  _T_1464; // @[MemPrimitives.scala 123:41:@10344.4]
  wire  _T_1465; // @[MemPrimitives.scala 123:41:@10345.4]
  wire  _T_1466; // @[MemPrimitives.scala 123:41:@10346.4]
  wire [2:0] _T_1468; // @[Cat.scala 30:58:@10348.4]
  wire [2:0] _T_1470; // @[Cat.scala 30:58:@10350.4]
  wire [2:0] _T_1472; // @[Cat.scala 30:58:@10352.4]
  wire [2:0] _T_1474; // @[Cat.scala 30:58:@10354.4]
  wire [2:0] _T_1476; // @[Cat.scala 30:58:@10356.4]
  wire [2:0] _T_1478; // @[Cat.scala 30:58:@10358.4]
  wire [2:0] _T_1479; // @[Mux.scala 31:69:@10359.4]
  wire [2:0] _T_1480; // @[Mux.scala 31:69:@10360.4]
  wire [2:0] _T_1481; // @[Mux.scala 31:69:@10361.4]
  wire [2:0] _T_1482; // @[Mux.scala 31:69:@10362.4]
  wire [2:0] _T_1483; // @[Mux.scala 31:69:@10363.4]
  wire  _T_1491; // @[MemPrimitives.scala 110:228:@10372.4]
  wire  _T_1497; // @[MemPrimitives.scala 110:228:@10376.4]
  wire  _T_1503; // @[MemPrimitives.scala 110:228:@10380.4]
  wire  _T_1509; // @[MemPrimitives.scala 110:228:@10384.4]
  wire  _T_1515; // @[MemPrimitives.scala 110:228:@10388.4]
  wire  _T_1521; // @[MemPrimitives.scala 110:228:@10392.4]
  wire  _T_1523; // @[MemPrimitives.scala 123:41:@10403.4]
  wire  _T_1524; // @[MemPrimitives.scala 123:41:@10404.4]
  wire  _T_1525; // @[MemPrimitives.scala 123:41:@10405.4]
  wire  _T_1526; // @[MemPrimitives.scala 123:41:@10406.4]
  wire  _T_1527; // @[MemPrimitives.scala 123:41:@10407.4]
  wire  _T_1528; // @[MemPrimitives.scala 123:41:@10408.4]
  wire [2:0] _T_1530; // @[Cat.scala 30:58:@10410.4]
  wire [2:0] _T_1532; // @[Cat.scala 30:58:@10412.4]
  wire [2:0] _T_1534; // @[Cat.scala 30:58:@10414.4]
  wire [2:0] _T_1536; // @[Cat.scala 30:58:@10416.4]
  wire [2:0] _T_1538; // @[Cat.scala 30:58:@10418.4]
  wire [2:0] _T_1540; // @[Cat.scala 30:58:@10420.4]
  wire [2:0] _T_1541; // @[Mux.scala 31:69:@10421.4]
  wire [2:0] _T_1542; // @[Mux.scala 31:69:@10422.4]
  wire [2:0] _T_1543; // @[Mux.scala 31:69:@10423.4]
  wire [2:0] _T_1544; // @[Mux.scala 31:69:@10424.4]
  wire [2:0] _T_1545; // @[Mux.scala 31:69:@10425.4]
  wire  _T_1553; // @[MemPrimitives.scala 110:228:@10434.4]
  wire  _T_1559; // @[MemPrimitives.scala 110:228:@10438.4]
  wire  _T_1565; // @[MemPrimitives.scala 110:228:@10442.4]
  wire  _T_1571; // @[MemPrimitives.scala 110:228:@10446.4]
  wire  _T_1577; // @[MemPrimitives.scala 110:228:@10450.4]
  wire  _T_1583; // @[MemPrimitives.scala 110:228:@10454.4]
  wire  _T_1585; // @[MemPrimitives.scala 123:41:@10465.4]
  wire  _T_1586; // @[MemPrimitives.scala 123:41:@10466.4]
  wire  _T_1587; // @[MemPrimitives.scala 123:41:@10467.4]
  wire  _T_1588; // @[MemPrimitives.scala 123:41:@10468.4]
  wire  _T_1589; // @[MemPrimitives.scala 123:41:@10469.4]
  wire  _T_1590; // @[MemPrimitives.scala 123:41:@10470.4]
  wire [2:0] _T_1592; // @[Cat.scala 30:58:@10472.4]
  wire [2:0] _T_1594; // @[Cat.scala 30:58:@10474.4]
  wire [2:0] _T_1596; // @[Cat.scala 30:58:@10476.4]
  wire [2:0] _T_1598; // @[Cat.scala 30:58:@10478.4]
  wire [2:0] _T_1600; // @[Cat.scala 30:58:@10480.4]
  wire [2:0] _T_1602; // @[Cat.scala 30:58:@10482.4]
  wire [2:0] _T_1603; // @[Mux.scala 31:69:@10483.4]
  wire [2:0] _T_1604; // @[Mux.scala 31:69:@10484.4]
  wire [2:0] _T_1605; // @[Mux.scala 31:69:@10485.4]
  wire [2:0] _T_1606; // @[Mux.scala 31:69:@10486.4]
  wire [2:0] _T_1607; // @[Mux.scala 31:69:@10487.4]
  wire  _T_1671; // @[package.scala 96:25:@10572.4 package.scala 96:25:@10573.4]
  wire [7:0] _T_1675; // @[Mux.scala 31:69:@10582.4]
  wire  _T_1668; // @[package.scala 96:25:@10564.4 package.scala 96:25:@10565.4]
  wire [7:0] _T_1676; // @[Mux.scala 31:69:@10583.4]
  wire  _T_1665; // @[package.scala 96:25:@10556.4 package.scala 96:25:@10557.4]
  wire [7:0] _T_1677; // @[Mux.scala 31:69:@10584.4]
  wire  _T_1662; // @[package.scala 96:25:@10548.4 package.scala 96:25:@10549.4]
  wire [7:0] _T_1678; // @[Mux.scala 31:69:@10585.4]
  wire  _T_1659; // @[package.scala 96:25:@10540.4 package.scala 96:25:@10541.4]
  wire [7:0] _T_1679; // @[Mux.scala 31:69:@10586.4]
  wire  _T_1656; // @[package.scala 96:25:@10532.4 package.scala 96:25:@10533.4]
  wire [7:0] _T_1680; // @[Mux.scala 31:69:@10587.4]
  wire  _T_1653; // @[package.scala 96:25:@10524.4 package.scala 96:25:@10525.4]
  wire  _T_1742; // @[package.scala 96:25:@10668.4 package.scala 96:25:@10669.4]
  wire [7:0] _T_1746; // @[Mux.scala 31:69:@10678.4]
  wire  _T_1739; // @[package.scala 96:25:@10660.4 package.scala 96:25:@10661.4]
  wire [7:0] _T_1747; // @[Mux.scala 31:69:@10679.4]
  wire  _T_1736; // @[package.scala 96:25:@10652.4 package.scala 96:25:@10653.4]
  wire [7:0] _T_1748; // @[Mux.scala 31:69:@10680.4]
  wire  _T_1733; // @[package.scala 96:25:@10644.4 package.scala 96:25:@10645.4]
  wire [7:0] _T_1749; // @[Mux.scala 31:69:@10681.4]
  wire  _T_1730; // @[package.scala 96:25:@10636.4 package.scala 96:25:@10637.4]
  wire [7:0] _T_1750; // @[Mux.scala 31:69:@10682.4]
  wire  _T_1727; // @[package.scala 96:25:@10628.4 package.scala 96:25:@10629.4]
  wire [7:0] _T_1751; // @[Mux.scala 31:69:@10683.4]
  wire  _T_1724; // @[package.scala 96:25:@10620.4 package.scala 96:25:@10621.4]
  wire  _T_1813; // @[package.scala 96:25:@10764.4 package.scala 96:25:@10765.4]
  wire [7:0] _T_1817; // @[Mux.scala 31:69:@10774.4]
  wire  _T_1810; // @[package.scala 96:25:@10756.4 package.scala 96:25:@10757.4]
  wire [7:0] _T_1818; // @[Mux.scala 31:69:@10775.4]
  wire  _T_1807; // @[package.scala 96:25:@10748.4 package.scala 96:25:@10749.4]
  wire [7:0] _T_1819; // @[Mux.scala 31:69:@10776.4]
  wire  _T_1804; // @[package.scala 96:25:@10740.4 package.scala 96:25:@10741.4]
  wire [7:0] _T_1820; // @[Mux.scala 31:69:@10777.4]
  wire  _T_1801; // @[package.scala 96:25:@10732.4 package.scala 96:25:@10733.4]
  wire [7:0] _T_1821; // @[Mux.scala 31:69:@10778.4]
  wire  _T_1798; // @[package.scala 96:25:@10724.4 package.scala 96:25:@10725.4]
  wire [7:0] _T_1822; // @[Mux.scala 31:69:@10779.4]
  wire  _T_1795; // @[package.scala 96:25:@10716.4 package.scala 96:25:@10717.4]
  wire  _T_1884; // @[package.scala 96:25:@10860.4 package.scala 96:25:@10861.4]
  wire [7:0] _T_1888; // @[Mux.scala 31:69:@10870.4]
  wire  _T_1881; // @[package.scala 96:25:@10852.4 package.scala 96:25:@10853.4]
  wire [7:0] _T_1889; // @[Mux.scala 31:69:@10871.4]
  wire  _T_1878; // @[package.scala 96:25:@10844.4 package.scala 96:25:@10845.4]
  wire [7:0] _T_1890; // @[Mux.scala 31:69:@10872.4]
  wire  _T_1875; // @[package.scala 96:25:@10836.4 package.scala 96:25:@10837.4]
  wire [7:0] _T_1891; // @[Mux.scala 31:69:@10873.4]
  wire  _T_1872; // @[package.scala 96:25:@10828.4 package.scala 96:25:@10829.4]
  wire [7:0] _T_1892; // @[Mux.scala 31:69:@10874.4]
  wire  _T_1869; // @[package.scala 96:25:@10820.4 package.scala 96:25:@10821.4]
  wire [7:0] _T_1893; // @[Mux.scala 31:69:@10875.4]
  wire  _T_1866; // @[package.scala 96:25:@10812.4 package.scala 96:25:@10813.4]
  wire  _T_1955; // @[package.scala 96:25:@10956.4 package.scala 96:25:@10957.4]
  wire [7:0] _T_1959; // @[Mux.scala 31:69:@10966.4]
  wire  _T_1952; // @[package.scala 96:25:@10948.4 package.scala 96:25:@10949.4]
  wire [7:0] _T_1960; // @[Mux.scala 31:69:@10967.4]
  wire  _T_1949; // @[package.scala 96:25:@10940.4 package.scala 96:25:@10941.4]
  wire [7:0] _T_1961; // @[Mux.scala 31:69:@10968.4]
  wire  _T_1946; // @[package.scala 96:25:@10932.4 package.scala 96:25:@10933.4]
  wire [7:0] _T_1962; // @[Mux.scala 31:69:@10969.4]
  wire  _T_1943; // @[package.scala 96:25:@10924.4 package.scala 96:25:@10925.4]
  wire [7:0] _T_1963; // @[Mux.scala 31:69:@10970.4]
  wire  _T_1940; // @[package.scala 96:25:@10916.4 package.scala 96:25:@10917.4]
  wire [7:0] _T_1964; // @[Mux.scala 31:69:@10971.4]
  wire  _T_1937; // @[package.scala 96:25:@10908.4 package.scala 96:25:@10909.4]
  wire  _T_2026; // @[package.scala 96:25:@11052.4 package.scala 96:25:@11053.4]
  wire [7:0] _T_2030; // @[Mux.scala 31:69:@11062.4]
  wire  _T_2023; // @[package.scala 96:25:@11044.4 package.scala 96:25:@11045.4]
  wire [7:0] _T_2031; // @[Mux.scala 31:69:@11063.4]
  wire  _T_2020; // @[package.scala 96:25:@11036.4 package.scala 96:25:@11037.4]
  wire [7:0] _T_2032; // @[Mux.scala 31:69:@11064.4]
  wire  _T_2017; // @[package.scala 96:25:@11028.4 package.scala 96:25:@11029.4]
  wire [7:0] _T_2033; // @[Mux.scala 31:69:@11065.4]
  wire  _T_2014; // @[package.scala 96:25:@11020.4 package.scala 96:25:@11021.4]
  wire [7:0] _T_2034; // @[Mux.scala 31:69:@11066.4]
  wire  _T_2011; // @[package.scala 96:25:@11012.4 package.scala 96:25:@11013.4]
  wire [7:0] _T_2035; // @[Mux.scala 31:69:@11067.4]
  wire  _T_2008; // @[package.scala 96:25:@11004.4 package.scala 96:25:@11005.4]
  wire  _T_2097; // @[package.scala 96:25:@11148.4 package.scala 96:25:@11149.4]
  wire [7:0] _T_2101; // @[Mux.scala 31:69:@11158.4]
  wire  _T_2094; // @[package.scala 96:25:@11140.4 package.scala 96:25:@11141.4]
  wire [7:0] _T_2102; // @[Mux.scala 31:69:@11159.4]
  wire  _T_2091; // @[package.scala 96:25:@11132.4 package.scala 96:25:@11133.4]
  wire [7:0] _T_2103; // @[Mux.scala 31:69:@11160.4]
  wire  _T_2088; // @[package.scala 96:25:@11124.4 package.scala 96:25:@11125.4]
  wire [7:0] _T_2104; // @[Mux.scala 31:69:@11161.4]
  wire  _T_2085; // @[package.scala 96:25:@11116.4 package.scala 96:25:@11117.4]
  wire [7:0] _T_2105; // @[Mux.scala 31:69:@11162.4]
  wire  _T_2082; // @[package.scala 96:25:@11108.4 package.scala 96:25:@11109.4]
  wire [7:0] _T_2106; // @[Mux.scala 31:69:@11163.4]
  wire  _T_2079; // @[package.scala 96:25:@11100.4 package.scala 96:25:@11101.4]
  wire  _T_2168; // @[package.scala 96:25:@11244.4 package.scala 96:25:@11245.4]
  wire [7:0] _T_2172; // @[Mux.scala 31:69:@11254.4]
  wire  _T_2165; // @[package.scala 96:25:@11236.4 package.scala 96:25:@11237.4]
  wire [7:0] _T_2173; // @[Mux.scala 31:69:@11255.4]
  wire  _T_2162; // @[package.scala 96:25:@11228.4 package.scala 96:25:@11229.4]
  wire [7:0] _T_2174; // @[Mux.scala 31:69:@11256.4]
  wire  _T_2159; // @[package.scala 96:25:@11220.4 package.scala 96:25:@11221.4]
  wire [7:0] _T_2175; // @[Mux.scala 31:69:@11257.4]
  wire  _T_2156; // @[package.scala 96:25:@11212.4 package.scala 96:25:@11213.4]
  wire [7:0] _T_2176; // @[Mux.scala 31:69:@11258.4]
  wire  _T_2153; // @[package.scala 96:25:@11204.4 package.scala 96:25:@11205.4]
  wire [7:0] _T_2177; // @[Mux.scala 31:69:@11259.4]
  wire  _T_2150; // @[package.scala 96:25:@11196.4 package.scala 96:25:@11197.4]
  wire  _T_2239; // @[package.scala 96:25:@11340.4 package.scala 96:25:@11341.4]
  wire [7:0] _T_2243; // @[Mux.scala 31:69:@11350.4]
  wire  _T_2236; // @[package.scala 96:25:@11332.4 package.scala 96:25:@11333.4]
  wire [7:0] _T_2244; // @[Mux.scala 31:69:@11351.4]
  wire  _T_2233; // @[package.scala 96:25:@11324.4 package.scala 96:25:@11325.4]
  wire [7:0] _T_2245; // @[Mux.scala 31:69:@11352.4]
  wire  _T_2230; // @[package.scala 96:25:@11316.4 package.scala 96:25:@11317.4]
  wire [7:0] _T_2246; // @[Mux.scala 31:69:@11353.4]
  wire  _T_2227; // @[package.scala 96:25:@11308.4 package.scala 96:25:@11309.4]
  wire [7:0] _T_2247; // @[Mux.scala 31:69:@11354.4]
  wire  _T_2224; // @[package.scala 96:25:@11300.4 package.scala 96:25:@11301.4]
  wire [7:0] _T_2248; // @[Mux.scala 31:69:@11355.4]
  wire  _T_2221; // @[package.scala 96:25:@11292.4 package.scala 96:25:@11293.4]
  wire  _T_2310; // @[package.scala 96:25:@11436.4 package.scala 96:25:@11437.4]
  wire [7:0] _T_2314; // @[Mux.scala 31:69:@11446.4]
  wire  _T_2307; // @[package.scala 96:25:@11428.4 package.scala 96:25:@11429.4]
  wire [7:0] _T_2315; // @[Mux.scala 31:69:@11447.4]
  wire  _T_2304; // @[package.scala 96:25:@11420.4 package.scala 96:25:@11421.4]
  wire [7:0] _T_2316; // @[Mux.scala 31:69:@11448.4]
  wire  _T_2301; // @[package.scala 96:25:@11412.4 package.scala 96:25:@11413.4]
  wire [7:0] _T_2317; // @[Mux.scala 31:69:@11449.4]
  wire  _T_2298; // @[package.scala 96:25:@11404.4 package.scala 96:25:@11405.4]
  wire [7:0] _T_2318; // @[Mux.scala 31:69:@11450.4]
  wire  _T_2295; // @[package.scala 96:25:@11396.4 package.scala 96:25:@11397.4]
  wire [7:0] _T_2319; // @[Mux.scala 31:69:@11451.4]
  wire  _T_2292; // @[package.scala 96:25:@11388.4 package.scala 96:25:@11389.4]
  wire  _T_2381; // @[package.scala 96:25:@11532.4 package.scala 96:25:@11533.4]
  wire [7:0] _T_2385; // @[Mux.scala 31:69:@11542.4]
  wire  _T_2378; // @[package.scala 96:25:@11524.4 package.scala 96:25:@11525.4]
  wire [7:0] _T_2386; // @[Mux.scala 31:69:@11543.4]
  wire  _T_2375; // @[package.scala 96:25:@11516.4 package.scala 96:25:@11517.4]
  wire [7:0] _T_2387; // @[Mux.scala 31:69:@11544.4]
  wire  _T_2372; // @[package.scala 96:25:@11508.4 package.scala 96:25:@11509.4]
  wire [7:0] _T_2388; // @[Mux.scala 31:69:@11545.4]
  wire  _T_2369; // @[package.scala 96:25:@11500.4 package.scala 96:25:@11501.4]
  wire [7:0] _T_2389; // @[Mux.scala 31:69:@11546.4]
  wire  _T_2366; // @[package.scala 96:25:@11492.4 package.scala 96:25:@11493.4]
  wire [7:0] _T_2390; // @[Mux.scala 31:69:@11547.4]
  wire  _T_2363; // @[package.scala 96:25:@11484.4 package.scala 96:25:@11485.4]
  wire  _T_2452; // @[package.scala 96:25:@11628.4 package.scala 96:25:@11629.4]
  wire [7:0] _T_2456; // @[Mux.scala 31:69:@11638.4]
  wire  _T_2449; // @[package.scala 96:25:@11620.4 package.scala 96:25:@11621.4]
  wire [7:0] _T_2457; // @[Mux.scala 31:69:@11639.4]
  wire  _T_2446; // @[package.scala 96:25:@11612.4 package.scala 96:25:@11613.4]
  wire [7:0] _T_2458; // @[Mux.scala 31:69:@11640.4]
  wire  _T_2443; // @[package.scala 96:25:@11604.4 package.scala 96:25:@11605.4]
  wire [7:0] _T_2459; // @[Mux.scala 31:69:@11641.4]
  wire  _T_2440; // @[package.scala 96:25:@11596.4 package.scala 96:25:@11597.4]
  wire [7:0] _T_2460; // @[Mux.scala 31:69:@11642.4]
  wire  _T_2437; // @[package.scala 96:25:@11588.4 package.scala 96:25:@11589.4]
  wire [7:0] _T_2461; // @[Mux.scala 31:69:@11643.4]
  wire  _T_2434; // @[package.scala 96:25:@11580.4 package.scala 96:25:@11581.4]
  Mem1D_4 Mem1D ( // @[MemPrimitives.scala 64:21:@9054.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  Mem1D_4 Mem1D_1 ( // @[MemPrimitives.scala 64:21:@9070.4]
    .clock(Mem1D_1_clock),
    .reset(Mem1D_1_reset),
    .io_r_ofs_0(Mem1D_1_io_r_ofs_0),
    .io_r_backpressure(Mem1D_1_io_r_backpressure),
    .io_w_ofs_0(Mem1D_1_io_w_ofs_0),
    .io_w_data_0(Mem1D_1_io_w_data_0),
    .io_w_en_0(Mem1D_1_io_w_en_0),
    .io_output(Mem1D_1_io_output)
  );
  Mem1D_4 Mem1D_2 ( // @[MemPrimitives.scala 64:21:@9086.4]
    .clock(Mem1D_2_clock),
    .reset(Mem1D_2_reset),
    .io_r_ofs_0(Mem1D_2_io_r_ofs_0),
    .io_r_backpressure(Mem1D_2_io_r_backpressure),
    .io_w_ofs_0(Mem1D_2_io_w_ofs_0),
    .io_w_data_0(Mem1D_2_io_w_data_0),
    .io_w_en_0(Mem1D_2_io_w_en_0),
    .io_output(Mem1D_2_io_output)
  );
  Mem1D_4 Mem1D_3 ( // @[MemPrimitives.scala 64:21:@9102.4]
    .clock(Mem1D_3_clock),
    .reset(Mem1D_3_reset),
    .io_r_ofs_0(Mem1D_3_io_r_ofs_0),
    .io_r_backpressure(Mem1D_3_io_r_backpressure),
    .io_w_ofs_0(Mem1D_3_io_w_ofs_0),
    .io_w_data_0(Mem1D_3_io_w_data_0),
    .io_w_en_0(Mem1D_3_io_w_en_0),
    .io_output(Mem1D_3_io_output)
  );
  Mem1D_4 Mem1D_4 ( // @[MemPrimitives.scala 64:21:@9118.4]
    .clock(Mem1D_4_clock),
    .reset(Mem1D_4_reset),
    .io_r_ofs_0(Mem1D_4_io_r_ofs_0),
    .io_r_backpressure(Mem1D_4_io_r_backpressure),
    .io_w_ofs_0(Mem1D_4_io_w_ofs_0),
    .io_w_data_0(Mem1D_4_io_w_data_0),
    .io_w_en_0(Mem1D_4_io_w_en_0),
    .io_output(Mem1D_4_io_output)
  );
  Mem1D_4 Mem1D_5 ( // @[MemPrimitives.scala 64:21:@9134.4]
    .clock(Mem1D_5_clock),
    .reset(Mem1D_5_reset),
    .io_r_ofs_0(Mem1D_5_io_r_ofs_0),
    .io_r_backpressure(Mem1D_5_io_r_backpressure),
    .io_w_ofs_0(Mem1D_5_io_w_ofs_0),
    .io_w_data_0(Mem1D_5_io_w_data_0),
    .io_w_en_0(Mem1D_5_io_w_en_0),
    .io_output(Mem1D_5_io_output)
  );
  Mem1D_4 Mem1D_6 ( // @[MemPrimitives.scala 64:21:@9150.4]
    .clock(Mem1D_6_clock),
    .reset(Mem1D_6_reset),
    .io_r_ofs_0(Mem1D_6_io_r_ofs_0),
    .io_r_backpressure(Mem1D_6_io_r_backpressure),
    .io_w_ofs_0(Mem1D_6_io_w_ofs_0),
    .io_w_data_0(Mem1D_6_io_w_data_0),
    .io_w_en_0(Mem1D_6_io_w_en_0),
    .io_output(Mem1D_6_io_output)
  );
  Mem1D_4 Mem1D_7 ( // @[MemPrimitives.scala 64:21:@9166.4]
    .clock(Mem1D_7_clock),
    .reset(Mem1D_7_reset),
    .io_r_ofs_0(Mem1D_7_io_r_ofs_0),
    .io_r_backpressure(Mem1D_7_io_r_backpressure),
    .io_w_ofs_0(Mem1D_7_io_w_ofs_0),
    .io_w_data_0(Mem1D_7_io_w_data_0),
    .io_w_en_0(Mem1D_7_io_w_en_0),
    .io_output(Mem1D_7_io_output)
  );
  Mem1D_4 Mem1D_8 ( // @[MemPrimitives.scala 64:21:@9182.4]
    .clock(Mem1D_8_clock),
    .reset(Mem1D_8_reset),
    .io_r_ofs_0(Mem1D_8_io_r_ofs_0),
    .io_r_backpressure(Mem1D_8_io_r_backpressure),
    .io_w_ofs_0(Mem1D_8_io_w_ofs_0),
    .io_w_data_0(Mem1D_8_io_w_data_0),
    .io_w_en_0(Mem1D_8_io_w_en_0),
    .io_output(Mem1D_8_io_output)
  );
  Mem1D_4 Mem1D_9 ( // @[MemPrimitives.scala 64:21:@9198.4]
    .clock(Mem1D_9_clock),
    .reset(Mem1D_9_reset),
    .io_r_ofs_0(Mem1D_9_io_r_ofs_0),
    .io_r_backpressure(Mem1D_9_io_r_backpressure),
    .io_w_ofs_0(Mem1D_9_io_w_ofs_0),
    .io_w_data_0(Mem1D_9_io_w_data_0),
    .io_w_en_0(Mem1D_9_io_w_en_0),
    .io_output(Mem1D_9_io_output)
  );
  Mem1D_4 Mem1D_10 ( // @[MemPrimitives.scala 64:21:@9214.4]
    .clock(Mem1D_10_clock),
    .reset(Mem1D_10_reset),
    .io_r_ofs_0(Mem1D_10_io_r_ofs_0),
    .io_r_backpressure(Mem1D_10_io_r_backpressure),
    .io_w_ofs_0(Mem1D_10_io_w_ofs_0),
    .io_w_data_0(Mem1D_10_io_w_data_0),
    .io_w_en_0(Mem1D_10_io_w_en_0),
    .io_output(Mem1D_10_io_output)
  );
  Mem1D_4 Mem1D_11 ( // @[MemPrimitives.scala 64:21:@9230.4]
    .clock(Mem1D_11_clock),
    .reset(Mem1D_11_reset),
    .io_r_ofs_0(Mem1D_11_io_r_ofs_0),
    .io_r_backpressure(Mem1D_11_io_r_backpressure),
    .io_w_ofs_0(Mem1D_11_io_w_ofs_0),
    .io_w_data_0(Mem1D_11_io_w_data_0),
    .io_w_en_0(Mem1D_11_io_w_en_0),
    .io_output(Mem1D_11_io_output)
  );
  Mem1D_4 Mem1D_12 ( // @[MemPrimitives.scala 64:21:@9246.4]
    .clock(Mem1D_12_clock),
    .reset(Mem1D_12_reset),
    .io_r_ofs_0(Mem1D_12_io_r_ofs_0),
    .io_r_backpressure(Mem1D_12_io_r_backpressure),
    .io_w_ofs_0(Mem1D_12_io_w_ofs_0),
    .io_w_data_0(Mem1D_12_io_w_data_0),
    .io_w_en_0(Mem1D_12_io_w_en_0),
    .io_output(Mem1D_12_io_output)
  );
  Mem1D_4 Mem1D_13 ( // @[MemPrimitives.scala 64:21:@9262.4]
    .clock(Mem1D_13_clock),
    .reset(Mem1D_13_reset),
    .io_r_ofs_0(Mem1D_13_io_r_ofs_0),
    .io_r_backpressure(Mem1D_13_io_r_backpressure),
    .io_w_ofs_0(Mem1D_13_io_w_ofs_0),
    .io_w_data_0(Mem1D_13_io_w_data_0),
    .io_w_en_0(Mem1D_13_io_w_en_0),
    .io_output(Mem1D_13_io_output)
  );
  Mem1D_4 Mem1D_14 ( // @[MemPrimitives.scala 64:21:@9278.4]
    .clock(Mem1D_14_clock),
    .reset(Mem1D_14_reset),
    .io_r_ofs_0(Mem1D_14_io_r_ofs_0),
    .io_r_backpressure(Mem1D_14_io_r_backpressure),
    .io_w_ofs_0(Mem1D_14_io_w_ofs_0),
    .io_w_data_0(Mem1D_14_io_w_data_0),
    .io_w_en_0(Mem1D_14_io_w_en_0),
    .io_output(Mem1D_14_io_output)
  );
  Mem1D_4 Mem1D_15 ( // @[MemPrimitives.scala 64:21:@9294.4]
    .clock(Mem1D_15_clock),
    .reset(Mem1D_15_reset),
    .io_r_ofs_0(Mem1D_15_io_r_ofs_0),
    .io_r_backpressure(Mem1D_15_io_r_backpressure),
    .io_w_ofs_0(Mem1D_15_io_w_ofs_0),
    .io_w_data_0(Mem1D_15_io_w_data_0),
    .io_w_en_0(Mem1D_15_io_w_en_0),
    .io_output(Mem1D_15_io_output)
  );
  StickySelects StickySelects ( // @[MemPrimitives.scala 121:29:@9526.4]
    .clock(StickySelects_clock),
    .reset(StickySelects_reset),
    .io_ins_0(StickySelects_io_ins_0),
    .io_ins_1(StickySelects_io_ins_1),
    .io_ins_2(StickySelects_io_ins_2),
    .io_ins_3(StickySelects_io_ins_3),
    .io_ins_4(StickySelects_io_ins_4),
    .io_ins_5(StickySelects_io_ins_5),
    .io_outs_0(StickySelects_io_outs_0),
    .io_outs_1(StickySelects_io_outs_1),
    .io_outs_2(StickySelects_io_outs_2),
    .io_outs_3(StickySelects_io_outs_3),
    .io_outs_4(StickySelects_io_outs_4),
    .io_outs_5(StickySelects_io_outs_5)
  );
  StickySelects StickySelects_1 ( // @[MemPrimitives.scala 121:29:@9588.4]
    .clock(StickySelects_1_clock),
    .reset(StickySelects_1_reset),
    .io_ins_0(StickySelects_1_io_ins_0),
    .io_ins_1(StickySelects_1_io_ins_1),
    .io_ins_2(StickySelects_1_io_ins_2),
    .io_ins_3(StickySelects_1_io_ins_3),
    .io_ins_4(StickySelects_1_io_ins_4),
    .io_ins_5(StickySelects_1_io_ins_5),
    .io_outs_0(StickySelects_1_io_outs_0),
    .io_outs_1(StickySelects_1_io_outs_1),
    .io_outs_2(StickySelects_1_io_outs_2),
    .io_outs_3(StickySelects_1_io_outs_3),
    .io_outs_4(StickySelects_1_io_outs_4),
    .io_outs_5(StickySelects_1_io_outs_5)
  );
  StickySelects StickySelects_2 ( // @[MemPrimitives.scala 121:29:@9650.4]
    .clock(StickySelects_2_clock),
    .reset(StickySelects_2_reset),
    .io_ins_0(StickySelects_2_io_ins_0),
    .io_ins_1(StickySelects_2_io_ins_1),
    .io_ins_2(StickySelects_2_io_ins_2),
    .io_ins_3(StickySelects_2_io_ins_3),
    .io_ins_4(StickySelects_2_io_ins_4),
    .io_ins_5(StickySelects_2_io_ins_5),
    .io_outs_0(StickySelects_2_io_outs_0),
    .io_outs_1(StickySelects_2_io_outs_1),
    .io_outs_2(StickySelects_2_io_outs_2),
    .io_outs_3(StickySelects_2_io_outs_3),
    .io_outs_4(StickySelects_2_io_outs_4),
    .io_outs_5(StickySelects_2_io_outs_5)
  );
  StickySelects StickySelects_3 ( // @[MemPrimitives.scala 121:29:@9712.4]
    .clock(StickySelects_3_clock),
    .reset(StickySelects_3_reset),
    .io_ins_0(StickySelects_3_io_ins_0),
    .io_ins_1(StickySelects_3_io_ins_1),
    .io_ins_2(StickySelects_3_io_ins_2),
    .io_ins_3(StickySelects_3_io_ins_3),
    .io_ins_4(StickySelects_3_io_ins_4),
    .io_ins_5(StickySelects_3_io_ins_5),
    .io_outs_0(StickySelects_3_io_outs_0),
    .io_outs_1(StickySelects_3_io_outs_1),
    .io_outs_2(StickySelects_3_io_outs_2),
    .io_outs_3(StickySelects_3_io_outs_3),
    .io_outs_4(StickySelects_3_io_outs_4),
    .io_outs_5(StickySelects_3_io_outs_5)
  );
  StickySelects StickySelects_4 ( // @[MemPrimitives.scala 121:29:@9774.4]
    .clock(StickySelects_4_clock),
    .reset(StickySelects_4_reset),
    .io_ins_0(StickySelects_4_io_ins_0),
    .io_ins_1(StickySelects_4_io_ins_1),
    .io_ins_2(StickySelects_4_io_ins_2),
    .io_ins_3(StickySelects_4_io_ins_3),
    .io_ins_4(StickySelects_4_io_ins_4),
    .io_ins_5(StickySelects_4_io_ins_5),
    .io_outs_0(StickySelects_4_io_outs_0),
    .io_outs_1(StickySelects_4_io_outs_1),
    .io_outs_2(StickySelects_4_io_outs_2),
    .io_outs_3(StickySelects_4_io_outs_3),
    .io_outs_4(StickySelects_4_io_outs_4),
    .io_outs_5(StickySelects_4_io_outs_5)
  );
  StickySelects StickySelects_5 ( // @[MemPrimitives.scala 121:29:@9836.4]
    .clock(StickySelects_5_clock),
    .reset(StickySelects_5_reset),
    .io_ins_0(StickySelects_5_io_ins_0),
    .io_ins_1(StickySelects_5_io_ins_1),
    .io_ins_2(StickySelects_5_io_ins_2),
    .io_ins_3(StickySelects_5_io_ins_3),
    .io_ins_4(StickySelects_5_io_ins_4),
    .io_ins_5(StickySelects_5_io_ins_5),
    .io_outs_0(StickySelects_5_io_outs_0),
    .io_outs_1(StickySelects_5_io_outs_1),
    .io_outs_2(StickySelects_5_io_outs_2),
    .io_outs_3(StickySelects_5_io_outs_3),
    .io_outs_4(StickySelects_5_io_outs_4),
    .io_outs_5(StickySelects_5_io_outs_5)
  );
  StickySelects StickySelects_6 ( // @[MemPrimitives.scala 121:29:@9898.4]
    .clock(StickySelects_6_clock),
    .reset(StickySelects_6_reset),
    .io_ins_0(StickySelects_6_io_ins_0),
    .io_ins_1(StickySelects_6_io_ins_1),
    .io_ins_2(StickySelects_6_io_ins_2),
    .io_ins_3(StickySelects_6_io_ins_3),
    .io_ins_4(StickySelects_6_io_ins_4),
    .io_ins_5(StickySelects_6_io_ins_5),
    .io_outs_0(StickySelects_6_io_outs_0),
    .io_outs_1(StickySelects_6_io_outs_1),
    .io_outs_2(StickySelects_6_io_outs_2),
    .io_outs_3(StickySelects_6_io_outs_3),
    .io_outs_4(StickySelects_6_io_outs_4),
    .io_outs_5(StickySelects_6_io_outs_5)
  );
  StickySelects StickySelects_7 ( // @[MemPrimitives.scala 121:29:@9960.4]
    .clock(StickySelects_7_clock),
    .reset(StickySelects_7_reset),
    .io_ins_0(StickySelects_7_io_ins_0),
    .io_ins_1(StickySelects_7_io_ins_1),
    .io_ins_2(StickySelects_7_io_ins_2),
    .io_ins_3(StickySelects_7_io_ins_3),
    .io_ins_4(StickySelects_7_io_ins_4),
    .io_ins_5(StickySelects_7_io_ins_5),
    .io_outs_0(StickySelects_7_io_outs_0),
    .io_outs_1(StickySelects_7_io_outs_1),
    .io_outs_2(StickySelects_7_io_outs_2),
    .io_outs_3(StickySelects_7_io_outs_3),
    .io_outs_4(StickySelects_7_io_outs_4),
    .io_outs_5(StickySelects_7_io_outs_5)
  );
  StickySelects StickySelects_8 ( // @[MemPrimitives.scala 121:29:@10022.4]
    .clock(StickySelects_8_clock),
    .reset(StickySelects_8_reset),
    .io_ins_0(StickySelects_8_io_ins_0),
    .io_ins_1(StickySelects_8_io_ins_1),
    .io_ins_2(StickySelects_8_io_ins_2),
    .io_ins_3(StickySelects_8_io_ins_3),
    .io_ins_4(StickySelects_8_io_ins_4),
    .io_ins_5(StickySelects_8_io_ins_5),
    .io_outs_0(StickySelects_8_io_outs_0),
    .io_outs_1(StickySelects_8_io_outs_1),
    .io_outs_2(StickySelects_8_io_outs_2),
    .io_outs_3(StickySelects_8_io_outs_3),
    .io_outs_4(StickySelects_8_io_outs_4),
    .io_outs_5(StickySelects_8_io_outs_5)
  );
  StickySelects StickySelects_9 ( // @[MemPrimitives.scala 121:29:@10084.4]
    .clock(StickySelects_9_clock),
    .reset(StickySelects_9_reset),
    .io_ins_0(StickySelects_9_io_ins_0),
    .io_ins_1(StickySelects_9_io_ins_1),
    .io_ins_2(StickySelects_9_io_ins_2),
    .io_ins_3(StickySelects_9_io_ins_3),
    .io_ins_4(StickySelects_9_io_ins_4),
    .io_ins_5(StickySelects_9_io_ins_5),
    .io_outs_0(StickySelects_9_io_outs_0),
    .io_outs_1(StickySelects_9_io_outs_1),
    .io_outs_2(StickySelects_9_io_outs_2),
    .io_outs_3(StickySelects_9_io_outs_3),
    .io_outs_4(StickySelects_9_io_outs_4),
    .io_outs_5(StickySelects_9_io_outs_5)
  );
  StickySelects StickySelects_10 ( // @[MemPrimitives.scala 121:29:@10146.4]
    .clock(StickySelects_10_clock),
    .reset(StickySelects_10_reset),
    .io_ins_0(StickySelects_10_io_ins_0),
    .io_ins_1(StickySelects_10_io_ins_1),
    .io_ins_2(StickySelects_10_io_ins_2),
    .io_ins_3(StickySelects_10_io_ins_3),
    .io_ins_4(StickySelects_10_io_ins_4),
    .io_ins_5(StickySelects_10_io_ins_5),
    .io_outs_0(StickySelects_10_io_outs_0),
    .io_outs_1(StickySelects_10_io_outs_1),
    .io_outs_2(StickySelects_10_io_outs_2),
    .io_outs_3(StickySelects_10_io_outs_3),
    .io_outs_4(StickySelects_10_io_outs_4),
    .io_outs_5(StickySelects_10_io_outs_5)
  );
  StickySelects StickySelects_11 ( // @[MemPrimitives.scala 121:29:@10208.4]
    .clock(StickySelects_11_clock),
    .reset(StickySelects_11_reset),
    .io_ins_0(StickySelects_11_io_ins_0),
    .io_ins_1(StickySelects_11_io_ins_1),
    .io_ins_2(StickySelects_11_io_ins_2),
    .io_ins_3(StickySelects_11_io_ins_3),
    .io_ins_4(StickySelects_11_io_ins_4),
    .io_ins_5(StickySelects_11_io_ins_5),
    .io_outs_0(StickySelects_11_io_outs_0),
    .io_outs_1(StickySelects_11_io_outs_1),
    .io_outs_2(StickySelects_11_io_outs_2),
    .io_outs_3(StickySelects_11_io_outs_3),
    .io_outs_4(StickySelects_11_io_outs_4),
    .io_outs_5(StickySelects_11_io_outs_5)
  );
  StickySelects StickySelects_12 ( // @[MemPrimitives.scala 121:29:@10270.4]
    .clock(StickySelects_12_clock),
    .reset(StickySelects_12_reset),
    .io_ins_0(StickySelects_12_io_ins_0),
    .io_ins_1(StickySelects_12_io_ins_1),
    .io_ins_2(StickySelects_12_io_ins_2),
    .io_ins_3(StickySelects_12_io_ins_3),
    .io_ins_4(StickySelects_12_io_ins_4),
    .io_ins_5(StickySelects_12_io_ins_5),
    .io_outs_0(StickySelects_12_io_outs_0),
    .io_outs_1(StickySelects_12_io_outs_1),
    .io_outs_2(StickySelects_12_io_outs_2),
    .io_outs_3(StickySelects_12_io_outs_3),
    .io_outs_4(StickySelects_12_io_outs_4),
    .io_outs_5(StickySelects_12_io_outs_5)
  );
  StickySelects StickySelects_13 ( // @[MemPrimitives.scala 121:29:@10332.4]
    .clock(StickySelects_13_clock),
    .reset(StickySelects_13_reset),
    .io_ins_0(StickySelects_13_io_ins_0),
    .io_ins_1(StickySelects_13_io_ins_1),
    .io_ins_2(StickySelects_13_io_ins_2),
    .io_ins_3(StickySelects_13_io_ins_3),
    .io_ins_4(StickySelects_13_io_ins_4),
    .io_ins_5(StickySelects_13_io_ins_5),
    .io_outs_0(StickySelects_13_io_outs_0),
    .io_outs_1(StickySelects_13_io_outs_1),
    .io_outs_2(StickySelects_13_io_outs_2),
    .io_outs_3(StickySelects_13_io_outs_3),
    .io_outs_4(StickySelects_13_io_outs_4),
    .io_outs_5(StickySelects_13_io_outs_5)
  );
  StickySelects StickySelects_14 ( // @[MemPrimitives.scala 121:29:@10394.4]
    .clock(StickySelects_14_clock),
    .reset(StickySelects_14_reset),
    .io_ins_0(StickySelects_14_io_ins_0),
    .io_ins_1(StickySelects_14_io_ins_1),
    .io_ins_2(StickySelects_14_io_ins_2),
    .io_ins_3(StickySelects_14_io_ins_3),
    .io_ins_4(StickySelects_14_io_ins_4),
    .io_ins_5(StickySelects_14_io_ins_5),
    .io_outs_0(StickySelects_14_io_outs_0),
    .io_outs_1(StickySelects_14_io_outs_1),
    .io_outs_2(StickySelects_14_io_outs_2),
    .io_outs_3(StickySelects_14_io_outs_3),
    .io_outs_4(StickySelects_14_io_outs_4),
    .io_outs_5(StickySelects_14_io_outs_5)
  );
  StickySelects StickySelects_15 ( // @[MemPrimitives.scala 121:29:@10456.4]
    .clock(StickySelects_15_clock),
    .reset(StickySelects_15_reset),
    .io_ins_0(StickySelects_15_io_ins_0),
    .io_ins_1(StickySelects_15_io_ins_1),
    .io_ins_2(StickySelects_15_io_ins_2),
    .io_ins_3(StickySelects_15_io_ins_3),
    .io_ins_4(StickySelects_15_io_ins_4),
    .io_ins_5(StickySelects_15_io_ins_5),
    .io_outs_0(StickySelects_15_io_outs_0),
    .io_outs_1(StickySelects_15_io_outs_1),
    .io_outs_2(StickySelects_15_io_outs_2),
    .io_outs_3(StickySelects_15_io_outs_3),
    .io_outs_4(StickySelects_15_io_outs_4),
    .io_outs_5(StickySelects_15_io_outs_5)
  );
  RetimeWrapper_52 RetimeWrapper ( // @[package.scala 93:22:@10519.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_1 ( // @[package.scala 93:22:@10527.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_2 ( // @[package.scala 93:22:@10535.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_3 ( // @[package.scala 93:22:@10543.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_4 ( // @[package.scala 93:22:@10551.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_5 ( // @[package.scala 93:22:@10559.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_6 ( // @[package.scala 93:22:@10567.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_7 ( // @[package.scala 93:22:@10575.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_8 ( // @[package.scala 93:22:@10615.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_9 ( // @[package.scala 93:22:@10623.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_10 ( // @[package.scala 93:22:@10631.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_11 ( // @[package.scala 93:22:@10639.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_12 ( // @[package.scala 93:22:@10647.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_13 ( // @[package.scala 93:22:@10655.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_14 ( // @[package.scala 93:22:@10663.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_15 ( // @[package.scala 93:22:@10671.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_16 ( // @[package.scala 93:22:@10711.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_17 ( // @[package.scala 93:22:@10719.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_18 ( // @[package.scala 93:22:@10727.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_19 ( // @[package.scala 93:22:@10735.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_20 ( // @[package.scala 93:22:@10743.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_21 ( // @[package.scala 93:22:@10751.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_22 ( // @[package.scala 93:22:@10759.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_23 ( // @[package.scala 93:22:@10767.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_24 ( // @[package.scala 93:22:@10807.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_25 ( // @[package.scala 93:22:@10815.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_26 ( // @[package.scala 93:22:@10823.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_27 ( // @[package.scala 93:22:@10831.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_28 ( // @[package.scala 93:22:@10839.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_29 ( // @[package.scala 93:22:@10847.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_30 ( // @[package.scala 93:22:@10855.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_31 ( // @[package.scala 93:22:@10863.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_32 ( // @[package.scala 93:22:@10903.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_33 ( // @[package.scala 93:22:@10911.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_34 ( // @[package.scala 93:22:@10919.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_35 ( // @[package.scala 93:22:@10927.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_36 ( // @[package.scala 93:22:@10935.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_37 ( // @[package.scala 93:22:@10943.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_38 ( // @[package.scala 93:22:@10951.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_39 ( // @[package.scala 93:22:@10959.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_40 ( // @[package.scala 93:22:@10999.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_41 ( // @[package.scala 93:22:@11007.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_42 ( // @[package.scala 93:22:@11015.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_43 ( // @[package.scala 93:22:@11023.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_44 ( // @[package.scala 93:22:@11031.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_45 ( // @[package.scala 93:22:@11039.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_46 ( // @[package.scala 93:22:@11047.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_47 ( // @[package.scala 93:22:@11055.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_48 ( // @[package.scala 93:22:@11095.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_49 ( // @[package.scala 93:22:@11103.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_50 ( // @[package.scala 93:22:@11111.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_51 ( // @[package.scala 93:22:@11119.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_52 ( // @[package.scala 93:22:@11127.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_53 ( // @[package.scala 93:22:@11135.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_54 ( // @[package.scala 93:22:@11143.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_55 ( // @[package.scala 93:22:@11151.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_56 ( // @[package.scala 93:22:@11191.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_57 ( // @[package.scala 93:22:@11199.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_58 ( // @[package.scala 93:22:@11207.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_59 ( // @[package.scala 93:22:@11215.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_60 ( // @[package.scala 93:22:@11223.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_61 ( // @[package.scala 93:22:@11231.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_62 ( // @[package.scala 93:22:@11239.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_63 ( // @[package.scala 93:22:@11247.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_64 ( // @[package.scala 93:22:@11287.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_65 ( // @[package.scala 93:22:@11295.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_66 ( // @[package.scala 93:22:@11303.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_67 ( // @[package.scala 93:22:@11311.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_68 ( // @[package.scala 93:22:@11319.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_69 ( // @[package.scala 93:22:@11327.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_70 ( // @[package.scala 93:22:@11335.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_71 ( // @[package.scala 93:22:@11343.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_72 ( // @[package.scala 93:22:@11383.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_73 ( // @[package.scala 93:22:@11391.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_74 ( // @[package.scala 93:22:@11399.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_75 ( // @[package.scala 93:22:@11407.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_76 ( // @[package.scala 93:22:@11415.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_77 ( // @[package.scala 93:22:@11423.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_78 ( // @[package.scala 93:22:@11431.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_79 ( // @[package.scala 93:22:@11439.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_80 ( // @[package.scala 93:22:@11479.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_81 ( // @[package.scala 93:22:@11487.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_82 ( // @[package.scala 93:22:@11495.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_83 ( // @[package.scala 93:22:@11503.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_84 ( // @[package.scala 93:22:@11511.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_85 ( // @[package.scala 93:22:@11519.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_86 ( // @[package.scala 93:22:@11527.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_87 ( // @[package.scala 93:22:@11535.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_88 ( // @[package.scala 93:22:@11575.4]
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_89 ( // @[package.scala 93:22:@11583.4]
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_90 ( // @[package.scala 93:22:@11591.4]
    .clock(RetimeWrapper_90_clock),
    .reset(RetimeWrapper_90_reset),
    .io_flow(RetimeWrapper_90_io_flow),
    .io_in(RetimeWrapper_90_io_in),
    .io_out(RetimeWrapper_90_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_91 ( // @[package.scala 93:22:@11599.4]
    .clock(RetimeWrapper_91_clock),
    .reset(RetimeWrapper_91_reset),
    .io_flow(RetimeWrapper_91_io_flow),
    .io_in(RetimeWrapper_91_io_in),
    .io_out(RetimeWrapper_91_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_92 ( // @[package.scala 93:22:@11607.4]
    .clock(RetimeWrapper_92_clock),
    .reset(RetimeWrapper_92_reset),
    .io_flow(RetimeWrapper_92_io_flow),
    .io_in(RetimeWrapper_92_io_in),
    .io_out(RetimeWrapper_92_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_93 ( // @[package.scala 93:22:@11615.4]
    .clock(RetimeWrapper_93_clock),
    .reset(RetimeWrapper_93_reset),
    .io_flow(RetimeWrapper_93_io_flow),
    .io_in(RetimeWrapper_93_io_in),
    .io_out(RetimeWrapper_93_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_94 ( // @[package.scala 93:22:@11623.4]
    .clock(RetimeWrapper_94_clock),
    .reset(RetimeWrapper_94_reset),
    .io_flow(RetimeWrapper_94_io_flow),
    .io_in(RetimeWrapper_94_io_in),
    .io_out(RetimeWrapper_94_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_95 ( // @[package.scala 93:22:@11631.4]
    .clock(RetimeWrapper_95_clock),
    .reset(RetimeWrapper_95_reset),
    .io_flow(RetimeWrapper_95_io_flow),
    .io_in(RetimeWrapper_95_io_in),
    .io_out(RetimeWrapper_95_io_out)
  );
  assign _T_444 = io_wPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@9310.4]
  assign _T_446 = io_wPort_0_banks_1 == 3'h0; // @[MemPrimitives.scala 82:210:@9311.4]
  assign _T_447 = _T_444 & _T_446; // @[MemPrimitives.scala 82:228:@9312.4]
  assign _T_448 = io_wPort_0_en_0 & _T_447; // @[MemPrimitives.scala 83:102:@9313.4]
  assign _T_450 = {_T_448,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9315.4]
  assign _T_455 = io_wPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@9322.4]
  assign _T_457 = io_wPort_1_banks_1 == 3'h1; // @[MemPrimitives.scala 82:210:@9323.4]
  assign _T_458 = _T_455 & _T_457; // @[MemPrimitives.scala 82:228:@9324.4]
  assign _T_459 = io_wPort_1_en_0 & _T_458; // @[MemPrimitives.scala 83:102:@9325.4]
  assign _T_461 = {_T_459,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@9327.4]
  assign _T_468 = io_wPort_0_banks_1 == 3'h2; // @[MemPrimitives.scala 82:210:@9335.4]
  assign _T_469 = _T_444 & _T_468; // @[MemPrimitives.scala 82:228:@9336.4]
  assign _T_470 = io_wPort_0_en_0 & _T_469; // @[MemPrimitives.scala 83:102:@9337.4]
  assign _T_472 = {_T_470,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9339.4]
  assign _T_479 = io_wPort_1_banks_1 == 3'h3; // @[MemPrimitives.scala 82:210:@9347.4]
  assign _T_480 = _T_455 & _T_479; // @[MemPrimitives.scala 82:228:@9348.4]
  assign _T_481 = io_wPort_1_en_0 & _T_480; // @[MemPrimitives.scala 83:102:@9349.4]
  assign _T_483 = {_T_481,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@9351.4]
  assign _T_488 = io_wPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@9358.4]
  assign _T_491 = _T_488 & _T_446; // @[MemPrimitives.scala 82:228:@9360.4]
  assign _T_492 = io_wPort_0_en_0 & _T_491; // @[MemPrimitives.scala 83:102:@9361.4]
  assign _T_494 = {_T_492,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9363.4]
  assign _T_499 = io_wPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@9370.4]
  assign _T_502 = _T_499 & _T_457; // @[MemPrimitives.scala 82:228:@9372.4]
  assign _T_503 = io_wPort_1_en_0 & _T_502; // @[MemPrimitives.scala 83:102:@9373.4]
  assign _T_505 = {_T_503,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@9375.4]
  assign _T_513 = _T_488 & _T_468; // @[MemPrimitives.scala 82:228:@9384.4]
  assign _T_514 = io_wPort_0_en_0 & _T_513; // @[MemPrimitives.scala 83:102:@9385.4]
  assign _T_516 = {_T_514,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9387.4]
  assign _T_524 = _T_499 & _T_479; // @[MemPrimitives.scala 82:228:@9396.4]
  assign _T_525 = io_wPort_1_en_0 & _T_524; // @[MemPrimitives.scala 83:102:@9397.4]
  assign _T_527 = {_T_525,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@9399.4]
  assign _T_532 = io_wPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@9406.4]
  assign _T_535 = _T_532 & _T_446; // @[MemPrimitives.scala 82:228:@9408.4]
  assign _T_536 = io_wPort_0_en_0 & _T_535; // @[MemPrimitives.scala 83:102:@9409.4]
  assign _T_538 = {_T_536,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9411.4]
  assign _T_543 = io_wPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@9418.4]
  assign _T_546 = _T_543 & _T_457; // @[MemPrimitives.scala 82:228:@9420.4]
  assign _T_547 = io_wPort_1_en_0 & _T_546; // @[MemPrimitives.scala 83:102:@9421.4]
  assign _T_549 = {_T_547,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@9423.4]
  assign _T_557 = _T_532 & _T_468; // @[MemPrimitives.scala 82:228:@9432.4]
  assign _T_558 = io_wPort_0_en_0 & _T_557; // @[MemPrimitives.scala 83:102:@9433.4]
  assign _T_560 = {_T_558,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9435.4]
  assign _T_568 = _T_543 & _T_479; // @[MemPrimitives.scala 82:228:@9444.4]
  assign _T_569 = io_wPort_1_en_0 & _T_568; // @[MemPrimitives.scala 83:102:@9445.4]
  assign _T_571 = {_T_569,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@9447.4]
  assign _T_576 = io_wPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@9454.4]
  assign _T_579 = _T_576 & _T_446; // @[MemPrimitives.scala 82:228:@9456.4]
  assign _T_580 = io_wPort_0_en_0 & _T_579; // @[MemPrimitives.scala 83:102:@9457.4]
  assign _T_582 = {_T_580,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9459.4]
  assign _T_587 = io_wPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@9466.4]
  assign _T_590 = _T_587 & _T_457; // @[MemPrimitives.scala 82:228:@9468.4]
  assign _T_591 = io_wPort_1_en_0 & _T_590; // @[MemPrimitives.scala 83:102:@9469.4]
  assign _T_593 = {_T_591,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@9471.4]
  assign _T_601 = _T_576 & _T_468; // @[MemPrimitives.scala 82:228:@9480.4]
  assign _T_602 = io_wPort_0_en_0 & _T_601; // @[MemPrimitives.scala 83:102:@9481.4]
  assign _T_604 = {_T_602,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9483.4]
  assign _T_612 = _T_587 & _T_479; // @[MemPrimitives.scala 82:228:@9492.4]
  assign _T_613 = io_wPort_1_en_0 & _T_612; // @[MemPrimitives.scala 83:102:@9493.4]
  assign _T_615 = {_T_613,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@9495.4]
  assign _T_620 = io_rPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9502.4]
  assign _T_622 = io_rPort_1_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@9503.4]
  assign _T_623 = _T_620 & _T_622; // @[MemPrimitives.scala 110:228:@9504.4]
  assign _T_626 = io_rPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9506.4]
  assign _T_628 = io_rPort_2_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@9507.4]
  assign _T_629 = _T_626 & _T_628; // @[MemPrimitives.scala 110:228:@9508.4]
  assign _T_632 = io_rPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9510.4]
  assign _T_634 = io_rPort_3_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@9511.4]
  assign _T_635 = _T_632 & _T_634; // @[MemPrimitives.scala 110:228:@9512.4]
  assign _T_638 = io_rPort_6_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9514.4]
  assign _T_640 = io_rPort_6_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@9515.4]
  assign _T_641 = _T_638 & _T_640; // @[MemPrimitives.scala 110:228:@9516.4]
  assign _T_644 = io_rPort_8_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9518.4]
  assign _T_646 = io_rPort_8_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@9519.4]
  assign _T_647 = _T_644 & _T_646; // @[MemPrimitives.scala 110:228:@9520.4]
  assign _T_650 = io_rPort_11_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9522.4]
  assign _T_652 = io_rPort_11_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@9523.4]
  assign _T_653 = _T_650 & _T_652; // @[MemPrimitives.scala 110:228:@9524.4]
  assign _T_655 = StickySelects_io_outs_0; // @[MemPrimitives.scala 123:41:@9535.4]
  assign _T_656 = StickySelects_io_outs_1; // @[MemPrimitives.scala 123:41:@9536.4]
  assign _T_657 = StickySelects_io_outs_2; // @[MemPrimitives.scala 123:41:@9537.4]
  assign _T_658 = StickySelects_io_outs_3; // @[MemPrimitives.scala 123:41:@9538.4]
  assign _T_659 = StickySelects_io_outs_4; // @[MemPrimitives.scala 123:41:@9539.4]
  assign _T_660 = StickySelects_io_outs_5; // @[MemPrimitives.scala 123:41:@9540.4]
  assign _T_662 = {_T_655,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@9542.4]
  assign _T_664 = {_T_656,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@9544.4]
  assign _T_666 = {_T_657,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@9546.4]
  assign _T_668 = {_T_658,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@9548.4]
  assign _T_670 = {_T_659,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@9550.4]
  assign _T_672 = {_T_660,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@9552.4]
  assign _T_673 = _T_659 ? _T_670 : _T_672; // @[Mux.scala 31:69:@9553.4]
  assign _T_674 = _T_658 ? _T_668 : _T_673; // @[Mux.scala 31:69:@9554.4]
  assign _T_675 = _T_657 ? _T_666 : _T_674; // @[Mux.scala 31:69:@9555.4]
  assign _T_676 = _T_656 ? _T_664 : _T_675; // @[Mux.scala 31:69:@9556.4]
  assign _T_677 = _T_655 ? _T_662 : _T_676; // @[Mux.scala 31:69:@9557.4]
  assign _T_682 = io_rPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9564.4]
  assign _T_684 = io_rPort_0_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@9565.4]
  assign _T_685 = _T_682 & _T_684; // @[MemPrimitives.scala 110:228:@9566.4]
  assign _T_688 = io_rPort_4_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9568.4]
  assign _T_690 = io_rPort_4_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@9569.4]
  assign _T_691 = _T_688 & _T_690; // @[MemPrimitives.scala 110:228:@9570.4]
  assign _T_694 = io_rPort_5_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9572.4]
  assign _T_696 = io_rPort_5_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@9573.4]
  assign _T_697 = _T_694 & _T_696; // @[MemPrimitives.scala 110:228:@9574.4]
  assign _T_700 = io_rPort_7_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9576.4]
  assign _T_702 = io_rPort_7_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@9577.4]
  assign _T_703 = _T_700 & _T_702; // @[MemPrimitives.scala 110:228:@9578.4]
  assign _T_706 = io_rPort_9_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9580.4]
  assign _T_708 = io_rPort_9_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@9581.4]
  assign _T_709 = _T_706 & _T_708; // @[MemPrimitives.scala 110:228:@9582.4]
  assign _T_712 = io_rPort_10_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9584.4]
  assign _T_714 = io_rPort_10_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@9585.4]
  assign _T_715 = _T_712 & _T_714; // @[MemPrimitives.scala 110:228:@9586.4]
  assign _T_717 = StickySelects_1_io_outs_0; // @[MemPrimitives.scala 123:41:@9597.4]
  assign _T_718 = StickySelects_1_io_outs_1; // @[MemPrimitives.scala 123:41:@9598.4]
  assign _T_719 = StickySelects_1_io_outs_2; // @[MemPrimitives.scala 123:41:@9599.4]
  assign _T_720 = StickySelects_1_io_outs_3; // @[MemPrimitives.scala 123:41:@9600.4]
  assign _T_721 = StickySelects_1_io_outs_4; // @[MemPrimitives.scala 123:41:@9601.4]
  assign _T_722 = StickySelects_1_io_outs_5; // @[MemPrimitives.scala 123:41:@9602.4]
  assign _T_724 = {_T_717,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@9604.4]
  assign _T_726 = {_T_718,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@9606.4]
  assign _T_728 = {_T_719,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@9608.4]
  assign _T_730 = {_T_720,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@9610.4]
  assign _T_732 = {_T_721,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@9612.4]
  assign _T_734 = {_T_722,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@9614.4]
  assign _T_735 = _T_721 ? _T_732 : _T_734; // @[Mux.scala 31:69:@9615.4]
  assign _T_736 = _T_720 ? _T_730 : _T_735; // @[Mux.scala 31:69:@9616.4]
  assign _T_737 = _T_719 ? _T_728 : _T_736; // @[Mux.scala 31:69:@9617.4]
  assign _T_738 = _T_718 ? _T_726 : _T_737; // @[Mux.scala 31:69:@9618.4]
  assign _T_739 = _T_717 ? _T_724 : _T_738; // @[Mux.scala 31:69:@9619.4]
  assign _T_746 = io_rPort_1_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@9627.4]
  assign _T_747 = _T_620 & _T_746; // @[MemPrimitives.scala 110:228:@9628.4]
  assign _T_752 = io_rPort_2_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@9631.4]
  assign _T_753 = _T_626 & _T_752; // @[MemPrimitives.scala 110:228:@9632.4]
  assign _T_758 = io_rPort_3_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@9635.4]
  assign _T_759 = _T_632 & _T_758; // @[MemPrimitives.scala 110:228:@9636.4]
  assign _T_764 = io_rPort_6_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@9639.4]
  assign _T_765 = _T_638 & _T_764; // @[MemPrimitives.scala 110:228:@9640.4]
  assign _T_770 = io_rPort_8_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@9643.4]
  assign _T_771 = _T_644 & _T_770; // @[MemPrimitives.scala 110:228:@9644.4]
  assign _T_776 = io_rPort_11_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@9647.4]
  assign _T_777 = _T_650 & _T_776; // @[MemPrimitives.scala 110:228:@9648.4]
  assign _T_779 = StickySelects_2_io_outs_0; // @[MemPrimitives.scala 123:41:@9659.4]
  assign _T_780 = StickySelects_2_io_outs_1; // @[MemPrimitives.scala 123:41:@9660.4]
  assign _T_781 = StickySelects_2_io_outs_2; // @[MemPrimitives.scala 123:41:@9661.4]
  assign _T_782 = StickySelects_2_io_outs_3; // @[MemPrimitives.scala 123:41:@9662.4]
  assign _T_783 = StickySelects_2_io_outs_4; // @[MemPrimitives.scala 123:41:@9663.4]
  assign _T_784 = StickySelects_2_io_outs_5; // @[MemPrimitives.scala 123:41:@9664.4]
  assign _T_786 = {_T_779,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@9666.4]
  assign _T_788 = {_T_780,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@9668.4]
  assign _T_790 = {_T_781,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@9670.4]
  assign _T_792 = {_T_782,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@9672.4]
  assign _T_794 = {_T_783,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@9674.4]
  assign _T_796 = {_T_784,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@9676.4]
  assign _T_797 = _T_783 ? _T_794 : _T_796; // @[Mux.scala 31:69:@9677.4]
  assign _T_798 = _T_782 ? _T_792 : _T_797; // @[Mux.scala 31:69:@9678.4]
  assign _T_799 = _T_781 ? _T_790 : _T_798; // @[Mux.scala 31:69:@9679.4]
  assign _T_800 = _T_780 ? _T_788 : _T_799; // @[Mux.scala 31:69:@9680.4]
  assign _T_801 = _T_779 ? _T_786 : _T_800; // @[Mux.scala 31:69:@9681.4]
  assign _T_808 = io_rPort_0_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@9689.4]
  assign _T_809 = _T_682 & _T_808; // @[MemPrimitives.scala 110:228:@9690.4]
  assign _T_814 = io_rPort_4_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@9693.4]
  assign _T_815 = _T_688 & _T_814; // @[MemPrimitives.scala 110:228:@9694.4]
  assign _T_820 = io_rPort_5_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@9697.4]
  assign _T_821 = _T_694 & _T_820; // @[MemPrimitives.scala 110:228:@9698.4]
  assign _T_826 = io_rPort_7_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@9701.4]
  assign _T_827 = _T_700 & _T_826; // @[MemPrimitives.scala 110:228:@9702.4]
  assign _T_832 = io_rPort_9_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@9705.4]
  assign _T_833 = _T_706 & _T_832; // @[MemPrimitives.scala 110:228:@9706.4]
  assign _T_838 = io_rPort_10_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@9709.4]
  assign _T_839 = _T_712 & _T_838; // @[MemPrimitives.scala 110:228:@9710.4]
  assign _T_841 = StickySelects_3_io_outs_0; // @[MemPrimitives.scala 123:41:@9721.4]
  assign _T_842 = StickySelects_3_io_outs_1; // @[MemPrimitives.scala 123:41:@9722.4]
  assign _T_843 = StickySelects_3_io_outs_2; // @[MemPrimitives.scala 123:41:@9723.4]
  assign _T_844 = StickySelects_3_io_outs_3; // @[MemPrimitives.scala 123:41:@9724.4]
  assign _T_845 = StickySelects_3_io_outs_4; // @[MemPrimitives.scala 123:41:@9725.4]
  assign _T_846 = StickySelects_3_io_outs_5; // @[MemPrimitives.scala 123:41:@9726.4]
  assign _T_848 = {_T_841,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@9728.4]
  assign _T_850 = {_T_842,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@9730.4]
  assign _T_852 = {_T_843,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@9732.4]
  assign _T_854 = {_T_844,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@9734.4]
  assign _T_856 = {_T_845,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@9736.4]
  assign _T_858 = {_T_846,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@9738.4]
  assign _T_859 = _T_845 ? _T_856 : _T_858; // @[Mux.scala 31:69:@9739.4]
  assign _T_860 = _T_844 ? _T_854 : _T_859; // @[Mux.scala 31:69:@9740.4]
  assign _T_861 = _T_843 ? _T_852 : _T_860; // @[Mux.scala 31:69:@9741.4]
  assign _T_862 = _T_842 ? _T_850 : _T_861; // @[Mux.scala 31:69:@9742.4]
  assign _T_863 = _T_841 ? _T_848 : _T_862; // @[Mux.scala 31:69:@9743.4]
  assign _T_868 = io_rPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9750.4]
  assign _T_871 = _T_868 & _T_622; // @[MemPrimitives.scala 110:228:@9752.4]
  assign _T_874 = io_rPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9754.4]
  assign _T_877 = _T_874 & _T_628; // @[MemPrimitives.scala 110:228:@9756.4]
  assign _T_880 = io_rPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9758.4]
  assign _T_883 = _T_880 & _T_634; // @[MemPrimitives.scala 110:228:@9760.4]
  assign _T_886 = io_rPort_6_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9762.4]
  assign _T_889 = _T_886 & _T_640; // @[MemPrimitives.scala 110:228:@9764.4]
  assign _T_892 = io_rPort_8_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9766.4]
  assign _T_895 = _T_892 & _T_646; // @[MemPrimitives.scala 110:228:@9768.4]
  assign _T_898 = io_rPort_11_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9770.4]
  assign _T_901 = _T_898 & _T_652; // @[MemPrimitives.scala 110:228:@9772.4]
  assign _T_903 = StickySelects_4_io_outs_0; // @[MemPrimitives.scala 123:41:@9783.4]
  assign _T_904 = StickySelects_4_io_outs_1; // @[MemPrimitives.scala 123:41:@9784.4]
  assign _T_905 = StickySelects_4_io_outs_2; // @[MemPrimitives.scala 123:41:@9785.4]
  assign _T_906 = StickySelects_4_io_outs_3; // @[MemPrimitives.scala 123:41:@9786.4]
  assign _T_907 = StickySelects_4_io_outs_4; // @[MemPrimitives.scala 123:41:@9787.4]
  assign _T_908 = StickySelects_4_io_outs_5; // @[MemPrimitives.scala 123:41:@9788.4]
  assign _T_910 = {_T_903,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@9790.4]
  assign _T_912 = {_T_904,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@9792.4]
  assign _T_914 = {_T_905,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@9794.4]
  assign _T_916 = {_T_906,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@9796.4]
  assign _T_918 = {_T_907,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@9798.4]
  assign _T_920 = {_T_908,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@9800.4]
  assign _T_921 = _T_907 ? _T_918 : _T_920; // @[Mux.scala 31:69:@9801.4]
  assign _T_922 = _T_906 ? _T_916 : _T_921; // @[Mux.scala 31:69:@9802.4]
  assign _T_923 = _T_905 ? _T_914 : _T_922; // @[Mux.scala 31:69:@9803.4]
  assign _T_924 = _T_904 ? _T_912 : _T_923; // @[Mux.scala 31:69:@9804.4]
  assign _T_925 = _T_903 ? _T_910 : _T_924; // @[Mux.scala 31:69:@9805.4]
  assign _T_930 = io_rPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9812.4]
  assign _T_933 = _T_930 & _T_684; // @[MemPrimitives.scala 110:228:@9814.4]
  assign _T_936 = io_rPort_4_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9816.4]
  assign _T_939 = _T_936 & _T_690; // @[MemPrimitives.scala 110:228:@9818.4]
  assign _T_942 = io_rPort_5_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9820.4]
  assign _T_945 = _T_942 & _T_696; // @[MemPrimitives.scala 110:228:@9822.4]
  assign _T_948 = io_rPort_7_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9824.4]
  assign _T_951 = _T_948 & _T_702; // @[MemPrimitives.scala 110:228:@9826.4]
  assign _T_954 = io_rPort_9_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9828.4]
  assign _T_957 = _T_954 & _T_708; // @[MemPrimitives.scala 110:228:@9830.4]
  assign _T_960 = io_rPort_10_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9832.4]
  assign _T_963 = _T_960 & _T_714; // @[MemPrimitives.scala 110:228:@9834.4]
  assign _T_965 = StickySelects_5_io_outs_0; // @[MemPrimitives.scala 123:41:@9845.4]
  assign _T_966 = StickySelects_5_io_outs_1; // @[MemPrimitives.scala 123:41:@9846.4]
  assign _T_967 = StickySelects_5_io_outs_2; // @[MemPrimitives.scala 123:41:@9847.4]
  assign _T_968 = StickySelects_5_io_outs_3; // @[MemPrimitives.scala 123:41:@9848.4]
  assign _T_969 = StickySelects_5_io_outs_4; // @[MemPrimitives.scala 123:41:@9849.4]
  assign _T_970 = StickySelects_5_io_outs_5; // @[MemPrimitives.scala 123:41:@9850.4]
  assign _T_972 = {_T_965,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@9852.4]
  assign _T_974 = {_T_966,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@9854.4]
  assign _T_976 = {_T_967,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@9856.4]
  assign _T_978 = {_T_968,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@9858.4]
  assign _T_980 = {_T_969,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@9860.4]
  assign _T_982 = {_T_970,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@9862.4]
  assign _T_983 = _T_969 ? _T_980 : _T_982; // @[Mux.scala 31:69:@9863.4]
  assign _T_984 = _T_968 ? _T_978 : _T_983; // @[Mux.scala 31:69:@9864.4]
  assign _T_985 = _T_967 ? _T_976 : _T_984; // @[Mux.scala 31:69:@9865.4]
  assign _T_986 = _T_966 ? _T_974 : _T_985; // @[Mux.scala 31:69:@9866.4]
  assign _T_987 = _T_965 ? _T_972 : _T_986; // @[Mux.scala 31:69:@9867.4]
  assign _T_995 = _T_868 & _T_746; // @[MemPrimitives.scala 110:228:@9876.4]
  assign _T_1001 = _T_874 & _T_752; // @[MemPrimitives.scala 110:228:@9880.4]
  assign _T_1007 = _T_880 & _T_758; // @[MemPrimitives.scala 110:228:@9884.4]
  assign _T_1013 = _T_886 & _T_764; // @[MemPrimitives.scala 110:228:@9888.4]
  assign _T_1019 = _T_892 & _T_770; // @[MemPrimitives.scala 110:228:@9892.4]
  assign _T_1025 = _T_898 & _T_776; // @[MemPrimitives.scala 110:228:@9896.4]
  assign _T_1027 = StickySelects_6_io_outs_0; // @[MemPrimitives.scala 123:41:@9907.4]
  assign _T_1028 = StickySelects_6_io_outs_1; // @[MemPrimitives.scala 123:41:@9908.4]
  assign _T_1029 = StickySelects_6_io_outs_2; // @[MemPrimitives.scala 123:41:@9909.4]
  assign _T_1030 = StickySelects_6_io_outs_3; // @[MemPrimitives.scala 123:41:@9910.4]
  assign _T_1031 = StickySelects_6_io_outs_4; // @[MemPrimitives.scala 123:41:@9911.4]
  assign _T_1032 = StickySelects_6_io_outs_5; // @[MemPrimitives.scala 123:41:@9912.4]
  assign _T_1034 = {_T_1027,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@9914.4]
  assign _T_1036 = {_T_1028,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@9916.4]
  assign _T_1038 = {_T_1029,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@9918.4]
  assign _T_1040 = {_T_1030,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@9920.4]
  assign _T_1042 = {_T_1031,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@9922.4]
  assign _T_1044 = {_T_1032,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@9924.4]
  assign _T_1045 = _T_1031 ? _T_1042 : _T_1044; // @[Mux.scala 31:69:@9925.4]
  assign _T_1046 = _T_1030 ? _T_1040 : _T_1045; // @[Mux.scala 31:69:@9926.4]
  assign _T_1047 = _T_1029 ? _T_1038 : _T_1046; // @[Mux.scala 31:69:@9927.4]
  assign _T_1048 = _T_1028 ? _T_1036 : _T_1047; // @[Mux.scala 31:69:@9928.4]
  assign _T_1049 = _T_1027 ? _T_1034 : _T_1048; // @[Mux.scala 31:69:@9929.4]
  assign _T_1057 = _T_930 & _T_808; // @[MemPrimitives.scala 110:228:@9938.4]
  assign _T_1063 = _T_936 & _T_814; // @[MemPrimitives.scala 110:228:@9942.4]
  assign _T_1069 = _T_942 & _T_820; // @[MemPrimitives.scala 110:228:@9946.4]
  assign _T_1075 = _T_948 & _T_826; // @[MemPrimitives.scala 110:228:@9950.4]
  assign _T_1081 = _T_954 & _T_832; // @[MemPrimitives.scala 110:228:@9954.4]
  assign _T_1087 = _T_960 & _T_838; // @[MemPrimitives.scala 110:228:@9958.4]
  assign _T_1089 = StickySelects_7_io_outs_0; // @[MemPrimitives.scala 123:41:@9969.4]
  assign _T_1090 = StickySelects_7_io_outs_1; // @[MemPrimitives.scala 123:41:@9970.4]
  assign _T_1091 = StickySelects_7_io_outs_2; // @[MemPrimitives.scala 123:41:@9971.4]
  assign _T_1092 = StickySelects_7_io_outs_3; // @[MemPrimitives.scala 123:41:@9972.4]
  assign _T_1093 = StickySelects_7_io_outs_4; // @[MemPrimitives.scala 123:41:@9973.4]
  assign _T_1094 = StickySelects_7_io_outs_5; // @[MemPrimitives.scala 123:41:@9974.4]
  assign _T_1096 = {_T_1089,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@9976.4]
  assign _T_1098 = {_T_1090,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@9978.4]
  assign _T_1100 = {_T_1091,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@9980.4]
  assign _T_1102 = {_T_1092,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@9982.4]
  assign _T_1104 = {_T_1093,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@9984.4]
  assign _T_1106 = {_T_1094,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@9986.4]
  assign _T_1107 = _T_1093 ? _T_1104 : _T_1106; // @[Mux.scala 31:69:@9987.4]
  assign _T_1108 = _T_1092 ? _T_1102 : _T_1107; // @[Mux.scala 31:69:@9988.4]
  assign _T_1109 = _T_1091 ? _T_1100 : _T_1108; // @[Mux.scala 31:69:@9989.4]
  assign _T_1110 = _T_1090 ? _T_1098 : _T_1109; // @[Mux.scala 31:69:@9990.4]
  assign _T_1111 = _T_1089 ? _T_1096 : _T_1110; // @[Mux.scala 31:69:@9991.4]
  assign _T_1116 = io_rPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@9998.4]
  assign _T_1119 = _T_1116 & _T_622; // @[MemPrimitives.scala 110:228:@10000.4]
  assign _T_1122 = io_rPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10002.4]
  assign _T_1125 = _T_1122 & _T_628; // @[MemPrimitives.scala 110:228:@10004.4]
  assign _T_1128 = io_rPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10006.4]
  assign _T_1131 = _T_1128 & _T_634; // @[MemPrimitives.scala 110:228:@10008.4]
  assign _T_1134 = io_rPort_6_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10010.4]
  assign _T_1137 = _T_1134 & _T_640; // @[MemPrimitives.scala 110:228:@10012.4]
  assign _T_1140 = io_rPort_8_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10014.4]
  assign _T_1143 = _T_1140 & _T_646; // @[MemPrimitives.scala 110:228:@10016.4]
  assign _T_1146 = io_rPort_11_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10018.4]
  assign _T_1149 = _T_1146 & _T_652; // @[MemPrimitives.scala 110:228:@10020.4]
  assign _T_1151 = StickySelects_8_io_outs_0; // @[MemPrimitives.scala 123:41:@10031.4]
  assign _T_1152 = StickySelects_8_io_outs_1; // @[MemPrimitives.scala 123:41:@10032.4]
  assign _T_1153 = StickySelects_8_io_outs_2; // @[MemPrimitives.scala 123:41:@10033.4]
  assign _T_1154 = StickySelects_8_io_outs_3; // @[MemPrimitives.scala 123:41:@10034.4]
  assign _T_1155 = StickySelects_8_io_outs_4; // @[MemPrimitives.scala 123:41:@10035.4]
  assign _T_1156 = StickySelects_8_io_outs_5; // @[MemPrimitives.scala 123:41:@10036.4]
  assign _T_1158 = {_T_1151,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@10038.4]
  assign _T_1160 = {_T_1152,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@10040.4]
  assign _T_1162 = {_T_1153,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@10042.4]
  assign _T_1164 = {_T_1154,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@10044.4]
  assign _T_1166 = {_T_1155,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@10046.4]
  assign _T_1168 = {_T_1156,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@10048.4]
  assign _T_1169 = _T_1155 ? _T_1166 : _T_1168; // @[Mux.scala 31:69:@10049.4]
  assign _T_1170 = _T_1154 ? _T_1164 : _T_1169; // @[Mux.scala 31:69:@10050.4]
  assign _T_1171 = _T_1153 ? _T_1162 : _T_1170; // @[Mux.scala 31:69:@10051.4]
  assign _T_1172 = _T_1152 ? _T_1160 : _T_1171; // @[Mux.scala 31:69:@10052.4]
  assign _T_1173 = _T_1151 ? _T_1158 : _T_1172; // @[Mux.scala 31:69:@10053.4]
  assign _T_1178 = io_rPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10060.4]
  assign _T_1181 = _T_1178 & _T_684; // @[MemPrimitives.scala 110:228:@10062.4]
  assign _T_1184 = io_rPort_4_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10064.4]
  assign _T_1187 = _T_1184 & _T_690; // @[MemPrimitives.scala 110:228:@10066.4]
  assign _T_1190 = io_rPort_5_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10068.4]
  assign _T_1193 = _T_1190 & _T_696; // @[MemPrimitives.scala 110:228:@10070.4]
  assign _T_1196 = io_rPort_7_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10072.4]
  assign _T_1199 = _T_1196 & _T_702; // @[MemPrimitives.scala 110:228:@10074.4]
  assign _T_1202 = io_rPort_9_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10076.4]
  assign _T_1205 = _T_1202 & _T_708; // @[MemPrimitives.scala 110:228:@10078.4]
  assign _T_1208 = io_rPort_10_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10080.4]
  assign _T_1211 = _T_1208 & _T_714; // @[MemPrimitives.scala 110:228:@10082.4]
  assign _T_1213 = StickySelects_9_io_outs_0; // @[MemPrimitives.scala 123:41:@10093.4]
  assign _T_1214 = StickySelects_9_io_outs_1; // @[MemPrimitives.scala 123:41:@10094.4]
  assign _T_1215 = StickySelects_9_io_outs_2; // @[MemPrimitives.scala 123:41:@10095.4]
  assign _T_1216 = StickySelects_9_io_outs_3; // @[MemPrimitives.scala 123:41:@10096.4]
  assign _T_1217 = StickySelects_9_io_outs_4; // @[MemPrimitives.scala 123:41:@10097.4]
  assign _T_1218 = StickySelects_9_io_outs_5; // @[MemPrimitives.scala 123:41:@10098.4]
  assign _T_1220 = {_T_1213,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@10100.4]
  assign _T_1222 = {_T_1214,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@10102.4]
  assign _T_1224 = {_T_1215,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@10104.4]
  assign _T_1226 = {_T_1216,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@10106.4]
  assign _T_1228 = {_T_1217,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@10108.4]
  assign _T_1230 = {_T_1218,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@10110.4]
  assign _T_1231 = _T_1217 ? _T_1228 : _T_1230; // @[Mux.scala 31:69:@10111.4]
  assign _T_1232 = _T_1216 ? _T_1226 : _T_1231; // @[Mux.scala 31:69:@10112.4]
  assign _T_1233 = _T_1215 ? _T_1224 : _T_1232; // @[Mux.scala 31:69:@10113.4]
  assign _T_1234 = _T_1214 ? _T_1222 : _T_1233; // @[Mux.scala 31:69:@10114.4]
  assign _T_1235 = _T_1213 ? _T_1220 : _T_1234; // @[Mux.scala 31:69:@10115.4]
  assign _T_1243 = _T_1116 & _T_746; // @[MemPrimitives.scala 110:228:@10124.4]
  assign _T_1249 = _T_1122 & _T_752; // @[MemPrimitives.scala 110:228:@10128.4]
  assign _T_1255 = _T_1128 & _T_758; // @[MemPrimitives.scala 110:228:@10132.4]
  assign _T_1261 = _T_1134 & _T_764; // @[MemPrimitives.scala 110:228:@10136.4]
  assign _T_1267 = _T_1140 & _T_770; // @[MemPrimitives.scala 110:228:@10140.4]
  assign _T_1273 = _T_1146 & _T_776; // @[MemPrimitives.scala 110:228:@10144.4]
  assign _T_1275 = StickySelects_10_io_outs_0; // @[MemPrimitives.scala 123:41:@10155.4]
  assign _T_1276 = StickySelects_10_io_outs_1; // @[MemPrimitives.scala 123:41:@10156.4]
  assign _T_1277 = StickySelects_10_io_outs_2; // @[MemPrimitives.scala 123:41:@10157.4]
  assign _T_1278 = StickySelects_10_io_outs_3; // @[MemPrimitives.scala 123:41:@10158.4]
  assign _T_1279 = StickySelects_10_io_outs_4; // @[MemPrimitives.scala 123:41:@10159.4]
  assign _T_1280 = StickySelects_10_io_outs_5; // @[MemPrimitives.scala 123:41:@10160.4]
  assign _T_1282 = {_T_1275,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@10162.4]
  assign _T_1284 = {_T_1276,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@10164.4]
  assign _T_1286 = {_T_1277,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@10166.4]
  assign _T_1288 = {_T_1278,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@10168.4]
  assign _T_1290 = {_T_1279,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@10170.4]
  assign _T_1292 = {_T_1280,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@10172.4]
  assign _T_1293 = _T_1279 ? _T_1290 : _T_1292; // @[Mux.scala 31:69:@10173.4]
  assign _T_1294 = _T_1278 ? _T_1288 : _T_1293; // @[Mux.scala 31:69:@10174.4]
  assign _T_1295 = _T_1277 ? _T_1286 : _T_1294; // @[Mux.scala 31:69:@10175.4]
  assign _T_1296 = _T_1276 ? _T_1284 : _T_1295; // @[Mux.scala 31:69:@10176.4]
  assign _T_1297 = _T_1275 ? _T_1282 : _T_1296; // @[Mux.scala 31:69:@10177.4]
  assign _T_1305 = _T_1178 & _T_808; // @[MemPrimitives.scala 110:228:@10186.4]
  assign _T_1311 = _T_1184 & _T_814; // @[MemPrimitives.scala 110:228:@10190.4]
  assign _T_1317 = _T_1190 & _T_820; // @[MemPrimitives.scala 110:228:@10194.4]
  assign _T_1323 = _T_1196 & _T_826; // @[MemPrimitives.scala 110:228:@10198.4]
  assign _T_1329 = _T_1202 & _T_832; // @[MemPrimitives.scala 110:228:@10202.4]
  assign _T_1335 = _T_1208 & _T_838; // @[MemPrimitives.scala 110:228:@10206.4]
  assign _T_1337 = StickySelects_11_io_outs_0; // @[MemPrimitives.scala 123:41:@10217.4]
  assign _T_1338 = StickySelects_11_io_outs_1; // @[MemPrimitives.scala 123:41:@10218.4]
  assign _T_1339 = StickySelects_11_io_outs_2; // @[MemPrimitives.scala 123:41:@10219.4]
  assign _T_1340 = StickySelects_11_io_outs_3; // @[MemPrimitives.scala 123:41:@10220.4]
  assign _T_1341 = StickySelects_11_io_outs_4; // @[MemPrimitives.scala 123:41:@10221.4]
  assign _T_1342 = StickySelects_11_io_outs_5; // @[MemPrimitives.scala 123:41:@10222.4]
  assign _T_1344 = {_T_1337,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@10224.4]
  assign _T_1346 = {_T_1338,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@10226.4]
  assign _T_1348 = {_T_1339,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@10228.4]
  assign _T_1350 = {_T_1340,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@10230.4]
  assign _T_1352 = {_T_1341,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@10232.4]
  assign _T_1354 = {_T_1342,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@10234.4]
  assign _T_1355 = _T_1341 ? _T_1352 : _T_1354; // @[Mux.scala 31:69:@10235.4]
  assign _T_1356 = _T_1340 ? _T_1350 : _T_1355; // @[Mux.scala 31:69:@10236.4]
  assign _T_1357 = _T_1339 ? _T_1348 : _T_1356; // @[Mux.scala 31:69:@10237.4]
  assign _T_1358 = _T_1338 ? _T_1346 : _T_1357; // @[Mux.scala 31:69:@10238.4]
  assign _T_1359 = _T_1337 ? _T_1344 : _T_1358; // @[Mux.scala 31:69:@10239.4]
  assign _T_1364 = io_rPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10246.4]
  assign _T_1367 = _T_1364 & _T_622; // @[MemPrimitives.scala 110:228:@10248.4]
  assign _T_1370 = io_rPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10250.4]
  assign _T_1373 = _T_1370 & _T_628; // @[MemPrimitives.scala 110:228:@10252.4]
  assign _T_1376 = io_rPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10254.4]
  assign _T_1379 = _T_1376 & _T_634; // @[MemPrimitives.scala 110:228:@10256.4]
  assign _T_1382 = io_rPort_6_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10258.4]
  assign _T_1385 = _T_1382 & _T_640; // @[MemPrimitives.scala 110:228:@10260.4]
  assign _T_1388 = io_rPort_8_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10262.4]
  assign _T_1391 = _T_1388 & _T_646; // @[MemPrimitives.scala 110:228:@10264.4]
  assign _T_1394 = io_rPort_11_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10266.4]
  assign _T_1397 = _T_1394 & _T_652; // @[MemPrimitives.scala 110:228:@10268.4]
  assign _T_1399 = StickySelects_12_io_outs_0; // @[MemPrimitives.scala 123:41:@10279.4]
  assign _T_1400 = StickySelects_12_io_outs_1; // @[MemPrimitives.scala 123:41:@10280.4]
  assign _T_1401 = StickySelects_12_io_outs_2; // @[MemPrimitives.scala 123:41:@10281.4]
  assign _T_1402 = StickySelects_12_io_outs_3; // @[MemPrimitives.scala 123:41:@10282.4]
  assign _T_1403 = StickySelects_12_io_outs_4; // @[MemPrimitives.scala 123:41:@10283.4]
  assign _T_1404 = StickySelects_12_io_outs_5; // @[MemPrimitives.scala 123:41:@10284.4]
  assign _T_1406 = {_T_1399,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@10286.4]
  assign _T_1408 = {_T_1400,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@10288.4]
  assign _T_1410 = {_T_1401,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@10290.4]
  assign _T_1412 = {_T_1402,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@10292.4]
  assign _T_1414 = {_T_1403,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@10294.4]
  assign _T_1416 = {_T_1404,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@10296.4]
  assign _T_1417 = _T_1403 ? _T_1414 : _T_1416; // @[Mux.scala 31:69:@10297.4]
  assign _T_1418 = _T_1402 ? _T_1412 : _T_1417; // @[Mux.scala 31:69:@10298.4]
  assign _T_1419 = _T_1401 ? _T_1410 : _T_1418; // @[Mux.scala 31:69:@10299.4]
  assign _T_1420 = _T_1400 ? _T_1408 : _T_1419; // @[Mux.scala 31:69:@10300.4]
  assign _T_1421 = _T_1399 ? _T_1406 : _T_1420; // @[Mux.scala 31:69:@10301.4]
  assign _T_1426 = io_rPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10308.4]
  assign _T_1429 = _T_1426 & _T_684; // @[MemPrimitives.scala 110:228:@10310.4]
  assign _T_1432 = io_rPort_4_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10312.4]
  assign _T_1435 = _T_1432 & _T_690; // @[MemPrimitives.scala 110:228:@10314.4]
  assign _T_1438 = io_rPort_5_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10316.4]
  assign _T_1441 = _T_1438 & _T_696; // @[MemPrimitives.scala 110:228:@10318.4]
  assign _T_1444 = io_rPort_7_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10320.4]
  assign _T_1447 = _T_1444 & _T_702; // @[MemPrimitives.scala 110:228:@10322.4]
  assign _T_1450 = io_rPort_9_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10324.4]
  assign _T_1453 = _T_1450 & _T_708; // @[MemPrimitives.scala 110:228:@10326.4]
  assign _T_1456 = io_rPort_10_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10328.4]
  assign _T_1459 = _T_1456 & _T_714; // @[MemPrimitives.scala 110:228:@10330.4]
  assign _T_1461 = StickySelects_13_io_outs_0; // @[MemPrimitives.scala 123:41:@10341.4]
  assign _T_1462 = StickySelects_13_io_outs_1; // @[MemPrimitives.scala 123:41:@10342.4]
  assign _T_1463 = StickySelects_13_io_outs_2; // @[MemPrimitives.scala 123:41:@10343.4]
  assign _T_1464 = StickySelects_13_io_outs_3; // @[MemPrimitives.scala 123:41:@10344.4]
  assign _T_1465 = StickySelects_13_io_outs_4; // @[MemPrimitives.scala 123:41:@10345.4]
  assign _T_1466 = StickySelects_13_io_outs_5; // @[MemPrimitives.scala 123:41:@10346.4]
  assign _T_1468 = {_T_1461,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@10348.4]
  assign _T_1470 = {_T_1462,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@10350.4]
  assign _T_1472 = {_T_1463,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@10352.4]
  assign _T_1474 = {_T_1464,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@10354.4]
  assign _T_1476 = {_T_1465,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@10356.4]
  assign _T_1478 = {_T_1466,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@10358.4]
  assign _T_1479 = _T_1465 ? _T_1476 : _T_1478; // @[Mux.scala 31:69:@10359.4]
  assign _T_1480 = _T_1464 ? _T_1474 : _T_1479; // @[Mux.scala 31:69:@10360.4]
  assign _T_1481 = _T_1463 ? _T_1472 : _T_1480; // @[Mux.scala 31:69:@10361.4]
  assign _T_1482 = _T_1462 ? _T_1470 : _T_1481; // @[Mux.scala 31:69:@10362.4]
  assign _T_1483 = _T_1461 ? _T_1468 : _T_1482; // @[Mux.scala 31:69:@10363.4]
  assign _T_1491 = _T_1364 & _T_746; // @[MemPrimitives.scala 110:228:@10372.4]
  assign _T_1497 = _T_1370 & _T_752; // @[MemPrimitives.scala 110:228:@10376.4]
  assign _T_1503 = _T_1376 & _T_758; // @[MemPrimitives.scala 110:228:@10380.4]
  assign _T_1509 = _T_1382 & _T_764; // @[MemPrimitives.scala 110:228:@10384.4]
  assign _T_1515 = _T_1388 & _T_770; // @[MemPrimitives.scala 110:228:@10388.4]
  assign _T_1521 = _T_1394 & _T_776; // @[MemPrimitives.scala 110:228:@10392.4]
  assign _T_1523 = StickySelects_14_io_outs_0; // @[MemPrimitives.scala 123:41:@10403.4]
  assign _T_1524 = StickySelects_14_io_outs_1; // @[MemPrimitives.scala 123:41:@10404.4]
  assign _T_1525 = StickySelects_14_io_outs_2; // @[MemPrimitives.scala 123:41:@10405.4]
  assign _T_1526 = StickySelects_14_io_outs_3; // @[MemPrimitives.scala 123:41:@10406.4]
  assign _T_1527 = StickySelects_14_io_outs_4; // @[MemPrimitives.scala 123:41:@10407.4]
  assign _T_1528 = StickySelects_14_io_outs_5; // @[MemPrimitives.scala 123:41:@10408.4]
  assign _T_1530 = {_T_1523,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@10410.4]
  assign _T_1532 = {_T_1524,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@10412.4]
  assign _T_1534 = {_T_1525,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@10414.4]
  assign _T_1536 = {_T_1526,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@10416.4]
  assign _T_1538 = {_T_1527,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@10418.4]
  assign _T_1540 = {_T_1528,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@10420.4]
  assign _T_1541 = _T_1527 ? _T_1538 : _T_1540; // @[Mux.scala 31:69:@10421.4]
  assign _T_1542 = _T_1526 ? _T_1536 : _T_1541; // @[Mux.scala 31:69:@10422.4]
  assign _T_1543 = _T_1525 ? _T_1534 : _T_1542; // @[Mux.scala 31:69:@10423.4]
  assign _T_1544 = _T_1524 ? _T_1532 : _T_1543; // @[Mux.scala 31:69:@10424.4]
  assign _T_1545 = _T_1523 ? _T_1530 : _T_1544; // @[Mux.scala 31:69:@10425.4]
  assign _T_1553 = _T_1426 & _T_808; // @[MemPrimitives.scala 110:228:@10434.4]
  assign _T_1559 = _T_1432 & _T_814; // @[MemPrimitives.scala 110:228:@10438.4]
  assign _T_1565 = _T_1438 & _T_820; // @[MemPrimitives.scala 110:228:@10442.4]
  assign _T_1571 = _T_1444 & _T_826; // @[MemPrimitives.scala 110:228:@10446.4]
  assign _T_1577 = _T_1450 & _T_832; // @[MemPrimitives.scala 110:228:@10450.4]
  assign _T_1583 = _T_1456 & _T_838; // @[MemPrimitives.scala 110:228:@10454.4]
  assign _T_1585 = StickySelects_15_io_outs_0; // @[MemPrimitives.scala 123:41:@10465.4]
  assign _T_1586 = StickySelects_15_io_outs_1; // @[MemPrimitives.scala 123:41:@10466.4]
  assign _T_1587 = StickySelects_15_io_outs_2; // @[MemPrimitives.scala 123:41:@10467.4]
  assign _T_1588 = StickySelects_15_io_outs_3; // @[MemPrimitives.scala 123:41:@10468.4]
  assign _T_1589 = StickySelects_15_io_outs_4; // @[MemPrimitives.scala 123:41:@10469.4]
  assign _T_1590 = StickySelects_15_io_outs_5; // @[MemPrimitives.scala 123:41:@10470.4]
  assign _T_1592 = {_T_1585,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@10472.4]
  assign _T_1594 = {_T_1586,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@10474.4]
  assign _T_1596 = {_T_1587,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@10476.4]
  assign _T_1598 = {_T_1588,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@10478.4]
  assign _T_1600 = {_T_1589,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@10480.4]
  assign _T_1602 = {_T_1590,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@10482.4]
  assign _T_1603 = _T_1589 ? _T_1600 : _T_1602; // @[Mux.scala 31:69:@10483.4]
  assign _T_1604 = _T_1588 ? _T_1598 : _T_1603; // @[Mux.scala 31:69:@10484.4]
  assign _T_1605 = _T_1587 ? _T_1596 : _T_1604; // @[Mux.scala 31:69:@10485.4]
  assign _T_1606 = _T_1586 ? _T_1594 : _T_1605; // @[Mux.scala 31:69:@10486.4]
  assign _T_1607 = _T_1585 ? _T_1592 : _T_1606; // @[Mux.scala 31:69:@10487.4]
  assign _T_1671 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@10572.4 package.scala 96:25:@10573.4]
  assign _T_1675 = _T_1671 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@10582.4]
  assign _T_1668 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@10564.4 package.scala 96:25:@10565.4]
  assign _T_1676 = _T_1668 ? Mem1D_11_io_output : _T_1675; // @[Mux.scala 31:69:@10583.4]
  assign _T_1665 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@10556.4 package.scala 96:25:@10557.4]
  assign _T_1677 = _T_1665 ? Mem1D_9_io_output : _T_1676; // @[Mux.scala 31:69:@10584.4]
  assign _T_1662 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@10548.4 package.scala 96:25:@10549.4]
  assign _T_1678 = _T_1662 ? Mem1D_7_io_output : _T_1677; // @[Mux.scala 31:69:@10585.4]
  assign _T_1659 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@10540.4 package.scala 96:25:@10541.4]
  assign _T_1679 = _T_1659 ? Mem1D_5_io_output : _T_1678; // @[Mux.scala 31:69:@10586.4]
  assign _T_1656 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@10532.4 package.scala 96:25:@10533.4]
  assign _T_1680 = _T_1656 ? Mem1D_3_io_output : _T_1679; // @[Mux.scala 31:69:@10587.4]
  assign _T_1653 = RetimeWrapper_io_out; // @[package.scala 96:25:@10524.4 package.scala 96:25:@10525.4]
  assign _T_1742 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@10668.4 package.scala 96:25:@10669.4]
  assign _T_1746 = _T_1742 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@10678.4]
  assign _T_1739 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@10660.4 package.scala 96:25:@10661.4]
  assign _T_1747 = _T_1739 ? Mem1D_10_io_output : _T_1746; // @[Mux.scala 31:69:@10679.4]
  assign _T_1736 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@10652.4 package.scala 96:25:@10653.4]
  assign _T_1748 = _T_1736 ? Mem1D_8_io_output : _T_1747; // @[Mux.scala 31:69:@10680.4]
  assign _T_1733 = RetimeWrapper_11_io_out; // @[package.scala 96:25:@10644.4 package.scala 96:25:@10645.4]
  assign _T_1749 = _T_1733 ? Mem1D_6_io_output : _T_1748; // @[Mux.scala 31:69:@10681.4]
  assign _T_1730 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@10636.4 package.scala 96:25:@10637.4]
  assign _T_1750 = _T_1730 ? Mem1D_4_io_output : _T_1749; // @[Mux.scala 31:69:@10682.4]
  assign _T_1727 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@10628.4 package.scala 96:25:@10629.4]
  assign _T_1751 = _T_1727 ? Mem1D_2_io_output : _T_1750; // @[Mux.scala 31:69:@10683.4]
  assign _T_1724 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@10620.4 package.scala 96:25:@10621.4]
  assign _T_1813 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@10764.4 package.scala 96:25:@10765.4]
  assign _T_1817 = _T_1813 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@10774.4]
  assign _T_1810 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@10756.4 package.scala 96:25:@10757.4]
  assign _T_1818 = _T_1810 ? Mem1D_10_io_output : _T_1817; // @[Mux.scala 31:69:@10775.4]
  assign _T_1807 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@10748.4 package.scala 96:25:@10749.4]
  assign _T_1819 = _T_1807 ? Mem1D_8_io_output : _T_1818; // @[Mux.scala 31:69:@10776.4]
  assign _T_1804 = RetimeWrapper_19_io_out; // @[package.scala 96:25:@10740.4 package.scala 96:25:@10741.4]
  assign _T_1820 = _T_1804 ? Mem1D_6_io_output : _T_1819; // @[Mux.scala 31:69:@10777.4]
  assign _T_1801 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@10732.4 package.scala 96:25:@10733.4]
  assign _T_1821 = _T_1801 ? Mem1D_4_io_output : _T_1820; // @[Mux.scala 31:69:@10778.4]
  assign _T_1798 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@10724.4 package.scala 96:25:@10725.4]
  assign _T_1822 = _T_1798 ? Mem1D_2_io_output : _T_1821; // @[Mux.scala 31:69:@10779.4]
  assign _T_1795 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@10716.4 package.scala 96:25:@10717.4]
  assign _T_1884 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@10860.4 package.scala 96:25:@10861.4]
  assign _T_1888 = _T_1884 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@10870.4]
  assign _T_1881 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@10852.4 package.scala 96:25:@10853.4]
  assign _T_1889 = _T_1881 ? Mem1D_10_io_output : _T_1888; // @[Mux.scala 31:69:@10871.4]
  assign _T_1878 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@10844.4 package.scala 96:25:@10845.4]
  assign _T_1890 = _T_1878 ? Mem1D_8_io_output : _T_1889; // @[Mux.scala 31:69:@10872.4]
  assign _T_1875 = RetimeWrapper_27_io_out; // @[package.scala 96:25:@10836.4 package.scala 96:25:@10837.4]
  assign _T_1891 = _T_1875 ? Mem1D_6_io_output : _T_1890; // @[Mux.scala 31:69:@10873.4]
  assign _T_1872 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@10828.4 package.scala 96:25:@10829.4]
  assign _T_1892 = _T_1872 ? Mem1D_4_io_output : _T_1891; // @[Mux.scala 31:69:@10874.4]
  assign _T_1869 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@10820.4 package.scala 96:25:@10821.4]
  assign _T_1893 = _T_1869 ? Mem1D_2_io_output : _T_1892; // @[Mux.scala 31:69:@10875.4]
  assign _T_1866 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@10812.4 package.scala 96:25:@10813.4]
  assign _T_1955 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@10956.4 package.scala 96:25:@10957.4]
  assign _T_1959 = _T_1955 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@10966.4]
  assign _T_1952 = RetimeWrapper_37_io_out; // @[package.scala 96:25:@10948.4 package.scala 96:25:@10949.4]
  assign _T_1960 = _T_1952 ? Mem1D_11_io_output : _T_1959; // @[Mux.scala 31:69:@10967.4]
  assign _T_1949 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@10940.4 package.scala 96:25:@10941.4]
  assign _T_1961 = _T_1949 ? Mem1D_9_io_output : _T_1960; // @[Mux.scala 31:69:@10968.4]
  assign _T_1946 = RetimeWrapper_35_io_out; // @[package.scala 96:25:@10932.4 package.scala 96:25:@10933.4]
  assign _T_1962 = _T_1946 ? Mem1D_7_io_output : _T_1961; // @[Mux.scala 31:69:@10969.4]
  assign _T_1943 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@10924.4 package.scala 96:25:@10925.4]
  assign _T_1963 = _T_1943 ? Mem1D_5_io_output : _T_1962; // @[Mux.scala 31:69:@10970.4]
  assign _T_1940 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@10916.4 package.scala 96:25:@10917.4]
  assign _T_1964 = _T_1940 ? Mem1D_3_io_output : _T_1963; // @[Mux.scala 31:69:@10971.4]
  assign _T_1937 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@10908.4 package.scala 96:25:@10909.4]
  assign _T_2026 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@11052.4 package.scala 96:25:@11053.4]
  assign _T_2030 = _T_2026 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@11062.4]
  assign _T_2023 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@11044.4 package.scala 96:25:@11045.4]
  assign _T_2031 = _T_2023 ? Mem1D_11_io_output : _T_2030; // @[Mux.scala 31:69:@11063.4]
  assign _T_2020 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@11036.4 package.scala 96:25:@11037.4]
  assign _T_2032 = _T_2020 ? Mem1D_9_io_output : _T_2031; // @[Mux.scala 31:69:@11064.4]
  assign _T_2017 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@11028.4 package.scala 96:25:@11029.4]
  assign _T_2033 = _T_2017 ? Mem1D_7_io_output : _T_2032; // @[Mux.scala 31:69:@11065.4]
  assign _T_2014 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@11020.4 package.scala 96:25:@11021.4]
  assign _T_2034 = _T_2014 ? Mem1D_5_io_output : _T_2033; // @[Mux.scala 31:69:@11066.4]
  assign _T_2011 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@11012.4 package.scala 96:25:@11013.4]
  assign _T_2035 = _T_2011 ? Mem1D_3_io_output : _T_2034; // @[Mux.scala 31:69:@11067.4]
  assign _T_2008 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@11004.4 package.scala 96:25:@11005.4]
  assign _T_2097 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@11148.4 package.scala 96:25:@11149.4]
  assign _T_2101 = _T_2097 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@11158.4]
  assign _T_2094 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@11140.4 package.scala 96:25:@11141.4]
  assign _T_2102 = _T_2094 ? Mem1D_10_io_output : _T_2101; // @[Mux.scala 31:69:@11159.4]
  assign _T_2091 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@11132.4 package.scala 96:25:@11133.4]
  assign _T_2103 = _T_2091 ? Mem1D_8_io_output : _T_2102; // @[Mux.scala 31:69:@11160.4]
  assign _T_2088 = RetimeWrapper_51_io_out; // @[package.scala 96:25:@11124.4 package.scala 96:25:@11125.4]
  assign _T_2104 = _T_2088 ? Mem1D_6_io_output : _T_2103; // @[Mux.scala 31:69:@11161.4]
  assign _T_2085 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@11116.4 package.scala 96:25:@11117.4]
  assign _T_2105 = _T_2085 ? Mem1D_4_io_output : _T_2104; // @[Mux.scala 31:69:@11162.4]
  assign _T_2082 = RetimeWrapper_49_io_out; // @[package.scala 96:25:@11108.4 package.scala 96:25:@11109.4]
  assign _T_2106 = _T_2082 ? Mem1D_2_io_output : _T_2105; // @[Mux.scala 31:69:@11163.4]
  assign _T_2079 = RetimeWrapper_48_io_out; // @[package.scala 96:25:@11100.4 package.scala 96:25:@11101.4]
  assign _T_2168 = RetimeWrapper_62_io_out; // @[package.scala 96:25:@11244.4 package.scala 96:25:@11245.4]
  assign _T_2172 = _T_2168 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@11254.4]
  assign _T_2165 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@11236.4 package.scala 96:25:@11237.4]
  assign _T_2173 = _T_2165 ? Mem1D_11_io_output : _T_2172; // @[Mux.scala 31:69:@11255.4]
  assign _T_2162 = RetimeWrapper_60_io_out; // @[package.scala 96:25:@11228.4 package.scala 96:25:@11229.4]
  assign _T_2174 = _T_2162 ? Mem1D_9_io_output : _T_2173; // @[Mux.scala 31:69:@11256.4]
  assign _T_2159 = RetimeWrapper_59_io_out; // @[package.scala 96:25:@11220.4 package.scala 96:25:@11221.4]
  assign _T_2175 = _T_2159 ? Mem1D_7_io_output : _T_2174; // @[Mux.scala 31:69:@11257.4]
  assign _T_2156 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@11212.4 package.scala 96:25:@11213.4]
  assign _T_2176 = _T_2156 ? Mem1D_5_io_output : _T_2175; // @[Mux.scala 31:69:@11258.4]
  assign _T_2153 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@11204.4 package.scala 96:25:@11205.4]
  assign _T_2177 = _T_2153 ? Mem1D_3_io_output : _T_2176; // @[Mux.scala 31:69:@11259.4]
  assign _T_2150 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@11196.4 package.scala 96:25:@11197.4]
  assign _T_2239 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@11340.4 package.scala 96:25:@11341.4]
  assign _T_2243 = _T_2239 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@11350.4]
  assign _T_2236 = RetimeWrapper_69_io_out; // @[package.scala 96:25:@11332.4 package.scala 96:25:@11333.4]
  assign _T_2244 = _T_2236 ? Mem1D_10_io_output : _T_2243; // @[Mux.scala 31:69:@11351.4]
  assign _T_2233 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@11324.4 package.scala 96:25:@11325.4]
  assign _T_2245 = _T_2233 ? Mem1D_8_io_output : _T_2244; // @[Mux.scala 31:69:@11352.4]
  assign _T_2230 = RetimeWrapper_67_io_out; // @[package.scala 96:25:@11316.4 package.scala 96:25:@11317.4]
  assign _T_2246 = _T_2230 ? Mem1D_6_io_output : _T_2245; // @[Mux.scala 31:69:@11353.4]
  assign _T_2227 = RetimeWrapper_66_io_out; // @[package.scala 96:25:@11308.4 package.scala 96:25:@11309.4]
  assign _T_2247 = _T_2227 ? Mem1D_4_io_output : _T_2246; // @[Mux.scala 31:69:@11354.4]
  assign _T_2224 = RetimeWrapper_65_io_out; // @[package.scala 96:25:@11300.4 package.scala 96:25:@11301.4]
  assign _T_2248 = _T_2224 ? Mem1D_2_io_output : _T_2247; // @[Mux.scala 31:69:@11355.4]
  assign _T_2221 = RetimeWrapper_64_io_out; // @[package.scala 96:25:@11292.4 package.scala 96:25:@11293.4]
  assign _T_2310 = RetimeWrapper_78_io_out; // @[package.scala 96:25:@11436.4 package.scala 96:25:@11437.4]
  assign _T_2314 = _T_2310 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@11446.4]
  assign _T_2307 = RetimeWrapper_77_io_out; // @[package.scala 96:25:@11428.4 package.scala 96:25:@11429.4]
  assign _T_2315 = _T_2307 ? Mem1D_11_io_output : _T_2314; // @[Mux.scala 31:69:@11447.4]
  assign _T_2304 = RetimeWrapper_76_io_out; // @[package.scala 96:25:@11420.4 package.scala 96:25:@11421.4]
  assign _T_2316 = _T_2304 ? Mem1D_9_io_output : _T_2315; // @[Mux.scala 31:69:@11448.4]
  assign _T_2301 = RetimeWrapper_75_io_out; // @[package.scala 96:25:@11412.4 package.scala 96:25:@11413.4]
  assign _T_2317 = _T_2301 ? Mem1D_7_io_output : _T_2316; // @[Mux.scala 31:69:@11449.4]
  assign _T_2298 = RetimeWrapper_74_io_out; // @[package.scala 96:25:@11404.4 package.scala 96:25:@11405.4]
  assign _T_2318 = _T_2298 ? Mem1D_5_io_output : _T_2317; // @[Mux.scala 31:69:@11450.4]
  assign _T_2295 = RetimeWrapper_73_io_out; // @[package.scala 96:25:@11396.4 package.scala 96:25:@11397.4]
  assign _T_2319 = _T_2295 ? Mem1D_3_io_output : _T_2318; // @[Mux.scala 31:69:@11451.4]
  assign _T_2292 = RetimeWrapper_72_io_out; // @[package.scala 96:25:@11388.4 package.scala 96:25:@11389.4]
  assign _T_2381 = RetimeWrapper_86_io_out; // @[package.scala 96:25:@11532.4 package.scala 96:25:@11533.4]
  assign _T_2385 = _T_2381 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@11542.4]
  assign _T_2378 = RetimeWrapper_85_io_out; // @[package.scala 96:25:@11524.4 package.scala 96:25:@11525.4]
  assign _T_2386 = _T_2378 ? Mem1D_11_io_output : _T_2385; // @[Mux.scala 31:69:@11543.4]
  assign _T_2375 = RetimeWrapper_84_io_out; // @[package.scala 96:25:@11516.4 package.scala 96:25:@11517.4]
  assign _T_2387 = _T_2375 ? Mem1D_9_io_output : _T_2386; // @[Mux.scala 31:69:@11544.4]
  assign _T_2372 = RetimeWrapper_83_io_out; // @[package.scala 96:25:@11508.4 package.scala 96:25:@11509.4]
  assign _T_2388 = _T_2372 ? Mem1D_7_io_output : _T_2387; // @[Mux.scala 31:69:@11545.4]
  assign _T_2369 = RetimeWrapper_82_io_out; // @[package.scala 96:25:@11500.4 package.scala 96:25:@11501.4]
  assign _T_2389 = _T_2369 ? Mem1D_5_io_output : _T_2388; // @[Mux.scala 31:69:@11546.4]
  assign _T_2366 = RetimeWrapper_81_io_out; // @[package.scala 96:25:@11492.4 package.scala 96:25:@11493.4]
  assign _T_2390 = _T_2366 ? Mem1D_3_io_output : _T_2389; // @[Mux.scala 31:69:@11547.4]
  assign _T_2363 = RetimeWrapper_80_io_out; // @[package.scala 96:25:@11484.4 package.scala 96:25:@11485.4]
  assign _T_2452 = RetimeWrapper_94_io_out; // @[package.scala 96:25:@11628.4 package.scala 96:25:@11629.4]
  assign _T_2456 = _T_2452 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@11638.4]
  assign _T_2449 = RetimeWrapper_93_io_out; // @[package.scala 96:25:@11620.4 package.scala 96:25:@11621.4]
  assign _T_2457 = _T_2449 ? Mem1D_10_io_output : _T_2456; // @[Mux.scala 31:69:@11639.4]
  assign _T_2446 = RetimeWrapper_92_io_out; // @[package.scala 96:25:@11612.4 package.scala 96:25:@11613.4]
  assign _T_2458 = _T_2446 ? Mem1D_8_io_output : _T_2457; // @[Mux.scala 31:69:@11640.4]
  assign _T_2443 = RetimeWrapper_91_io_out; // @[package.scala 96:25:@11604.4 package.scala 96:25:@11605.4]
  assign _T_2459 = _T_2443 ? Mem1D_6_io_output : _T_2458; // @[Mux.scala 31:69:@11641.4]
  assign _T_2440 = RetimeWrapper_90_io_out; // @[package.scala 96:25:@11596.4 package.scala 96:25:@11597.4]
  assign _T_2460 = _T_2440 ? Mem1D_4_io_output : _T_2459; // @[Mux.scala 31:69:@11642.4]
  assign _T_2437 = RetimeWrapper_89_io_out; // @[package.scala 96:25:@11588.4 package.scala 96:25:@11589.4]
  assign _T_2461 = _T_2437 ? Mem1D_2_io_output : _T_2460; // @[Mux.scala 31:69:@11643.4]
  assign _T_2434 = RetimeWrapper_88_io_out; // @[package.scala 96:25:@11580.4 package.scala 96:25:@11581.4]
  assign io_rPort_11_output_0 = _T_2434 ? Mem1D_io_output : _T_2461; // @[MemPrimitives.scala 148:13:@11645.4]
  assign io_rPort_10_output_0 = _T_2363 ? Mem1D_1_io_output : _T_2390; // @[MemPrimitives.scala 148:13:@11549.4]
  assign io_rPort_9_output_0 = _T_2292 ? Mem1D_1_io_output : _T_2319; // @[MemPrimitives.scala 148:13:@11453.4]
  assign io_rPort_8_output_0 = _T_2221 ? Mem1D_io_output : _T_2248; // @[MemPrimitives.scala 148:13:@11357.4]
  assign io_rPort_7_output_0 = _T_2150 ? Mem1D_1_io_output : _T_2177; // @[MemPrimitives.scala 148:13:@11261.4]
  assign io_rPort_6_output_0 = _T_2079 ? Mem1D_io_output : _T_2106; // @[MemPrimitives.scala 148:13:@11165.4]
  assign io_rPort_5_output_0 = _T_2008 ? Mem1D_1_io_output : _T_2035; // @[MemPrimitives.scala 148:13:@11069.4]
  assign io_rPort_4_output_0 = _T_1937 ? Mem1D_1_io_output : _T_1964; // @[MemPrimitives.scala 148:13:@10973.4]
  assign io_rPort_3_output_0 = _T_1866 ? Mem1D_io_output : _T_1893; // @[MemPrimitives.scala 148:13:@10877.4]
  assign io_rPort_2_output_0 = _T_1795 ? Mem1D_io_output : _T_1822; // @[MemPrimitives.scala 148:13:@10781.4]
  assign io_rPort_1_output_0 = _T_1724 ? Mem1D_io_output : _T_1751; // @[MemPrimitives.scala 148:13:@10685.4]
  assign io_rPort_0_output_0 = _T_1653 ? Mem1D_1_io_output : _T_1680; // @[MemPrimitives.scala 148:13:@10589.4]
  assign Mem1D_clock = clock; // @[:@9055.4]
  assign Mem1D_reset = reset; // @[:@9056.4]
  assign Mem1D_io_r_ofs_0 = _T_677[0]; // @[MemPrimitives.scala 127:28:@9561.4]
  assign Mem1D_io_r_backpressure = _T_677[1]; // @[MemPrimitives.scala 128:32:@9562.4]
  assign Mem1D_io_w_ofs_0 = _T_450[0]; // @[MemPrimitives.scala 94:28:@9319.4]
  assign Mem1D_io_w_data_0 = _T_450[8:1]; // @[MemPrimitives.scala 95:29:@9320.4]
  assign Mem1D_io_w_en_0 = _T_450[9]; // @[MemPrimitives.scala 96:27:@9321.4]
  assign Mem1D_1_clock = clock; // @[:@9071.4]
  assign Mem1D_1_reset = reset; // @[:@9072.4]
  assign Mem1D_1_io_r_ofs_0 = _T_739[0]; // @[MemPrimitives.scala 127:28:@9623.4]
  assign Mem1D_1_io_r_backpressure = _T_739[1]; // @[MemPrimitives.scala 128:32:@9624.4]
  assign Mem1D_1_io_w_ofs_0 = _T_461[0]; // @[MemPrimitives.scala 94:28:@9331.4]
  assign Mem1D_1_io_w_data_0 = _T_461[8:1]; // @[MemPrimitives.scala 95:29:@9332.4]
  assign Mem1D_1_io_w_en_0 = _T_461[9]; // @[MemPrimitives.scala 96:27:@9333.4]
  assign Mem1D_2_clock = clock; // @[:@9087.4]
  assign Mem1D_2_reset = reset; // @[:@9088.4]
  assign Mem1D_2_io_r_ofs_0 = _T_801[0]; // @[MemPrimitives.scala 127:28:@9685.4]
  assign Mem1D_2_io_r_backpressure = _T_801[1]; // @[MemPrimitives.scala 128:32:@9686.4]
  assign Mem1D_2_io_w_ofs_0 = _T_472[0]; // @[MemPrimitives.scala 94:28:@9343.4]
  assign Mem1D_2_io_w_data_0 = _T_472[8:1]; // @[MemPrimitives.scala 95:29:@9344.4]
  assign Mem1D_2_io_w_en_0 = _T_472[9]; // @[MemPrimitives.scala 96:27:@9345.4]
  assign Mem1D_3_clock = clock; // @[:@9103.4]
  assign Mem1D_3_reset = reset; // @[:@9104.4]
  assign Mem1D_3_io_r_ofs_0 = _T_863[0]; // @[MemPrimitives.scala 127:28:@9747.4]
  assign Mem1D_3_io_r_backpressure = _T_863[1]; // @[MemPrimitives.scala 128:32:@9748.4]
  assign Mem1D_3_io_w_ofs_0 = _T_483[0]; // @[MemPrimitives.scala 94:28:@9355.4]
  assign Mem1D_3_io_w_data_0 = _T_483[8:1]; // @[MemPrimitives.scala 95:29:@9356.4]
  assign Mem1D_3_io_w_en_0 = _T_483[9]; // @[MemPrimitives.scala 96:27:@9357.4]
  assign Mem1D_4_clock = clock; // @[:@9119.4]
  assign Mem1D_4_reset = reset; // @[:@9120.4]
  assign Mem1D_4_io_r_ofs_0 = _T_925[0]; // @[MemPrimitives.scala 127:28:@9809.4]
  assign Mem1D_4_io_r_backpressure = _T_925[1]; // @[MemPrimitives.scala 128:32:@9810.4]
  assign Mem1D_4_io_w_ofs_0 = _T_494[0]; // @[MemPrimitives.scala 94:28:@9367.4]
  assign Mem1D_4_io_w_data_0 = _T_494[8:1]; // @[MemPrimitives.scala 95:29:@9368.4]
  assign Mem1D_4_io_w_en_0 = _T_494[9]; // @[MemPrimitives.scala 96:27:@9369.4]
  assign Mem1D_5_clock = clock; // @[:@9135.4]
  assign Mem1D_5_reset = reset; // @[:@9136.4]
  assign Mem1D_5_io_r_ofs_0 = _T_987[0]; // @[MemPrimitives.scala 127:28:@9871.4]
  assign Mem1D_5_io_r_backpressure = _T_987[1]; // @[MemPrimitives.scala 128:32:@9872.4]
  assign Mem1D_5_io_w_ofs_0 = _T_505[0]; // @[MemPrimitives.scala 94:28:@9379.4]
  assign Mem1D_5_io_w_data_0 = _T_505[8:1]; // @[MemPrimitives.scala 95:29:@9380.4]
  assign Mem1D_5_io_w_en_0 = _T_505[9]; // @[MemPrimitives.scala 96:27:@9381.4]
  assign Mem1D_6_clock = clock; // @[:@9151.4]
  assign Mem1D_6_reset = reset; // @[:@9152.4]
  assign Mem1D_6_io_r_ofs_0 = _T_1049[0]; // @[MemPrimitives.scala 127:28:@9933.4]
  assign Mem1D_6_io_r_backpressure = _T_1049[1]; // @[MemPrimitives.scala 128:32:@9934.4]
  assign Mem1D_6_io_w_ofs_0 = _T_516[0]; // @[MemPrimitives.scala 94:28:@9391.4]
  assign Mem1D_6_io_w_data_0 = _T_516[8:1]; // @[MemPrimitives.scala 95:29:@9392.4]
  assign Mem1D_6_io_w_en_0 = _T_516[9]; // @[MemPrimitives.scala 96:27:@9393.4]
  assign Mem1D_7_clock = clock; // @[:@9167.4]
  assign Mem1D_7_reset = reset; // @[:@9168.4]
  assign Mem1D_7_io_r_ofs_0 = _T_1111[0]; // @[MemPrimitives.scala 127:28:@9995.4]
  assign Mem1D_7_io_r_backpressure = _T_1111[1]; // @[MemPrimitives.scala 128:32:@9996.4]
  assign Mem1D_7_io_w_ofs_0 = _T_527[0]; // @[MemPrimitives.scala 94:28:@9403.4]
  assign Mem1D_7_io_w_data_0 = _T_527[8:1]; // @[MemPrimitives.scala 95:29:@9404.4]
  assign Mem1D_7_io_w_en_0 = _T_527[9]; // @[MemPrimitives.scala 96:27:@9405.4]
  assign Mem1D_8_clock = clock; // @[:@9183.4]
  assign Mem1D_8_reset = reset; // @[:@9184.4]
  assign Mem1D_8_io_r_ofs_0 = _T_1173[0]; // @[MemPrimitives.scala 127:28:@10057.4]
  assign Mem1D_8_io_r_backpressure = _T_1173[1]; // @[MemPrimitives.scala 128:32:@10058.4]
  assign Mem1D_8_io_w_ofs_0 = _T_538[0]; // @[MemPrimitives.scala 94:28:@9415.4]
  assign Mem1D_8_io_w_data_0 = _T_538[8:1]; // @[MemPrimitives.scala 95:29:@9416.4]
  assign Mem1D_8_io_w_en_0 = _T_538[9]; // @[MemPrimitives.scala 96:27:@9417.4]
  assign Mem1D_9_clock = clock; // @[:@9199.4]
  assign Mem1D_9_reset = reset; // @[:@9200.4]
  assign Mem1D_9_io_r_ofs_0 = _T_1235[0]; // @[MemPrimitives.scala 127:28:@10119.4]
  assign Mem1D_9_io_r_backpressure = _T_1235[1]; // @[MemPrimitives.scala 128:32:@10120.4]
  assign Mem1D_9_io_w_ofs_0 = _T_549[0]; // @[MemPrimitives.scala 94:28:@9427.4]
  assign Mem1D_9_io_w_data_0 = _T_549[8:1]; // @[MemPrimitives.scala 95:29:@9428.4]
  assign Mem1D_9_io_w_en_0 = _T_549[9]; // @[MemPrimitives.scala 96:27:@9429.4]
  assign Mem1D_10_clock = clock; // @[:@9215.4]
  assign Mem1D_10_reset = reset; // @[:@9216.4]
  assign Mem1D_10_io_r_ofs_0 = _T_1297[0]; // @[MemPrimitives.scala 127:28:@10181.4]
  assign Mem1D_10_io_r_backpressure = _T_1297[1]; // @[MemPrimitives.scala 128:32:@10182.4]
  assign Mem1D_10_io_w_ofs_0 = _T_560[0]; // @[MemPrimitives.scala 94:28:@9439.4]
  assign Mem1D_10_io_w_data_0 = _T_560[8:1]; // @[MemPrimitives.scala 95:29:@9440.4]
  assign Mem1D_10_io_w_en_0 = _T_560[9]; // @[MemPrimitives.scala 96:27:@9441.4]
  assign Mem1D_11_clock = clock; // @[:@9231.4]
  assign Mem1D_11_reset = reset; // @[:@9232.4]
  assign Mem1D_11_io_r_ofs_0 = _T_1359[0]; // @[MemPrimitives.scala 127:28:@10243.4]
  assign Mem1D_11_io_r_backpressure = _T_1359[1]; // @[MemPrimitives.scala 128:32:@10244.4]
  assign Mem1D_11_io_w_ofs_0 = _T_571[0]; // @[MemPrimitives.scala 94:28:@9451.4]
  assign Mem1D_11_io_w_data_0 = _T_571[8:1]; // @[MemPrimitives.scala 95:29:@9452.4]
  assign Mem1D_11_io_w_en_0 = _T_571[9]; // @[MemPrimitives.scala 96:27:@9453.4]
  assign Mem1D_12_clock = clock; // @[:@9247.4]
  assign Mem1D_12_reset = reset; // @[:@9248.4]
  assign Mem1D_12_io_r_ofs_0 = _T_1421[0]; // @[MemPrimitives.scala 127:28:@10305.4]
  assign Mem1D_12_io_r_backpressure = _T_1421[1]; // @[MemPrimitives.scala 128:32:@10306.4]
  assign Mem1D_12_io_w_ofs_0 = _T_582[0]; // @[MemPrimitives.scala 94:28:@9463.4]
  assign Mem1D_12_io_w_data_0 = _T_582[8:1]; // @[MemPrimitives.scala 95:29:@9464.4]
  assign Mem1D_12_io_w_en_0 = _T_582[9]; // @[MemPrimitives.scala 96:27:@9465.4]
  assign Mem1D_13_clock = clock; // @[:@9263.4]
  assign Mem1D_13_reset = reset; // @[:@9264.4]
  assign Mem1D_13_io_r_ofs_0 = _T_1483[0]; // @[MemPrimitives.scala 127:28:@10367.4]
  assign Mem1D_13_io_r_backpressure = _T_1483[1]; // @[MemPrimitives.scala 128:32:@10368.4]
  assign Mem1D_13_io_w_ofs_0 = _T_593[0]; // @[MemPrimitives.scala 94:28:@9475.4]
  assign Mem1D_13_io_w_data_0 = _T_593[8:1]; // @[MemPrimitives.scala 95:29:@9476.4]
  assign Mem1D_13_io_w_en_0 = _T_593[9]; // @[MemPrimitives.scala 96:27:@9477.4]
  assign Mem1D_14_clock = clock; // @[:@9279.4]
  assign Mem1D_14_reset = reset; // @[:@9280.4]
  assign Mem1D_14_io_r_ofs_0 = _T_1545[0]; // @[MemPrimitives.scala 127:28:@10429.4]
  assign Mem1D_14_io_r_backpressure = _T_1545[1]; // @[MemPrimitives.scala 128:32:@10430.4]
  assign Mem1D_14_io_w_ofs_0 = _T_604[0]; // @[MemPrimitives.scala 94:28:@9487.4]
  assign Mem1D_14_io_w_data_0 = _T_604[8:1]; // @[MemPrimitives.scala 95:29:@9488.4]
  assign Mem1D_14_io_w_en_0 = _T_604[9]; // @[MemPrimitives.scala 96:27:@9489.4]
  assign Mem1D_15_clock = clock; // @[:@9295.4]
  assign Mem1D_15_reset = reset; // @[:@9296.4]
  assign Mem1D_15_io_r_ofs_0 = _T_1607[0]; // @[MemPrimitives.scala 127:28:@10491.4]
  assign Mem1D_15_io_r_backpressure = _T_1607[1]; // @[MemPrimitives.scala 128:32:@10492.4]
  assign Mem1D_15_io_w_ofs_0 = _T_615[0]; // @[MemPrimitives.scala 94:28:@9499.4]
  assign Mem1D_15_io_w_data_0 = _T_615[8:1]; // @[MemPrimitives.scala 95:29:@9500.4]
  assign Mem1D_15_io_w_en_0 = _T_615[9]; // @[MemPrimitives.scala 96:27:@9501.4]
  assign StickySelects_clock = clock; // @[:@9527.4]
  assign StickySelects_reset = reset; // @[:@9528.4]
  assign StickySelects_io_ins_0 = io_rPort_1_en_0 & _T_623; // @[MemPrimitives.scala 122:60:@9529.4]
  assign StickySelects_io_ins_1 = io_rPort_2_en_0 & _T_629; // @[MemPrimitives.scala 122:60:@9530.4]
  assign StickySelects_io_ins_2 = io_rPort_3_en_0 & _T_635; // @[MemPrimitives.scala 122:60:@9531.4]
  assign StickySelects_io_ins_3 = io_rPort_6_en_0 & _T_641; // @[MemPrimitives.scala 122:60:@9532.4]
  assign StickySelects_io_ins_4 = io_rPort_8_en_0 & _T_647; // @[MemPrimitives.scala 122:60:@9533.4]
  assign StickySelects_io_ins_5 = io_rPort_11_en_0 & _T_653; // @[MemPrimitives.scala 122:60:@9534.4]
  assign StickySelects_1_clock = clock; // @[:@9589.4]
  assign StickySelects_1_reset = reset; // @[:@9590.4]
  assign StickySelects_1_io_ins_0 = io_rPort_0_en_0 & _T_685; // @[MemPrimitives.scala 122:60:@9591.4]
  assign StickySelects_1_io_ins_1 = io_rPort_4_en_0 & _T_691; // @[MemPrimitives.scala 122:60:@9592.4]
  assign StickySelects_1_io_ins_2 = io_rPort_5_en_0 & _T_697; // @[MemPrimitives.scala 122:60:@9593.4]
  assign StickySelects_1_io_ins_3 = io_rPort_7_en_0 & _T_703; // @[MemPrimitives.scala 122:60:@9594.4]
  assign StickySelects_1_io_ins_4 = io_rPort_9_en_0 & _T_709; // @[MemPrimitives.scala 122:60:@9595.4]
  assign StickySelects_1_io_ins_5 = io_rPort_10_en_0 & _T_715; // @[MemPrimitives.scala 122:60:@9596.4]
  assign StickySelects_2_clock = clock; // @[:@9651.4]
  assign StickySelects_2_reset = reset; // @[:@9652.4]
  assign StickySelects_2_io_ins_0 = io_rPort_1_en_0 & _T_747; // @[MemPrimitives.scala 122:60:@9653.4]
  assign StickySelects_2_io_ins_1 = io_rPort_2_en_0 & _T_753; // @[MemPrimitives.scala 122:60:@9654.4]
  assign StickySelects_2_io_ins_2 = io_rPort_3_en_0 & _T_759; // @[MemPrimitives.scala 122:60:@9655.4]
  assign StickySelects_2_io_ins_3 = io_rPort_6_en_0 & _T_765; // @[MemPrimitives.scala 122:60:@9656.4]
  assign StickySelects_2_io_ins_4 = io_rPort_8_en_0 & _T_771; // @[MemPrimitives.scala 122:60:@9657.4]
  assign StickySelects_2_io_ins_5 = io_rPort_11_en_0 & _T_777; // @[MemPrimitives.scala 122:60:@9658.4]
  assign StickySelects_3_clock = clock; // @[:@9713.4]
  assign StickySelects_3_reset = reset; // @[:@9714.4]
  assign StickySelects_3_io_ins_0 = io_rPort_0_en_0 & _T_809; // @[MemPrimitives.scala 122:60:@9715.4]
  assign StickySelects_3_io_ins_1 = io_rPort_4_en_0 & _T_815; // @[MemPrimitives.scala 122:60:@9716.4]
  assign StickySelects_3_io_ins_2 = io_rPort_5_en_0 & _T_821; // @[MemPrimitives.scala 122:60:@9717.4]
  assign StickySelects_3_io_ins_3 = io_rPort_7_en_0 & _T_827; // @[MemPrimitives.scala 122:60:@9718.4]
  assign StickySelects_3_io_ins_4 = io_rPort_9_en_0 & _T_833; // @[MemPrimitives.scala 122:60:@9719.4]
  assign StickySelects_3_io_ins_5 = io_rPort_10_en_0 & _T_839; // @[MemPrimitives.scala 122:60:@9720.4]
  assign StickySelects_4_clock = clock; // @[:@9775.4]
  assign StickySelects_4_reset = reset; // @[:@9776.4]
  assign StickySelects_4_io_ins_0 = io_rPort_1_en_0 & _T_871; // @[MemPrimitives.scala 122:60:@9777.4]
  assign StickySelects_4_io_ins_1 = io_rPort_2_en_0 & _T_877; // @[MemPrimitives.scala 122:60:@9778.4]
  assign StickySelects_4_io_ins_2 = io_rPort_3_en_0 & _T_883; // @[MemPrimitives.scala 122:60:@9779.4]
  assign StickySelects_4_io_ins_3 = io_rPort_6_en_0 & _T_889; // @[MemPrimitives.scala 122:60:@9780.4]
  assign StickySelects_4_io_ins_4 = io_rPort_8_en_0 & _T_895; // @[MemPrimitives.scala 122:60:@9781.4]
  assign StickySelects_4_io_ins_5 = io_rPort_11_en_0 & _T_901; // @[MemPrimitives.scala 122:60:@9782.4]
  assign StickySelects_5_clock = clock; // @[:@9837.4]
  assign StickySelects_5_reset = reset; // @[:@9838.4]
  assign StickySelects_5_io_ins_0 = io_rPort_0_en_0 & _T_933; // @[MemPrimitives.scala 122:60:@9839.4]
  assign StickySelects_5_io_ins_1 = io_rPort_4_en_0 & _T_939; // @[MemPrimitives.scala 122:60:@9840.4]
  assign StickySelects_5_io_ins_2 = io_rPort_5_en_0 & _T_945; // @[MemPrimitives.scala 122:60:@9841.4]
  assign StickySelects_5_io_ins_3 = io_rPort_7_en_0 & _T_951; // @[MemPrimitives.scala 122:60:@9842.4]
  assign StickySelects_5_io_ins_4 = io_rPort_9_en_0 & _T_957; // @[MemPrimitives.scala 122:60:@9843.4]
  assign StickySelects_5_io_ins_5 = io_rPort_10_en_0 & _T_963; // @[MemPrimitives.scala 122:60:@9844.4]
  assign StickySelects_6_clock = clock; // @[:@9899.4]
  assign StickySelects_6_reset = reset; // @[:@9900.4]
  assign StickySelects_6_io_ins_0 = io_rPort_1_en_0 & _T_995; // @[MemPrimitives.scala 122:60:@9901.4]
  assign StickySelects_6_io_ins_1 = io_rPort_2_en_0 & _T_1001; // @[MemPrimitives.scala 122:60:@9902.4]
  assign StickySelects_6_io_ins_2 = io_rPort_3_en_0 & _T_1007; // @[MemPrimitives.scala 122:60:@9903.4]
  assign StickySelects_6_io_ins_3 = io_rPort_6_en_0 & _T_1013; // @[MemPrimitives.scala 122:60:@9904.4]
  assign StickySelects_6_io_ins_4 = io_rPort_8_en_0 & _T_1019; // @[MemPrimitives.scala 122:60:@9905.4]
  assign StickySelects_6_io_ins_5 = io_rPort_11_en_0 & _T_1025; // @[MemPrimitives.scala 122:60:@9906.4]
  assign StickySelects_7_clock = clock; // @[:@9961.4]
  assign StickySelects_7_reset = reset; // @[:@9962.4]
  assign StickySelects_7_io_ins_0 = io_rPort_0_en_0 & _T_1057; // @[MemPrimitives.scala 122:60:@9963.4]
  assign StickySelects_7_io_ins_1 = io_rPort_4_en_0 & _T_1063; // @[MemPrimitives.scala 122:60:@9964.4]
  assign StickySelects_7_io_ins_2 = io_rPort_5_en_0 & _T_1069; // @[MemPrimitives.scala 122:60:@9965.4]
  assign StickySelects_7_io_ins_3 = io_rPort_7_en_0 & _T_1075; // @[MemPrimitives.scala 122:60:@9966.4]
  assign StickySelects_7_io_ins_4 = io_rPort_9_en_0 & _T_1081; // @[MemPrimitives.scala 122:60:@9967.4]
  assign StickySelects_7_io_ins_5 = io_rPort_10_en_0 & _T_1087; // @[MemPrimitives.scala 122:60:@9968.4]
  assign StickySelects_8_clock = clock; // @[:@10023.4]
  assign StickySelects_8_reset = reset; // @[:@10024.4]
  assign StickySelects_8_io_ins_0 = io_rPort_1_en_0 & _T_1119; // @[MemPrimitives.scala 122:60:@10025.4]
  assign StickySelects_8_io_ins_1 = io_rPort_2_en_0 & _T_1125; // @[MemPrimitives.scala 122:60:@10026.4]
  assign StickySelects_8_io_ins_2 = io_rPort_3_en_0 & _T_1131; // @[MemPrimitives.scala 122:60:@10027.4]
  assign StickySelects_8_io_ins_3 = io_rPort_6_en_0 & _T_1137; // @[MemPrimitives.scala 122:60:@10028.4]
  assign StickySelects_8_io_ins_4 = io_rPort_8_en_0 & _T_1143; // @[MemPrimitives.scala 122:60:@10029.4]
  assign StickySelects_8_io_ins_5 = io_rPort_11_en_0 & _T_1149; // @[MemPrimitives.scala 122:60:@10030.4]
  assign StickySelects_9_clock = clock; // @[:@10085.4]
  assign StickySelects_9_reset = reset; // @[:@10086.4]
  assign StickySelects_9_io_ins_0 = io_rPort_0_en_0 & _T_1181; // @[MemPrimitives.scala 122:60:@10087.4]
  assign StickySelects_9_io_ins_1 = io_rPort_4_en_0 & _T_1187; // @[MemPrimitives.scala 122:60:@10088.4]
  assign StickySelects_9_io_ins_2 = io_rPort_5_en_0 & _T_1193; // @[MemPrimitives.scala 122:60:@10089.4]
  assign StickySelects_9_io_ins_3 = io_rPort_7_en_0 & _T_1199; // @[MemPrimitives.scala 122:60:@10090.4]
  assign StickySelects_9_io_ins_4 = io_rPort_9_en_0 & _T_1205; // @[MemPrimitives.scala 122:60:@10091.4]
  assign StickySelects_9_io_ins_5 = io_rPort_10_en_0 & _T_1211; // @[MemPrimitives.scala 122:60:@10092.4]
  assign StickySelects_10_clock = clock; // @[:@10147.4]
  assign StickySelects_10_reset = reset; // @[:@10148.4]
  assign StickySelects_10_io_ins_0 = io_rPort_1_en_0 & _T_1243; // @[MemPrimitives.scala 122:60:@10149.4]
  assign StickySelects_10_io_ins_1 = io_rPort_2_en_0 & _T_1249; // @[MemPrimitives.scala 122:60:@10150.4]
  assign StickySelects_10_io_ins_2 = io_rPort_3_en_0 & _T_1255; // @[MemPrimitives.scala 122:60:@10151.4]
  assign StickySelects_10_io_ins_3 = io_rPort_6_en_0 & _T_1261; // @[MemPrimitives.scala 122:60:@10152.4]
  assign StickySelects_10_io_ins_4 = io_rPort_8_en_0 & _T_1267; // @[MemPrimitives.scala 122:60:@10153.4]
  assign StickySelects_10_io_ins_5 = io_rPort_11_en_0 & _T_1273; // @[MemPrimitives.scala 122:60:@10154.4]
  assign StickySelects_11_clock = clock; // @[:@10209.4]
  assign StickySelects_11_reset = reset; // @[:@10210.4]
  assign StickySelects_11_io_ins_0 = io_rPort_0_en_0 & _T_1305; // @[MemPrimitives.scala 122:60:@10211.4]
  assign StickySelects_11_io_ins_1 = io_rPort_4_en_0 & _T_1311; // @[MemPrimitives.scala 122:60:@10212.4]
  assign StickySelects_11_io_ins_2 = io_rPort_5_en_0 & _T_1317; // @[MemPrimitives.scala 122:60:@10213.4]
  assign StickySelects_11_io_ins_3 = io_rPort_7_en_0 & _T_1323; // @[MemPrimitives.scala 122:60:@10214.4]
  assign StickySelects_11_io_ins_4 = io_rPort_9_en_0 & _T_1329; // @[MemPrimitives.scala 122:60:@10215.4]
  assign StickySelects_11_io_ins_5 = io_rPort_10_en_0 & _T_1335; // @[MemPrimitives.scala 122:60:@10216.4]
  assign StickySelects_12_clock = clock; // @[:@10271.4]
  assign StickySelects_12_reset = reset; // @[:@10272.4]
  assign StickySelects_12_io_ins_0 = io_rPort_1_en_0 & _T_1367; // @[MemPrimitives.scala 122:60:@10273.4]
  assign StickySelects_12_io_ins_1 = io_rPort_2_en_0 & _T_1373; // @[MemPrimitives.scala 122:60:@10274.4]
  assign StickySelects_12_io_ins_2 = io_rPort_3_en_0 & _T_1379; // @[MemPrimitives.scala 122:60:@10275.4]
  assign StickySelects_12_io_ins_3 = io_rPort_6_en_0 & _T_1385; // @[MemPrimitives.scala 122:60:@10276.4]
  assign StickySelects_12_io_ins_4 = io_rPort_8_en_0 & _T_1391; // @[MemPrimitives.scala 122:60:@10277.4]
  assign StickySelects_12_io_ins_5 = io_rPort_11_en_0 & _T_1397; // @[MemPrimitives.scala 122:60:@10278.4]
  assign StickySelects_13_clock = clock; // @[:@10333.4]
  assign StickySelects_13_reset = reset; // @[:@10334.4]
  assign StickySelects_13_io_ins_0 = io_rPort_0_en_0 & _T_1429; // @[MemPrimitives.scala 122:60:@10335.4]
  assign StickySelects_13_io_ins_1 = io_rPort_4_en_0 & _T_1435; // @[MemPrimitives.scala 122:60:@10336.4]
  assign StickySelects_13_io_ins_2 = io_rPort_5_en_0 & _T_1441; // @[MemPrimitives.scala 122:60:@10337.4]
  assign StickySelects_13_io_ins_3 = io_rPort_7_en_0 & _T_1447; // @[MemPrimitives.scala 122:60:@10338.4]
  assign StickySelects_13_io_ins_4 = io_rPort_9_en_0 & _T_1453; // @[MemPrimitives.scala 122:60:@10339.4]
  assign StickySelects_13_io_ins_5 = io_rPort_10_en_0 & _T_1459; // @[MemPrimitives.scala 122:60:@10340.4]
  assign StickySelects_14_clock = clock; // @[:@10395.4]
  assign StickySelects_14_reset = reset; // @[:@10396.4]
  assign StickySelects_14_io_ins_0 = io_rPort_1_en_0 & _T_1491; // @[MemPrimitives.scala 122:60:@10397.4]
  assign StickySelects_14_io_ins_1 = io_rPort_2_en_0 & _T_1497; // @[MemPrimitives.scala 122:60:@10398.4]
  assign StickySelects_14_io_ins_2 = io_rPort_3_en_0 & _T_1503; // @[MemPrimitives.scala 122:60:@10399.4]
  assign StickySelects_14_io_ins_3 = io_rPort_6_en_0 & _T_1509; // @[MemPrimitives.scala 122:60:@10400.4]
  assign StickySelects_14_io_ins_4 = io_rPort_8_en_0 & _T_1515; // @[MemPrimitives.scala 122:60:@10401.4]
  assign StickySelects_14_io_ins_5 = io_rPort_11_en_0 & _T_1521; // @[MemPrimitives.scala 122:60:@10402.4]
  assign StickySelects_15_clock = clock; // @[:@10457.4]
  assign StickySelects_15_reset = reset; // @[:@10458.4]
  assign StickySelects_15_io_ins_0 = io_rPort_0_en_0 & _T_1553; // @[MemPrimitives.scala 122:60:@10459.4]
  assign StickySelects_15_io_ins_1 = io_rPort_4_en_0 & _T_1559; // @[MemPrimitives.scala 122:60:@10460.4]
  assign StickySelects_15_io_ins_2 = io_rPort_5_en_0 & _T_1565; // @[MemPrimitives.scala 122:60:@10461.4]
  assign StickySelects_15_io_ins_3 = io_rPort_7_en_0 & _T_1571; // @[MemPrimitives.scala 122:60:@10462.4]
  assign StickySelects_15_io_ins_4 = io_rPort_9_en_0 & _T_1577; // @[MemPrimitives.scala 122:60:@10463.4]
  assign StickySelects_15_io_ins_5 = io_rPort_10_en_0 & _T_1583; // @[MemPrimitives.scala 122:60:@10464.4]
  assign RetimeWrapper_clock = clock; // @[:@10520.4]
  assign RetimeWrapper_reset = reset; // @[:@10521.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@10523.4]
  assign RetimeWrapper_io_in = _T_685 & io_rPort_0_en_0; // @[package.scala 94:16:@10522.4]
  assign RetimeWrapper_1_clock = clock; // @[:@10528.4]
  assign RetimeWrapper_1_reset = reset; // @[:@10529.4]
  assign RetimeWrapper_1_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@10531.4]
  assign RetimeWrapper_1_io_in = _T_809 & io_rPort_0_en_0; // @[package.scala 94:16:@10530.4]
  assign RetimeWrapper_2_clock = clock; // @[:@10536.4]
  assign RetimeWrapper_2_reset = reset; // @[:@10537.4]
  assign RetimeWrapper_2_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@10539.4]
  assign RetimeWrapper_2_io_in = _T_933 & io_rPort_0_en_0; // @[package.scala 94:16:@10538.4]
  assign RetimeWrapper_3_clock = clock; // @[:@10544.4]
  assign RetimeWrapper_3_reset = reset; // @[:@10545.4]
  assign RetimeWrapper_3_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@10547.4]
  assign RetimeWrapper_3_io_in = _T_1057 & io_rPort_0_en_0; // @[package.scala 94:16:@10546.4]
  assign RetimeWrapper_4_clock = clock; // @[:@10552.4]
  assign RetimeWrapper_4_reset = reset; // @[:@10553.4]
  assign RetimeWrapper_4_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@10555.4]
  assign RetimeWrapper_4_io_in = _T_1181 & io_rPort_0_en_0; // @[package.scala 94:16:@10554.4]
  assign RetimeWrapper_5_clock = clock; // @[:@10560.4]
  assign RetimeWrapper_5_reset = reset; // @[:@10561.4]
  assign RetimeWrapper_5_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@10563.4]
  assign RetimeWrapper_5_io_in = _T_1305 & io_rPort_0_en_0; // @[package.scala 94:16:@10562.4]
  assign RetimeWrapper_6_clock = clock; // @[:@10568.4]
  assign RetimeWrapper_6_reset = reset; // @[:@10569.4]
  assign RetimeWrapper_6_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@10571.4]
  assign RetimeWrapper_6_io_in = _T_1429 & io_rPort_0_en_0; // @[package.scala 94:16:@10570.4]
  assign RetimeWrapper_7_clock = clock; // @[:@10576.4]
  assign RetimeWrapper_7_reset = reset; // @[:@10577.4]
  assign RetimeWrapper_7_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@10579.4]
  assign RetimeWrapper_7_io_in = _T_1553 & io_rPort_0_en_0; // @[package.scala 94:16:@10578.4]
  assign RetimeWrapper_8_clock = clock; // @[:@10616.4]
  assign RetimeWrapper_8_reset = reset; // @[:@10617.4]
  assign RetimeWrapper_8_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@10619.4]
  assign RetimeWrapper_8_io_in = _T_623 & io_rPort_1_en_0; // @[package.scala 94:16:@10618.4]
  assign RetimeWrapper_9_clock = clock; // @[:@10624.4]
  assign RetimeWrapper_9_reset = reset; // @[:@10625.4]
  assign RetimeWrapper_9_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@10627.4]
  assign RetimeWrapper_9_io_in = _T_747 & io_rPort_1_en_0; // @[package.scala 94:16:@10626.4]
  assign RetimeWrapper_10_clock = clock; // @[:@10632.4]
  assign RetimeWrapper_10_reset = reset; // @[:@10633.4]
  assign RetimeWrapper_10_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@10635.4]
  assign RetimeWrapper_10_io_in = _T_871 & io_rPort_1_en_0; // @[package.scala 94:16:@10634.4]
  assign RetimeWrapper_11_clock = clock; // @[:@10640.4]
  assign RetimeWrapper_11_reset = reset; // @[:@10641.4]
  assign RetimeWrapper_11_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@10643.4]
  assign RetimeWrapper_11_io_in = _T_995 & io_rPort_1_en_0; // @[package.scala 94:16:@10642.4]
  assign RetimeWrapper_12_clock = clock; // @[:@10648.4]
  assign RetimeWrapper_12_reset = reset; // @[:@10649.4]
  assign RetimeWrapper_12_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@10651.4]
  assign RetimeWrapper_12_io_in = _T_1119 & io_rPort_1_en_0; // @[package.scala 94:16:@10650.4]
  assign RetimeWrapper_13_clock = clock; // @[:@10656.4]
  assign RetimeWrapper_13_reset = reset; // @[:@10657.4]
  assign RetimeWrapper_13_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@10659.4]
  assign RetimeWrapper_13_io_in = _T_1243 & io_rPort_1_en_0; // @[package.scala 94:16:@10658.4]
  assign RetimeWrapper_14_clock = clock; // @[:@10664.4]
  assign RetimeWrapper_14_reset = reset; // @[:@10665.4]
  assign RetimeWrapper_14_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@10667.4]
  assign RetimeWrapper_14_io_in = _T_1367 & io_rPort_1_en_0; // @[package.scala 94:16:@10666.4]
  assign RetimeWrapper_15_clock = clock; // @[:@10672.4]
  assign RetimeWrapper_15_reset = reset; // @[:@10673.4]
  assign RetimeWrapper_15_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@10675.4]
  assign RetimeWrapper_15_io_in = _T_1491 & io_rPort_1_en_0; // @[package.scala 94:16:@10674.4]
  assign RetimeWrapper_16_clock = clock; // @[:@10712.4]
  assign RetimeWrapper_16_reset = reset; // @[:@10713.4]
  assign RetimeWrapper_16_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@10715.4]
  assign RetimeWrapper_16_io_in = _T_629 & io_rPort_2_en_0; // @[package.scala 94:16:@10714.4]
  assign RetimeWrapper_17_clock = clock; // @[:@10720.4]
  assign RetimeWrapper_17_reset = reset; // @[:@10721.4]
  assign RetimeWrapper_17_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@10723.4]
  assign RetimeWrapper_17_io_in = _T_753 & io_rPort_2_en_0; // @[package.scala 94:16:@10722.4]
  assign RetimeWrapper_18_clock = clock; // @[:@10728.4]
  assign RetimeWrapper_18_reset = reset; // @[:@10729.4]
  assign RetimeWrapper_18_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@10731.4]
  assign RetimeWrapper_18_io_in = _T_877 & io_rPort_2_en_0; // @[package.scala 94:16:@10730.4]
  assign RetimeWrapper_19_clock = clock; // @[:@10736.4]
  assign RetimeWrapper_19_reset = reset; // @[:@10737.4]
  assign RetimeWrapper_19_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@10739.4]
  assign RetimeWrapper_19_io_in = _T_1001 & io_rPort_2_en_0; // @[package.scala 94:16:@10738.4]
  assign RetimeWrapper_20_clock = clock; // @[:@10744.4]
  assign RetimeWrapper_20_reset = reset; // @[:@10745.4]
  assign RetimeWrapper_20_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@10747.4]
  assign RetimeWrapper_20_io_in = _T_1125 & io_rPort_2_en_0; // @[package.scala 94:16:@10746.4]
  assign RetimeWrapper_21_clock = clock; // @[:@10752.4]
  assign RetimeWrapper_21_reset = reset; // @[:@10753.4]
  assign RetimeWrapper_21_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@10755.4]
  assign RetimeWrapper_21_io_in = _T_1249 & io_rPort_2_en_0; // @[package.scala 94:16:@10754.4]
  assign RetimeWrapper_22_clock = clock; // @[:@10760.4]
  assign RetimeWrapper_22_reset = reset; // @[:@10761.4]
  assign RetimeWrapper_22_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@10763.4]
  assign RetimeWrapper_22_io_in = _T_1373 & io_rPort_2_en_0; // @[package.scala 94:16:@10762.4]
  assign RetimeWrapper_23_clock = clock; // @[:@10768.4]
  assign RetimeWrapper_23_reset = reset; // @[:@10769.4]
  assign RetimeWrapper_23_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@10771.4]
  assign RetimeWrapper_23_io_in = _T_1497 & io_rPort_2_en_0; // @[package.scala 94:16:@10770.4]
  assign RetimeWrapper_24_clock = clock; // @[:@10808.4]
  assign RetimeWrapper_24_reset = reset; // @[:@10809.4]
  assign RetimeWrapper_24_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@10811.4]
  assign RetimeWrapper_24_io_in = _T_635 & io_rPort_3_en_0; // @[package.scala 94:16:@10810.4]
  assign RetimeWrapper_25_clock = clock; // @[:@10816.4]
  assign RetimeWrapper_25_reset = reset; // @[:@10817.4]
  assign RetimeWrapper_25_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@10819.4]
  assign RetimeWrapper_25_io_in = _T_759 & io_rPort_3_en_0; // @[package.scala 94:16:@10818.4]
  assign RetimeWrapper_26_clock = clock; // @[:@10824.4]
  assign RetimeWrapper_26_reset = reset; // @[:@10825.4]
  assign RetimeWrapper_26_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@10827.4]
  assign RetimeWrapper_26_io_in = _T_883 & io_rPort_3_en_0; // @[package.scala 94:16:@10826.4]
  assign RetimeWrapper_27_clock = clock; // @[:@10832.4]
  assign RetimeWrapper_27_reset = reset; // @[:@10833.4]
  assign RetimeWrapper_27_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@10835.4]
  assign RetimeWrapper_27_io_in = _T_1007 & io_rPort_3_en_0; // @[package.scala 94:16:@10834.4]
  assign RetimeWrapper_28_clock = clock; // @[:@10840.4]
  assign RetimeWrapper_28_reset = reset; // @[:@10841.4]
  assign RetimeWrapper_28_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@10843.4]
  assign RetimeWrapper_28_io_in = _T_1131 & io_rPort_3_en_0; // @[package.scala 94:16:@10842.4]
  assign RetimeWrapper_29_clock = clock; // @[:@10848.4]
  assign RetimeWrapper_29_reset = reset; // @[:@10849.4]
  assign RetimeWrapper_29_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@10851.4]
  assign RetimeWrapper_29_io_in = _T_1255 & io_rPort_3_en_0; // @[package.scala 94:16:@10850.4]
  assign RetimeWrapper_30_clock = clock; // @[:@10856.4]
  assign RetimeWrapper_30_reset = reset; // @[:@10857.4]
  assign RetimeWrapper_30_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@10859.4]
  assign RetimeWrapper_30_io_in = _T_1379 & io_rPort_3_en_0; // @[package.scala 94:16:@10858.4]
  assign RetimeWrapper_31_clock = clock; // @[:@10864.4]
  assign RetimeWrapper_31_reset = reset; // @[:@10865.4]
  assign RetimeWrapper_31_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@10867.4]
  assign RetimeWrapper_31_io_in = _T_1503 & io_rPort_3_en_0; // @[package.scala 94:16:@10866.4]
  assign RetimeWrapper_32_clock = clock; // @[:@10904.4]
  assign RetimeWrapper_32_reset = reset; // @[:@10905.4]
  assign RetimeWrapper_32_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@10907.4]
  assign RetimeWrapper_32_io_in = _T_691 & io_rPort_4_en_0; // @[package.scala 94:16:@10906.4]
  assign RetimeWrapper_33_clock = clock; // @[:@10912.4]
  assign RetimeWrapper_33_reset = reset; // @[:@10913.4]
  assign RetimeWrapper_33_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@10915.4]
  assign RetimeWrapper_33_io_in = _T_815 & io_rPort_4_en_0; // @[package.scala 94:16:@10914.4]
  assign RetimeWrapper_34_clock = clock; // @[:@10920.4]
  assign RetimeWrapper_34_reset = reset; // @[:@10921.4]
  assign RetimeWrapper_34_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@10923.4]
  assign RetimeWrapper_34_io_in = _T_939 & io_rPort_4_en_0; // @[package.scala 94:16:@10922.4]
  assign RetimeWrapper_35_clock = clock; // @[:@10928.4]
  assign RetimeWrapper_35_reset = reset; // @[:@10929.4]
  assign RetimeWrapper_35_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@10931.4]
  assign RetimeWrapper_35_io_in = _T_1063 & io_rPort_4_en_0; // @[package.scala 94:16:@10930.4]
  assign RetimeWrapper_36_clock = clock; // @[:@10936.4]
  assign RetimeWrapper_36_reset = reset; // @[:@10937.4]
  assign RetimeWrapper_36_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@10939.4]
  assign RetimeWrapper_36_io_in = _T_1187 & io_rPort_4_en_0; // @[package.scala 94:16:@10938.4]
  assign RetimeWrapper_37_clock = clock; // @[:@10944.4]
  assign RetimeWrapper_37_reset = reset; // @[:@10945.4]
  assign RetimeWrapper_37_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@10947.4]
  assign RetimeWrapper_37_io_in = _T_1311 & io_rPort_4_en_0; // @[package.scala 94:16:@10946.4]
  assign RetimeWrapper_38_clock = clock; // @[:@10952.4]
  assign RetimeWrapper_38_reset = reset; // @[:@10953.4]
  assign RetimeWrapper_38_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@10955.4]
  assign RetimeWrapper_38_io_in = _T_1435 & io_rPort_4_en_0; // @[package.scala 94:16:@10954.4]
  assign RetimeWrapper_39_clock = clock; // @[:@10960.4]
  assign RetimeWrapper_39_reset = reset; // @[:@10961.4]
  assign RetimeWrapper_39_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@10963.4]
  assign RetimeWrapper_39_io_in = _T_1559 & io_rPort_4_en_0; // @[package.scala 94:16:@10962.4]
  assign RetimeWrapper_40_clock = clock; // @[:@11000.4]
  assign RetimeWrapper_40_reset = reset; // @[:@11001.4]
  assign RetimeWrapper_40_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@11003.4]
  assign RetimeWrapper_40_io_in = _T_697 & io_rPort_5_en_0; // @[package.scala 94:16:@11002.4]
  assign RetimeWrapper_41_clock = clock; // @[:@11008.4]
  assign RetimeWrapper_41_reset = reset; // @[:@11009.4]
  assign RetimeWrapper_41_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@11011.4]
  assign RetimeWrapper_41_io_in = _T_821 & io_rPort_5_en_0; // @[package.scala 94:16:@11010.4]
  assign RetimeWrapper_42_clock = clock; // @[:@11016.4]
  assign RetimeWrapper_42_reset = reset; // @[:@11017.4]
  assign RetimeWrapper_42_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@11019.4]
  assign RetimeWrapper_42_io_in = _T_945 & io_rPort_5_en_0; // @[package.scala 94:16:@11018.4]
  assign RetimeWrapper_43_clock = clock; // @[:@11024.4]
  assign RetimeWrapper_43_reset = reset; // @[:@11025.4]
  assign RetimeWrapper_43_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@11027.4]
  assign RetimeWrapper_43_io_in = _T_1069 & io_rPort_5_en_0; // @[package.scala 94:16:@11026.4]
  assign RetimeWrapper_44_clock = clock; // @[:@11032.4]
  assign RetimeWrapper_44_reset = reset; // @[:@11033.4]
  assign RetimeWrapper_44_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@11035.4]
  assign RetimeWrapper_44_io_in = _T_1193 & io_rPort_5_en_0; // @[package.scala 94:16:@11034.4]
  assign RetimeWrapper_45_clock = clock; // @[:@11040.4]
  assign RetimeWrapper_45_reset = reset; // @[:@11041.4]
  assign RetimeWrapper_45_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@11043.4]
  assign RetimeWrapper_45_io_in = _T_1317 & io_rPort_5_en_0; // @[package.scala 94:16:@11042.4]
  assign RetimeWrapper_46_clock = clock; // @[:@11048.4]
  assign RetimeWrapper_46_reset = reset; // @[:@11049.4]
  assign RetimeWrapper_46_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@11051.4]
  assign RetimeWrapper_46_io_in = _T_1441 & io_rPort_5_en_0; // @[package.scala 94:16:@11050.4]
  assign RetimeWrapper_47_clock = clock; // @[:@11056.4]
  assign RetimeWrapper_47_reset = reset; // @[:@11057.4]
  assign RetimeWrapper_47_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@11059.4]
  assign RetimeWrapper_47_io_in = _T_1565 & io_rPort_5_en_0; // @[package.scala 94:16:@11058.4]
  assign RetimeWrapper_48_clock = clock; // @[:@11096.4]
  assign RetimeWrapper_48_reset = reset; // @[:@11097.4]
  assign RetimeWrapper_48_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@11099.4]
  assign RetimeWrapper_48_io_in = _T_641 & io_rPort_6_en_0; // @[package.scala 94:16:@11098.4]
  assign RetimeWrapper_49_clock = clock; // @[:@11104.4]
  assign RetimeWrapper_49_reset = reset; // @[:@11105.4]
  assign RetimeWrapper_49_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@11107.4]
  assign RetimeWrapper_49_io_in = _T_765 & io_rPort_6_en_0; // @[package.scala 94:16:@11106.4]
  assign RetimeWrapper_50_clock = clock; // @[:@11112.4]
  assign RetimeWrapper_50_reset = reset; // @[:@11113.4]
  assign RetimeWrapper_50_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@11115.4]
  assign RetimeWrapper_50_io_in = _T_889 & io_rPort_6_en_0; // @[package.scala 94:16:@11114.4]
  assign RetimeWrapper_51_clock = clock; // @[:@11120.4]
  assign RetimeWrapper_51_reset = reset; // @[:@11121.4]
  assign RetimeWrapper_51_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@11123.4]
  assign RetimeWrapper_51_io_in = _T_1013 & io_rPort_6_en_0; // @[package.scala 94:16:@11122.4]
  assign RetimeWrapper_52_clock = clock; // @[:@11128.4]
  assign RetimeWrapper_52_reset = reset; // @[:@11129.4]
  assign RetimeWrapper_52_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@11131.4]
  assign RetimeWrapper_52_io_in = _T_1137 & io_rPort_6_en_0; // @[package.scala 94:16:@11130.4]
  assign RetimeWrapper_53_clock = clock; // @[:@11136.4]
  assign RetimeWrapper_53_reset = reset; // @[:@11137.4]
  assign RetimeWrapper_53_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@11139.4]
  assign RetimeWrapper_53_io_in = _T_1261 & io_rPort_6_en_0; // @[package.scala 94:16:@11138.4]
  assign RetimeWrapper_54_clock = clock; // @[:@11144.4]
  assign RetimeWrapper_54_reset = reset; // @[:@11145.4]
  assign RetimeWrapper_54_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@11147.4]
  assign RetimeWrapper_54_io_in = _T_1385 & io_rPort_6_en_0; // @[package.scala 94:16:@11146.4]
  assign RetimeWrapper_55_clock = clock; // @[:@11152.4]
  assign RetimeWrapper_55_reset = reset; // @[:@11153.4]
  assign RetimeWrapper_55_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@11155.4]
  assign RetimeWrapper_55_io_in = _T_1509 & io_rPort_6_en_0; // @[package.scala 94:16:@11154.4]
  assign RetimeWrapper_56_clock = clock; // @[:@11192.4]
  assign RetimeWrapper_56_reset = reset; // @[:@11193.4]
  assign RetimeWrapper_56_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@11195.4]
  assign RetimeWrapper_56_io_in = _T_703 & io_rPort_7_en_0; // @[package.scala 94:16:@11194.4]
  assign RetimeWrapper_57_clock = clock; // @[:@11200.4]
  assign RetimeWrapper_57_reset = reset; // @[:@11201.4]
  assign RetimeWrapper_57_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@11203.4]
  assign RetimeWrapper_57_io_in = _T_827 & io_rPort_7_en_0; // @[package.scala 94:16:@11202.4]
  assign RetimeWrapper_58_clock = clock; // @[:@11208.4]
  assign RetimeWrapper_58_reset = reset; // @[:@11209.4]
  assign RetimeWrapper_58_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@11211.4]
  assign RetimeWrapper_58_io_in = _T_951 & io_rPort_7_en_0; // @[package.scala 94:16:@11210.4]
  assign RetimeWrapper_59_clock = clock; // @[:@11216.4]
  assign RetimeWrapper_59_reset = reset; // @[:@11217.4]
  assign RetimeWrapper_59_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@11219.4]
  assign RetimeWrapper_59_io_in = _T_1075 & io_rPort_7_en_0; // @[package.scala 94:16:@11218.4]
  assign RetimeWrapper_60_clock = clock; // @[:@11224.4]
  assign RetimeWrapper_60_reset = reset; // @[:@11225.4]
  assign RetimeWrapper_60_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@11227.4]
  assign RetimeWrapper_60_io_in = _T_1199 & io_rPort_7_en_0; // @[package.scala 94:16:@11226.4]
  assign RetimeWrapper_61_clock = clock; // @[:@11232.4]
  assign RetimeWrapper_61_reset = reset; // @[:@11233.4]
  assign RetimeWrapper_61_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@11235.4]
  assign RetimeWrapper_61_io_in = _T_1323 & io_rPort_7_en_0; // @[package.scala 94:16:@11234.4]
  assign RetimeWrapper_62_clock = clock; // @[:@11240.4]
  assign RetimeWrapper_62_reset = reset; // @[:@11241.4]
  assign RetimeWrapper_62_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@11243.4]
  assign RetimeWrapper_62_io_in = _T_1447 & io_rPort_7_en_0; // @[package.scala 94:16:@11242.4]
  assign RetimeWrapper_63_clock = clock; // @[:@11248.4]
  assign RetimeWrapper_63_reset = reset; // @[:@11249.4]
  assign RetimeWrapper_63_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@11251.4]
  assign RetimeWrapper_63_io_in = _T_1571 & io_rPort_7_en_0; // @[package.scala 94:16:@11250.4]
  assign RetimeWrapper_64_clock = clock; // @[:@11288.4]
  assign RetimeWrapper_64_reset = reset; // @[:@11289.4]
  assign RetimeWrapper_64_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@11291.4]
  assign RetimeWrapper_64_io_in = _T_647 & io_rPort_8_en_0; // @[package.scala 94:16:@11290.4]
  assign RetimeWrapper_65_clock = clock; // @[:@11296.4]
  assign RetimeWrapper_65_reset = reset; // @[:@11297.4]
  assign RetimeWrapper_65_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@11299.4]
  assign RetimeWrapper_65_io_in = _T_771 & io_rPort_8_en_0; // @[package.scala 94:16:@11298.4]
  assign RetimeWrapper_66_clock = clock; // @[:@11304.4]
  assign RetimeWrapper_66_reset = reset; // @[:@11305.4]
  assign RetimeWrapper_66_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@11307.4]
  assign RetimeWrapper_66_io_in = _T_895 & io_rPort_8_en_0; // @[package.scala 94:16:@11306.4]
  assign RetimeWrapper_67_clock = clock; // @[:@11312.4]
  assign RetimeWrapper_67_reset = reset; // @[:@11313.4]
  assign RetimeWrapper_67_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@11315.4]
  assign RetimeWrapper_67_io_in = _T_1019 & io_rPort_8_en_0; // @[package.scala 94:16:@11314.4]
  assign RetimeWrapper_68_clock = clock; // @[:@11320.4]
  assign RetimeWrapper_68_reset = reset; // @[:@11321.4]
  assign RetimeWrapper_68_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@11323.4]
  assign RetimeWrapper_68_io_in = _T_1143 & io_rPort_8_en_0; // @[package.scala 94:16:@11322.4]
  assign RetimeWrapper_69_clock = clock; // @[:@11328.4]
  assign RetimeWrapper_69_reset = reset; // @[:@11329.4]
  assign RetimeWrapper_69_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@11331.4]
  assign RetimeWrapper_69_io_in = _T_1267 & io_rPort_8_en_0; // @[package.scala 94:16:@11330.4]
  assign RetimeWrapper_70_clock = clock; // @[:@11336.4]
  assign RetimeWrapper_70_reset = reset; // @[:@11337.4]
  assign RetimeWrapper_70_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@11339.4]
  assign RetimeWrapper_70_io_in = _T_1391 & io_rPort_8_en_0; // @[package.scala 94:16:@11338.4]
  assign RetimeWrapper_71_clock = clock; // @[:@11344.4]
  assign RetimeWrapper_71_reset = reset; // @[:@11345.4]
  assign RetimeWrapper_71_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@11347.4]
  assign RetimeWrapper_71_io_in = _T_1515 & io_rPort_8_en_0; // @[package.scala 94:16:@11346.4]
  assign RetimeWrapper_72_clock = clock; // @[:@11384.4]
  assign RetimeWrapper_72_reset = reset; // @[:@11385.4]
  assign RetimeWrapper_72_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@11387.4]
  assign RetimeWrapper_72_io_in = _T_709 & io_rPort_9_en_0; // @[package.scala 94:16:@11386.4]
  assign RetimeWrapper_73_clock = clock; // @[:@11392.4]
  assign RetimeWrapper_73_reset = reset; // @[:@11393.4]
  assign RetimeWrapper_73_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@11395.4]
  assign RetimeWrapper_73_io_in = _T_833 & io_rPort_9_en_0; // @[package.scala 94:16:@11394.4]
  assign RetimeWrapper_74_clock = clock; // @[:@11400.4]
  assign RetimeWrapper_74_reset = reset; // @[:@11401.4]
  assign RetimeWrapper_74_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@11403.4]
  assign RetimeWrapper_74_io_in = _T_957 & io_rPort_9_en_0; // @[package.scala 94:16:@11402.4]
  assign RetimeWrapper_75_clock = clock; // @[:@11408.4]
  assign RetimeWrapper_75_reset = reset; // @[:@11409.4]
  assign RetimeWrapper_75_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@11411.4]
  assign RetimeWrapper_75_io_in = _T_1081 & io_rPort_9_en_0; // @[package.scala 94:16:@11410.4]
  assign RetimeWrapper_76_clock = clock; // @[:@11416.4]
  assign RetimeWrapper_76_reset = reset; // @[:@11417.4]
  assign RetimeWrapper_76_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@11419.4]
  assign RetimeWrapper_76_io_in = _T_1205 & io_rPort_9_en_0; // @[package.scala 94:16:@11418.4]
  assign RetimeWrapper_77_clock = clock; // @[:@11424.4]
  assign RetimeWrapper_77_reset = reset; // @[:@11425.4]
  assign RetimeWrapper_77_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@11427.4]
  assign RetimeWrapper_77_io_in = _T_1329 & io_rPort_9_en_0; // @[package.scala 94:16:@11426.4]
  assign RetimeWrapper_78_clock = clock; // @[:@11432.4]
  assign RetimeWrapper_78_reset = reset; // @[:@11433.4]
  assign RetimeWrapper_78_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@11435.4]
  assign RetimeWrapper_78_io_in = _T_1453 & io_rPort_9_en_0; // @[package.scala 94:16:@11434.4]
  assign RetimeWrapper_79_clock = clock; // @[:@11440.4]
  assign RetimeWrapper_79_reset = reset; // @[:@11441.4]
  assign RetimeWrapper_79_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@11443.4]
  assign RetimeWrapper_79_io_in = _T_1577 & io_rPort_9_en_0; // @[package.scala 94:16:@11442.4]
  assign RetimeWrapper_80_clock = clock; // @[:@11480.4]
  assign RetimeWrapper_80_reset = reset; // @[:@11481.4]
  assign RetimeWrapper_80_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@11483.4]
  assign RetimeWrapper_80_io_in = _T_715 & io_rPort_10_en_0; // @[package.scala 94:16:@11482.4]
  assign RetimeWrapper_81_clock = clock; // @[:@11488.4]
  assign RetimeWrapper_81_reset = reset; // @[:@11489.4]
  assign RetimeWrapper_81_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@11491.4]
  assign RetimeWrapper_81_io_in = _T_839 & io_rPort_10_en_0; // @[package.scala 94:16:@11490.4]
  assign RetimeWrapper_82_clock = clock; // @[:@11496.4]
  assign RetimeWrapper_82_reset = reset; // @[:@11497.4]
  assign RetimeWrapper_82_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@11499.4]
  assign RetimeWrapper_82_io_in = _T_963 & io_rPort_10_en_0; // @[package.scala 94:16:@11498.4]
  assign RetimeWrapper_83_clock = clock; // @[:@11504.4]
  assign RetimeWrapper_83_reset = reset; // @[:@11505.4]
  assign RetimeWrapper_83_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@11507.4]
  assign RetimeWrapper_83_io_in = _T_1087 & io_rPort_10_en_0; // @[package.scala 94:16:@11506.4]
  assign RetimeWrapper_84_clock = clock; // @[:@11512.4]
  assign RetimeWrapper_84_reset = reset; // @[:@11513.4]
  assign RetimeWrapper_84_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@11515.4]
  assign RetimeWrapper_84_io_in = _T_1211 & io_rPort_10_en_0; // @[package.scala 94:16:@11514.4]
  assign RetimeWrapper_85_clock = clock; // @[:@11520.4]
  assign RetimeWrapper_85_reset = reset; // @[:@11521.4]
  assign RetimeWrapper_85_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@11523.4]
  assign RetimeWrapper_85_io_in = _T_1335 & io_rPort_10_en_0; // @[package.scala 94:16:@11522.4]
  assign RetimeWrapper_86_clock = clock; // @[:@11528.4]
  assign RetimeWrapper_86_reset = reset; // @[:@11529.4]
  assign RetimeWrapper_86_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@11531.4]
  assign RetimeWrapper_86_io_in = _T_1459 & io_rPort_10_en_0; // @[package.scala 94:16:@11530.4]
  assign RetimeWrapper_87_clock = clock; // @[:@11536.4]
  assign RetimeWrapper_87_reset = reset; // @[:@11537.4]
  assign RetimeWrapper_87_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@11539.4]
  assign RetimeWrapper_87_io_in = _T_1583 & io_rPort_10_en_0; // @[package.scala 94:16:@11538.4]
  assign RetimeWrapper_88_clock = clock; // @[:@11576.4]
  assign RetimeWrapper_88_reset = reset; // @[:@11577.4]
  assign RetimeWrapper_88_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@11579.4]
  assign RetimeWrapper_88_io_in = _T_653 & io_rPort_11_en_0; // @[package.scala 94:16:@11578.4]
  assign RetimeWrapper_89_clock = clock; // @[:@11584.4]
  assign RetimeWrapper_89_reset = reset; // @[:@11585.4]
  assign RetimeWrapper_89_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@11587.4]
  assign RetimeWrapper_89_io_in = _T_777 & io_rPort_11_en_0; // @[package.scala 94:16:@11586.4]
  assign RetimeWrapper_90_clock = clock; // @[:@11592.4]
  assign RetimeWrapper_90_reset = reset; // @[:@11593.4]
  assign RetimeWrapper_90_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@11595.4]
  assign RetimeWrapper_90_io_in = _T_901 & io_rPort_11_en_0; // @[package.scala 94:16:@11594.4]
  assign RetimeWrapper_91_clock = clock; // @[:@11600.4]
  assign RetimeWrapper_91_reset = reset; // @[:@11601.4]
  assign RetimeWrapper_91_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@11603.4]
  assign RetimeWrapper_91_io_in = _T_1025 & io_rPort_11_en_0; // @[package.scala 94:16:@11602.4]
  assign RetimeWrapper_92_clock = clock; // @[:@11608.4]
  assign RetimeWrapper_92_reset = reset; // @[:@11609.4]
  assign RetimeWrapper_92_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@11611.4]
  assign RetimeWrapper_92_io_in = _T_1149 & io_rPort_11_en_0; // @[package.scala 94:16:@11610.4]
  assign RetimeWrapper_93_clock = clock; // @[:@11616.4]
  assign RetimeWrapper_93_reset = reset; // @[:@11617.4]
  assign RetimeWrapper_93_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@11619.4]
  assign RetimeWrapper_93_io_in = _T_1273 & io_rPort_11_en_0; // @[package.scala 94:16:@11618.4]
  assign RetimeWrapper_94_clock = clock; // @[:@11624.4]
  assign RetimeWrapper_94_reset = reset; // @[:@11625.4]
  assign RetimeWrapper_94_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@11627.4]
  assign RetimeWrapper_94_io_in = _T_1397 & io_rPort_11_en_0; // @[package.scala 94:16:@11626.4]
  assign RetimeWrapper_95_clock = clock; // @[:@11632.4]
  assign RetimeWrapper_95_reset = reset; // @[:@11633.4]
  assign RetimeWrapper_95_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@11635.4]
  assign RetimeWrapper_95_io_in = _T_1521 & io_rPort_11_en_0; // @[package.scala 94:16:@11634.4]
endmodule
module StickySelects_16( // @[:@13167.2]
  input   clock, // @[:@13168.4]
  input   reset, // @[:@13169.4]
  input   io_ins_0, // @[:@13170.4]
  input   io_ins_1, // @[:@13170.4]
  output  io_outs_0, // @[:@13170.4]
  output  io_outs_1 // @[:@13170.4]
);
  reg  _T_19; // @[StickySelects.scala 21:22:@13172.4]
  reg [31:0] _RAND_0;
  wire  _T_21; // @[StickySelects.scala 24:52:@13173.4]
  wire  _T_22; // @[StickySelects.scala 24:21:@13174.4]
  reg  _T_25; // @[StickySelects.scala 21:22:@13176.4]
  reg [31:0] _RAND_1;
  wire  _T_27; // @[StickySelects.scala 24:52:@13177.4]
  wire  _T_28; // @[StickySelects.scala 24:21:@13178.4]
  assign _T_21 = io_ins_0 | _T_19; // @[StickySelects.scala 24:52:@13173.4]
  assign _T_22 = io_ins_1 ? 1'h0 : _T_21; // @[StickySelects.scala 24:21:@13174.4]
  assign _T_27 = io_ins_1 | _T_25; // @[StickySelects.scala 24:52:@13177.4]
  assign _T_28 = io_ins_0 ? 1'h0 : _T_27; // @[StickySelects.scala 24:21:@13178.4]
  assign io_outs_0 = io_ins_1 ? 1'h0 : _T_21; // @[StickySelects.scala 28:52:@13180.4]
  assign io_outs_1 = io_ins_0 ? 1'h0 : _T_27; // @[StickySelects.scala 28:52:@13181.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_25 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (io_ins_1) begin
        _T_19 <= 1'h0;
      end else begin
        _T_19 <= _T_21;
      end
    end
    if (reset) begin
      _T_25 <= 1'h0;
    end else begin
      if (io_ins_0) begin
        _T_25 <= 1'h0;
      end else begin
        _T_25 <= _T_27;
      end
    end
  end
endmodule
module StickySelects_17( // @[:@13183.2]
  input   clock, // @[:@13184.4]
  input   reset, // @[:@13185.4]
  input   io_ins_0, // @[:@13186.4]
  input   io_ins_1, // @[:@13186.4]
  input   io_ins_2, // @[:@13186.4]
  input   io_ins_3, // @[:@13186.4]
  output  io_outs_0, // @[:@13186.4]
  output  io_outs_1, // @[:@13186.4]
  output  io_outs_2, // @[:@13186.4]
  output  io_outs_3 // @[:@13186.4]
);
  reg  _T_19; // @[StickySelects.scala 21:22:@13188.4]
  reg [31:0] _RAND_0;
  wire  _T_20; // @[StickySelects.scala 22:54:@13189.4]
  wire  _T_21; // @[StickySelects.scala 22:54:@13190.4]
  wire  _T_23; // @[StickySelects.scala 24:52:@13191.4]
  wire  _T_24; // @[StickySelects.scala 24:21:@13192.4]
  reg  _T_27; // @[StickySelects.scala 21:22:@13194.4]
  reg [31:0] _RAND_1;
  wire  _T_28; // @[StickySelects.scala 22:54:@13195.4]
  wire  _T_29; // @[StickySelects.scala 22:54:@13196.4]
  wire  _T_31; // @[StickySelects.scala 24:52:@13197.4]
  wire  _T_32; // @[StickySelects.scala 24:21:@13198.4]
  reg  _T_35; // @[StickySelects.scala 21:22:@13200.4]
  reg [31:0] _RAND_2;
  wire  _T_36; // @[StickySelects.scala 22:54:@13201.4]
  wire  _T_37; // @[StickySelects.scala 22:54:@13202.4]
  wire  _T_39; // @[StickySelects.scala 24:52:@13203.4]
  wire  _T_40; // @[StickySelects.scala 24:21:@13204.4]
  reg  _T_43; // @[StickySelects.scala 21:22:@13206.4]
  reg [31:0] _RAND_3;
  wire  _T_45; // @[StickySelects.scala 22:54:@13208.4]
  wire  _T_47; // @[StickySelects.scala 24:52:@13209.4]
  wire  _T_48; // @[StickySelects.scala 24:21:@13210.4]
  assign _T_20 = io_ins_1 | io_ins_2; // @[StickySelects.scala 22:54:@13189.4]
  assign _T_21 = _T_20 | io_ins_3; // @[StickySelects.scala 22:54:@13190.4]
  assign _T_23 = io_ins_0 | _T_19; // @[StickySelects.scala 24:52:@13191.4]
  assign _T_24 = _T_21 ? 1'h0 : _T_23; // @[StickySelects.scala 24:21:@13192.4]
  assign _T_28 = io_ins_0 | io_ins_2; // @[StickySelects.scala 22:54:@13195.4]
  assign _T_29 = _T_28 | io_ins_3; // @[StickySelects.scala 22:54:@13196.4]
  assign _T_31 = io_ins_1 | _T_27; // @[StickySelects.scala 24:52:@13197.4]
  assign _T_32 = _T_29 ? 1'h0 : _T_31; // @[StickySelects.scala 24:21:@13198.4]
  assign _T_36 = io_ins_0 | io_ins_1; // @[StickySelects.scala 22:54:@13201.4]
  assign _T_37 = _T_36 | io_ins_3; // @[StickySelects.scala 22:54:@13202.4]
  assign _T_39 = io_ins_2 | _T_35; // @[StickySelects.scala 24:52:@13203.4]
  assign _T_40 = _T_37 ? 1'h0 : _T_39; // @[StickySelects.scala 24:21:@13204.4]
  assign _T_45 = _T_36 | io_ins_2; // @[StickySelects.scala 22:54:@13208.4]
  assign _T_47 = io_ins_3 | _T_43; // @[StickySelects.scala 24:52:@13209.4]
  assign _T_48 = _T_45 ? 1'h0 : _T_47; // @[StickySelects.scala 24:21:@13210.4]
  assign io_outs_0 = _T_21 ? 1'h0 : _T_23; // @[StickySelects.scala 28:52:@13212.4]
  assign io_outs_1 = _T_29 ? 1'h0 : _T_31; // @[StickySelects.scala 28:52:@13213.4]
  assign io_outs_2 = _T_37 ? 1'h0 : _T_39; // @[StickySelects.scala 28:52:@13214.4]
  assign io_outs_3 = _T_45 ? 1'h0 : _T_47; // @[StickySelects.scala 28:52:@13215.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_27 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_35 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_43 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (_T_21) begin
        _T_19 <= 1'h0;
      end else begin
        _T_19 <= _T_23;
      end
    end
    if (reset) begin
      _T_27 <= 1'h0;
    end else begin
      if (_T_29) begin
        _T_27 <= 1'h0;
      end else begin
        _T_27 <= _T_31;
      end
    end
    if (reset) begin
      _T_35 <= 1'h0;
    end else begin
      if (_T_37) begin
        _T_35 <= 1'h0;
      end else begin
        _T_35 <= _T_39;
      end
    end
    if (reset) begin
      _T_43 <= 1'h0;
    end else begin
      if (_T_45) begin
        _T_43 <= 1'h0;
      end else begin
        _T_43 <= _T_47;
      end
    end
  end
endmodule
module x289_lb2_0( // @[:@15103.2]
  input        clock, // @[:@15104.4]
  input        reset, // @[:@15105.4]
  input  [2:0] io_rPort_5_banks_1, // @[:@15106.4]
  input  [2:0] io_rPort_5_banks_0, // @[:@15106.4]
  input        io_rPort_5_ofs_0, // @[:@15106.4]
  input        io_rPort_5_en_0, // @[:@15106.4]
  input        io_rPort_5_backpressure, // @[:@15106.4]
  output [7:0] io_rPort_5_output_0, // @[:@15106.4]
  input  [2:0] io_rPort_4_banks_1, // @[:@15106.4]
  input  [2:0] io_rPort_4_banks_0, // @[:@15106.4]
  input        io_rPort_4_ofs_0, // @[:@15106.4]
  input        io_rPort_4_en_0, // @[:@15106.4]
  input        io_rPort_4_backpressure, // @[:@15106.4]
  output [7:0] io_rPort_4_output_0, // @[:@15106.4]
  input  [2:0] io_rPort_3_banks_1, // @[:@15106.4]
  input  [2:0] io_rPort_3_banks_0, // @[:@15106.4]
  input        io_rPort_3_ofs_0, // @[:@15106.4]
  input        io_rPort_3_en_0, // @[:@15106.4]
  input        io_rPort_3_backpressure, // @[:@15106.4]
  output [7:0] io_rPort_3_output_0, // @[:@15106.4]
  input  [2:0] io_rPort_2_banks_1, // @[:@15106.4]
  input  [2:0] io_rPort_2_banks_0, // @[:@15106.4]
  input        io_rPort_2_ofs_0, // @[:@15106.4]
  input        io_rPort_2_en_0, // @[:@15106.4]
  input        io_rPort_2_backpressure, // @[:@15106.4]
  output [7:0] io_rPort_2_output_0, // @[:@15106.4]
  input  [2:0] io_rPort_1_banks_1, // @[:@15106.4]
  input  [2:0] io_rPort_1_banks_0, // @[:@15106.4]
  input        io_rPort_1_ofs_0, // @[:@15106.4]
  input        io_rPort_1_en_0, // @[:@15106.4]
  input        io_rPort_1_backpressure, // @[:@15106.4]
  output [7:0] io_rPort_1_output_0, // @[:@15106.4]
  input  [2:0] io_rPort_0_banks_1, // @[:@15106.4]
  input  [2:0] io_rPort_0_banks_0, // @[:@15106.4]
  input        io_rPort_0_ofs_0, // @[:@15106.4]
  input        io_rPort_0_en_0, // @[:@15106.4]
  input        io_rPort_0_backpressure, // @[:@15106.4]
  output [7:0] io_rPort_0_output_0, // @[:@15106.4]
  input  [2:0] io_wPort_1_banks_1, // @[:@15106.4]
  input  [2:0] io_wPort_1_banks_0, // @[:@15106.4]
  input        io_wPort_1_ofs_0, // @[:@15106.4]
  input  [7:0] io_wPort_1_data_0, // @[:@15106.4]
  input        io_wPort_1_en_0, // @[:@15106.4]
  input  [2:0] io_wPort_0_banks_1, // @[:@15106.4]
  input  [2:0] io_wPort_0_banks_0, // @[:@15106.4]
  input        io_wPort_0_ofs_0, // @[:@15106.4]
  input  [7:0] io_wPort_0_data_0, // @[:@15106.4]
  input        io_wPort_0_en_0 // @[:@15106.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@15161.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@15161.4]
  wire  Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15161.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15161.4]
  wire  Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15161.4]
  wire [7:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@15161.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@15161.4]
  wire [7:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@15161.4]
  wire  Mem1D_1_clock; // @[MemPrimitives.scala 64:21:@15177.4]
  wire  Mem1D_1_reset; // @[MemPrimitives.scala 64:21:@15177.4]
  wire  Mem1D_1_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15177.4]
  wire  Mem1D_1_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15177.4]
  wire  Mem1D_1_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15177.4]
  wire [7:0] Mem1D_1_io_w_data_0; // @[MemPrimitives.scala 64:21:@15177.4]
  wire  Mem1D_1_io_w_en_0; // @[MemPrimitives.scala 64:21:@15177.4]
  wire [7:0] Mem1D_1_io_output; // @[MemPrimitives.scala 64:21:@15177.4]
  wire  Mem1D_2_clock; // @[MemPrimitives.scala 64:21:@15193.4]
  wire  Mem1D_2_reset; // @[MemPrimitives.scala 64:21:@15193.4]
  wire  Mem1D_2_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15193.4]
  wire  Mem1D_2_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15193.4]
  wire  Mem1D_2_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15193.4]
  wire [7:0] Mem1D_2_io_w_data_0; // @[MemPrimitives.scala 64:21:@15193.4]
  wire  Mem1D_2_io_w_en_0; // @[MemPrimitives.scala 64:21:@15193.4]
  wire [7:0] Mem1D_2_io_output; // @[MemPrimitives.scala 64:21:@15193.4]
  wire  Mem1D_3_clock; // @[MemPrimitives.scala 64:21:@15209.4]
  wire  Mem1D_3_reset; // @[MemPrimitives.scala 64:21:@15209.4]
  wire  Mem1D_3_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15209.4]
  wire  Mem1D_3_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15209.4]
  wire  Mem1D_3_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15209.4]
  wire [7:0] Mem1D_3_io_w_data_0; // @[MemPrimitives.scala 64:21:@15209.4]
  wire  Mem1D_3_io_w_en_0; // @[MemPrimitives.scala 64:21:@15209.4]
  wire [7:0] Mem1D_3_io_output; // @[MemPrimitives.scala 64:21:@15209.4]
  wire  Mem1D_4_clock; // @[MemPrimitives.scala 64:21:@15225.4]
  wire  Mem1D_4_reset; // @[MemPrimitives.scala 64:21:@15225.4]
  wire  Mem1D_4_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15225.4]
  wire  Mem1D_4_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15225.4]
  wire  Mem1D_4_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15225.4]
  wire [7:0] Mem1D_4_io_w_data_0; // @[MemPrimitives.scala 64:21:@15225.4]
  wire  Mem1D_4_io_w_en_0; // @[MemPrimitives.scala 64:21:@15225.4]
  wire [7:0] Mem1D_4_io_output; // @[MemPrimitives.scala 64:21:@15225.4]
  wire  Mem1D_5_clock; // @[MemPrimitives.scala 64:21:@15241.4]
  wire  Mem1D_5_reset; // @[MemPrimitives.scala 64:21:@15241.4]
  wire  Mem1D_5_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15241.4]
  wire  Mem1D_5_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15241.4]
  wire  Mem1D_5_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15241.4]
  wire [7:0] Mem1D_5_io_w_data_0; // @[MemPrimitives.scala 64:21:@15241.4]
  wire  Mem1D_5_io_w_en_0; // @[MemPrimitives.scala 64:21:@15241.4]
  wire [7:0] Mem1D_5_io_output; // @[MemPrimitives.scala 64:21:@15241.4]
  wire  Mem1D_6_clock; // @[MemPrimitives.scala 64:21:@15257.4]
  wire  Mem1D_6_reset; // @[MemPrimitives.scala 64:21:@15257.4]
  wire  Mem1D_6_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15257.4]
  wire  Mem1D_6_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15257.4]
  wire  Mem1D_6_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15257.4]
  wire [7:0] Mem1D_6_io_w_data_0; // @[MemPrimitives.scala 64:21:@15257.4]
  wire  Mem1D_6_io_w_en_0; // @[MemPrimitives.scala 64:21:@15257.4]
  wire [7:0] Mem1D_6_io_output; // @[MemPrimitives.scala 64:21:@15257.4]
  wire  Mem1D_7_clock; // @[MemPrimitives.scala 64:21:@15273.4]
  wire  Mem1D_7_reset; // @[MemPrimitives.scala 64:21:@15273.4]
  wire  Mem1D_7_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15273.4]
  wire  Mem1D_7_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15273.4]
  wire  Mem1D_7_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15273.4]
  wire [7:0] Mem1D_7_io_w_data_0; // @[MemPrimitives.scala 64:21:@15273.4]
  wire  Mem1D_7_io_w_en_0; // @[MemPrimitives.scala 64:21:@15273.4]
  wire [7:0] Mem1D_7_io_output; // @[MemPrimitives.scala 64:21:@15273.4]
  wire  Mem1D_8_clock; // @[MemPrimitives.scala 64:21:@15289.4]
  wire  Mem1D_8_reset; // @[MemPrimitives.scala 64:21:@15289.4]
  wire  Mem1D_8_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15289.4]
  wire  Mem1D_8_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15289.4]
  wire  Mem1D_8_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15289.4]
  wire [7:0] Mem1D_8_io_w_data_0; // @[MemPrimitives.scala 64:21:@15289.4]
  wire  Mem1D_8_io_w_en_0; // @[MemPrimitives.scala 64:21:@15289.4]
  wire [7:0] Mem1D_8_io_output; // @[MemPrimitives.scala 64:21:@15289.4]
  wire  Mem1D_9_clock; // @[MemPrimitives.scala 64:21:@15305.4]
  wire  Mem1D_9_reset; // @[MemPrimitives.scala 64:21:@15305.4]
  wire  Mem1D_9_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15305.4]
  wire  Mem1D_9_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15305.4]
  wire  Mem1D_9_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15305.4]
  wire [7:0] Mem1D_9_io_w_data_0; // @[MemPrimitives.scala 64:21:@15305.4]
  wire  Mem1D_9_io_w_en_0; // @[MemPrimitives.scala 64:21:@15305.4]
  wire [7:0] Mem1D_9_io_output; // @[MemPrimitives.scala 64:21:@15305.4]
  wire  Mem1D_10_clock; // @[MemPrimitives.scala 64:21:@15321.4]
  wire  Mem1D_10_reset; // @[MemPrimitives.scala 64:21:@15321.4]
  wire  Mem1D_10_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15321.4]
  wire  Mem1D_10_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15321.4]
  wire  Mem1D_10_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15321.4]
  wire [7:0] Mem1D_10_io_w_data_0; // @[MemPrimitives.scala 64:21:@15321.4]
  wire  Mem1D_10_io_w_en_0; // @[MemPrimitives.scala 64:21:@15321.4]
  wire [7:0] Mem1D_10_io_output; // @[MemPrimitives.scala 64:21:@15321.4]
  wire  Mem1D_11_clock; // @[MemPrimitives.scala 64:21:@15337.4]
  wire  Mem1D_11_reset; // @[MemPrimitives.scala 64:21:@15337.4]
  wire  Mem1D_11_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15337.4]
  wire  Mem1D_11_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15337.4]
  wire  Mem1D_11_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15337.4]
  wire [7:0] Mem1D_11_io_w_data_0; // @[MemPrimitives.scala 64:21:@15337.4]
  wire  Mem1D_11_io_w_en_0; // @[MemPrimitives.scala 64:21:@15337.4]
  wire [7:0] Mem1D_11_io_output; // @[MemPrimitives.scala 64:21:@15337.4]
  wire  Mem1D_12_clock; // @[MemPrimitives.scala 64:21:@15353.4]
  wire  Mem1D_12_reset; // @[MemPrimitives.scala 64:21:@15353.4]
  wire  Mem1D_12_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15353.4]
  wire  Mem1D_12_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15353.4]
  wire  Mem1D_12_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15353.4]
  wire [7:0] Mem1D_12_io_w_data_0; // @[MemPrimitives.scala 64:21:@15353.4]
  wire  Mem1D_12_io_w_en_0; // @[MemPrimitives.scala 64:21:@15353.4]
  wire [7:0] Mem1D_12_io_output; // @[MemPrimitives.scala 64:21:@15353.4]
  wire  Mem1D_13_clock; // @[MemPrimitives.scala 64:21:@15369.4]
  wire  Mem1D_13_reset; // @[MemPrimitives.scala 64:21:@15369.4]
  wire  Mem1D_13_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15369.4]
  wire  Mem1D_13_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15369.4]
  wire  Mem1D_13_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15369.4]
  wire [7:0] Mem1D_13_io_w_data_0; // @[MemPrimitives.scala 64:21:@15369.4]
  wire  Mem1D_13_io_w_en_0; // @[MemPrimitives.scala 64:21:@15369.4]
  wire [7:0] Mem1D_13_io_output; // @[MemPrimitives.scala 64:21:@15369.4]
  wire  Mem1D_14_clock; // @[MemPrimitives.scala 64:21:@15385.4]
  wire  Mem1D_14_reset; // @[MemPrimitives.scala 64:21:@15385.4]
  wire  Mem1D_14_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15385.4]
  wire  Mem1D_14_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15385.4]
  wire  Mem1D_14_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15385.4]
  wire [7:0] Mem1D_14_io_w_data_0; // @[MemPrimitives.scala 64:21:@15385.4]
  wire  Mem1D_14_io_w_en_0; // @[MemPrimitives.scala 64:21:@15385.4]
  wire [7:0] Mem1D_14_io_output; // @[MemPrimitives.scala 64:21:@15385.4]
  wire  Mem1D_15_clock; // @[MemPrimitives.scala 64:21:@15401.4]
  wire  Mem1D_15_reset; // @[MemPrimitives.scala 64:21:@15401.4]
  wire  Mem1D_15_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15401.4]
  wire  Mem1D_15_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15401.4]
  wire  Mem1D_15_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15401.4]
  wire [7:0] Mem1D_15_io_w_data_0; // @[MemPrimitives.scala 64:21:@15401.4]
  wire  Mem1D_15_io_w_en_0; // @[MemPrimitives.scala 64:21:@15401.4]
  wire [7:0] Mem1D_15_io_output; // @[MemPrimitives.scala 64:21:@15401.4]
  wire  StickySelects_clock; // @[MemPrimitives.scala 121:29:@15617.4]
  wire  StickySelects_reset; // @[MemPrimitives.scala 121:29:@15617.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 121:29:@15617.4]
  wire  StickySelects_io_ins_1; // @[MemPrimitives.scala 121:29:@15617.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 121:29:@15617.4]
  wire  StickySelects_io_outs_1; // @[MemPrimitives.scala 121:29:@15617.4]
  wire  StickySelects_1_clock; // @[MemPrimitives.scala 121:29:@15651.4]
  wire  StickySelects_1_reset; // @[MemPrimitives.scala 121:29:@15651.4]
  wire  StickySelects_1_io_ins_0; // @[MemPrimitives.scala 121:29:@15651.4]
  wire  StickySelects_1_io_ins_1; // @[MemPrimitives.scala 121:29:@15651.4]
  wire  StickySelects_1_io_ins_2; // @[MemPrimitives.scala 121:29:@15651.4]
  wire  StickySelects_1_io_ins_3; // @[MemPrimitives.scala 121:29:@15651.4]
  wire  StickySelects_1_io_outs_0; // @[MemPrimitives.scala 121:29:@15651.4]
  wire  StickySelects_1_io_outs_1; // @[MemPrimitives.scala 121:29:@15651.4]
  wire  StickySelects_1_io_outs_2; // @[MemPrimitives.scala 121:29:@15651.4]
  wire  StickySelects_1_io_outs_3; // @[MemPrimitives.scala 121:29:@15651.4]
  wire  StickySelects_2_clock; // @[MemPrimitives.scala 121:29:@15687.4]
  wire  StickySelects_2_reset; // @[MemPrimitives.scala 121:29:@15687.4]
  wire  StickySelects_2_io_ins_0; // @[MemPrimitives.scala 121:29:@15687.4]
  wire  StickySelects_2_io_ins_1; // @[MemPrimitives.scala 121:29:@15687.4]
  wire  StickySelects_2_io_outs_0; // @[MemPrimitives.scala 121:29:@15687.4]
  wire  StickySelects_2_io_outs_1; // @[MemPrimitives.scala 121:29:@15687.4]
  wire  StickySelects_3_clock; // @[MemPrimitives.scala 121:29:@15721.4]
  wire  StickySelects_3_reset; // @[MemPrimitives.scala 121:29:@15721.4]
  wire  StickySelects_3_io_ins_0; // @[MemPrimitives.scala 121:29:@15721.4]
  wire  StickySelects_3_io_ins_1; // @[MemPrimitives.scala 121:29:@15721.4]
  wire  StickySelects_3_io_ins_2; // @[MemPrimitives.scala 121:29:@15721.4]
  wire  StickySelects_3_io_ins_3; // @[MemPrimitives.scala 121:29:@15721.4]
  wire  StickySelects_3_io_outs_0; // @[MemPrimitives.scala 121:29:@15721.4]
  wire  StickySelects_3_io_outs_1; // @[MemPrimitives.scala 121:29:@15721.4]
  wire  StickySelects_3_io_outs_2; // @[MemPrimitives.scala 121:29:@15721.4]
  wire  StickySelects_3_io_outs_3; // @[MemPrimitives.scala 121:29:@15721.4]
  wire  StickySelects_4_clock; // @[MemPrimitives.scala 121:29:@15757.4]
  wire  StickySelects_4_reset; // @[MemPrimitives.scala 121:29:@15757.4]
  wire  StickySelects_4_io_ins_0; // @[MemPrimitives.scala 121:29:@15757.4]
  wire  StickySelects_4_io_ins_1; // @[MemPrimitives.scala 121:29:@15757.4]
  wire  StickySelects_4_io_outs_0; // @[MemPrimitives.scala 121:29:@15757.4]
  wire  StickySelects_4_io_outs_1; // @[MemPrimitives.scala 121:29:@15757.4]
  wire  StickySelects_5_clock; // @[MemPrimitives.scala 121:29:@15791.4]
  wire  StickySelects_5_reset; // @[MemPrimitives.scala 121:29:@15791.4]
  wire  StickySelects_5_io_ins_0; // @[MemPrimitives.scala 121:29:@15791.4]
  wire  StickySelects_5_io_ins_1; // @[MemPrimitives.scala 121:29:@15791.4]
  wire  StickySelects_5_io_ins_2; // @[MemPrimitives.scala 121:29:@15791.4]
  wire  StickySelects_5_io_ins_3; // @[MemPrimitives.scala 121:29:@15791.4]
  wire  StickySelects_5_io_outs_0; // @[MemPrimitives.scala 121:29:@15791.4]
  wire  StickySelects_5_io_outs_1; // @[MemPrimitives.scala 121:29:@15791.4]
  wire  StickySelects_5_io_outs_2; // @[MemPrimitives.scala 121:29:@15791.4]
  wire  StickySelects_5_io_outs_3; // @[MemPrimitives.scala 121:29:@15791.4]
  wire  StickySelects_6_clock; // @[MemPrimitives.scala 121:29:@15827.4]
  wire  StickySelects_6_reset; // @[MemPrimitives.scala 121:29:@15827.4]
  wire  StickySelects_6_io_ins_0; // @[MemPrimitives.scala 121:29:@15827.4]
  wire  StickySelects_6_io_ins_1; // @[MemPrimitives.scala 121:29:@15827.4]
  wire  StickySelects_6_io_outs_0; // @[MemPrimitives.scala 121:29:@15827.4]
  wire  StickySelects_6_io_outs_1; // @[MemPrimitives.scala 121:29:@15827.4]
  wire  StickySelects_7_clock; // @[MemPrimitives.scala 121:29:@15861.4]
  wire  StickySelects_7_reset; // @[MemPrimitives.scala 121:29:@15861.4]
  wire  StickySelects_7_io_ins_0; // @[MemPrimitives.scala 121:29:@15861.4]
  wire  StickySelects_7_io_ins_1; // @[MemPrimitives.scala 121:29:@15861.4]
  wire  StickySelects_7_io_ins_2; // @[MemPrimitives.scala 121:29:@15861.4]
  wire  StickySelects_7_io_ins_3; // @[MemPrimitives.scala 121:29:@15861.4]
  wire  StickySelects_7_io_outs_0; // @[MemPrimitives.scala 121:29:@15861.4]
  wire  StickySelects_7_io_outs_1; // @[MemPrimitives.scala 121:29:@15861.4]
  wire  StickySelects_7_io_outs_2; // @[MemPrimitives.scala 121:29:@15861.4]
  wire  StickySelects_7_io_outs_3; // @[MemPrimitives.scala 121:29:@15861.4]
  wire  StickySelects_8_clock; // @[MemPrimitives.scala 121:29:@15897.4]
  wire  StickySelects_8_reset; // @[MemPrimitives.scala 121:29:@15897.4]
  wire  StickySelects_8_io_ins_0; // @[MemPrimitives.scala 121:29:@15897.4]
  wire  StickySelects_8_io_ins_1; // @[MemPrimitives.scala 121:29:@15897.4]
  wire  StickySelects_8_io_outs_0; // @[MemPrimitives.scala 121:29:@15897.4]
  wire  StickySelects_8_io_outs_1; // @[MemPrimitives.scala 121:29:@15897.4]
  wire  StickySelects_9_clock; // @[MemPrimitives.scala 121:29:@15931.4]
  wire  StickySelects_9_reset; // @[MemPrimitives.scala 121:29:@15931.4]
  wire  StickySelects_9_io_ins_0; // @[MemPrimitives.scala 121:29:@15931.4]
  wire  StickySelects_9_io_ins_1; // @[MemPrimitives.scala 121:29:@15931.4]
  wire  StickySelects_9_io_ins_2; // @[MemPrimitives.scala 121:29:@15931.4]
  wire  StickySelects_9_io_ins_3; // @[MemPrimitives.scala 121:29:@15931.4]
  wire  StickySelects_9_io_outs_0; // @[MemPrimitives.scala 121:29:@15931.4]
  wire  StickySelects_9_io_outs_1; // @[MemPrimitives.scala 121:29:@15931.4]
  wire  StickySelects_9_io_outs_2; // @[MemPrimitives.scala 121:29:@15931.4]
  wire  StickySelects_9_io_outs_3; // @[MemPrimitives.scala 121:29:@15931.4]
  wire  StickySelects_10_clock; // @[MemPrimitives.scala 121:29:@15967.4]
  wire  StickySelects_10_reset; // @[MemPrimitives.scala 121:29:@15967.4]
  wire  StickySelects_10_io_ins_0; // @[MemPrimitives.scala 121:29:@15967.4]
  wire  StickySelects_10_io_ins_1; // @[MemPrimitives.scala 121:29:@15967.4]
  wire  StickySelects_10_io_outs_0; // @[MemPrimitives.scala 121:29:@15967.4]
  wire  StickySelects_10_io_outs_1; // @[MemPrimitives.scala 121:29:@15967.4]
  wire  StickySelects_11_clock; // @[MemPrimitives.scala 121:29:@16001.4]
  wire  StickySelects_11_reset; // @[MemPrimitives.scala 121:29:@16001.4]
  wire  StickySelects_11_io_ins_0; // @[MemPrimitives.scala 121:29:@16001.4]
  wire  StickySelects_11_io_ins_1; // @[MemPrimitives.scala 121:29:@16001.4]
  wire  StickySelects_11_io_ins_2; // @[MemPrimitives.scala 121:29:@16001.4]
  wire  StickySelects_11_io_ins_3; // @[MemPrimitives.scala 121:29:@16001.4]
  wire  StickySelects_11_io_outs_0; // @[MemPrimitives.scala 121:29:@16001.4]
  wire  StickySelects_11_io_outs_1; // @[MemPrimitives.scala 121:29:@16001.4]
  wire  StickySelects_11_io_outs_2; // @[MemPrimitives.scala 121:29:@16001.4]
  wire  StickySelects_11_io_outs_3; // @[MemPrimitives.scala 121:29:@16001.4]
  wire  StickySelects_12_clock; // @[MemPrimitives.scala 121:29:@16037.4]
  wire  StickySelects_12_reset; // @[MemPrimitives.scala 121:29:@16037.4]
  wire  StickySelects_12_io_ins_0; // @[MemPrimitives.scala 121:29:@16037.4]
  wire  StickySelects_12_io_ins_1; // @[MemPrimitives.scala 121:29:@16037.4]
  wire  StickySelects_12_io_outs_0; // @[MemPrimitives.scala 121:29:@16037.4]
  wire  StickySelects_12_io_outs_1; // @[MemPrimitives.scala 121:29:@16037.4]
  wire  StickySelects_13_clock; // @[MemPrimitives.scala 121:29:@16071.4]
  wire  StickySelects_13_reset; // @[MemPrimitives.scala 121:29:@16071.4]
  wire  StickySelects_13_io_ins_0; // @[MemPrimitives.scala 121:29:@16071.4]
  wire  StickySelects_13_io_ins_1; // @[MemPrimitives.scala 121:29:@16071.4]
  wire  StickySelects_13_io_ins_2; // @[MemPrimitives.scala 121:29:@16071.4]
  wire  StickySelects_13_io_ins_3; // @[MemPrimitives.scala 121:29:@16071.4]
  wire  StickySelects_13_io_outs_0; // @[MemPrimitives.scala 121:29:@16071.4]
  wire  StickySelects_13_io_outs_1; // @[MemPrimitives.scala 121:29:@16071.4]
  wire  StickySelects_13_io_outs_2; // @[MemPrimitives.scala 121:29:@16071.4]
  wire  StickySelects_13_io_outs_3; // @[MemPrimitives.scala 121:29:@16071.4]
  wire  StickySelects_14_clock; // @[MemPrimitives.scala 121:29:@16107.4]
  wire  StickySelects_14_reset; // @[MemPrimitives.scala 121:29:@16107.4]
  wire  StickySelects_14_io_ins_0; // @[MemPrimitives.scala 121:29:@16107.4]
  wire  StickySelects_14_io_ins_1; // @[MemPrimitives.scala 121:29:@16107.4]
  wire  StickySelects_14_io_outs_0; // @[MemPrimitives.scala 121:29:@16107.4]
  wire  StickySelects_14_io_outs_1; // @[MemPrimitives.scala 121:29:@16107.4]
  wire  StickySelects_15_clock; // @[MemPrimitives.scala 121:29:@16141.4]
  wire  StickySelects_15_reset; // @[MemPrimitives.scala 121:29:@16141.4]
  wire  StickySelects_15_io_ins_0; // @[MemPrimitives.scala 121:29:@16141.4]
  wire  StickySelects_15_io_ins_1; // @[MemPrimitives.scala 121:29:@16141.4]
  wire  StickySelects_15_io_ins_2; // @[MemPrimitives.scala 121:29:@16141.4]
  wire  StickySelects_15_io_ins_3; // @[MemPrimitives.scala 121:29:@16141.4]
  wire  StickySelects_15_io_outs_0; // @[MemPrimitives.scala 121:29:@16141.4]
  wire  StickySelects_15_io_outs_1; // @[MemPrimitives.scala 121:29:@16141.4]
  wire  StickySelects_15_io_outs_2; // @[MemPrimitives.scala 121:29:@16141.4]
  wire  StickySelects_15_io_outs_3; // @[MemPrimitives.scala 121:29:@16141.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@16194.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@16194.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@16194.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@16194.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@16194.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@16202.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@16202.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@16202.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@16202.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@16202.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@16210.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@16210.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@16210.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@16210.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@16210.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@16218.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@16218.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@16218.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@16218.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@16218.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@16226.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@16226.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@16226.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@16226.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@16226.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@16234.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@16234.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@16234.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@16234.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@16234.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@16242.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@16242.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@16242.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@16242.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@16242.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@16250.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@16250.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@16250.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@16250.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@16250.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@16290.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@16290.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@16290.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@16290.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@16290.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@16298.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@16298.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@16298.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@16298.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@16298.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@16306.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@16306.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@16306.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@16306.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@16306.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@16314.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@16314.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@16314.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@16314.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@16314.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@16322.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@16322.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@16322.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@16322.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@16322.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@16330.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@16330.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@16330.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@16330.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@16330.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@16338.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@16338.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@16338.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@16338.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@16338.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@16346.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@16346.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@16346.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@16346.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@16346.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@16386.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@16386.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@16386.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@16386.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@16386.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@16394.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@16394.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@16394.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@16394.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@16394.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@16402.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@16402.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@16402.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@16402.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@16402.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@16410.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@16410.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@16410.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@16410.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@16410.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@16418.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@16418.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@16418.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@16418.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@16418.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@16426.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@16426.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@16426.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@16426.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@16426.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@16434.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@16434.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@16434.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@16434.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@16434.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@16442.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@16442.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@16442.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@16442.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@16442.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@16482.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@16482.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@16482.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@16482.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@16482.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@16490.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@16490.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@16490.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@16490.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@16490.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@16498.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@16498.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@16498.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@16498.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@16498.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@16506.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@16506.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@16506.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@16506.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@16506.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@16514.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@16514.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@16514.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@16514.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@16514.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@16522.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@16522.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@16522.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@16522.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@16522.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@16530.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@16530.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@16530.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@16530.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@16530.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@16538.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@16538.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@16538.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@16538.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@16538.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@16578.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@16578.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@16578.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@16578.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@16578.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@16586.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@16586.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@16586.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@16586.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@16586.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@16594.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@16594.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@16594.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@16594.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@16594.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@16602.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@16602.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@16602.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@16602.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@16602.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@16610.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@16610.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@16610.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@16610.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@16610.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@16618.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@16618.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@16618.4]
  wire  RetimeWrapper_37_io_in; // @[package.scala 93:22:@16618.4]
  wire  RetimeWrapper_37_io_out; // @[package.scala 93:22:@16618.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@16626.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@16626.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@16626.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@16626.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@16626.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@16634.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@16634.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@16634.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@16634.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@16634.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@16674.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@16674.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@16674.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@16674.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@16674.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@16682.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@16682.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@16682.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@16682.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@16682.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@16690.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@16690.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@16690.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@16690.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@16690.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@16698.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@16698.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@16698.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@16698.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@16698.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@16706.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@16706.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@16706.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@16706.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@16706.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@16714.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@16714.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@16714.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@16714.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@16714.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@16722.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@16722.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@16722.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@16722.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@16722.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@16730.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@16730.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@16730.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@16730.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@16730.4]
  wire  _T_264; // @[MemPrimitives.scala 82:210:@15417.4]
  wire  _T_266; // @[MemPrimitives.scala 82:210:@15418.4]
  wire  _T_267; // @[MemPrimitives.scala 82:228:@15419.4]
  wire  _T_268; // @[MemPrimitives.scala 83:102:@15420.4]
  wire [9:0] _T_270; // @[Cat.scala 30:58:@15422.4]
  wire  _T_275; // @[MemPrimitives.scala 82:210:@15429.4]
  wire  _T_277; // @[MemPrimitives.scala 82:210:@15430.4]
  wire  _T_278; // @[MemPrimitives.scala 82:228:@15431.4]
  wire  _T_279; // @[MemPrimitives.scala 83:102:@15432.4]
  wire [9:0] _T_281; // @[Cat.scala 30:58:@15434.4]
  wire  _T_288; // @[MemPrimitives.scala 82:210:@15442.4]
  wire  _T_289; // @[MemPrimitives.scala 82:228:@15443.4]
  wire  _T_290; // @[MemPrimitives.scala 83:102:@15444.4]
  wire [9:0] _T_292; // @[Cat.scala 30:58:@15446.4]
  wire  _T_299; // @[MemPrimitives.scala 82:210:@15454.4]
  wire  _T_300; // @[MemPrimitives.scala 82:228:@15455.4]
  wire  _T_301; // @[MemPrimitives.scala 83:102:@15456.4]
  wire [9:0] _T_303; // @[Cat.scala 30:58:@15458.4]
  wire  _T_308; // @[MemPrimitives.scala 82:210:@15465.4]
  wire  _T_311; // @[MemPrimitives.scala 82:228:@15467.4]
  wire  _T_312; // @[MemPrimitives.scala 83:102:@15468.4]
  wire [9:0] _T_314; // @[Cat.scala 30:58:@15470.4]
  wire  _T_319; // @[MemPrimitives.scala 82:210:@15477.4]
  wire  _T_322; // @[MemPrimitives.scala 82:228:@15479.4]
  wire  _T_323; // @[MemPrimitives.scala 83:102:@15480.4]
  wire [9:0] _T_325; // @[Cat.scala 30:58:@15482.4]
  wire  _T_333; // @[MemPrimitives.scala 82:228:@15491.4]
  wire  _T_334; // @[MemPrimitives.scala 83:102:@15492.4]
  wire [9:0] _T_336; // @[Cat.scala 30:58:@15494.4]
  wire  _T_344; // @[MemPrimitives.scala 82:228:@15503.4]
  wire  _T_345; // @[MemPrimitives.scala 83:102:@15504.4]
  wire [9:0] _T_347; // @[Cat.scala 30:58:@15506.4]
  wire  _T_352; // @[MemPrimitives.scala 82:210:@15513.4]
  wire  _T_355; // @[MemPrimitives.scala 82:228:@15515.4]
  wire  _T_356; // @[MemPrimitives.scala 83:102:@15516.4]
  wire [9:0] _T_358; // @[Cat.scala 30:58:@15518.4]
  wire  _T_363; // @[MemPrimitives.scala 82:210:@15525.4]
  wire  _T_366; // @[MemPrimitives.scala 82:228:@15527.4]
  wire  _T_367; // @[MemPrimitives.scala 83:102:@15528.4]
  wire [9:0] _T_369; // @[Cat.scala 30:58:@15530.4]
  wire  _T_377; // @[MemPrimitives.scala 82:228:@15539.4]
  wire  _T_378; // @[MemPrimitives.scala 83:102:@15540.4]
  wire [9:0] _T_380; // @[Cat.scala 30:58:@15542.4]
  wire  _T_388; // @[MemPrimitives.scala 82:228:@15551.4]
  wire  _T_389; // @[MemPrimitives.scala 83:102:@15552.4]
  wire [9:0] _T_391; // @[Cat.scala 30:58:@15554.4]
  wire  _T_396; // @[MemPrimitives.scala 82:210:@15561.4]
  wire  _T_399; // @[MemPrimitives.scala 82:228:@15563.4]
  wire  _T_400; // @[MemPrimitives.scala 83:102:@15564.4]
  wire [9:0] _T_402; // @[Cat.scala 30:58:@15566.4]
  wire  _T_407; // @[MemPrimitives.scala 82:210:@15573.4]
  wire  _T_410; // @[MemPrimitives.scala 82:228:@15575.4]
  wire  _T_411; // @[MemPrimitives.scala 83:102:@15576.4]
  wire [9:0] _T_413; // @[Cat.scala 30:58:@15578.4]
  wire  _T_421; // @[MemPrimitives.scala 82:228:@15587.4]
  wire  _T_422; // @[MemPrimitives.scala 83:102:@15588.4]
  wire [9:0] _T_424; // @[Cat.scala 30:58:@15590.4]
  wire  _T_432; // @[MemPrimitives.scala 82:228:@15599.4]
  wire  _T_433; // @[MemPrimitives.scala 83:102:@15600.4]
  wire [9:0] _T_435; // @[Cat.scala 30:58:@15602.4]
  wire  _T_440; // @[MemPrimitives.scala 110:210:@15609.4]
  wire  _T_442; // @[MemPrimitives.scala 110:210:@15610.4]
  wire  _T_443; // @[MemPrimitives.scala 110:228:@15611.4]
  wire  _T_446; // @[MemPrimitives.scala 110:210:@15613.4]
  wire  _T_448; // @[MemPrimitives.scala 110:210:@15614.4]
  wire  _T_449; // @[MemPrimitives.scala 110:228:@15615.4]
  wire  _T_451; // @[MemPrimitives.scala 123:41:@15622.4]
  wire  _T_452; // @[MemPrimitives.scala 123:41:@15623.4]
  wire [2:0] _T_454; // @[Cat.scala 30:58:@15625.4]
  wire [2:0] _T_456; // @[Cat.scala 30:58:@15627.4]
  wire [2:0] _T_457; // @[Mux.scala 31:69:@15628.4]
  wire  _T_462; // @[MemPrimitives.scala 110:210:@15635.4]
  wire  _T_464; // @[MemPrimitives.scala 110:210:@15636.4]
  wire  _T_465; // @[MemPrimitives.scala 110:228:@15637.4]
  wire  _T_468; // @[MemPrimitives.scala 110:210:@15639.4]
  wire  _T_470; // @[MemPrimitives.scala 110:210:@15640.4]
  wire  _T_471; // @[MemPrimitives.scala 110:228:@15641.4]
  wire  _T_474; // @[MemPrimitives.scala 110:210:@15643.4]
  wire  _T_476; // @[MemPrimitives.scala 110:210:@15644.4]
  wire  _T_477; // @[MemPrimitives.scala 110:228:@15645.4]
  wire  _T_480; // @[MemPrimitives.scala 110:210:@15647.4]
  wire  _T_482; // @[MemPrimitives.scala 110:210:@15648.4]
  wire  _T_483; // @[MemPrimitives.scala 110:228:@15649.4]
  wire  _T_485; // @[MemPrimitives.scala 123:41:@15658.4]
  wire  _T_486; // @[MemPrimitives.scala 123:41:@15659.4]
  wire  _T_487; // @[MemPrimitives.scala 123:41:@15660.4]
  wire  _T_488; // @[MemPrimitives.scala 123:41:@15661.4]
  wire [2:0] _T_490; // @[Cat.scala 30:58:@15663.4]
  wire [2:0] _T_492; // @[Cat.scala 30:58:@15665.4]
  wire [2:0] _T_494; // @[Cat.scala 30:58:@15667.4]
  wire [2:0] _T_496; // @[Cat.scala 30:58:@15669.4]
  wire [2:0] _T_497; // @[Mux.scala 31:69:@15670.4]
  wire [2:0] _T_498; // @[Mux.scala 31:69:@15671.4]
  wire [2:0] _T_499; // @[Mux.scala 31:69:@15672.4]
  wire  _T_506; // @[MemPrimitives.scala 110:210:@15680.4]
  wire  _T_507; // @[MemPrimitives.scala 110:228:@15681.4]
  wire  _T_512; // @[MemPrimitives.scala 110:210:@15684.4]
  wire  _T_513; // @[MemPrimitives.scala 110:228:@15685.4]
  wire  _T_515; // @[MemPrimitives.scala 123:41:@15692.4]
  wire  _T_516; // @[MemPrimitives.scala 123:41:@15693.4]
  wire [2:0] _T_518; // @[Cat.scala 30:58:@15695.4]
  wire [2:0] _T_520; // @[Cat.scala 30:58:@15697.4]
  wire [2:0] _T_521; // @[Mux.scala 31:69:@15698.4]
  wire  _T_528; // @[MemPrimitives.scala 110:210:@15706.4]
  wire  _T_529; // @[MemPrimitives.scala 110:228:@15707.4]
  wire  _T_534; // @[MemPrimitives.scala 110:210:@15710.4]
  wire  _T_535; // @[MemPrimitives.scala 110:228:@15711.4]
  wire  _T_540; // @[MemPrimitives.scala 110:210:@15714.4]
  wire  _T_541; // @[MemPrimitives.scala 110:228:@15715.4]
  wire  _T_546; // @[MemPrimitives.scala 110:210:@15718.4]
  wire  _T_547; // @[MemPrimitives.scala 110:228:@15719.4]
  wire  _T_549; // @[MemPrimitives.scala 123:41:@15728.4]
  wire  _T_550; // @[MemPrimitives.scala 123:41:@15729.4]
  wire  _T_551; // @[MemPrimitives.scala 123:41:@15730.4]
  wire  _T_552; // @[MemPrimitives.scala 123:41:@15731.4]
  wire [2:0] _T_554; // @[Cat.scala 30:58:@15733.4]
  wire [2:0] _T_556; // @[Cat.scala 30:58:@15735.4]
  wire [2:0] _T_558; // @[Cat.scala 30:58:@15737.4]
  wire [2:0] _T_560; // @[Cat.scala 30:58:@15739.4]
  wire [2:0] _T_561; // @[Mux.scala 31:69:@15740.4]
  wire [2:0] _T_562; // @[Mux.scala 31:69:@15741.4]
  wire [2:0] _T_563; // @[Mux.scala 31:69:@15742.4]
  wire  _T_568; // @[MemPrimitives.scala 110:210:@15749.4]
  wire  _T_571; // @[MemPrimitives.scala 110:228:@15751.4]
  wire  _T_574; // @[MemPrimitives.scala 110:210:@15753.4]
  wire  _T_577; // @[MemPrimitives.scala 110:228:@15755.4]
  wire  _T_579; // @[MemPrimitives.scala 123:41:@15762.4]
  wire  _T_580; // @[MemPrimitives.scala 123:41:@15763.4]
  wire [2:0] _T_582; // @[Cat.scala 30:58:@15765.4]
  wire [2:0] _T_584; // @[Cat.scala 30:58:@15767.4]
  wire [2:0] _T_585; // @[Mux.scala 31:69:@15768.4]
  wire  _T_590; // @[MemPrimitives.scala 110:210:@15775.4]
  wire  _T_593; // @[MemPrimitives.scala 110:228:@15777.4]
  wire  _T_596; // @[MemPrimitives.scala 110:210:@15779.4]
  wire  _T_599; // @[MemPrimitives.scala 110:228:@15781.4]
  wire  _T_602; // @[MemPrimitives.scala 110:210:@15783.4]
  wire  _T_605; // @[MemPrimitives.scala 110:228:@15785.4]
  wire  _T_608; // @[MemPrimitives.scala 110:210:@15787.4]
  wire  _T_611; // @[MemPrimitives.scala 110:228:@15789.4]
  wire  _T_613; // @[MemPrimitives.scala 123:41:@15798.4]
  wire  _T_614; // @[MemPrimitives.scala 123:41:@15799.4]
  wire  _T_615; // @[MemPrimitives.scala 123:41:@15800.4]
  wire  _T_616; // @[MemPrimitives.scala 123:41:@15801.4]
  wire [2:0] _T_618; // @[Cat.scala 30:58:@15803.4]
  wire [2:0] _T_620; // @[Cat.scala 30:58:@15805.4]
  wire [2:0] _T_622; // @[Cat.scala 30:58:@15807.4]
  wire [2:0] _T_624; // @[Cat.scala 30:58:@15809.4]
  wire [2:0] _T_625; // @[Mux.scala 31:69:@15810.4]
  wire [2:0] _T_626; // @[Mux.scala 31:69:@15811.4]
  wire [2:0] _T_627; // @[Mux.scala 31:69:@15812.4]
  wire  _T_635; // @[MemPrimitives.scala 110:228:@15821.4]
  wire  _T_641; // @[MemPrimitives.scala 110:228:@15825.4]
  wire  _T_643; // @[MemPrimitives.scala 123:41:@15832.4]
  wire  _T_644; // @[MemPrimitives.scala 123:41:@15833.4]
  wire [2:0] _T_646; // @[Cat.scala 30:58:@15835.4]
  wire [2:0] _T_648; // @[Cat.scala 30:58:@15837.4]
  wire [2:0] _T_649; // @[Mux.scala 31:69:@15838.4]
  wire  _T_657; // @[MemPrimitives.scala 110:228:@15847.4]
  wire  _T_663; // @[MemPrimitives.scala 110:228:@15851.4]
  wire  _T_669; // @[MemPrimitives.scala 110:228:@15855.4]
  wire  _T_675; // @[MemPrimitives.scala 110:228:@15859.4]
  wire  _T_677; // @[MemPrimitives.scala 123:41:@15868.4]
  wire  _T_678; // @[MemPrimitives.scala 123:41:@15869.4]
  wire  _T_679; // @[MemPrimitives.scala 123:41:@15870.4]
  wire  _T_680; // @[MemPrimitives.scala 123:41:@15871.4]
  wire [2:0] _T_682; // @[Cat.scala 30:58:@15873.4]
  wire [2:0] _T_684; // @[Cat.scala 30:58:@15875.4]
  wire [2:0] _T_686; // @[Cat.scala 30:58:@15877.4]
  wire [2:0] _T_688; // @[Cat.scala 30:58:@15879.4]
  wire [2:0] _T_689; // @[Mux.scala 31:69:@15880.4]
  wire [2:0] _T_690; // @[Mux.scala 31:69:@15881.4]
  wire [2:0] _T_691; // @[Mux.scala 31:69:@15882.4]
  wire  _T_696; // @[MemPrimitives.scala 110:210:@15889.4]
  wire  _T_699; // @[MemPrimitives.scala 110:228:@15891.4]
  wire  _T_702; // @[MemPrimitives.scala 110:210:@15893.4]
  wire  _T_705; // @[MemPrimitives.scala 110:228:@15895.4]
  wire  _T_707; // @[MemPrimitives.scala 123:41:@15902.4]
  wire  _T_708; // @[MemPrimitives.scala 123:41:@15903.4]
  wire [2:0] _T_710; // @[Cat.scala 30:58:@15905.4]
  wire [2:0] _T_712; // @[Cat.scala 30:58:@15907.4]
  wire [2:0] _T_713; // @[Mux.scala 31:69:@15908.4]
  wire  _T_718; // @[MemPrimitives.scala 110:210:@15915.4]
  wire  _T_721; // @[MemPrimitives.scala 110:228:@15917.4]
  wire  _T_724; // @[MemPrimitives.scala 110:210:@15919.4]
  wire  _T_727; // @[MemPrimitives.scala 110:228:@15921.4]
  wire  _T_730; // @[MemPrimitives.scala 110:210:@15923.4]
  wire  _T_733; // @[MemPrimitives.scala 110:228:@15925.4]
  wire  _T_736; // @[MemPrimitives.scala 110:210:@15927.4]
  wire  _T_739; // @[MemPrimitives.scala 110:228:@15929.4]
  wire  _T_741; // @[MemPrimitives.scala 123:41:@15938.4]
  wire  _T_742; // @[MemPrimitives.scala 123:41:@15939.4]
  wire  _T_743; // @[MemPrimitives.scala 123:41:@15940.4]
  wire  _T_744; // @[MemPrimitives.scala 123:41:@15941.4]
  wire [2:0] _T_746; // @[Cat.scala 30:58:@15943.4]
  wire [2:0] _T_748; // @[Cat.scala 30:58:@15945.4]
  wire [2:0] _T_750; // @[Cat.scala 30:58:@15947.4]
  wire [2:0] _T_752; // @[Cat.scala 30:58:@15949.4]
  wire [2:0] _T_753; // @[Mux.scala 31:69:@15950.4]
  wire [2:0] _T_754; // @[Mux.scala 31:69:@15951.4]
  wire [2:0] _T_755; // @[Mux.scala 31:69:@15952.4]
  wire  _T_763; // @[MemPrimitives.scala 110:228:@15961.4]
  wire  _T_769; // @[MemPrimitives.scala 110:228:@15965.4]
  wire  _T_771; // @[MemPrimitives.scala 123:41:@15972.4]
  wire  _T_772; // @[MemPrimitives.scala 123:41:@15973.4]
  wire [2:0] _T_774; // @[Cat.scala 30:58:@15975.4]
  wire [2:0] _T_776; // @[Cat.scala 30:58:@15977.4]
  wire [2:0] _T_777; // @[Mux.scala 31:69:@15978.4]
  wire  _T_785; // @[MemPrimitives.scala 110:228:@15987.4]
  wire  _T_791; // @[MemPrimitives.scala 110:228:@15991.4]
  wire  _T_797; // @[MemPrimitives.scala 110:228:@15995.4]
  wire  _T_803; // @[MemPrimitives.scala 110:228:@15999.4]
  wire  _T_805; // @[MemPrimitives.scala 123:41:@16008.4]
  wire  _T_806; // @[MemPrimitives.scala 123:41:@16009.4]
  wire  _T_807; // @[MemPrimitives.scala 123:41:@16010.4]
  wire  _T_808; // @[MemPrimitives.scala 123:41:@16011.4]
  wire [2:0] _T_810; // @[Cat.scala 30:58:@16013.4]
  wire [2:0] _T_812; // @[Cat.scala 30:58:@16015.4]
  wire [2:0] _T_814; // @[Cat.scala 30:58:@16017.4]
  wire [2:0] _T_816; // @[Cat.scala 30:58:@16019.4]
  wire [2:0] _T_817; // @[Mux.scala 31:69:@16020.4]
  wire [2:0] _T_818; // @[Mux.scala 31:69:@16021.4]
  wire [2:0] _T_819; // @[Mux.scala 31:69:@16022.4]
  wire  _T_824; // @[MemPrimitives.scala 110:210:@16029.4]
  wire  _T_827; // @[MemPrimitives.scala 110:228:@16031.4]
  wire  _T_830; // @[MemPrimitives.scala 110:210:@16033.4]
  wire  _T_833; // @[MemPrimitives.scala 110:228:@16035.4]
  wire  _T_835; // @[MemPrimitives.scala 123:41:@16042.4]
  wire  _T_836; // @[MemPrimitives.scala 123:41:@16043.4]
  wire [2:0] _T_838; // @[Cat.scala 30:58:@16045.4]
  wire [2:0] _T_840; // @[Cat.scala 30:58:@16047.4]
  wire [2:0] _T_841; // @[Mux.scala 31:69:@16048.4]
  wire  _T_846; // @[MemPrimitives.scala 110:210:@16055.4]
  wire  _T_849; // @[MemPrimitives.scala 110:228:@16057.4]
  wire  _T_852; // @[MemPrimitives.scala 110:210:@16059.4]
  wire  _T_855; // @[MemPrimitives.scala 110:228:@16061.4]
  wire  _T_858; // @[MemPrimitives.scala 110:210:@16063.4]
  wire  _T_861; // @[MemPrimitives.scala 110:228:@16065.4]
  wire  _T_864; // @[MemPrimitives.scala 110:210:@16067.4]
  wire  _T_867; // @[MemPrimitives.scala 110:228:@16069.4]
  wire  _T_869; // @[MemPrimitives.scala 123:41:@16078.4]
  wire  _T_870; // @[MemPrimitives.scala 123:41:@16079.4]
  wire  _T_871; // @[MemPrimitives.scala 123:41:@16080.4]
  wire  _T_872; // @[MemPrimitives.scala 123:41:@16081.4]
  wire [2:0] _T_874; // @[Cat.scala 30:58:@16083.4]
  wire [2:0] _T_876; // @[Cat.scala 30:58:@16085.4]
  wire [2:0] _T_878; // @[Cat.scala 30:58:@16087.4]
  wire [2:0] _T_880; // @[Cat.scala 30:58:@16089.4]
  wire [2:0] _T_881; // @[Mux.scala 31:69:@16090.4]
  wire [2:0] _T_882; // @[Mux.scala 31:69:@16091.4]
  wire [2:0] _T_883; // @[Mux.scala 31:69:@16092.4]
  wire  _T_891; // @[MemPrimitives.scala 110:228:@16101.4]
  wire  _T_897; // @[MemPrimitives.scala 110:228:@16105.4]
  wire  _T_899; // @[MemPrimitives.scala 123:41:@16112.4]
  wire  _T_900; // @[MemPrimitives.scala 123:41:@16113.4]
  wire [2:0] _T_902; // @[Cat.scala 30:58:@16115.4]
  wire [2:0] _T_904; // @[Cat.scala 30:58:@16117.4]
  wire [2:0] _T_905; // @[Mux.scala 31:69:@16118.4]
  wire  _T_913; // @[MemPrimitives.scala 110:228:@16127.4]
  wire  _T_919; // @[MemPrimitives.scala 110:228:@16131.4]
  wire  _T_925; // @[MemPrimitives.scala 110:228:@16135.4]
  wire  _T_931; // @[MemPrimitives.scala 110:228:@16139.4]
  wire  _T_933; // @[MemPrimitives.scala 123:41:@16148.4]
  wire  _T_934; // @[MemPrimitives.scala 123:41:@16149.4]
  wire  _T_935; // @[MemPrimitives.scala 123:41:@16150.4]
  wire  _T_936; // @[MemPrimitives.scala 123:41:@16151.4]
  wire [2:0] _T_938; // @[Cat.scala 30:58:@16153.4]
  wire [2:0] _T_940; // @[Cat.scala 30:58:@16155.4]
  wire [2:0] _T_942; // @[Cat.scala 30:58:@16157.4]
  wire [2:0] _T_944; // @[Cat.scala 30:58:@16159.4]
  wire [2:0] _T_945; // @[Mux.scala 31:69:@16160.4]
  wire [2:0] _T_946; // @[Mux.scala 31:69:@16161.4]
  wire [2:0] _T_947; // @[Mux.scala 31:69:@16162.4]
  wire  _T_1011; // @[package.scala 96:25:@16247.4 package.scala 96:25:@16248.4]
  wire [7:0] _T_1015; // @[Mux.scala 31:69:@16257.4]
  wire  _T_1008; // @[package.scala 96:25:@16239.4 package.scala 96:25:@16240.4]
  wire [7:0] _T_1016; // @[Mux.scala 31:69:@16258.4]
  wire  _T_1005; // @[package.scala 96:25:@16231.4 package.scala 96:25:@16232.4]
  wire [7:0] _T_1017; // @[Mux.scala 31:69:@16259.4]
  wire  _T_1002; // @[package.scala 96:25:@16223.4 package.scala 96:25:@16224.4]
  wire [7:0] _T_1018; // @[Mux.scala 31:69:@16260.4]
  wire  _T_999; // @[package.scala 96:25:@16215.4 package.scala 96:25:@16216.4]
  wire [7:0] _T_1019; // @[Mux.scala 31:69:@16261.4]
  wire  _T_996; // @[package.scala 96:25:@16207.4 package.scala 96:25:@16208.4]
  wire [7:0] _T_1020; // @[Mux.scala 31:69:@16262.4]
  wire  _T_993; // @[package.scala 96:25:@16199.4 package.scala 96:25:@16200.4]
  wire  _T_1082; // @[package.scala 96:25:@16343.4 package.scala 96:25:@16344.4]
  wire [7:0] _T_1086; // @[Mux.scala 31:69:@16353.4]
  wire  _T_1079; // @[package.scala 96:25:@16335.4 package.scala 96:25:@16336.4]
  wire [7:0] _T_1087; // @[Mux.scala 31:69:@16354.4]
  wire  _T_1076; // @[package.scala 96:25:@16327.4 package.scala 96:25:@16328.4]
  wire [7:0] _T_1088; // @[Mux.scala 31:69:@16355.4]
  wire  _T_1073; // @[package.scala 96:25:@16319.4 package.scala 96:25:@16320.4]
  wire [7:0] _T_1089; // @[Mux.scala 31:69:@16356.4]
  wire  _T_1070; // @[package.scala 96:25:@16311.4 package.scala 96:25:@16312.4]
  wire [7:0] _T_1090; // @[Mux.scala 31:69:@16357.4]
  wire  _T_1067; // @[package.scala 96:25:@16303.4 package.scala 96:25:@16304.4]
  wire [7:0] _T_1091; // @[Mux.scala 31:69:@16358.4]
  wire  _T_1064; // @[package.scala 96:25:@16295.4 package.scala 96:25:@16296.4]
  wire  _T_1153; // @[package.scala 96:25:@16439.4 package.scala 96:25:@16440.4]
  wire [7:0] _T_1157; // @[Mux.scala 31:69:@16449.4]
  wire  _T_1150; // @[package.scala 96:25:@16431.4 package.scala 96:25:@16432.4]
  wire [7:0] _T_1158; // @[Mux.scala 31:69:@16450.4]
  wire  _T_1147; // @[package.scala 96:25:@16423.4 package.scala 96:25:@16424.4]
  wire [7:0] _T_1159; // @[Mux.scala 31:69:@16451.4]
  wire  _T_1144; // @[package.scala 96:25:@16415.4 package.scala 96:25:@16416.4]
  wire [7:0] _T_1160; // @[Mux.scala 31:69:@16452.4]
  wire  _T_1141; // @[package.scala 96:25:@16407.4 package.scala 96:25:@16408.4]
  wire [7:0] _T_1161; // @[Mux.scala 31:69:@16453.4]
  wire  _T_1138; // @[package.scala 96:25:@16399.4 package.scala 96:25:@16400.4]
  wire [7:0] _T_1162; // @[Mux.scala 31:69:@16454.4]
  wire  _T_1135; // @[package.scala 96:25:@16391.4 package.scala 96:25:@16392.4]
  wire  _T_1224; // @[package.scala 96:25:@16535.4 package.scala 96:25:@16536.4]
  wire [7:0] _T_1228; // @[Mux.scala 31:69:@16545.4]
  wire  _T_1221; // @[package.scala 96:25:@16527.4 package.scala 96:25:@16528.4]
  wire [7:0] _T_1229; // @[Mux.scala 31:69:@16546.4]
  wire  _T_1218; // @[package.scala 96:25:@16519.4 package.scala 96:25:@16520.4]
  wire [7:0] _T_1230; // @[Mux.scala 31:69:@16547.4]
  wire  _T_1215; // @[package.scala 96:25:@16511.4 package.scala 96:25:@16512.4]
  wire [7:0] _T_1231; // @[Mux.scala 31:69:@16548.4]
  wire  _T_1212; // @[package.scala 96:25:@16503.4 package.scala 96:25:@16504.4]
  wire [7:0] _T_1232; // @[Mux.scala 31:69:@16549.4]
  wire  _T_1209; // @[package.scala 96:25:@16495.4 package.scala 96:25:@16496.4]
  wire [7:0] _T_1233; // @[Mux.scala 31:69:@16550.4]
  wire  _T_1206; // @[package.scala 96:25:@16487.4 package.scala 96:25:@16488.4]
  wire  _T_1295; // @[package.scala 96:25:@16631.4 package.scala 96:25:@16632.4]
  wire [7:0] _T_1299; // @[Mux.scala 31:69:@16641.4]
  wire  _T_1292; // @[package.scala 96:25:@16623.4 package.scala 96:25:@16624.4]
  wire [7:0] _T_1300; // @[Mux.scala 31:69:@16642.4]
  wire  _T_1289; // @[package.scala 96:25:@16615.4 package.scala 96:25:@16616.4]
  wire [7:0] _T_1301; // @[Mux.scala 31:69:@16643.4]
  wire  _T_1286; // @[package.scala 96:25:@16607.4 package.scala 96:25:@16608.4]
  wire [7:0] _T_1302; // @[Mux.scala 31:69:@16644.4]
  wire  _T_1283; // @[package.scala 96:25:@16599.4 package.scala 96:25:@16600.4]
  wire [7:0] _T_1303; // @[Mux.scala 31:69:@16645.4]
  wire  _T_1280; // @[package.scala 96:25:@16591.4 package.scala 96:25:@16592.4]
  wire [7:0] _T_1304; // @[Mux.scala 31:69:@16646.4]
  wire  _T_1277; // @[package.scala 96:25:@16583.4 package.scala 96:25:@16584.4]
  wire  _T_1366; // @[package.scala 96:25:@16727.4 package.scala 96:25:@16728.4]
  wire [7:0] _T_1370; // @[Mux.scala 31:69:@16737.4]
  wire  _T_1363; // @[package.scala 96:25:@16719.4 package.scala 96:25:@16720.4]
  wire [7:0] _T_1371; // @[Mux.scala 31:69:@16738.4]
  wire  _T_1360; // @[package.scala 96:25:@16711.4 package.scala 96:25:@16712.4]
  wire [7:0] _T_1372; // @[Mux.scala 31:69:@16739.4]
  wire  _T_1357; // @[package.scala 96:25:@16703.4 package.scala 96:25:@16704.4]
  wire [7:0] _T_1373; // @[Mux.scala 31:69:@16740.4]
  wire  _T_1354; // @[package.scala 96:25:@16695.4 package.scala 96:25:@16696.4]
  wire [7:0] _T_1374; // @[Mux.scala 31:69:@16741.4]
  wire  _T_1351; // @[package.scala 96:25:@16687.4 package.scala 96:25:@16688.4]
  wire [7:0] _T_1375; // @[Mux.scala 31:69:@16742.4]
  wire  _T_1348; // @[package.scala 96:25:@16679.4 package.scala 96:25:@16680.4]
  Mem1D_4 Mem1D ( // @[MemPrimitives.scala 64:21:@15161.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  Mem1D_4 Mem1D_1 ( // @[MemPrimitives.scala 64:21:@15177.4]
    .clock(Mem1D_1_clock),
    .reset(Mem1D_1_reset),
    .io_r_ofs_0(Mem1D_1_io_r_ofs_0),
    .io_r_backpressure(Mem1D_1_io_r_backpressure),
    .io_w_ofs_0(Mem1D_1_io_w_ofs_0),
    .io_w_data_0(Mem1D_1_io_w_data_0),
    .io_w_en_0(Mem1D_1_io_w_en_0),
    .io_output(Mem1D_1_io_output)
  );
  Mem1D_4 Mem1D_2 ( // @[MemPrimitives.scala 64:21:@15193.4]
    .clock(Mem1D_2_clock),
    .reset(Mem1D_2_reset),
    .io_r_ofs_0(Mem1D_2_io_r_ofs_0),
    .io_r_backpressure(Mem1D_2_io_r_backpressure),
    .io_w_ofs_0(Mem1D_2_io_w_ofs_0),
    .io_w_data_0(Mem1D_2_io_w_data_0),
    .io_w_en_0(Mem1D_2_io_w_en_0),
    .io_output(Mem1D_2_io_output)
  );
  Mem1D_4 Mem1D_3 ( // @[MemPrimitives.scala 64:21:@15209.4]
    .clock(Mem1D_3_clock),
    .reset(Mem1D_3_reset),
    .io_r_ofs_0(Mem1D_3_io_r_ofs_0),
    .io_r_backpressure(Mem1D_3_io_r_backpressure),
    .io_w_ofs_0(Mem1D_3_io_w_ofs_0),
    .io_w_data_0(Mem1D_3_io_w_data_0),
    .io_w_en_0(Mem1D_3_io_w_en_0),
    .io_output(Mem1D_3_io_output)
  );
  Mem1D_4 Mem1D_4 ( // @[MemPrimitives.scala 64:21:@15225.4]
    .clock(Mem1D_4_clock),
    .reset(Mem1D_4_reset),
    .io_r_ofs_0(Mem1D_4_io_r_ofs_0),
    .io_r_backpressure(Mem1D_4_io_r_backpressure),
    .io_w_ofs_0(Mem1D_4_io_w_ofs_0),
    .io_w_data_0(Mem1D_4_io_w_data_0),
    .io_w_en_0(Mem1D_4_io_w_en_0),
    .io_output(Mem1D_4_io_output)
  );
  Mem1D_4 Mem1D_5 ( // @[MemPrimitives.scala 64:21:@15241.4]
    .clock(Mem1D_5_clock),
    .reset(Mem1D_5_reset),
    .io_r_ofs_0(Mem1D_5_io_r_ofs_0),
    .io_r_backpressure(Mem1D_5_io_r_backpressure),
    .io_w_ofs_0(Mem1D_5_io_w_ofs_0),
    .io_w_data_0(Mem1D_5_io_w_data_0),
    .io_w_en_0(Mem1D_5_io_w_en_0),
    .io_output(Mem1D_5_io_output)
  );
  Mem1D_4 Mem1D_6 ( // @[MemPrimitives.scala 64:21:@15257.4]
    .clock(Mem1D_6_clock),
    .reset(Mem1D_6_reset),
    .io_r_ofs_0(Mem1D_6_io_r_ofs_0),
    .io_r_backpressure(Mem1D_6_io_r_backpressure),
    .io_w_ofs_0(Mem1D_6_io_w_ofs_0),
    .io_w_data_0(Mem1D_6_io_w_data_0),
    .io_w_en_0(Mem1D_6_io_w_en_0),
    .io_output(Mem1D_6_io_output)
  );
  Mem1D_4 Mem1D_7 ( // @[MemPrimitives.scala 64:21:@15273.4]
    .clock(Mem1D_7_clock),
    .reset(Mem1D_7_reset),
    .io_r_ofs_0(Mem1D_7_io_r_ofs_0),
    .io_r_backpressure(Mem1D_7_io_r_backpressure),
    .io_w_ofs_0(Mem1D_7_io_w_ofs_0),
    .io_w_data_0(Mem1D_7_io_w_data_0),
    .io_w_en_0(Mem1D_7_io_w_en_0),
    .io_output(Mem1D_7_io_output)
  );
  Mem1D_4 Mem1D_8 ( // @[MemPrimitives.scala 64:21:@15289.4]
    .clock(Mem1D_8_clock),
    .reset(Mem1D_8_reset),
    .io_r_ofs_0(Mem1D_8_io_r_ofs_0),
    .io_r_backpressure(Mem1D_8_io_r_backpressure),
    .io_w_ofs_0(Mem1D_8_io_w_ofs_0),
    .io_w_data_0(Mem1D_8_io_w_data_0),
    .io_w_en_0(Mem1D_8_io_w_en_0),
    .io_output(Mem1D_8_io_output)
  );
  Mem1D_4 Mem1D_9 ( // @[MemPrimitives.scala 64:21:@15305.4]
    .clock(Mem1D_9_clock),
    .reset(Mem1D_9_reset),
    .io_r_ofs_0(Mem1D_9_io_r_ofs_0),
    .io_r_backpressure(Mem1D_9_io_r_backpressure),
    .io_w_ofs_0(Mem1D_9_io_w_ofs_0),
    .io_w_data_0(Mem1D_9_io_w_data_0),
    .io_w_en_0(Mem1D_9_io_w_en_0),
    .io_output(Mem1D_9_io_output)
  );
  Mem1D_4 Mem1D_10 ( // @[MemPrimitives.scala 64:21:@15321.4]
    .clock(Mem1D_10_clock),
    .reset(Mem1D_10_reset),
    .io_r_ofs_0(Mem1D_10_io_r_ofs_0),
    .io_r_backpressure(Mem1D_10_io_r_backpressure),
    .io_w_ofs_0(Mem1D_10_io_w_ofs_0),
    .io_w_data_0(Mem1D_10_io_w_data_0),
    .io_w_en_0(Mem1D_10_io_w_en_0),
    .io_output(Mem1D_10_io_output)
  );
  Mem1D_4 Mem1D_11 ( // @[MemPrimitives.scala 64:21:@15337.4]
    .clock(Mem1D_11_clock),
    .reset(Mem1D_11_reset),
    .io_r_ofs_0(Mem1D_11_io_r_ofs_0),
    .io_r_backpressure(Mem1D_11_io_r_backpressure),
    .io_w_ofs_0(Mem1D_11_io_w_ofs_0),
    .io_w_data_0(Mem1D_11_io_w_data_0),
    .io_w_en_0(Mem1D_11_io_w_en_0),
    .io_output(Mem1D_11_io_output)
  );
  Mem1D_4 Mem1D_12 ( // @[MemPrimitives.scala 64:21:@15353.4]
    .clock(Mem1D_12_clock),
    .reset(Mem1D_12_reset),
    .io_r_ofs_0(Mem1D_12_io_r_ofs_0),
    .io_r_backpressure(Mem1D_12_io_r_backpressure),
    .io_w_ofs_0(Mem1D_12_io_w_ofs_0),
    .io_w_data_0(Mem1D_12_io_w_data_0),
    .io_w_en_0(Mem1D_12_io_w_en_0),
    .io_output(Mem1D_12_io_output)
  );
  Mem1D_4 Mem1D_13 ( // @[MemPrimitives.scala 64:21:@15369.4]
    .clock(Mem1D_13_clock),
    .reset(Mem1D_13_reset),
    .io_r_ofs_0(Mem1D_13_io_r_ofs_0),
    .io_r_backpressure(Mem1D_13_io_r_backpressure),
    .io_w_ofs_0(Mem1D_13_io_w_ofs_0),
    .io_w_data_0(Mem1D_13_io_w_data_0),
    .io_w_en_0(Mem1D_13_io_w_en_0),
    .io_output(Mem1D_13_io_output)
  );
  Mem1D_4 Mem1D_14 ( // @[MemPrimitives.scala 64:21:@15385.4]
    .clock(Mem1D_14_clock),
    .reset(Mem1D_14_reset),
    .io_r_ofs_0(Mem1D_14_io_r_ofs_0),
    .io_r_backpressure(Mem1D_14_io_r_backpressure),
    .io_w_ofs_0(Mem1D_14_io_w_ofs_0),
    .io_w_data_0(Mem1D_14_io_w_data_0),
    .io_w_en_0(Mem1D_14_io_w_en_0),
    .io_output(Mem1D_14_io_output)
  );
  Mem1D_4 Mem1D_15 ( // @[MemPrimitives.scala 64:21:@15401.4]
    .clock(Mem1D_15_clock),
    .reset(Mem1D_15_reset),
    .io_r_ofs_0(Mem1D_15_io_r_ofs_0),
    .io_r_backpressure(Mem1D_15_io_r_backpressure),
    .io_w_ofs_0(Mem1D_15_io_w_ofs_0),
    .io_w_data_0(Mem1D_15_io_w_data_0),
    .io_w_en_0(Mem1D_15_io_w_en_0),
    .io_output(Mem1D_15_io_output)
  );
  StickySelects_16 StickySelects ( // @[MemPrimitives.scala 121:29:@15617.4]
    .clock(StickySelects_clock),
    .reset(StickySelects_reset),
    .io_ins_0(StickySelects_io_ins_0),
    .io_ins_1(StickySelects_io_ins_1),
    .io_outs_0(StickySelects_io_outs_0),
    .io_outs_1(StickySelects_io_outs_1)
  );
  StickySelects_17 StickySelects_1 ( // @[MemPrimitives.scala 121:29:@15651.4]
    .clock(StickySelects_1_clock),
    .reset(StickySelects_1_reset),
    .io_ins_0(StickySelects_1_io_ins_0),
    .io_ins_1(StickySelects_1_io_ins_1),
    .io_ins_2(StickySelects_1_io_ins_2),
    .io_ins_3(StickySelects_1_io_ins_3),
    .io_outs_0(StickySelects_1_io_outs_0),
    .io_outs_1(StickySelects_1_io_outs_1),
    .io_outs_2(StickySelects_1_io_outs_2),
    .io_outs_3(StickySelects_1_io_outs_3)
  );
  StickySelects_16 StickySelects_2 ( // @[MemPrimitives.scala 121:29:@15687.4]
    .clock(StickySelects_2_clock),
    .reset(StickySelects_2_reset),
    .io_ins_0(StickySelects_2_io_ins_0),
    .io_ins_1(StickySelects_2_io_ins_1),
    .io_outs_0(StickySelects_2_io_outs_0),
    .io_outs_1(StickySelects_2_io_outs_1)
  );
  StickySelects_17 StickySelects_3 ( // @[MemPrimitives.scala 121:29:@15721.4]
    .clock(StickySelects_3_clock),
    .reset(StickySelects_3_reset),
    .io_ins_0(StickySelects_3_io_ins_0),
    .io_ins_1(StickySelects_3_io_ins_1),
    .io_ins_2(StickySelects_3_io_ins_2),
    .io_ins_3(StickySelects_3_io_ins_3),
    .io_outs_0(StickySelects_3_io_outs_0),
    .io_outs_1(StickySelects_3_io_outs_1),
    .io_outs_2(StickySelects_3_io_outs_2),
    .io_outs_3(StickySelects_3_io_outs_3)
  );
  StickySelects_16 StickySelects_4 ( // @[MemPrimitives.scala 121:29:@15757.4]
    .clock(StickySelects_4_clock),
    .reset(StickySelects_4_reset),
    .io_ins_0(StickySelects_4_io_ins_0),
    .io_ins_1(StickySelects_4_io_ins_1),
    .io_outs_0(StickySelects_4_io_outs_0),
    .io_outs_1(StickySelects_4_io_outs_1)
  );
  StickySelects_17 StickySelects_5 ( // @[MemPrimitives.scala 121:29:@15791.4]
    .clock(StickySelects_5_clock),
    .reset(StickySelects_5_reset),
    .io_ins_0(StickySelects_5_io_ins_0),
    .io_ins_1(StickySelects_5_io_ins_1),
    .io_ins_2(StickySelects_5_io_ins_2),
    .io_ins_3(StickySelects_5_io_ins_3),
    .io_outs_0(StickySelects_5_io_outs_0),
    .io_outs_1(StickySelects_5_io_outs_1),
    .io_outs_2(StickySelects_5_io_outs_2),
    .io_outs_3(StickySelects_5_io_outs_3)
  );
  StickySelects_16 StickySelects_6 ( // @[MemPrimitives.scala 121:29:@15827.4]
    .clock(StickySelects_6_clock),
    .reset(StickySelects_6_reset),
    .io_ins_0(StickySelects_6_io_ins_0),
    .io_ins_1(StickySelects_6_io_ins_1),
    .io_outs_0(StickySelects_6_io_outs_0),
    .io_outs_1(StickySelects_6_io_outs_1)
  );
  StickySelects_17 StickySelects_7 ( // @[MemPrimitives.scala 121:29:@15861.4]
    .clock(StickySelects_7_clock),
    .reset(StickySelects_7_reset),
    .io_ins_0(StickySelects_7_io_ins_0),
    .io_ins_1(StickySelects_7_io_ins_1),
    .io_ins_2(StickySelects_7_io_ins_2),
    .io_ins_3(StickySelects_7_io_ins_3),
    .io_outs_0(StickySelects_7_io_outs_0),
    .io_outs_1(StickySelects_7_io_outs_1),
    .io_outs_2(StickySelects_7_io_outs_2),
    .io_outs_3(StickySelects_7_io_outs_3)
  );
  StickySelects_16 StickySelects_8 ( // @[MemPrimitives.scala 121:29:@15897.4]
    .clock(StickySelects_8_clock),
    .reset(StickySelects_8_reset),
    .io_ins_0(StickySelects_8_io_ins_0),
    .io_ins_1(StickySelects_8_io_ins_1),
    .io_outs_0(StickySelects_8_io_outs_0),
    .io_outs_1(StickySelects_8_io_outs_1)
  );
  StickySelects_17 StickySelects_9 ( // @[MemPrimitives.scala 121:29:@15931.4]
    .clock(StickySelects_9_clock),
    .reset(StickySelects_9_reset),
    .io_ins_0(StickySelects_9_io_ins_0),
    .io_ins_1(StickySelects_9_io_ins_1),
    .io_ins_2(StickySelects_9_io_ins_2),
    .io_ins_3(StickySelects_9_io_ins_3),
    .io_outs_0(StickySelects_9_io_outs_0),
    .io_outs_1(StickySelects_9_io_outs_1),
    .io_outs_2(StickySelects_9_io_outs_2),
    .io_outs_3(StickySelects_9_io_outs_3)
  );
  StickySelects_16 StickySelects_10 ( // @[MemPrimitives.scala 121:29:@15967.4]
    .clock(StickySelects_10_clock),
    .reset(StickySelects_10_reset),
    .io_ins_0(StickySelects_10_io_ins_0),
    .io_ins_1(StickySelects_10_io_ins_1),
    .io_outs_0(StickySelects_10_io_outs_0),
    .io_outs_1(StickySelects_10_io_outs_1)
  );
  StickySelects_17 StickySelects_11 ( // @[MemPrimitives.scala 121:29:@16001.4]
    .clock(StickySelects_11_clock),
    .reset(StickySelects_11_reset),
    .io_ins_0(StickySelects_11_io_ins_0),
    .io_ins_1(StickySelects_11_io_ins_1),
    .io_ins_2(StickySelects_11_io_ins_2),
    .io_ins_3(StickySelects_11_io_ins_3),
    .io_outs_0(StickySelects_11_io_outs_0),
    .io_outs_1(StickySelects_11_io_outs_1),
    .io_outs_2(StickySelects_11_io_outs_2),
    .io_outs_3(StickySelects_11_io_outs_3)
  );
  StickySelects_16 StickySelects_12 ( // @[MemPrimitives.scala 121:29:@16037.4]
    .clock(StickySelects_12_clock),
    .reset(StickySelects_12_reset),
    .io_ins_0(StickySelects_12_io_ins_0),
    .io_ins_1(StickySelects_12_io_ins_1),
    .io_outs_0(StickySelects_12_io_outs_0),
    .io_outs_1(StickySelects_12_io_outs_1)
  );
  StickySelects_17 StickySelects_13 ( // @[MemPrimitives.scala 121:29:@16071.4]
    .clock(StickySelects_13_clock),
    .reset(StickySelects_13_reset),
    .io_ins_0(StickySelects_13_io_ins_0),
    .io_ins_1(StickySelects_13_io_ins_1),
    .io_ins_2(StickySelects_13_io_ins_2),
    .io_ins_3(StickySelects_13_io_ins_3),
    .io_outs_0(StickySelects_13_io_outs_0),
    .io_outs_1(StickySelects_13_io_outs_1),
    .io_outs_2(StickySelects_13_io_outs_2),
    .io_outs_3(StickySelects_13_io_outs_3)
  );
  StickySelects_16 StickySelects_14 ( // @[MemPrimitives.scala 121:29:@16107.4]
    .clock(StickySelects_14_clock),
    .reset(StickySelects_14_reset),
    .io_ins_0(StickySelects_14_io_ins_0),
    .io_ins_1(StickySelects_14_io_ins_1),
    .io_outs_0(StickySelects_14_io_outs_0),
    .io_outs_1(StickySelects_14_io_outs_1)
  );
  StickySelects_17 StickySelects_15 ( // @[MemPrimitives.scala 121:29:@16141.4]
    .clock(StickySelects_15_clock),
    .reset(StickySelects_15_reset),
    .io_ins_0(StickySelects_15_io_ins_0),
    .io_ins_1(StickySelects_15_io_ins_1),
    .io_ins_2(StickySelects_15_io_ins_2),
    .io_ins_3(StickySelects_15_io_ins_3),
    .io_outs_0(StickySelects_15_io_outs_0),
    .io_outs_1(StickySelects_15_io_outs_1),
    .io_outs_2(StickySelects_15_io_outs_2),
    .io_outs_3(StickySelects_15_io_outs_3)
  );
  RetimeWrapper_52 RetimeWrapper ( // @[package.scala 93:22:@16194.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_1 ( // @[package.scala 93:22:@16202.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_2 ( // @[package.scala 93:22:@16210.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_3 ( // @[package.scala 93:22:@16218.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_4 ( // @[package.scala 93:22:@16226.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_5 ( // @[package.scala 93:22:@16234.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_6 ( // @[package.scala 93:22:@16242.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_7 ( // @[package.scala 93:22:@16250.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_8 ( // @[package.scala 93:22:@16290.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_9 ( // @[package.scala 93:22:@16298.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_10 ( // @[package.scala 93:22:@16306.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_11 ( // @[package.scala 93:22:@16314.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_12 ( // @[package.scala 93:22:@16322.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_13 ( // @[package.scala 93:22:@16330.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_14 ( // @[package.scala 93:22:@16338.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_15 ( // @[package.scala 93:22:@16346.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_16 ( // @[package.scala 93:22:@16386.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_17 ( // @[package.scala 93:22:@16394.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_18 ( // @[package.scala 93:22:@16402.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_19 ( // @[package.scala 93:22:@16410.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_20 ( // @[package.scala 93:22:@16418.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_21 ( // @[package.scala 93:22:@16426.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_22 ( // @[package.scala 93:22:@16434.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_23 ( // @[package.scala 93:22:@16442.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_24 ( // @[package.scala 93:22:@16482.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_25 ( // @[package.scala 93:22:@16490.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_26 ( // @[package.scala 93:22:@16498.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_27 ( // @[package.scala 93:22:@16506.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_28 ( // @[package.scala 93:22:@16514.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_29 ( // @[package.scala 93:22:@16522.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_30 ( // @[package.scala 93:22:@16530.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_31 ( // @[package.scala 93:22:@16538.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_32 ( // @[package.scala 93:22:@16578.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_33 ( // @[package.scala 93:22:@16586.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_34 ( // @[package.scala 93:22:@16594.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_35 ( // @[package.scala 93:22:@16602.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_36 ( // @[package.scala 93:22:@16610.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_37 ( // @[package.scala 93:22:@16618.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_38 ( // @[package.scala 93:22:@16626.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_39 ( // @[package.scala 93:22:@16634.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_40 ( // @[package.scala 93:22:@16674.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_41 ( // @[package.scala 93:22:@16682.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_42 ( // @[package.scala 93:22:@16690.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_43 ( // @[package.scala 93:22:@16698.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_44 ( // @[package.scala 93:22:@16706.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_45 ( // @[package.scala 93:22:@16714.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_46 ( // @[package.scala 93:22:@16722.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_47 ( // @[package.scala 93:22:@16730.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  assign _T_264 = io_wPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@15417.4]
  assign _T_266 = io_wPort_0_banks_1 == 3'h0; // @[MemPrimitives.scala 82:210:@15418.4]
  assign _T_267 = _T_264 & _T_266; // @[MemPrimitives.scala 82:228:@15419.4]
  assign _T_268 = io_wPort_0_en_0 & _T_267; // @[MemPrimitives.scala 83:102:@15420.4]
  assign _T_270 = {_T_268,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@15422.4]
  assign _T_275 = io_wPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@15429.4]
  assign _T_277 = io_wPort_1_banks_1 == 3'h1; // @[MemPrimitives.scala 82:210:@15430.4]
  assign _T_278 = _T_275 & _T_277; // @[MemPrimitives.scala 82:228:@15431.4]
  assign _T_279 = io_wPort_1_en_0 & _T_278; // @[MemPrimitives.scala 83:102:@15432.4]
  assign _T_281 = {_T_279,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@15434.4]
  assign _T_288 = io_wPort_0_banks_1 == 3'h2; // @[MemPrimitives.scala 82:210:@15442.4]
  assign _T_289 = _T_264 & _T_288; // @[MemPrimitives.scala 82:228:@15443.4]
  assign _T_290 = io_wPort_0_en_0 & _T_289; // @[MemPrimitives.scala 83:102:@15444.4]
  assign _T_292 = {_T_290,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@15446.4]
  assign _T_299 = io_wPort_1_banks_1 == 3'h3; // @[MemPrimitives.scala 82:210:@15454.4]
  assign _T_300 = _T_275 & _T_299; // @[MemPrimitives.scala 82:228:@15455.4]
  assign _T_301 = io_wPort_1_en_0 & _T_300; // @[MemPrimitives.scala 83:102:@15456.4]
  assign _T_303 = {_T_301,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@15458.4]
  assign _T_308 = io_wPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@15465.4]
  assign _T_311 = _T_308 & _T_266; // @[MemPrimitives.scala 82:228:@15467.4]
  assign _T_312 = io_wPort_0_en_0 & _T_311; // @[MemPrimitives.scala 83:102:@15468.4]
  assign _T_314 = {_T_312,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@15470.4]
  assign _T_319 = io_wPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@15477.4]
  assign _T_322 = _T_319 & _T_277; // @[MemPrimitives.scala 82:228:@15479.4]
  assign _T_323 = io_wPort_1_en_0 & _T_322; // @[MemPrimitives.scala 83:102:@15480.4]
  assign _T_325 = {_T_323,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@15482.4]
  assign _T_333 = _T_308 & _T_288; // @[MemPrimitives.scala 82:228:@15491.4]
  assign _T_334 = io_wPort_0_en_0 & _T_333; // @[MemPrimitives.scala 83:102:@15492.4]
  assign _T_336 = {_T_334,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@15494.4]
  assign _T_344 = _T_319 & _T_299; // @[MemPrimitives.scala 82:228:@15503.4]
  assign _T_345 = io_wPort_1_en_0 & _T_344; // @[MemPrimitives.scala 83:102:@15504.4]
  assign _T_347 = {_T_345,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@15506.4]
  assign _T_352 = io_wPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@15513.4]
  assign _T_355 = _T_352 & _T_266; // @[MemPrimitives.scala 82:228:@15515.4]
  assign _T_356 = io_wPort_0_en_0 & _T_355; // @[MemPrimitives.scala 83:102:@15516.4]
  assign _T_358 = {_T_356,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@15518.4]
  assign _T_363 = io_wPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@15525.4]
  assign _T_366 = _T_363 & _T_277; // @[MemPrimitives.scala 82:228:@15527.4]
  assign _T_367 = io_wPort_1_en_0 & _T_366; // @[MemPrimitives.scala 83:102:@15528.4]
  assign _T_369 = {_T_367,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@15530.4]
  assign _T_377 = _T_352 & _T_288; // @[MemPrimitives.scala 82:228:@15539.4]
  assign _T_378 = io_wPort_0_en_0 & _T_377; // @[MemPrimitives.scala 83:102:@15540.4]
  assign _T_380 = {_T_378,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@15542.4]
  assign _T_388 = _T_363 & _T_299; // @[MemPrimitives.scala 82:228:@15551.4]
  assign _T_389 = io_wPort_1_en_0 & _T_388; // @[MemPrimitives.scala 83:102:@15552.4]
  assign _T_391 = {_T_389,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@15554.4]
  assign _T_396 = io_wPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@15561.4]
  assign _T_399 = _T_396 & _T_266; // @[MemPrimitives.scala 82:228:@15563.4]
  assign _T_400 = io_wPort_0_en_0 & _T_399; // @[MemPrimitives.scala 83:102:@15564.4]
  assign _T_402 = {_T_400,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@15566.4]
  assign _T_407 = io_wPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@15573.4]
  assign _T_410 = _T_407 & _T_277; // @[MemPrimitives.scala 82:228:@15575.4]
  assign _T_411 = io_wPort_1_en_0 & _T_410; // @[MemPrimitives.scala 83:102:@15576.4]
  assign _T_413 = {_T_411,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@15578.4]
  assign _T_421 = _T_396 & _T_288; // @[MemPrimitives.scala 82:228:@15587.4]
  assign _T_422 = io_wPort_0_en_0 & _T_421; // @[MemPrimitives.scala 83:102:@15588.4]
  assign _T_424 = {_T_422,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@15590.4]
  assign _T_432 = _T_407 & _T_299; // @[MemPrimitives.scala 82:228:@15599.4]
  assign _T_433 = io_wPort_1_en_0 & _T_432; // @[MemPrimitives.scala 83:102:@15600.4]
  assign _T_435 = {_T_433,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@15602.4]
  assign _T_440 = io_rPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@15609.4]
  assign _T_442 = io_rPort_1_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@15610.4]
  assign _T_443 = _T_440 & _T_442; // @[MemPrimitives.scala 110:228:@15611.4]
  assign _T_446 = io_rPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@15613.4]
  assign _T_448 = io_rPort_2_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@15614.4]
  assign _T_449 = _T_446 & _T_448; // @[MemPrimitives.scala 110:228:@15615.4]
  assign _T_451 = StickySelects_io_outs_0; // @[MemPrimitives.scala 123:41:@15622.4]
  assign _T_452 = StickySelects_io_outs_1; // @[MemPrimitives.scala 123:41:@15623.4]
  assign _T_454 = {_T_451,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@15625.4]
  assign _T_456 = {_T_452,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@15627.4]
  assign _T_457 = _T_451 ? _T_454 : _T_456; // @[Mux.scala 31:69:@15628.4]
  assign _T_462 = io_rPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@15635.4]
  assign _T_464 = io_rPort_0_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@15636.4]
  assign _T_465 = _T_462 & _T_464; // @[MemPrimitives.scala 110:228:@15637.4]
  assign _T_468 = io_rPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@15639.4]
  assign _T_470 = io_rPort_3_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@15640.4]
  assign _T_471 = _T_468 & _T_470; // @[MemPrimitives.scala 110:228:@15641.4]
  assign _T_474 = io_rPort_4_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@15643.4]
  assign _T_476 = io_rPort_4_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@15644.4]
  assign _T_477 = _T_474 & _T_476; // @[MemPrimitives.scala 110:228:@15645.4]
  assign _T_480 = io_rPort_5_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@15647.4]
  assign _T_482 = io_rPort_5_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@15648.4]
  assign _T_483 = _T_480 & _T_482; // @[MemPrimitives.scala 110:228:@15649.4]
  assign _T_485 = StickySelects_1_io_outs_0; // @[MemPrimitives.scala 123:41:@15658.4]
  assign _T_486 = StickySelects_1_io_outs_1; // @[MemPrimitives.scala 123:41:@15659.4]
  assign _T_487 = StickySelects_1_io_outs_2; // @[MemPrimitives.scala 123:41:@15660.4]
  assign _T_488 = StickySelects_1_io_outs_3; // @[MemPrimitives.scala 123:41:@15661.4]
  assign _T_490 = {_T_485,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@15663.4]
  assign _T_492 = {_T_486,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@15665.4]
  assign _T_494 = {_T_487,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@15667.4]
  assign _T_496 = {_T_488,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@15669.4]
  assign _T_497 = _T_487 ? _T_494 : _T_496; // @[Mux.scala 31:69:@15670.4]
  assign _T_498 = _T_486 ? _T_492 : _T_497; // @[Mux.scala 31:69:@15671.4]
  assign _T_499 = _T_485 ? _T_490 : _T_498; // @[Mux.scala 31:69:@15672.4]
  assign _T_506 = io_rPort_1_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@15680.4]
  assign _T_507 = _T_440 & _T_506; // @[MemPrimitives.scala 110:228:@15681.4]
  assign _T_512 = io_rPort_2_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@15684.4]
  assign _T_513 = _T_446 & _T_512; // @[MemPrimitives.scala 110:228:@15685.4]
  assign _T_515 = StickySelects_2_io_outs_0; // @[MemPrimitives.scala 123:41:@15692.4]
  assign _T_516 = StickySelects_2_io_outs_1; // @[MemPrimitives.scala 123:41:@15693.4]
  assign _T_518 = {_T_515,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@15695.4]
  assign _T_520 = {_T_516,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@15697.4]
  assign _T_521 = _T_515 ? _T_518 : _T_520; // @[Mux.scala 31:69:@15698.4]
  assign _T_528 = io_rPort_0_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@15706.4]
  assign _T_529 = _T_462 & _T_528; // @[MemPrimitives.scala 110:228:@15707.4]
  assign _T_534 = io_rPort_3_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@15710.4]
  assign _T_535 = _T_468 & _T_534; // @[MemPrimitives.scala 110:228:@15711.4]
  assign _T_540 = io_rPort_4_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@15714.4]
  assign _T_541 = _T_474 & _T_540; // @[MemPrimitives.scala 110:228:@15715.4]
  assign _T_546 = io_rPort_5_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@15718.4]
  assign _T_547 = _T_480 & _T_546; // @[MemPrimitives.scala 110:228:@15719.4]
  assign _T_549 = StickySelects_3_io_outs_0; // @[MemPrimitives.scala 123:41:@15728.4]
  assign _T_550 = StickySelects_3_io_outs_1; // @[MemPrimitives.scala 123:41:@15729.4]
  assign _T_551 = StickySelects_3_io_outs_2; // @[MemPrimitives.scala 123:41:@15730.4]
  assign _T_552 = StickySelects_3_io_outs_3; // @[MemPrimitives.scala 123:41:@15731.4]
  assign _T_554 = {_T_549,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@15733.4]
  assign _T_556 = {_T_550,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@15735.4]
  assign _T_558 = {_T_551,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@15737.4]
  assign _T_560 = {_T_552,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@15739.4]
  assign _T_561 = _T_551 ? _T_558 : _T_560; // @[Mux.scala 31:69:@15740.4]
  assign _T_562 = _T_550 ? _T_556 : _T_561; // @[Mux.scala 31:69:@15741.4]
  assign _T_563 = _T_549 ? _T_554 : _T_562; // @[Mux.scala 31:69:@15742.4]
  assign _T_568 = io_rPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@15749.4]
  assign _T_571 = _T_568 & _T_442; // @[MemPrimitives.scala 110:228:@15751.4]
  assign _T_574 = io_rPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@15753.4]
  assign _T_577 = _T_574 & _T_448; // @[MemPrimitives.scala 110:228:@15755.4]
  assign _T_579 = StickySelects_4_io_outs_0; // @[MemPrimitives.scala 123:41:@15762.4]
  assign _T_580 = StickySelects_4_io_outs_1; // @[MemPrimitives.scala 123:41:@15763.4]
  assign _T_582 = {_T_579,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@15765.4]
  assign _T_584 = {_T_580,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@15767.4]
  assign _T_585 = _T_579 ? _T_582 : _T_584; // @[Mux.scala 31:69:@15768.4]
  assign _T_590 = io_rPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@15775.4]
  assign _T_593 = _T_590 & _T_464; // @[MemPrimitives.scala 110:228:@15777.4]
  assign _T_596 = io_rPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@15779.4]
  assign _T_599 = _T_596 & _T_470; // @[MemPrimitives.scala 110:228:@15781.4]
  assign _T_602 = io_rPort_4_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@15783.4]
  assign _T_605 = _T_602 & _T_476; // @[MemPrimitives.scala 110:228:@15785.4]
  assign _T_608 = io_rPort_5_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@15787.4]
  assign _T_611 = _T_608 & _T_482; // @[MemPrimitives.scala 110:228:@15789.4]
  assign _T_613 = StickySelects_5_io_outs_0; // @[MemPrimitives.scala 123:41:@15798.4]
  assign _T_614 = StickySelects_5_io_outs_1; // @[MemPrimitives.scala 123:41:@15799.4]
  assign _T_615 = StickySelects_5_io_outs_2; // @[MemPrimitives.scala 123:41:@15800.4]
  assign _T_616 = StickySelects_5_io_outs_3; // @[MemPrimitives.scala 123:41:@15801.4]
  assign _T_618 = {_T_613,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@15803.4]
  assign _T_620 = {_T_614,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@15805.4]
  assign _T_622 = {_T_615,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@15807.4]
  assign _T_624 = {_T_616,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@15809.4]
  assign _T_625 = _T_615 ? _T_622 : _T_624; // @[Mux.scala 31:69:@15810.4]
  assign _T_626 = _T_614 ? _T_620 : _T_625; // @[Mux.scala 31:69:@15811.4]
  assign _T_627 = _T_613 ? _T_618 : _T_626; // @[Mux.scala 31:69:@15812.4]
  assign _T_635 = _T_568 & _T_506; // @[MemPrimitives.scala 110:228:@15821.4]
  assign _T_641 = _T_574 & _T_512; // @[MemPrimitives.scala 110:228:@15825.4]
  assign _T_643 = StickySelects_6_io_outs_0; // @[MemPrimitives.scala 123:41:@15832.4]
  assign _T_644 = StickySelects_6_io_outs_1; // @[MemPrimitives.scala 123:41:@15833.4]
  assign _T_646 = {_T_643,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@15835.4]
  assign _T_648 = {_T_644,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@15837.4]
  assign _T_649 = _T_643 ? _T_646 : _T_648; // @[Mux.scala 31:69:@15838.4]
  assign _T_657 = _T_590 & _T_528; // @[MemPrimitives.scala 110:228:@15847.4]
  assign _T_663 = _T_596 & _T_534; // @[MemPrimitives.scala 110:228:@15851.4]
  assign _T_669 = _T_602 & _T_540; // @[MemPrimitives.scala 110:228:@15855.4]
  assign _T_675 = _T_608 & _T_546; // @[MemPrimitives.scala 110:228:@15859.4]
  assign _T_677 = StickySelects_7_io_outs_0; // @[MemPrimitives.scala 123:41:@15868.4]
  assign _T_678 = StickySelects_7_io_outs_1; // @[MemPrimitives.scala 123:41:@15869.4]
  assign _T_679 = StickySelects_7_io_outs_2; // @[MemPrimitives.scala 123:41:@15870.4]
  assign _T_680 = StickySelects_7_io_outs_3; // @[MemPrimitives.scala 123:41:@15871.4]
  assign _T_682 = {_T_677,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@15873.4]
  assign _T_684 = {_T_678,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@15875.4]
  assign _T_686 = {_T_679,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@15877.4]
  assign _T_688 = {_T_680,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@15879.4]
  assign _T_689 = _T_679 ? _T_686 : _T_688; // @[Mux.scala 31:69:@15880.4]
  assign _T_690 = _T_678 ? _T_684 : _T_689; // @[Mux.scala 31:69:@15881.4]
  assign _T_691 = _T_677 ? _T_682 : _T_690; // @[Mux.scala 31:69:@15882.4]
  assign _T_696 = io_rPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@15889.4]
  assign _T_699 = _T_696 & _T_442; // @[MemPrimitives.scala 110:228:@15891.4]
  assign _T_702 = io_rPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@15893.4]
  assign _T_705 = _T_702 & _T_448; // @[MemPrimitives.scala 110:228:@15895.4]
  assign _T_707 = StickySelects_8_io_outs_0; // @[MemPrimitives.scala 123:41:@15902.4]
  assign _T_708 = StickySelects_8_io_outs_1; // @[MemPrimitives.scala 123:41:@15903.4]
  assign _T_710 = {_T_707,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@15905.4]
  assign _T_712 = {_T_708,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@15907.4]
  assign _T_713 = _T_707 ? _T_710 : _T_712; // @[Mux.scala 31:69:@15908.4]
  assign _T_718 = io_rPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@15915.4]
  assign _T_721 = _T_718 & _T_464; // @[MemPrimitives.scala 110:228:@15917.4]
  assign _T_724 = io_rPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@15919.4]
  assign _T_727 = _T_724 & _T_470; // @[MemPrimitives.scala 110:228:@15921.4]
  assign _T_730 = io_rPort_4_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@15923.4]
  assign _T_733 = _T_730 & _T_476; // @[MemPrimitives.scala 110:228:@15925.4]
  assign _T_736 = io_rPort_5_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@15927.4]
  assign _T_739 = _T_736 & _T_482; // @[MemPrimitives.scala 110:228:@15929.4]
  assign _T_741 = StickySelects_9_io_outs_0; // @[MemPrimitives.scala 123:41:@15938.4]
  assign _T_742 = StickySelects_9_io_outs_1; // @[MemPrimitives.scala 123:41:@15939.4]
  assign _T_743 = StickySelects_9_io_outs_2; // @[MemPrimitives.scala 123:41:@15940.4]
  assign _T_744 = StickySelects_9_io_outs_3; // @[MemPrimitives.scala 123:41:@15941.4]
  assign _T_746 = {_T_741,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@15943.4]
  assign _T_748 = {_T_742,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@15945.4]
  assign _T_750 = {_T_743,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@15947.4]
  assign _T_752 = {_T_744,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@15949.4]
  assign _T_753 = _T_743 ? _T_750 : _T_752; // @[Mux.scala 31:69:@15950.4]
  assign _T_754 = _T_742 ? _T_748 : _T_753; // @[Mux.scala 31:69:@15951.4]
  assign _T_755 = _T_741 ? _T_746 : _T_754; // @[Mux.scala 31:69:@15952.4]
  assign _T_763 = _T_696 & _T_506; // @[MemPrimitives.scala 110:228:@15961.4]
  assign _T_769 = _T_702 & _T_512; // @[MemPrimitives.scala 110:228:@15965.4]
  assign _T_771 = StickySelects_10_io_outs_0; // @[MemPrimitives.scala 123:41:@15972.4]
  assign _T_772 = StickySelects_10_io_outs_1; // @[MemPrimitives.scala 123:41:@15973.4]
  assign _T_774 = {_T_771,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@15975.4]
  assign _T_776 = {_T_772,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@15977.4]
  assign _T_777 = _T_771 ? _T_774 : _T_776; // @[Mux.scala 31:69:@15978.4]
  assign _T_785 = _T_718 & _T_528; // @[MemPrimitives.scala 110:228:@15987.4]
  assign _T_791 = _T_724 & _T_534; // @[MemPrimitives.scala 110:228:@15991.4]
  assign _T_797 = _T_730 & _T_540; // @[MemPrimitives.scala 110:228:@15995.4]
  assign _T_803 = _T_736 & _T_546; // @[MemPrimitives.scala 110:228:@15999.4]
  assign _T_805 = StickySelects_11_io_outs_0; // @[MemPrimitives.scala 123:41:@16008.4]
  assign _T_806 = StickySelects_11_io_outs_1; // @[MemPrimitives.scala 123:41:@16009.4]
  assign _T_807 = StickySelects_11_io_outs_2; // @[MemPrimitives.scala 123:41:@16010.4]
  assign _T_808 = StickySelects_11_io_outs_3; // @[MemPrimitives.scala 123:41:@16011.4]
  assign _T_810 = {_T_805,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@16013.4]
  assign _T_812 = {_T_806,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@16015.4]
  assign _T_814 = {_T_807,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@16017.4]
  assign _T_816 = {_T_808,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@16019.4]
  assign _T_817 = _T_807 ? _T_814 : _T_816; // @[Mux.scala 31:69:@16020.4]
  assign _T_818 = _T_806 ? _T_812 : _T_817; // @[Mux.scala 31:69:@16021.4]
  assign _T_819 = _T_805 ? _T_810 : _T_818; // @[Mux.scala 31:69:@16022.4]
  assign _T_824 = io_rPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@16029.4]
  assign _T_827 = _T_824 & _T_442; // @[MemPrimitives.scala 110:228:@16031.4]
  assign _T_830 = io_rPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@16033.4]
  assign _T_833 = _T_830 & _T_448; // @[MemPrimitives.scala 110:228:@16035.4]
  assign _T_835 = StickySelects_12_io_outs_0; // @[MemPrimitives.scala 123:41:@16042.4]
  assign _T_836 = StickySelects_12_io_outs_1; // @[MemPrimitives.scala 123:41:@16043.4]
  assign _T_838 = {_T_835,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@16045.4]
  assign _T_840 = {_T_836,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@16047.4]
  assign _T_841 = _T_835 ? _T_838 : _T_840; // @[Mux.scala 31:69:@16048.4]
  assign _T_846 = io_rPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@16055.4]
  assign _T_849 = _T_846 & _T_464; // @[MemPrimitives.scala 110:228:@16057.4]
  assign _T_852 = io_rPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@16059.4]
  assign _T_855 = _T_852 & _T_470; // @[MemPrimitives.scala 110:228:@16061.4]
  assign _T_858 = io_rPort_4_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@16063.4]
  assign _T_861 = _T_858 & _T_476; // @[MemPrimitives.scala 110:228:@16065.4]
  assign _T_864 = io_rPort_5_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@16067.4]
  assign _T_867 = _T_864 & _T_482; // @[MemPrimitives.scala 110:228:@16069.4]
  assign _T_869 = StickySelects_13_io_outs_0; // @[MemPrimitives.scala 123:41:@16078.4]
  assign _T_870 = StickySelects_13_io_outs_1; // @[MemPrimitives.scala 123:41:@16079.4]
  assign _T_871 = StickySelects_13_io_outs_2; // @[MemPrimitives.scala 123:41:@16080.4]
  assign _T_872 = StickySelects_13_io_outs_3; // @[MemPrimitives.scala 123:41:@16081.4]
  assign _T_874 = {_T_869,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@16083.4]
  assign _T_876 = {_T_870,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@16085.4]
  assign _T_878 = {_T_871,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@16087.4]
  assign _T_880 = {_T_872,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@16089.4]
  assign _T_881 = _T_871 ? _T_878 : _T_880; // @[Mux.scala 31:69:@16090.4]
  assign _T_882 = _T_870 ? _T_876 : _T_881; // @[Mux.scala 31:69:@16091.4]
  assign _T_883 = _T_869 ? _T_874 : _T_882; // @[Mux.scala 31:69:@16092.4]
  assign _T_891 = _T_824 & _T_506; // @[MemPrimitives.scala 110:228:@16101.4]
  assign _T_897 = _T_830 & _T_512; // @[MemPrimitives.scala 110:228:@16105.4]
  assign _T_899 = StickySelects_14_io_outs_0; // @[MemPrimitives.scala 123:41:@16112.4]
  assign _T_900 = StickySelects_14_io_outs_1; // @[MemPrimitives.scala 123:41:@16113.4]
  assign _T_902 = {_T_899,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@16115.4]
  assign _T_904 = {_T_900,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@16117.4]
  assign _T_905 = _T_899 ? _T_902 : _T_904; // @[Mux.scala 31:69:@16118.4]
  assign _T_913 = _T_846 & _T_528; // @[MemPrimitives.scala 110:228:@16127.4]
  assign _T_919 = _T_852 & _T_534; // @[MemPrimitives.scala 110:228:@16131.4]
  assign _T_925 = _T_858 & _T_540; // @[MemPrimitives.scala 110:228:@16135.4]
  assign _T_931 = _T_864 & _T_546; // @[MemPrimitives.scala 110:228:@16139.4]
  assign _T_933 = StickySelects_15_io_outs_0; // @[MemPrimitives.scala 123:41:@16148.4]
  assign _T_934 = StickySelects_15_io_outs_1; // @[MemPrimitives.scala 123:41:@16149.4]
  assign _T_935 = StickySelects_15_io_outs_2; // @[MemPrimitives.scala 123:41:@16150.4]
  assign _T_936 = StickySelects_15_io_outs_3; // @[MemPrimitives.scala 123:41:@16151.4]
  assign _T_938 = {_T_933,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@16153.4]
  assign _T_940 = {_T_934,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@16155.4]
  assign _T_942 = {_T_935,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@16157.4]
  assign _T_944 = {_T_936,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@16159.4]
  assign _T_945 = _T_935 ? _T_942 : _T_944; // @[Mux.scala 31:69:@16160.4]
  assign _T_946 = _T_934 ? _T_940 : _T_945; // @[Mux.scala 31:69:@16161.4]
  assign _T_947 = _T_933 ? _T_938 : _T_946; // @[Mux.scala 31:69:@16162.4]
  assign _T_1011 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@16247.4 package.scala 96:25:@16248.4]
  assign _T_1015 = _T_1011 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@16257.4]
  assign _T_1008 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@16239.4 package.scala 96:25:@16240.4]
  assign _T_1016 = _T_1008 ? Mem1D_11_io_output : _T_1015; // @[Mux.scala 31:69:@16258.4]
  assign _T_1005 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@16231.4 package.scala 96:25:@16232.4]
  assign _T_1017 = _T_1005 ? Mem1D_9_io_output : _T_1016; // @[Mux.scala 31:69:@16259.4]
  assign _T_1002 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@16223.4 package.scala 96:25:@16224.4]
  assign _T_1018 = _T_1002 ? Mem1D_7_io_output : _T_1017; // @[Mux.scala 31:69:@16260.4]
  assign _T_999 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@16215.4 package.scala 96:25:@16216.4]
  assign _T_1019 = _T_999 ? Mem1D_5_io_output : _T_1018; // @[Mux.scala 31:69:@16261.4]
  assign _T_996 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@16207.4 package.scala 96:25:@16208.4]
  assign _T_1020 = _T_996 ? Mem1D_3_io_output : _T_1019; // @[Mux.scala 31:69:@16262.4]
  assign _T_993 = RetimeWrapper_io_out; // @[package.scala 96:25:@16199.4 package.scala 96:25:@16200.4]
  assign _T_1082 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@16343.4 package.scala 96:25:@16344.4]
  assign _T_1086 = _T_1082 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@16353.4]
  assign _T_1079 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@16335.4 package.scala 96:25:@16336.4]
  assign _T_1087 = _T_1079 ? Mem1D_10_io_output : _T_1086; // @[Mux.scala 31:69:@16354.4]
  assign _T_1076 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@16327.4 package.scala 96:25:@16328.4]
  assign _T_1088 = _T_1076 ? Mem1D_8_io_output : _T_1087; // @[Mux.scala 31:69:@16355.4]
  assign _T_1073 = RetimeWrapper_11_io_out; // @[package.scala 96:25:@16319.4 package.scala 96:25:@16320.4]
  assign _T_1089 = _T_1073 ? Mem1D_6_io_output : _T_1088; // @[Mux.scala 31:69:@16356.4]
  assign _T_1070 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@16311.4 package.scala 96:25:@16312.4]
  assign _T_1090 = _T_1070 ? Mem1D_4_io_output : _T_1089; // @[Mux.scala 31:69:@16357.4]
  assign _T_1067 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@16303.4 package.scala 96:25:@16304.4]
  assign _T_1091 = _T_1067 ? Mem1D_2_io_output : _T_1090; // @[Mux.scala 31:69:@16358.4]
  assign _T_1064 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@16295.4 package.scala 96:25:@16296.4]
  assign _T_1153 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@16439.4 package.scala 96:25:@16440.4]
  assign _T_1157 = _T_1153 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@16449.4]
  assign _T_1150 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@16431.4 package.scala 96:25:@16432.4]
  assign _T_1158 = _T_1150 ? Mem1D_10_io_output : _T_1157; // @[Mux.scala 31:69:@16450.4]
  assign _T_1147 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@16423.4 package.scala 96:25:@16424.4]
  assign _T_1159 = _T_1147 ? Mem1D_8_io_output : _T_1158; // @[Mux.scala 31:69:@16451.4]
  assign _T_1144 = RetimeWrapper_19_io_out; // @[package.scala 96:25:@16415.4 package.scala 96:25:@16416.4]
  assign _T_1160 = _T_1144 ? Mem1D_6_io_output : _T_1159; // @[Mux.scala 31:69:@16452.4]
  assign _T_1141 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@16407.4 package.scala 96:25:@16408.4]
  assign _T_1161 = _T_1141 ? Mem1D_4_io_output : _T_1160; // @[Mux.scala 31:69:@16453.4]
  assign _T_1138 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@16399.4 package.scala 96:25:@16400.4]
  assign _T_1162 = _T_1138 ? Mem1D_2_io_output : _T_1161; // @[Mux.scala 31:69:@16454.4]
  assign _T_1135 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@16391.4 package.scala 96:25:@16392.4]
  assign _T_1224 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@16535.4 package.scala 96:25:@16536.4]
  assign _T_1228 = _T_1224 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@16545.4]
  assign _T_1221 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@16527.4 package.scala 96:25:@16528.4]
  assign _T_1229 = _T_1221 ? Mem1D_11_io_output : _T_1228; // @[Mux.scala 31:69:@16546.4]
  assign _T_1218 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@16519.4 package.scala 96:25:@16520.4]
  assign _T_1230 = _T_1218 ? Mem1D_9_io_output : _T_1229; // @[Mux.scala 31:69:@16547.4]
  assign _T_1215 = RetimeWrapper_27_io_out; // @[package.scala 96:25:@16511.4 package.scala 96:25:@16512.4]
  assign _T_1231 = _T_1215 ? Mem1D_7_io_output : _T_1230; // @[Mux.scala 31:69:@16548.4]
  assign _T_1212 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@16503.4 package.scala 96:25:@16504.4]
  assign _T_1232 = _T_1212 ? Mem1D_5_io_output : _T_1231; // @[Mux.scala 31:69:@16549.4]
  assign _T_1209 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@16495.4 package.scala 96:25:@16496.4]
  assign _T_1233 = _T_1209 ? Mem1D_3_io_output : _T_1232; // @[Mux.scala 31:69:@16550.4]
  assign _T_1206 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@16487.4 package.scala 96:25:@16488.4]
  assign _T_1295 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@16631.4 package.scala 96:25:@16632.4]
  assign _T_1299 = _T_1295 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@16641.4]
  assign _T_1292 = RetimeWrapper_37_io_out; // @[package.scala 96:25:@16623.4 package.scala 96:25:@16624.4]
  assign _T_1300 = _T_1292 ? Mem1D_11_io_output : _T_1299; // @[Mux.scala 31:69:@16642.4]
  assign _T_1289 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@16615.4 package.scala 96:25:@16616.4]
  assign _T_1301 = _T_1289 ? Mem1D_9_io_output : _T_1300; // @[Mux.scala 31:69:@16643.4]
  assign _T_1286 = RetimeWrapper_35_io_out; // @[package.scala 96:25:@16607.4 package.scala 96:25:@16608.4]
  assign _T_1302 = _T_1286 ? Mem1D_7_io_output : _T_1301; // @[Mux.scala 31:69:@16644.4]
  assign _T_1283 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@16599.4 package.scala 96:25:@16600.4]
  assign _T_1303 = _T_1283 ? Mem1D_5_io_output : _T_1302; // @[Mux.scala 31:69:@16645.4]
  assign _T_1280 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@16591.4 package.scala 96:25:@16592.4]
  assign _T_1304 = _T_1280 ? Mem1D_3_io_output : _T_1303; // @[Mux.scala 31:69:@16646.4]
  assign _T_1277 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@16583.4 package.scala 96:25:@16584.4]
  assign _T_1366 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@16727.4 package.scala 96:25:@16728.4]
  assign _T_1370 = _T_1366 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@16737.4]
  assign _T_1363 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@16719.4 package.scala 96:25:@16720.4]
  assign _T_1371 = _T_1363 ? Mem1D_11_io_output : _T_1370; // @[Mux.scala 31:69:@16738.4]
  assign _T_1360 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@16711.4 package.scala 96:25:@16712.4]
  assign _T_1372 = _T_1360 ? Mem1D_9_io_output : _T_1371; // @[Mux.scala 31:69:@16739.4]
  assign _T_1357 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@16703.4 package.scala 96:25:@16704.4]
  assign _T_1373 = _T_1357 ? Mem1D_7_io_output : _T_1372; // @[Mux.scala 31:69:@16740.4]
  assign _T_1354 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@16695.4 package.scala 96:25:@16696.4]
  assign _T_1374 = _T_1354 ? Mem1D_5_io_output : _T_1373; // @[Mux.scala 31:69:@16741.4]
  assign _T_1351 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@16687.4 package.scala 96:25:@16688.4]
  assign _T_1375 = _T_1351 ? Mem1D_3_io_output : _T_1374; // @[Mux.scala 31:69:@16742.4]
  assign _T_1348 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@16679.4 package.scala 96:25:@16680.4]
  assign io_rPort_5_output_0 = _T_1348 ? Mem1D_1_io_output : _T_1375; // @[MemPrimitives.scala 148:13:@16744.4]
  assign io_rPort_4_output_0 = _T_1277 ? Mem1D_1_io_output : _T_1304; // @[MemPrimitives.scala 148:13:@16648.4]
  assign io_rPort_3_output_0 = _T_1206 ? Mem1D_1_io_output : _T_1233; // @[MemPrimitives.scala 148:13:@16552.4]
  assign io_rPort_2_output_0 = _T_1135 ? Mem1D_io_output : _T_1162; // @[MemPrimitives.scala 148:13:@16456.4]
  assign io_rPort_1_output_0 = _T_1064 ? Mem1D_io_output : _T_1091; // @[MemPrimitives.scala 148:13:@16360.4]
  assign io_rPort_0_output_0 = _T_993 ? Mem1D_1_io_output : _T_1020; // @[MemPrimitives.scala 148:13:@16264.4]
  assign Mem1D_clock = clock; // @[:@15162.4]
  assign Mem1D_reset = reset; // @[:@15163.4]
  assign Mem1D_io_r_ofs_0 = _T_457[0]; // @[MemPrimitives.scala 127:28:@15632.4]
  assign Mem1D_io_r_backpressure = _T_457[1]; // @[MemPrimitives.scala 128:32:@15633.4]
  assign Mem1D_io_w_ofs_0 = _T_270[0]; // @[MemPrimitives.scala 94:28:@15426.4]
  assign Mem1D_io_w_data_0 = _T_270[8:1]; // @[MemPrimitives.scala 95:29:@15427.4]
  assign Mem1D_io_w_en_0 = _T_270[9]; // @[MemPrimitives.scala 96:27:@15428.4]
  assign Mem1D_1_clock = clock; // @[:@15178.4]
  assign Mem1D_1_reset = reset; // @[:@15179.4]
  assign Mem1D_1_io_r_ofs_0 = _T_499[0]; // @[MemPrimitives.scala 127:28:@15676.4]
  assign Mem1D_1_io_r_backpressure = _T_499[1]; // @[MemPrimitives.scala 128:32:@15677.4]
  assign Mem1D_1_io_w_ofs_0 = _T_281[0]; // @[MemPrimitives.scala 94:28:@15438.4]
  assign Mem1D_1_io_w_data_0 = _T_281[8:1]; // @[MemPrimitives.scala 95:29:@15439.4]
  assign Mem1D_1_io_w_en_0 = _T_281[9]; // @[MemPrimitives.scala 96:27:@15440.4]
  assign Mem1D_2_clock = clock; // @[:@15194.4]
  assign Mem1D_2_reset = reset; // @[:@15195.4]
  assign Mem1D_2_io_r_ofs_0 = _T_521[0]; // @[MemPrimitives.scala 127:28:@15702.4]
  assign Mem1D_2_io_r_backpressure = _T_521[1]; // @[MemPrimitives.scala 128:32:@15703.4]
  assign Mem1D_2_io_w_ofs_0 = _T_292[0]; // @[MemPrimitives.scala 94:28:@15450.4]
  assign Mem1D_2_io_w_data_0 = _T_292[8:1]; // @[MemPrimitives.scala 95:29:@15451.4]
  assign Mem1D_2_io_w_en_0 = _T_292[9]; // @[MemPrimitives.scala 96:27:@15452.4]
  assign Mem1D_3_clock = clock; // @[:@15210.4]
  assign Mem1D_3_reset = reset; // @[:@15211.4]
  assign Mem1D_3_io_r_ofs_0 = _T_563[0]; // @[MemPrimitives.scala 127:28:@15746.4]
  assign Mem1D_3_io_r_backpressure = _T_563[1]; // @[MemPrimitives.scala 128:32:@15747.4]
  assign Mem1D_3_io_w_ofs_0 = _T_303[0]; // @[MemPrimitives.scala 94:28:@15462.4]
  assign Mem1D_3_io_w_data_0 = _T_303[8:1]; // @[MemPrimitives.scala 95:29:@15463.4]
  assign Mem1D_3_io_w_en_0 = _T_303[9]; // @[MemPrimitives.scala 96:27:@15464.4]
  assign Mem1D_4_clock = clock; // @[:@15226.4]
  assign Mem1D_4_reset = reset; // @[:@15227.4]
  assign Mem1D_4_io_r_ofs_0 = _T_585[0]; // @[MemPrimitives.scala 127:28:@15772.4]
  assign Mem1D_4_io_r_backpressure = _T_585[1]; // @[MemPrimitives.scala 128:32:@15773.4]
  assign Mem1D_4_io_w_ofs_0 = _T_314[0]; // @[MemPrimitives.scala 94:28:@15474.4]
  assign Mem1D_4_io_w_data_0 = _T_314[8:1]; // @[MemPrimitives.scala 95:29:@15475.4]
  assign Mem1D_4_io_w_en_0 = _T_314[9]; // @[MemPrimitives.scala 96:27:@15476.4]
  assign Mem1D_5_clock = clock; // @[:@15242.4]
  assign Mem1D_5_reset = reset; // @[:@15243.4]
  assign Mem1D_5_io_r_ofs_0 = _T_627[0]; // @[MemPrimitives.scala 127:28:@15816.4]
  assign Mem1D_5_io_r_backpressure = _T_627[1]; // @[MemPrimitives.scala 128:32:@15817.4]
  assign Mem1D_5_io_w_ofs_0 = _T_325[0]; // @[MemPrimitives.scala 94:28:@15486.4]
  assign Mem1D_5_io_w_data_0 = _T_325[8:1]; // @[MemPrimitives.scala 95:29:@15487.4]
  assign Mem1D_5_io_w_en_0 = _T_325[9]; // @[MemPrimitives.scala 96:27:@15488.4]
  assign Mem1D_6_clock = clock; // @[:@15258.4]
  assign Mem1D_6_reset = reset; // @[:@15259.4]
  assign Mem1D_6_io_r_ofs_0 = _T_649[0]; // @[MemPrimitives.scala 127:28:@15842.4]
  assign Mem1D_6_io_r_backpressure = _T_649[1]; // @[MemPrimitives.scala 128:32:@15843.4]
  assign Mem1D_6_io_w_ofs_0 = _T_336[0]; // @[MemPrimitives.scala 94:28:@15498.4]
  assign Mem1D_6_io_w_data_0 = _T_336[8:1]; // @[MemPrimitives.scala 95:29:@15499.4]
  assign Mem1D_6_io_w_en_0 = _T_336[9]; // @[MemPrimitives.scala 96:27:@15500.4]
  assign Mem1D_7_clock = clock; // @[:@15274.4]
  assign Mem1D_7_reset = reset; // @[:@15275.4]
  assign Mem1D_7_io_r_ofs_0 = _T_691[0]; // @[MemPrimitives.scala 127:28:@15886.4]
  assign Mem1D_7_io_r_backpressure = _T_691[1]; // @[MemPrimitives.scala 128:32:@15887.4]
  assign Mem1D_7_io_w_ofs_0 = _T_347[0]; // @[MemPrimitives.scala 94:28:@15510.4]
  assign Mem1D_7_io_w_data_0 = _T_347[8:1]; // @[MemPrimitives.scala 95:29:@15511.4]
  assign Mem1D_7_io_w_en_0 = _T_347[9]; // @[MemPrimitives.scala 96:27:@15512.4]
  assign Mem1D_8_clock = clock; // @[:@15290.4]
  assign Mem1D_8_reset = reset; // @[:@15291.4]
  assign Mem1D_8_io_r_ofs_0 = _T_713[0]; // @[MemPrimitives.scala 127:28:@15912.4]
  assign Mem1D_8_io_r_backpressure = _T_713[1]; // @[MemPrimitives.scala 128:32:@15913.4]
  assign Mem1D_8_io_w_ofs_0 = _T_358[0]; // @[MemPrimitives.scala 94:28:@15522.4]
  assign Mem1D_8_io_w_data_0 = _T_358[8:1]; // @[MemPrimitives.scala 95:29:@15523.4]
  assign Mem1D_8_io_w_en_0 = _T_358[9]; // @[MemPrimitives.scala 96:27:@15524.4]
  assign Mem1D_9_clock = clock; // @[:@15306.4]
  assign Mem1D_9_reset = reset; // @[:@15307.4]
  assign Mem1D_9_io_r_ofs_0 = _T_755[0]; // @[MemPrimitives.scala 127:28:@15956.4]
  assign Mem1D_9_io_r_backpressure = _T_755[1]; // @[MemPrimitives.scala 128:32:@15957.4]
  assign Mem1D_9_io_w_ofs_0 = _T_369[0]; // @[MemPrimitives.scala 94:28:@15534.4]
  assign Mem1D_9_io_w_data_0 = _T_369[8:1]; // @[MemPrimitives.scala 95:29:@15535.4]
  assign Mem1D_9_io_w_en_0 = _T_369[9]; // @[MemPrimitives.scala 96:27:@15536.4]
  assign Mem1D_10_clock = clock; // @[:@15322.4]
  assign Mem1D_10_reset = reset; // @[:@15323.4]
  assign Mem1D_10_io_r_ofs_0 = _T_777[0]; // @[MemPrimitives.scala 127:28:@15982.4]
  assign Mem1D_10_io_r_backpressure = _T_777[1]; // @[MemPrimitives.scala 128:32:@15983.4]
  assign Mem1D_10_io_w_ofs_0 = _T_380[0]; // @[MemPrimitives.scala 94:28:@15546.4]
  assign Mem1D_10_io_w_data_0 = _T_380[8:1]; // @[MemPrimitives.scala 95:29:@15547.4]
  assign Mem1D_10_io_w_en_0 = _T_380[9]; // @[MemPrimitives.scala 96:27:@15548.4]
  assign Mem1D_11_clock = clock; // @[:@15338.4]
  assign Mem1D_11_reset = reset; // @[:@15339.4]
  assign Mem1D_11_io_r_ofs_0 = _T_819[0]; // @[MemPrimitives.scala 127:28:@16026.4]
  assign Mem1D_11_io_r_backpressure = _T_819[1]; // @[MemPrimitives.scala 128:32:@16027.4]
  assign Mem1D_11_io_w_ofs_0 = _T_391[0]; // @[MemPrimitives.scala 94:28:@15558.4]
  assign Mem1D_11_io_w_data_0 = _T_391[8:1]; // @[MemPrimitives.scala 95:29:@15559.4]
  assign Mem1D_11_io_w_en_0 = _T_391[9]; // @[MemPrimitives.scala 96:27:@15560.4]
  assign Mem1D_12_clock = clock; // @[:@15354.4]
  assign Mem1D_12_reset = reset; // @[:@15355.4]
  assign Mem1D_12_io_r_ofs_0 = _T_841[0]; // @[MemPrimitives.scala 127:28:@16052.4]
  assign Mem1D_12_io_r_backpressure = _T_841[1]; // @[MemPrimitives.scala 128:32:@16053.4]
  assign Mem1D_12_io_w_ofs_0 = _T_402[0]; // @[MemPrimitives.scala 94:28:@15570.4]
  assign Mem1D_12_io_w_data_0 = _T_402[8:1]; // @[MemPrimitives.scala 95:29:@15571.4]
  assign Mem1D_12_io_w_en_0 = _T_402[9]; // @[MemPrimitives.scala 96:27:@15572.4]
  assign Mem1D_13_clock = clock; // @[:@15370.4]
  assign Mem1D_13_reset = reset; // @[:@15371.4]
  assign Mem1D_13_io_r_ofs_0 = _T_883[0]; // @[MemPrimitives.scala 127:28:@16096.4]
  assign Mem1D_13_io_r_backpressure = _T_883[1]; // @[MemPrimitives.scala 128:32:@16097.4]
  assign Mem1D_13_io_w_ofs_0 = _T_413[0]; // @[MemPrimitives.scala 94:28:@15582.4]
  assign Mem1D_13_io_w_data_0 = _T_413[8:1]; // @[MemPrimitives.scala 95:29:@15583.4]
  assign Mem1D_13_io_w_en_0 = _T_413[9]; // @[MemPrimitives.scala 96:27:@15584.4]
  assign Mem1D_14_clock = clock; // @[:@15386.4]
  assign Mem1D_14_reset = reset; // @[:@15387.4]
  assign Mem1D_14_io_r_ofs_0 = _T_905[0]; // @[MemPrimitives.scala 127:28:@16122.4]
  assign Mem1D_14_io_r_backpressure = _T_905[1]; // @[MemPrimitives.scala 128:32:@16123.4]
  assign Mem1D_14_io_w_ofs_0 = _T_424[0]; // @[MemPrimitives.scala 94:28:@15594.4]
  assign Mem1D_14_io_w_data_0 = _T_424[8:1]; // @[MemPrimitives.scala 95:29:@15595.4]
  assign Mem1D_14_io_w_en_0 = _T_424[9]; // @[MemPrimitives.scala 96:27:@15596.4]
  assign Mem1D_15_clock = clock; // @[:@15402.4]
  assign Mem1D_15_reset = reset; // @[:@15403.4]
  assign Mem1D_15_io_r_ofs_0 = _T_947[0]; // @[MemPrimitives.scala 127:28:@16166.4]
  assign Mem1D_15_io_r_backpressure = _T_947[1]; // @[MemPrimitives.scala 128:32:@16167.4]
  assign Mem1D_15_io_w_ofs_0 = _T_435[0]; // @[MemPrimitives.scala 94:28:@15606.4]
  assign Mem1D_15_io_w_data_0 = _T_435[8:1]; // @[MemPrimitives.scala 95:29:@15607.4]
  assign Mem1D_15_io_w_en_0 = _T_435[9]; // @[MemPrimitives.scala 96:27:@15608.4]
  assign StickySelects_clock = clock; // @[:@15618.4]
  assign StickySelects_reset = reset; // @[:@15619.4]
  assign StickySelects_io_ins_0 = io_rPort_1_en_0 & _T_443; // @[MemPrimitives.scala 122:60:@15620.4]
  assign StickySelects_io_ins_1 = io_rPort_2_en_0 & _T_449; // @[MemPrimitives.scala 122:60:@15621.4]
  assign StickySelects_1_clock = clock; // @[:@15652.4]
  assign StickySelects_1_reset = reset; // @[:@15653.4]
  assign StickySelects_1_io_ins_0 = io_rPort_0_en_0 & _T_465; // @[MemPrimitives.scala 122:60:@15654.4]
  assign StickySelects_1_io_ins_1 = io_rPort_3_en_0 & _T_471; // @[MemPrimitives.scala 122:60:@15655.4]
  assign StickySelects_1_io_ins_2 = io_rPort_4_en_0 & _T_477; // @[MemPrimitives.scala 122:60:@15656.4]
  assign StickySelects_1_io_ins_3 = io_rPort_5_en_0 & _T_483; // @[MemPrimitives.scala 122:60:@15657.4]
  assign StickySelects_2_clock = clock; // @[:@15688.4]
  assign StickySelects_2_reset = reset; // @[:@15689.4]
  assign StickySelects_2_io_ins_0 = io_rPort_1_en_0 & _T_507; // @[MemPrimitives.scala 122:60:@15690.4]
  assign StickySelects_2_io_ins_1 = io_rPort_2_en_0 & _T_513; // @[MemPrimitives.scala 122:60:@15691.4]
  assign StickySelects_3_clock = clock; // @[:@15722.4]
  assign StickySelects_3_reset = reset; // @[:@15723.4]
  assign StickySelects_3_io_ins_0 = io_rPort_0_en_0 & _T_529; // @[MemPrimitives.scala 122:60:@15724.4]
  assign StickySelects_3_io_ins_1 = io_rPort_3_en_0 & _T_535; // @[MemPrimitives.scala 122:60:@15725.4]
  assign StickySelects_3_io_ins_2 = io_rPort_4_en_0 & _T_541; // @[MemPrimitives.scala 122:60:@15726.4]
  assign StickySelects_3_io_ins_3 = io_rPort_5_en_0 & _T_547; // @[MemPrimitives.scala 122:60:@15727.4]
  assign StickySelects_4_clock = clock; // @[:@15758.4]
  assign StickySelects_4_reset = reset; // @[:@15759.4]
  assign StickySelects_4_io_ins_0 = io_rPort_1_en_0 & _T_571; // @[MemPrimitives.scala 122:60:@15760.4]
  assign StickySelects_4_io_ins_1 = io_rPort_2_en_0 & _T_577; // @[MemPrimitives.scala 122:60:@15761.4]
  assign StickySelects_5_clock = clock; // @[:@15792.4]
  assign StickySelects_5_reset = reset; // @[:@15793.4]
  assign StickySelects_5_io_ins_0 = io_rPort_0_en_0 & _T_593; // @[MemPrimitives.scala 122:60:@15794.4]
  assign StickySelects_5_io_ins_1 = io_rPort_3_en_0 & _T_599; // @[MemPrimitives.scala 122:60:@15795.4]
  assign StickySelects_5_io_ins_2 = io_rPort_4_en_0 & _T_605; // @[MemPrimitives.scala 122:60:@15796.4]
  assign StickySelects_5_io_ins_3 = io_rPort_5_en_0 & _T_611; // @[MemPrimitives.scala 122:60:@15797.4]
  assign StickySelects_6_clock = clock; // @[:@15828.4]
  assign StickySelects_6_reset = reset; // @[:@15829.4]
  assign StickySelects_6_io_ins_0 = io_rPort_1_en_0 & _T_635; // @[MemPrimitives.scala 122:60:@15830.4]
  assign StickySelects_6_io_ins_1 = io_rPort_2_en_0 & _T_641; // @[MemPrimitives.scala 122:60:@15831.4]
  assign StickySelects_7_clock = clock; // @[:@15862.4]
  assign StickySelects_7_reset = reset; // @[:@15863.4]
  assign StickySelects_7_io_ins_0 = io_rPort_0_en_0 & _T_657; // @[MemPrimitives.scala 122:60:@15864.4]
  assign StickySelects_7_io_ins_1 = io_rPort_3_en_0 & _T_663; // @[MemPrimitives.scala 122:60:@15865.4]
  assign StickySelects_7_io_ins_2 = io_rPort_4_en_0 & _T_669; // @[MemPrimitives.scala 122:60:@15866.4]
  assign StickySelects_7_io_ins_3 = io_rPort_5_en_0 & _T_675; // @[MemPrimitives.scala 122:60:@15867.4]
  assign StickySelects_8_clock = clock; // @[:@15898.4]
  assign StickySelects_8_reset = reset; // @[:@15899.4]
  assign StickySelects_8_io_ins_0 = io_rPort_1_en_0 & _T_699; // @[MemPrimitives.scala 122:60:@15900.4]
  assign StickySelects_8_io_ins_1 = io_rPort_2_en_0 & _T_705; // @[MemPrimitives.scala 122:60:@15901.4]
  assign StickySelects_9_clock = clock; // @[:@15932.4]
  assign StickySelects_9_reset = reset; // @[:@15933.4]
  assign StickySelects_9_io_ins_0 = io_rPort_0_en_0 & _T_721; // @[MemPrimitives.scala 122:60:@15934.4]
  assign StickySelects_9_io_ins_1 = io_rPort_3_en_0 & _T_727; // @[MemPrimitives.scala 122:60:@15935.4]
  assign StickySelects_9_io_ins_2 = io_rPort_4_en_0 & _T_733; // @[MemPrimitives.scala 122:60:@15936.4]
  assign StickySelects_9_io_ins_3 = io_rPort_5_en_0 & _T_739; // @[MemPrimitives.scala 122:60:@15937.4]
  assign StickySelects_10_clock = clock; // @[:@15968.4]
  assign StickySelects_10_reset = reset; // @[:@15969.4]
  assign StickySelects_10_io_ins_0 = io_rPort_1_en_0 & _T_763; // @[MemPrimitives.scala 122:60:@15970.4]
  assign StickySelects_10_io_ins_1 = io_rPort_2_en_0 & _T_769; // @[MemPrimitives.scala 122:60:@15971.4]
  assign StickySelects_11_clock = clock; // @[:@16002.4]
  assign StickySelects_11_reset = reset; // @[:@16003.4]
  assign StickySelects_11_io_ins_0 = io_rPort_0_en_0 & _T_785; // @[MemPrimitives.scala 122:60:@16004.4]
  assign StickySelects_11_io_ins_1 = io_rPort_3_en_0 & _T_791; // @[MemPrimitives.scala 122:60:@16005.4]
  assign StickySelects_11_io_ins_2 = io_rPort_4_en_0 & _T_797; // @[MemPrimitives.scala 122:60:@16006.4]
  assign StickySelects_11_io_ins_3 = io_rPort_5_en_0 & _T_803; // @[MemPrimitives.scala 122:60:@16007.4]
  assign StickySelects_12_clock = clock; // @[:@16038.4]
  assign StickySelects_12_reset = reset; // @[:@16039.4]
  assign StickySelects_12_io_ins_0 = io_rPort_1_en_0 & _T_827; // @[MemPrimitives.scala 122:60:@16040.4]
  assign StickySelects_12_io_ins_1 = io_rPort_2_en_0 & _T_833; // @[MemPrimitives.scala 122:60:@16041.4]
  assign StickySelects_13_clock = clock; // @[:@16072.4]
  assign StickySelects_13_reset = reset; // @[:@16073.4]
  assign StickySelects_13_io_ins_0 = io_rPort_0_en_0 & _T_849; // @[MemPrimitives.scala 122:60:@16074.4]
  assign StickySelects_13_io_ins_1 = io_rPort_3_en_0 & _T_855; // @[MemPrimitives.scala 122:60:@16075.4]
  assign StickySelects_13_io_ins_2 = io_rPort_4_en_0 & _T_861; // @[MemPrimitives.scala 122:60:@16076.4]
  assign StickySelects_13_io_ins_3 = io_rPort_5_en_0 & _T_867; // @[MemPrimitives.scala 122:60:@16077.4]
  assign StickySelects_14_clock = clock; // @[:@16108.4]
  assign StickySelects_14_reset = reset; // @[:@16109.4]
  assign StickySelects_14_io_ins_0 = io_rPort_1_en_0 & _T_891; // @[MemPrimitives.scala 122:60:@16110.4]
  assign StickySelects_14_io_ins_1 = io_rPort_2_en_0 & _T_897; // @[MemPrimitives.scala 122:60:@16111.4]
  assign StickySelects_15_clock = clock; // @[:@16142.4]
  assign StickySelects_15_reset = reset; // @[:@16143.4]
  assign StickySelects_15_io_ins_0 = io_rPort_0_en_0 & _T_913; // @[MemPrimitives.scala 122:60:@16144.4]
  assign StickySelects_15_io_ins_1 = io_rPort_3_en_0 & _T_919; // @[MemPrimitives.scala 122:60:@16145.4]
  assign StickySelects_15_io_ins_2 = io_rPort_4_en_0 & _T_925; // @[MemPrimitives.scala 122:60:@16146.4]
  assign StickySelects_15_io_ins_3 = io_rPort_5_en_0 & _T_931; // @[MemPrimitives.scala 122:60:@16147.4]
  assign RetimeWrapper_clock = clock; // @[:@16195.4]
  assign RetimeWrapper_reset = reset; // @[:@16196.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@16198.4]
  assign RetimeWrapper_io_in = _T_465 & io_rPort_0_en_0; // @[package.scala 94:16:@16197.4]
  assign RetimeWrapper_1_clock = clock; // @[:@16203.4]
  assign RetimeWrapper_1_reset = reset; // @[:@16204.4]
  assign RetimeWrapper_1_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@16206.4]
  assign RetimeWrapper_1_io_in = _T_529 & io_rPort_0_en_0; // @[package.scala 94:16:@16205.4]
  assign RetimeWrapper_2_clock = clock; // @[:@16211.4]
  assign RetimeWrapper_2_reset = reset; // @[:@16212.4]
  assign RetimeWrapper_2_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@16214.4]
  assign RetimeWrapper_2_io_in = _T_593 & io_rPort_0_en_0; // @[package.scala 94:16:@16213.4]
  assign RetimeWrapper_3_clock = clock; // @[:@16219.4]
  assign RetimeWrapper_3_reset = reset; // @[:@16220.4]
  assign RetimeWrapper_3_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@16222.4]
  assign RetimeWrapper_3_io_in = _T_657 & io_rPort_0_en_0; // @[package.scala 94:16:@16221.4]
  assign RetimeWrapper_4_clock = clock; // @[:@16227.4]
  assign RetimeWrapper_4_reset = reset; // @[:@16228.4]
  assign RetimeWrapper_4_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@16230.4]
  assign RetimeWrapper_4_io_in = _T_721 & io_rPort_0_en_0; // @[package.scala 94:16:@16229.4]
  assign RetimeWrapper_5_clock = clock; // @[:@16235.4]
  assign RetimeWrapper_5_reset = reset; // @[:@16236.4]
  assign RetimeWrapper_5_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@16238.4]
  assign RetimeWrapper_5_io_in = _T_785 & io_rPort_0_en_0; // @[package.scala 94:16:@16237.4]
  assign RetimeWrapper_6_clock = clock; // @[:@16243.4]
  assign RetimeWrapper_6_reset = reset; // @[:@16244.4]
  assign RetimeWrapper_6_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@16246.4]
  assign RetimeWrapper_6_io_in = _T_849 & io_rPort_0_en_0; // @[package.scala 94:16:@16245.4]
  assign RetimeWrapper_7_clock = clock; // @[:@16251.4]
  assign RetimeWrapper_7_reset = reset; // @[:@16252.4]
  assign RetimeWrapper_7_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@16254.4]
  assign RetimeWrapper_7_io_in = _T_913 & io_rPort_0_en_0; // @[package.scala 94:16:@16253.4]
  assign RetimeWrapper_8_clock = clock; // @[:@16291.4]
  assign RetimeWrapper_8_reset = reset; // @[:@16292.4]
  assign RetimeWrapper_8_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@16294.4]
  assign RetimeWrapper_8_io_in = _T_443 & io_rPort_1_en_0; // @[package.scala 94:16:@16293.4]
  assign RetimeWrapper_9_clock = clock; // @[:@16299.4]
  assign RetimeWrapper_9_reset = reset; // @[:@16300.4]
  assign RetimeWrapper_9_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@16302.4]
  assign RetimeWrapper_9_io_in = _T_507 & io_rPort_1_en_0; // @[package.scala 94:16:@16301.4]
  assign RetimeWrapper_10_clock = clock; // @[:@16307.4]
  assign RetimeWrapper_10_reset = reset; // @[:@16308.4]
  assign RetimeWrapper_10_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@16310.4]
  assign RetimeWrapper_10_io_in = _T_571 & io_rPort_1_en_0; // @[package.scala 94:16:@16309.4]
  assign RetimeWrapper_11_clock = clock; // @[:@16315.4]
  assign RetimeWrapper_11_reset = reset; // @[:@16316.4]
  assign RetimeWrapper_11_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@16318.4]
  assign RetimeWrapper_11_io_in = _T_635 & io_rPort_1_en_0; // @[package.scala 94:16:@16317.4]
  assign RetimeWrapper_12_clock = clock; // @[:@16323.4]
  assign RetimeWrapper_12_reset = reset; // @[:@16324.4]
  assign RetimeWrapper_12_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@16326.4]
  assign RetimeWrapper_12_io_in = _T_699 & io_rPort_1_en_0; // @[package.scala 94:16:@16325.4]
  assign RetimeWrapper_13_clock = clock; // @[:@16331.4]
  assign RetimeWrapper_13_reset = reset; // @[:@16332.4]
  assign RetimeWrapper_13_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@16334.4]
  assign RetimeWrapper_13_io_in = _T_763 & io_rPort_1_en_0; // @[package.scala 94:16:@16333.4]
  assign RetimeWrapper_14_clock = clock; // @[:@16339.4]
  assign RetimeWrapper_14_reset = reset; // @[:@16340.4]
  assign RetimeWrapper_14_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@16342.4]
  assign RetimeWrapper_14_io_in = _T_827 & io_rPort_1_en_0; // @[package.scala 94:16:@16341.4]
  assign RetimeWrapper_15_clock = clock; // @[:@16347.4]
  assign RetimeWrapper_15_reset = reset; // @[:@16348.4]
  assign RetimeWrapper_15_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@16350.4]
  assign RetimeWrapper_15_io_in = _T_891 & io_rPort_1_en_0; // @[package.scala 94:16:@16349.4]
  assign RetimeWrapper_16_clock = clock; // @[:@16387.4]
  assign RetimeWrapper_16_reset = reset; // @[:@16388.4]
  assign RetimeWrapper_16_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@16390.4]
  assign RetimeWrapper_16_io_in = _T_449 & io_rPort_2_en_0; // @[package.scala 94:16:@16389.4]
  assign RetimeWrapper_17_clock = clock; // @[:@16395.4]
  assign RetimeWrapper_17_reset = reset; // @[:@16396.4]
  assign RetimeWrapper_17_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@16398.4]
  assign RetimeWrapper_17_io_in = _T_513 & io_rPort_2_en_0; // @[package.scala 94:16:@16397.4]
  assign RetimeWrapper_18_clock = clock; // @[:@16403.4]
  assign RetimeWrapper_18_reset = reset; // @[:@16404.4]
  assign RetimeWrapper_18_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@16406.4]
  assign RetimeWrapper_18_io_in = _T_577 & io_rPort_2_en_0; // @[package.scala 94:16:@16405.4]
  assign RetimeWrapper_19_clock = clock; // @[:@16411.4]
  assign RetimeWrapper_19_reset = reset; // @[:@16412.4]
  assign RetimeWrapper_19_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@16414.4]
  assign RetimeWrapper_19_io_in = _T_641 & io_rPort_2_en_0; // @[package.scala 94:16:@16413.4]
  assign RetimeWrapper_20_clock = clock; // @[:@16419.4]
  assign RetimeWrapper_20_reset = reset; // @[:@16420.4]
  assign RetimeWrapper_20_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@16422.4]
  assign RetimeWrapper_20_io_in = _T_705 & io_rPort_2_en_0; // @[package.scala 94:16:@16421.4]
  assign RetimeWrapper_21_clock = clock; // @[:@16427.4]
  assign RetimeWrapper_21_reset = reset; // @[:@16428.4]
  assign RetimeWrapper_21_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@16430.4]
  assign RetimeWrapper_21_io_in = _T_769 & io_rPort_2_en_0; // @[package.scala 94:16:@16429.4]
  assign RetimeWrapper_22_clock = clock; // @[:@16435.4]
  assign RetimeWrapper_22_reset = reset; // @[:@16436.4]
  assign RetimeWrapper_22_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@16438.4]
  assign RetimeWrapper_22_io_in = _T_833 & io_rPort_2_en_0; // @[package.scala 94:16:@16437.4]
  assign RetimeWrapper_23_clock = clock; // @[:@16443.4]
  assign RetimeWrapper_23_reset = reset; // @[:@16444.4]
  assign RetimeWrapper_23_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@16446.4]
  assign RetimeWrapper_23_io_in = _T_897 & io_rPort_2_en_0; // @[package.scala 94:16:@16445.4]
  assign RetimeWrapper_24_clock = clock; // @[:@16483.4]
  assign RetimeWrapper_24_reset = reset; // @[:@16484.4]
  assign RetimeWrapper_24_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@16486.4]
  assign RetimeWrapper_24_io_in = _T_471 & io_rPort_3_en_0; // @[package.scala 94:16:@16485.4]
  assign RetimeWrapper_25_clock = clock; // @[:@16491.4]
  assign RetimeWrapper_25_reset = reset; // @[:@16492.4]
  assign RetimeWrapper_25_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@16494.4]
  assign RetimeWrapper_25_io_in = _T_535 & io_rPort_3_en_0; // @[package.scala 94:16:@16493.4]
  assign RetimeWrapper_26_clock = clock; // @[:@16499.4]
  assign RetimeWrapper_26_reset = reset; // @[:@16500.4]
  assign RetimeWrapper_26_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@16502.4]
  assign RetimeWrapper_26_io_in = _T_599 & io_rPort_3_en_0; // @[package.scala 94:16:@16501.4]
  assign RetimeWrapper_27_clock = clock; // @[:@16507.4]
  assign RetimeWrapper_27_reset = reset; // @[:@16508.4]
  assign RetimeWrapper_27_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@16510.4]
  assign RetimeWrapper_27_io_in = _T_663 & io_rPort_3_en_0; // @[package.scala 94:16:@16509.4]
  assign RetimeWrapper_28_clock = clock; // @[:@16515.4]
  assign RetimeWrapper_28_reset = reset; // @[:@16516.4]
  assign RetimeWrapper_28_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@16518.4]
  assign RetimeWrapper_28_io_in = _T_727 & io_rPort_3_en_0; // @[package.scala 94:16:@16517.4]
  assign RetimeWrapper_29_clock = clock; // @[:@16523.4]
  assign RetimeWrapper_29_reset = reset; // @[:@16524.4]
  assign RetimeWrapper_29_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@16526.4]
  assign RetimeWrapper_29_io_in = _T_791 & io_rPort_3_en_0; // @[package.scala 94:16:@16525.4]
  assign RetimeWrapper_30_clock = clock; // @[:@16531.4]
  assign RetimeWrapper_30_reset = reset; // @[:@16532.4]
  assign RetimeWrapper_30_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@16534.4]
  assign RetimeWrapper_30_io_in = _T_855 & io_rPort_3_en_0; // @[package.scala 94:16:@16533.4]
  assign RetimeWrapper_31_clock = clock; // @[:@16539.4]
  assign RetimeWrapper_31_reset = reset; // @[:@16540.4]
  assign RetimeWrapper_31_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@16542.4]
  assign RetimeWrapper_31_io_in = _T_919 & io_rPort_3_en_0; // @[package.scala 94:16:@16541.4]
  assign RetimeWrapper_32_clock = clock; // @[:@16579.4]
  assign RetimeWrapper_32_reset = reset; // @[:@16580.4]
  assign RetimeWrapper_32_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@16582.4]
  assign RetimeWrapper_32_io_in = _T_477 & io_rPort_4_en_0; // @[package.scala 94:16:@16581.4]
  assign RetimeWrapper_33_clock = clock; // @[:@16587.4]
  assign RetimeWrapper_33_reset = reset; // @[:@16588.4]
  assign RetimeWrapper_33_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@16590.4]
  assign RetimeWrapper_33_io_in = _T_541 & io_rPort_4_en_0; // @[package.scala 94:16:@16589.4]
  assign RetimeWrapper_34_clock = clock; // @[:@16595.4]
  assign RetimeWrapper_34_reset = reset; // @[:@16596.4]
  assign RetimeWrapper_34_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@16598.4]
  assign RetimeWrapper_34_io_in = _T_605 & io_rPort_4_en_0; // @[package.scala 94:16:@16597.4]
  assign RetimeWrapper_35_clock = clock; // @[:@16603.4]
  assign RetimeWrapper_35_reset = reset; // @[:@16604.4]
  assign RetimeWrapper_35_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@16606.4]
  assign RetimeWrapper_35_io_in = _T_669 & io_rPort_4_en_0; // @[package.scala 94:16:@16605.4]
  assign RetimeWrapper_36_clock = clock; // @[:@16611.4]
  assign RetimeWrapper_36_reset = reset; // @[:@16612.4]
  assign RetimeWrapper_36_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@16614.4]
  assign RetimeWrapper_36_io_in = _T_733 & io_rPort_4_en_0; // @[package.scala 94:16:@16613.4]
  assign RetimeWrapper_37_clock = clock; // @[:@16619.4]
  assign RetimeWrapper_37_reset = reset; // @[:@16620.4]
  assign RetimeWrapper_37_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@16622.4]
  assign RetimeWrapper_37_io_in = _T_797 & io_rPort_4_en_0; // @[package.scala 94:16:@16621.4]
  assign RetimeWrapper_38_clock = clock; // @[:@16627.4]
  assign RetimeWrapper_38_reset = reset; // @[:@16628.4]
  assign RetimeWrapper_38_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@16630.4]
  assign RetimeWrapper_38_io_in = _T_861 & io_rPort_4_en_0; // @[package.scala 94:16:@16629.4]
  assign RetimeWrapper_39_clock = clock; // @[:@16635.4]
  assign RetimeWrapper_39_reset = reset; // @[:@16636.4]
  assign RetimeWrapper_39_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@16638.4]
  assign RetimeWrapper_39_io_in = _T_925 & io_rPort_4_en_0; // @[package.scala 94:16:@16637.4]
  assign RetimeWrapper_40_clock = clock; // @[:@16675.4]
  assign RetimeWrapper_40_reset = reset; // @[:@16676.4]
  assign RetimeWrapper_40_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@16678.4]
  assign RetimeWrapper_40_io_in = _T_483 & io_rPort_5_en_0; // @[package.scala 94:16:@16677.4]
  assign RetimeWrapper_41_clock = clock; // @[:@16683.4]
  assign RetimeWrapper_41_reset = reset; // @[:@16684.4]
  assign RetimeWrapper_41_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@16686.4]
  assign RetimeWrapper_41_io_in = _T_547 & io_rPort_5_en_0; // @[package.scala 94:16:@16685.4]
  assign RetimeWrapper_42_clock = clock; // @[:@16691.4]
  assign RetimeWrapper_42_reset = reset; // @[:@16692.4]
  assign RetimeWrapper_42_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@16694.4]
  assign RetimeWrapper_42_io_in = _T_611 & io_rPort_5_en_0; // @[package.scala 94:16:@16693.4]
  assign RetimeWrapper_43_clock = clock; // @[:@16699.4]
  assign RetimeWrapper_43_reset = reset; // @[:@16700.4]
  assign RetimeWrapper_43_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@16702.4]
  assign RetimeWrapper_43_io_in = _T_675 & io_rPort_5_en_0; // @[package.scala 94:16:@16701.4]
  assign RetimeWrapper_44_clock = clock; // @[:@16707.4]
  assign RetimeWrapper_44_reset = reset; // @[:@16708.4]
  assign RetimeWrapper_44_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@16710.4]
  assign RetimeWrapper_44_io_in = _T_739 & io_rPort_5_en_0; // @[package.scala 94:16:@16709.4]
  assign RetimeWrapper_45_clock = clock; // @[:@16715.4]
  assign RetimeWrapper_45_reset = reset; // @[:@16716.4]
  assign RetimeWrapper_45_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@16718.4]
  assign RetimeWrapper_45_io_in = _T_803 & io_rPort_5_en_0; // @[package.scala 94:16:@16717.4]
  assign RetimeWrapper_46_clock = clock; // @[:@16723.4]
  assign RetimeWrapper_46_reset = reset; // @[:@16724.4]
  assign RetimeWrapper_46_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@16726.4]
  assign RetimeWrapper_46_io_in = _T_867 & io_rPort_5_en_0; // @[package.scala 94:16:@16725.4]
  assign RetimeWrapper_47_clock = clock; // @[:@16731.4]
  assign RetimeWrapper_47_reset = reset; // @[:@16732.4]
  assign RetimeWrapper_47_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@16734.4]
  assign RetimeWrapper_47_io_in = _T_931 & io_rPort_5_en_0; // @[package.scala 94:16:@16733.4]
endmodule
module RetimeWrapper_228( // @[:@16758.2]
  input         clock, // @[:@16759.4]
  input         reset, // @[:@16760.4]
  input         io_flow, // @[:@16761.4]
  input  [15:0] io_in, // @[:@16761.4]
  output [15:0] io_out // @[:@16761.4]
);
  wire [15:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@16763.4]
  wire [15:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@16763.4]
  wire [15:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@16763.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@16763.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@16763.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@16763.4]
  RetimeShiftRegister #(.WIDTH(16), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@16763.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@16776.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@16775.4]
  assign sr_init = 16'h0; // @[RetimeShiftRegister.scala 19:16:@16774.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@16773.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@16772.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@16770.4]
endmodule
module SimBlackBoxesfix2fixBox_2( // @[:@16778.2]
  input  [31:0] io_a, // @[:@16781.4]
  output [32:0] io_b // @[:@16781.4]
);
  wire  _T_20; // @[implicits.scala 69:16:@16788.4]
  assign _T_20 = io_a[31]; // @[implicits.scala 69:16:@16788.4]
  assign io_b = {_T_20,io_a}; // @[SimBlackBoxes.scala 99:40:@16793.4]
endmodule
module __2( // @[:@16795.2]
  input  [31:0] io_b, // @[:@16798.4]
  output [32:0] io_result // @[:@16798.4]
);
  wire [31:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@16803.4]
  wire [32:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@16803.4]
  SimBlackBoxesfix2fixBox_2 SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@16803.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@16816.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@16811.4]
endmodule
module RetimeWrapper_229( // @[:@16870.2]
  input         clock, // @[:@16871.4]
  input         reset, // @[:@16872.4]
  input         io_flow, // @[:@16873.4]
  input  [31:0] io_in, // @[:@16873.4]
  output [31:0] io_out // @[:@16873.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@16875.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@16875.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@16875.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@16875.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@16875.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@16875.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@16875.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@16888.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@16887.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@16886.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@16885.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@16884.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@16882.4]
endmodule
module fix2fixBox( // @[:@16890.2]
  input         clock, // @[:@16891.4]
  input         reset, // @[:@16892.4]
  input  [32:0] io_a, // @[:@16893.4]
  input         io_flow, // @[:@16893.4]
  output [31:0] io_b // @[:@16893.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@16903.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@16903.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@16903.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@16903.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@16903.4]
  RetimeWrapper_229 RetimeWrapper ( // @[package.scala 93:22:@16903.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@16910.4]
  assign RetimeWrapper_clock = clock; // @[:@16904.4]
  assign RetimeWrapper_reset = reset; // @[:@16905.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@16907.4]
  assign RetimeWrapper_io_in = io_a[31:0]; // @[package.scala 94:16:@16906.4]
endmodule
module x303_sum( // @[:@16912.2]
  input         clock, // @[:@16913.4]
  input         reset, // @[:@16914.4]
  input  [31:0] io_a, // @[:@16915.4]
  input  [31:0] io_b, // @[:@16915.4]
  input         io_flow, // @[:@16915.4]
  output [31:0] io_result // @[:@16915.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@16923.4]
  wire [32:0] __io_result; // @[Math.scala 709:24:@16923.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@16930.4]
  wire [32:0] __1_io_result; // @[Math.scala 709:24:@16930.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@16948.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@16948.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@16948.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@16948.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@16948.4]
  wire [32:0] a_upcast_number; // @[Math.scala 712:22:@16928.4 Math.scala 713:14:@16929.4]
  wire [32:0] b_upcast_number; // @[Math.scala 712:22:@16935.4 Math.scala 713:14:@16936.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@16937.4]
  __2 _ ( // @[Math.scala 709:24:@16923.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 709:24:@16930.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox fix2fixBox ( // @[Math.scala 141:30:@16948.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@16928.4 Math.scala 713:14:@16929.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@16935.4 Math.scala 713:14:@16936.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@16937.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@16956.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@16926.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@16933.4]
  assign fix2fixBox_clock = clock; // @[:@16949.4]
  assign fix2fixBox_reset = reset; // @[:@16950.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@16951.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@16954.4]
endmodule
module RetimeWrapper_230( // @[:@16970.2]
  input         clock, // @[:@16971.4]
  input         reset, // @[:@16972.4]
  input         io_flow, // @[:@16973.4]
  input  [31:0] io_in, // @[:@16973.4]
  output [31:0] io_out // @[:@16973.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@16975.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@16975.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@16975.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@16975.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@16975.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@16975.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@16975.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@16988.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@16987.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@16986.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@16985.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@16984.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@16982.4]
endmodule
module RetimeWrapper_243( // @[:@17682.2]
  input         clock, // @[:@17683.4]
  input         reset, // @[:@17684.4]
  input         io_flow, // @[:@17685.4]
  input  [31:0] io_in, // @[:@17685.4]
  output [31:0] io_out // @[:@17685.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@17687.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@17687.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@17687.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@17687.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@17687.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@17687.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(4)) sr ( // @[RetimeShiftRegister.scala 15:20:@17687.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@17700.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@17699.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@17698.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@17697.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@17696.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@17694.4]
endmodule
module RetimeWrapper_249( // @[:@18022.2]
  input         clock, // @[:@18023.4]
  input         reset, // @[:@18024.4]
  input         io_flow, // @[:@18025.4]
  input  [31:0] io_in, // @[:@18025.4]
  output [31:0] io_out // @[:@18025.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@18027.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@18027.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@18027.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@18027.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@18027.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@18027.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(5)) sr ( // @[RetimeShiftRegister.scala 15:20:@18027.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@18040.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@18039.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@18038.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@18037.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@18036.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@18034.4]
endmodule
module RetimeWrapper_250( // @[:@18054.2]
  input   clock, // @[:@18055.4]
  input   reset, // @[:@18056.4]
  input   io_flow, // @[:@18057.4]
  input   io_in, // @[:@18057.4]
  output  io_out // @[:@18057.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@18059.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@18059.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@18059.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@18059.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@18059.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@18059.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(6)) sr ( // @[RetimeShiftRegister.scala 15:20:@18059.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@18072.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@18071.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@18070.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@18069.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@18068.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@18066.4]
endmodule
module RetimeWrapper_259( // @[:@18490.2]
  input         clock, // @[:@18491.4]
  input         reset, // @[:@18492.4]
  input         io_flow, // @[:@18493.4]
  input  [31:0] io_in, // @[:@18493.4]
  output [31:0] io_out // @[:@18493.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@18495.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@18495.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@18495.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@18495.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@18495.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@18495.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(6)) sr ( // @[RetimeShiftRegister.scala 15:20:@18495.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@18508.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@18507.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@18506.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@18505.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@18504.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@18502.4]
endmodule
module x364_rdrow( // @[:@19620.2]
  input         clock, // @[:@19621.4]
  input         reset, // @[:@19622.4]
  input  [31:0] io_a, // @[:@19623.4]
  input  [31:0] io_b, // @[:@19623.4]
  input         io_flow, // @[:@19623.4]
  output [31:0] io_result // @[:@19623.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@19631.4]
  wire [32:0] __io_result; // @[Math.scala 709:24:@19631.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@19638.4]
  wire [32:0] __1_io_result; // @[Math.scala 709:24:@19638.4]
  wire  fix2fixBox_clock; // @[Math.scala 182:30:@19657.4]
  wire  fix2fixBox_reset; // @[Math.scala 182:30:@19657.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 182:30:@19657.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 182:30:@19657.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 182:30:@19657.4]
  wire [32:0] a_upcast_number; // @[Math.scala 712:22:@19636.4 Math.scala 713:14:@19637.4]
  wire [32:0] b_upcast_number; // @[Math.scala 712:22:@19643.4 Math.scala 713:14:@19644.4]
  wire [33:0] _T_21; // @[Math.scala 177:37:@19645.4]
  wire [33:0] _T_22; // @[Math.scala 177:37:@19646.4]
  __2 _ ( // @[Math.scala 709:24:@19631.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 709:24:@19638.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox fix2fixBox ( // @[Math.scala 182:30:@19657.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@19636.4 Math.scala 713:14:@19637.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@19643.4 Math.scala 713:14:@19644.4]
  assign _T_21 = a_upcast_number - b_upcast_number; // @[Math.scala 177:37:@19645.4]
  assign _T_22 = $unsigned(_T_21); // @[Math.scala 177:37:@19646.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 188:17:@19665.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@19634.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@19641.4]
  assign fix2fixBox_clock = clock; // @[:@19658.4]
  assign fix2fixBox_reset = reset; // @[:@19659.4]
  assign fix2fixBox_io_a = _T_22[32:0]; // @[Math.scala 183:23:@19660.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 186:26:@19663.4]
endmodule
module SimBlackBoxesfix2fixBox_40( // @[:@21928.2]
  input  [7:0] io_a, // @[:@21931.4]
  output [8:0] io_b // @[:@21931.4]
);
  assign io_b = {1'h0,io_a}; // @[SimBlackBoxes.scala 99:40:@21942.4]
endmodule
module __40( // @[:@21944.2]
  input  [7:0] io_b, // @[:@21947.4]
  output [8:0] io_result // @[:@21947.4]
);
  wire [7:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@21952.4]
  wire [8:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@21952.4]
  SimBlackBoxesfix2fixBox_40 SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@21952.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@21965.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@21960.4]
endmodule
module fix2fixBox_19( // @[:@22038.2]
  input        clock, // @[:@22039.4]
  input        reset, // @[:@22040.4]
  input  [8:0] io_a, // @[:@22041.4]
  input        io_flow, // @[:@22041.4]
  output [7:0] io_b // @[:@22041.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@22051.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@22051.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@22051.4]
  wire [7:0] RetimeWrapper_io_in; // @[package.scala 93:22:@22051.4]
  wire [7:0] RetimeWrapper_io_out; // @[package.scala 93:22:@22051.4]
  RetimeWrapper_21 RetimeWrapper ( // @[package.scala 93:22:@22051.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@22058.4]
  assign RetimeWrapper_clock = clock; // @[:@22052.4]
  assign RetimeWrapper_reset = reset; // @[:@22053.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@22055.4]
  assign RetimeWrapper_io_in = io_a[7:0]; // @[package.scala 94:16:@22054.4]
endmodule
module x437_x23( // @[:@22060.2]
  input        clock, // @[:@22061.4]
  input        reset, // @[:@22062.4]
  input  [7:0] io_a, // @[:@22063.4]
  input  [7:0] io_b, // @[:@22063.4]
  input        io_flow, // @[:@22063.4]
  output [7:0] io_result // @[:@22063.4]
);
  wire [7:0] __io_b; // @[Math.scala 709:24:@22071.4]
  wire [8:0] __io_result; // @[Math.scala 709:24:@22071.4]
  wire [7:0] __1_io_b; // @[Math.scala 709:24:@22078.4]
  wire [8:0] __1_io_result; // @[Math.scala 709:24:@22078.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@22088.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@22088.4]
  wire [8:0] fix2fixBox_io_a; // @[Math.scala 141:30:@22088.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@22088.4]
  wire [7:0] fix2fixBox_io_b; // @[Math.scala 141:30:@22088.4]
  wire [8:0] a_upcast_number; // @[Math.scala 712:22:@22076.4 Math.scala 713:14:@22077.4]
  wire [8:0] b_upcast_number; // @[Math.scala 712:22:@22083.4 Math.scala 713:14:@22084.4]
  wire [9:0] _T_21; // @[Math.scala 136:37:@22085.4]
  __40 _ ( // @[Math.scala 709:24:@22071.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __40 __1 ( // @[Math.scala 709:24:@22078.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_19 fix2fixBox ( // @[Math.scala 141:30:@22088.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@22076.4 Math.scala 713:14:@22077.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@22083.4 Math.scala 713:14:@22084.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@22085.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@22096.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@22074.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@22081.4]
  assign fix2fixBox_clock = clock; // @[:@22089.4]
  assign fix2fixBox_reset = reset; // @[:@22090.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@22091.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@22094.4]
endmodule
module fix2fixBox_23( // @[:@22686.2]
  input  [8:0] io_a, // @[:@22689.4]
  output [7:0] io_b // @[:@22689.4]
);
  assign io_b = io_a[7:0]; // @[Converter.scala 95:38:@22699.4]
endmodule
module x441_x23( // @[:@22701.2]
  input  [7:0] io_a, // @[:@22704.4]
  input  [7:0] io_b, // @[:@22704.4]
  output [7:0] io_result // @[:@22704.4]
);
  wire [7:0] __io_b; // @[Math.scala 709:24:@22712.4]
  wire [8:0] __io_result; // @[Math.scala 709:24:@22712.4]
  wire [7:0] __1_io_b; // @[Math.scala 709:24:@22719.4]
  wire [8:0] __1_io_result; // @[Math.scala 709:24:@22719.4]
  wire [8:0] fix2fixBox_io_a; // @[Math.scala 141:30:@22729.4]
  wire [7:0] fix2fixBox_io_b; // @[Math.scala 141:30:@22729.4]
  wire [8:0] a_upcast_number; // @[Math.scala 712:22:@22717.4 Math.scala 713:14:@22718.4]
  wire [8:0] b_upcast_number; // @[Math.scala 712:22:@22724.4 Math.scala 713:14:@22725.4]
  wire [9:0] _T_21; // @[Math.scala 136:37:@22726.4]
  __40 _ ( // @[Math.scala 709:24:@22712.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __40 __1 ( // @[Math.scala 709:24:@22719.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_23 fix2fixBox ( // @[Math.scala 141:30:@22729.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@22717.4 Math.scala 713:14:@22718.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@22724.4 Math.scala 713:14:@22725.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@22726.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@22737.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@22715.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@22722.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@22732.4]
endmodule
module RetimeWrapper_314( // @[:@24476.2]
  input         clock, // @[:@24477.4]
  input         reset, // @[:@24478.4]
  input         io_flow, // @[:@24479.4]
  input  [31:0] io_in, // @[:@24479.4]
  output [31:0] io_out // @[:@24479.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@24481.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@24481.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@24481.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@24481.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@24481.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@24481.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(10)) sr ( // @[RetimeShiftRegister.scala 15:20:@24481.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@24494.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@24493.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@24492.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@24491.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@24490.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@24488.4]
endmodule
module RetimeWrapper_315( // @[:@24508.2]
  input   clock, // @[:@24509.4]
  input   reset, // @[:@24510.4]
  input   io_flow, // @[:@24511.4]
  input   io_in, // @[:@24511.4]
  output  io_out // @[:@24511.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@24513.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@24513.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@24513.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@24513.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@24513.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@24513.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(10)) sr ( // @[RetimeShiftRegister.scala 15:20:@24513.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@24526.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@24525.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@24524.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@24523.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@24522.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@24520.4]
endmodule
module RetimeWrapper_316( // @[:@24540.2]
  input         clock, // @[:@24541.4]
  input         reset, // @[:@24542.4]
  input         io_flow, // @[:@24543.4]
  input  [31:0] io_in, // @[:@24543.4]
  output [31:0] io_out // @[:@24543.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@24545.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@24545.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@24545.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@24545.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@24545.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@24545.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(9)) sr ( // @[RetimeShiftRegister.scala 15:20:@24545.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@24558.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@24557.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@24556.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@24555.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@24554.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@24552.4]
endmodule
module RetimeWrapper_321( // @[:@24700.2]
  input         clock, // @[:@24701.4]
  input         reset, // @[:@24702.4]
  input         io_flow, // @[:@24703.4]
  input  [31:0] io_in, // @[:@24703.4]
  output [31:0] io_out // @[:@24703.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@24705.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@24705.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@24705.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@24705.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@24705.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@24705.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(8)) sr ( // @[RetimeShiftRegister.scala 15:20:@24705.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@24718.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@24717.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@24716.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@24715.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@24714.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@24712.4]
endmodule
module RetimeWrapper_323( // @[:@24764.2]
  input   clock, // @[:@24765.4]
  input   reset, // @[:@24766.4]
  input   io_flow, // @[:@24767.4]
  input   io_in, // @[:@24767.4]
  output  io_out // @[:@24767.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@24769.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@24769.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@24769.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@24769.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@24769.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@24769.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(5)) sr ( // @[RetimeShiftRegister.scala 15:20:@24769.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@24782.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@24781.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@24780.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@24779.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@24778.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@24776.4]
endmodule
module RetimeWrapper_344( // @[:@25829.2]
  input        clock, // @[:@25830.4]
  input        reset, // @[:@25831.4]
  input        io_flow, // @[:@25832.4]
  input  [7:0] io_in, // @[:@25832.4]
  output [7:0] io_out // @[:@25832.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@25834.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@25834.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@25834.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@25834.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@25834.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@25834.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(5)) sr ( // @[RetimeShiftRegister.scala 15:20:@25834.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@25847.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@25846.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@25845.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@25844.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@25843.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@25841.4]
endmodule
module SimBlackBoxesfix2fixBox_78( // @[:@25849.2]
  input  [7:0] io_a, // @[:@25852.4]
  output [7:0] io_b // @[:@25852.4]
);
  assign io_b = io_a; // @[SimBlackBoxes.scala 99:40:@25862.4]
endmodule
module __78( // @[:@25864.2]
  input  [7:0] io_b, // @[:@25867.4]
  output [7:0] io_result // @[:@25867.4]
);
  wire [7:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@25872.4]
  wire [7:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@25872.4]
  SimBlackBoxesfix2fixBox_78 SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@25872.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@25885.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@25880.4]
endmodule
module x481_div( // @[:@25887.2]
  input        clock, // @[:@25888.4]
  input        reset, // @[:@25889.4]
  input  [7:0] io_a, // @[:@25890.4]
  input        io_flow, // @[:@25890.4]
  output [7:0] io_result // @[:@25890.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@25897.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@25897.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@25897.4]
  wire [7:0] RetimeWrapper_io_in; // @[package.scala 93:22:@25897.4]
  wire [7:0] RetimeWrapper_io_out; // @[package.scala 93:22:@25897.4]
  wire [7:0] __io_b; // @[Math.scala 709:24:@25907.4]
  wire [7:0] __io_result; // @[Math.scala 709:24:@25907.4]
  RetimeWrapper_344 RetimeWrapper ( // @[package.scala 93:22:@25897.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  __78 _ ( // @[Math.scala 709:24:@25907.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  assign io_result = __io_result; // @[Math.scala 291:34:@25915.4]
  assign RetimeWrapper_clock = clock; // @[:@25898.4]
  assign RetimeWrapper_reset = reset; // @[:@25899.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@25901.4]
  assign RetimeWrapper_io_in = io_a / 8'h6; // @[package.scala 94:16:@25900.4]
  assign __io_b = RetimeWrapper_io_out; // @[Math.scala 710:17:@25910.4]
endmodule
module RetimeWrapper_346( // @[:@26422.2]
  input         clock, // @[:@26423.4]
  input         reset, // @[:@26424.4]
  input         io_flow, // @[:@26425.4]
  input  [15:0] io_in, // @[:@26425.4]
  output [15:0] io_out // @[:@26425.4]
);
  wire [15:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@26427.4]
  wire [15:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@26427.4]
  wire [15:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@26427.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@26427.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@26427.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@26427.4]
  RetimeShiftRegister #(.WIDTH(16), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@26427.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@26440.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@26439.4]
  assign sr_init = 16'h0; // @[RetimeShiftRegister.scala 19:16:@26438.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@26437.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@26436.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@26434.4]
endmodule
module RetimeWrapper_347( // @[:@26454.2]
  input   clock, // @[:@26455.4]
  input   reset, // @[:@26456.4]
  input   io_flow, // @[:@26457.4]
  input   io_in, // @[:@26457.4]
  output  io_out // @[:@26457.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@26459.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@26459.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@26459.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@26459.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@26459.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@26459.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(20)) sr ( // @[RetimeShiftRegister.scala 15:20:@26459.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@26472.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@26471.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@26470.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@26469.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@26468.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@26466.4]
endmodule
module x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1( // @[:@26538.2]
  input          clock, // @[:@26539.4]
  input          reset, // @[:@26540.4]
  output         io_in_x276_TVALID, // @[:@26541.4]
  input          io_in_x276_TREADY, // @[:@26541.4]
  output [255:0] io_in_x276_TDATA, // @[:@26541.4]
  output         io_in_x275_TREADY, // @[:@26541.4]
  input  [255:0] io_in_x275_TDATA, // @[:@26541.4]
  input  [7:0]   io_in_x275_TID, // @[:@26541.4]
  input  [7:0]   io_in_x275_TDEST, // @[:@26541.4]
  input          io_sigsIn_backpressure, // @[:@26541.4]
  input          io_sigsIn_datapathEn, // @[:@26541.4]
  input          io_sigsIn_break, // @[:@26541.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_1, // @[:@26541.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_0, // @[:@26541.4]
  input          io_sigsIn_cchainOutputs_0_oobs_0, // @[:@26541.4]
  input          io_sigsIn_cchainOutputs_0_oobs_1, // @[:@26541.4]
  input          io_rr // @[:@26541.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@26555.4]
  wire [31:0] __io_result; // @[Math.scala 709:24:@26555.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@26567.4]
  wire [31:0] __1_io_result; // @[Math.scala 709:24:@26567.4]
  wire  x288_lb_0_clock; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire  x288_lb_0_reset; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire [2:0] x288_lb_0_io_rPort_11_banks_1; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire [2:0] x288_lb_0_io_rPort_11_banks_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire  x288_lb_0_io_rPort_11_ofs_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire  x288_lb_0_io_rPort_11_en_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire  x288_lb_0_io_rPort_11_backpressure; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire [7:0] x288_lb_0_io_rPort_11_output_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire [2:0] x288_lb_0_io_rPort_10_banks_1; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire [2:0] x288_lb_0_io_rPort_10_banks_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire  x288_lb_0_io_rPort_10_ofs_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire  x288_lb_0_io_rPort_10_en_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire  x288_lb_0_io_rPort_10_backpressure; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire [7:0] x288_lb_0_io_rPort_10_output_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire [2:0] x288_lb_0_io_rPort_9_banks_1; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire [2:0] x288_lb_0_io_rPort_9_banks_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire  x288_lb_0_io_rPort_9_ofs_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire  x288_lb_0_io_rPort_9_en_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire  x288_lb_0_io_rPort_9_backpressure; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire [7:0] x288_lb_0_io_rPort_9_output_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire [2:0] x288_lb_0_io_rPort_8_banks_1; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire [2:0] x288_lb_0_io_rPort_8_banks_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire  x288_lb_0_io_rPort_8_ofs_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire  x288_lb_0_io_rPort_8_en_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire  x288_lb_0_io_rPort_8_backpressure; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire [7:0] x288_lb_0_io_rPort_8_output_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire [2:0] x288_lb_0_io_rPort_7_banks_1; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire [2:0] x288_lb_0_io_rPort_7_banks_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire  x288_lb_0_io_rPort_7_ofs_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire  x288_lb_0_io_rPort_7_en_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire  x288_lb_0_io_rPort_7_backpressure; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire [7:0] x288_lb_0_io_rPort_7_output_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire [2:0] x288_lb_0_io_rPort_6_banks_1; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire [2:0] x288_lb_0_io_rPort_6_banks_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire  x288_lb_0_io_rPort_6_ofs_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire  x288_lb_0_io_rPort_6_en_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire  x288_lb_0_io_rPort_6_backpressure; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire [7:0] x288_lb_0_io_rPort_6_output_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire [2:0] x288_lb_0_io_rPort_5_banks_1; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire [2:0] x288_lb_0_io_rPort_5_banks_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire  x288_lb_0_io_rPort_5_ofs_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire  x288_lb_0_io_rPort_5_en_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire  x288_lb_0_io_rPort_5_backpressure; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire [7:0] x288_lb_0_io_rPort_5_output_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire [2:0] x288_lb_0_io_rPort_4_banks_1; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire [2:0] x288_lb_0_io_rPort_4_banks_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire  x288_lb_0_io_rPort_4_ofs_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire  x288_lb_0_io_rPort_4_en_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire  x288_lb_0_io_rPort_4_backpressure; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire [7:0] x288_lb_0_io_rPort_4_output_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire [2:0] x288_lb_0_io_rPort_3_banks_1; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire [2:0] x288_lb_0_io_rPort_3_banks_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire  x288_lb_0_io_rPort_3_ofs_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire  x288_lb_0_io_rPort_3_en_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire  x288_lb_0_io_rPort_3_backpressure; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire [7:0] x288_lb_0_io_rPort_3_output_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire [2:0] x288_lb_0_io_rPort_2_banks_1; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire [2:0] x288_lb_0_io_rPort_2_banks_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire  x288_lb_0_io_rPort_2_ofs_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire  x288_lb_0_io_rPort_2_en_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire  x288_lb_0_io_rPort_2_backpressure; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire [7:0] x288_lb_0_io_rPort_2_output_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire [2:0] x288_lb_0_io_rPort_1_banks_1; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire [2:0] x288_lb_0_io_rPort_1_banks_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire  x288_lb_0_io_rPort_1_ofs_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire  x288_lb_0_io_rPort_1_en_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire  x288_lb_0_io_rPort_1_backpressure; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire [7:0] x288_lb_0_io_rPort_1_output_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire [2:0] x288_lb_0_io_rPort_0_banks_1; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire [2:0] x288_lb_0_io_rPort_0_banks_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire  x288_lb_0_io_rPort_0_ofs_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire  x288_lb_0_io_rPort_0_en_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire  x288_lb_0_io_rPort_0_backpressure; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire [7:0] x288_lb_0_io_rPort_0_output_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire [2:0] x288_lb_0_io_wPort_1_banks_1; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire [2:0] x288_lb_0_io_wPort_1_banks_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire  x288_lb_0_io_wPort_1_ofs_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire [7:0] x288_lb_0_io_wPort_1_data_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire  x288_lb_0_io_wPort_1_en_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire [2:0] x288_lb_0_io_wPort_0_banks_1; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire [2:0] x288_lb_0_io_wPort_0_banks_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire  x288_lb_0_io_wPort_0_ofs_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire [7:0] x288_lb_0_io_wPort_0_data_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire  x288_lb_0_io_wPort_0_en_0; // @[m_x288_lb_0.scala 39:17:@26577.4]
  wire  x289_lb2_0_clock; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire  x289_lb2_0_reset; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire [2:0] x289_lb2_0_io_rPort_5_banks_1; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire [2:0] x289_lb2_0_io_rPort_5_banks_0; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire  x289_lb2_0_io_rPort_5_ofs_0; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire  x289_lb2_0_io_rPort_5_en_0; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire  x289_lb2_0_io_rPort_5_backpressure; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire [7:0] x289_lb2_0_io_rPort_5_output_0; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire [2:0] x289_lb2_0_io_rPort_4_banks_1; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire [2:0] x289_lb2_0_io_rPort_4_banks_0; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire  x289_lb2_0_io_rPort_4_ofs_0; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire  x289_lb2_0_io_rPort_4_en_0; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire  x289_lb2_0_io_rPort_4_backpressure; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire [7:0] x289_lb2_0_io_rPort_4_output_0; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire [2:0] x289_lb2_0_io_rPort_3_banks_1; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire [2:0] x289_lb2_0_io_rPort_3_banks_0; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire  x289_lb2_0_io_rPort_3_ofs_0; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire  x289_lb2_0_io_rPort_3_en_0; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire  x289_lb2_0_io_rPort_3_backpressure; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire [7:0] x289_lb2_0_io_rPort_3_output_0; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire [2:0] x289_lb2_0_io_rPort_2_banks_1; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire [2:0] x289_lb2_0_io_rPort_2_banks_0; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire  x289_lb2_0_io_rPort_2_ofs_0; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire  x289_lb2_0_io_rPort_2_en_0; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire  x289_lb2_0_io_rPort_2_backpressure; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire [7:0] x289_lb2_0_io_rPort_2_output_0; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire [2:0] x289_lb2_0_io_rPort_1_banks_1; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire [2:0] x289_lb2_0_io_rPort_1_banks_0; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire  x289_lb2_0_io_rPort_1_ofs_0; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire  x289_lb2_0_io_rPort_1_en_0; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire  x289_lb2_0_io_rPort_1_backpressure; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire [7:0] x289_lb2_0_io_rPort_1_output_0; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire [2:0] x289_lb2_0_io_rPort_0_banks_1; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire [2:0] x289_lb2_0_io_rPort_0_banks_0; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire  x289_lb2_0_io_rPort_0_ofs_0; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire  x289_lb2_0_io_rPort_0_en_0; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire  x289_lb2_0_io_rPort_0_backpressure; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire [7:0] x289_lb2_0_io_rPort_0_output_0; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire [2:0] x289_lb2_0_io_wPort_1_banks_1; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire [2:0] x289_lb2_0_io_wPort_1_banks_0; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire  x289_lb2_0_io_wPort_1_ofs_0; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire [7:0] x289_lb2_0_io_wPort_1_data_0; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire  x289_lb2_0_io_wPort_1_en_0; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire [2:0] x289_lb2_0_io_wPort_0_banks_1; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire [2:0] x289_lb2_0_io_wPort_0_banks_0; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire  x289_lb2_0_io_wPort_0_ofs_0; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire [7:0] x289_lb2_0_io_wPort_0_data_0; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire  x289_lb2_0_io_wPort_0_en_0; // @[m_x289_lb2_0.scala 33:17:@26670.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@26740.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@26740.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@26740.4]
  wire [15:0] RetimeWrapper_io_in; // @[package.scala 93:22:@26740.4]
  wire [15:0] RetimeWrapper_io_out; // @[package.scala 93:22:@26740.4]
  wire  x303_sum_1_clock; // @[Math.scala 150:24:@26847.4]
  wire  x303_sum_1_reset; // @[Math.scala 150:24:@26847.4]
  wire [31:0] x303_sum_1_io_a; // @[Math.scala 150:24:@26847.4]
  wire [31:0] x303_sum_1_io_b; // @[Math.scala 150:24:@26847.4]
  wire  x303_sum_1_io_flow; // @[Math.scala 150:24:@26847.4]
  wire [31:0] x303_sum_1_io_result; // @[Math.scala 150:24:@26847.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@26857.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@26857.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@26857.4]
  wire [31:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@26857.4]
  wire [31:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@26857.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@26866.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@26866.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@26866.4]
  wire [7:0] RetimeWrapper_2_io_in; // @[package.scala 93:22:@26866.4]
  wire [7:0] RetimeWrapper_2_io_out; // @[package.scala 93:22:@26866.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@26875.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@26875.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@26875.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@26875.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@26875.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@26884.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@26884.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@26884.4]
  wire [31:0] RetimeWrapper_4_io_in; // @[package.scala 93:22:@26884.4]
  wire [31:0] RetimeWrapper_4_io_out; // @[package.scala 93:22:@26884.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@26893.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@26893.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@26893.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@26893.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@26893.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@26902.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@26902.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@26902.4]
  wire [31:0] RetimeWrapper_6_io_in; // @[package.scala 93:22:@26902.4]
  wire [31:0] RetimeWrapper_6_io_out; // @[package.scala 93:22:@26902.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@26913.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@26913.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@26913.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@26913.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@26913.4]
  wire  x309_rdcol_1_clock; // @[Math.scala 150:24:@26936.4]
  wire  x309_rdcol_1_reset; // @[Math.scala 150:24:@26936.4]
  wire [31:0] x309_rdcol_1_io_a; // @[Math.scala 150:24:@26936.4]
  wire [31:0] x309_rdcol_1_io_b; // @[Math.scala 150:24:@26936.4]
  wire  x309_rdcol_1_io_flow; // @[Math.scala 150:24:@26936.4]
  wire [31:0] x309_rdcol_1_io_result; // @[Math.scala 150:24:@26936.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@26968.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@26968.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@26968.4]
  wire [31:0] RetimeWrapper_8_io_in; // @[package.scala 93:22:@26968.4]
  wire [31:0] RetimeWrapper_8_io_out; // @[package.scala 93:22:@26968.4]
  wire  x313_sum_1_clock; // @[Math.scala 150:24:@26977.4]
  wire  x313_sum_1_reset; // @[Math.scala 150:24:@26977.4]
  wire [31:0] x313_sum_1_io_a; // @[Math.scala 150:24:@26977.4]
  wire [31:0] x313_sum_1_io_b; // @[Math.scala 150:24:@26977.4]
  wire  x313_sum_1_io_flow; // @[Math.scala 150:24:@26977.4]
  wire [31:0] x313_sum_1_io_result; // @[Math.scala 150:24:@26977.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@26987.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@26987.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@26987.4]
  wire [31:0] RetimeWrapper_9_io_in; // @[package.scala 93:22:@26987.4]
  wire [31:0] RetimeWrapper_9_io_out; // @[package.scala 93:22:@26987.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@26996.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@26996.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@26996.4]
  wire [7:0] RetimeWrapper_10_io_in; // @[package.scala 93:22:@26996.4]
  wire [7:0] RetimeWrapper_10_io_out; // @[package.scala 93:22:@26996.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@27007.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@27007.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@27007.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@27007.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@27007.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@27028.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@27028.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@27028.4]
  wire [31:0] RetimeWrapper_12_io_in; // @[package.scala 93:22:@27028.4]
  wire [31:0] RetimeWrapper_12_io_out; // @[package.scala 93:22:@27028.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@27055.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@27055.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@27055.4]
  wire [31:0] RetimeWrapper_13_io_in; // @[package.scala 93:22:@27055.4]
  wire [31:0] RetimeWrapper_13_io_out; // @[package.scala 93:22:@27055.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@27071.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@27071.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@27071.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@27071.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@27071.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@27106.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@27106.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@27106.4]
  wire [31:0] RetimeWrapper_15_io_in; // @[package.scala 93:22:@27106.4]
  wire [31:0] RetimeWrapper_15_io_out; // @[package.scala 93:22:@27106.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@27115.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@27115.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@27115.4]
  wire [31:0] RetimeWrapper_16_io_in; // @[package.scala 93:22:@27115.4]
  wire [31:0] RetimeWrapper_16_io_out; // @[package.scala 93:22:@27115.4]
  wire  x326_sum_1_clock; // @[Math.scala 150:24:@27124.4]
  wire  x326_sum_1_reset; // @[Math.scala 150:24:@27124.4]
  wire [31:0] x326_sum_1_io_a; // @[Math.scala 150:24:@27124.4]
  wire [31:0] x326_sum_1_io_b; // @[Math.scala 150:24:@27124.4]
  wire  x326_sum_1_io_flow; // @[Math.scala 150:24:@27124.4]
  wire [31:0] x326_sum_1_io_result; // @[Math.scala 150:24:@27124.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@27134.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@27134.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@27134.4]
  wire [31:0] RetimeWrapper_17_io_in; // @[package.scala 93:22:@27134.4]
  wire [31:0] RetimeWrapper_17_io_out; // @[package.scala 93:22:@27134.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@27143.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@27143.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@27143.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@27143.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@27143.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@27152.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@27152.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@27152.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@27152.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@27152.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@27161.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@27161.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@27161.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@27161.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@27161.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@27170.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@27170.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@27170.4]
  wire [31:0] RetimeWrapper_21_io_in; // @[package.scala 93:22:@27170.4]
  wire [31:0] RetimeWrapper_21_io_out; // @[package.scala 93:22:@27170.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@27182.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@27182.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@27182.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@27182.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@27182.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@27203.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@27203.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@27203.4]
  wire [31:0] RetimeWrapper_23_io_in; // @[package.scala 93:22:@27203.4]
  wire [31:0] RetimeWrapper_23_io_out; // @[package.scala 93:22:@27203.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@27227.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@27227.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@27227.4]
  wire [31:0] RetimeWrapper_24_io_in; // @[package.scala 93:22:@27227.4]
  wire [31:0] RetimeWrapper_24_io_out; // @[package.scala 93:22:@27227.4]
  wire  x335_sum_1_clock; // @[Math.scala 150:24:@27236.4]
  wire  x335_sum_1_reset; // @[Math.scala 150:24:@27236.4]
  wire [31:0] x335_sum_1_io_a; // @[Math.scala 150:24:@27236.4]
  wire [31:0] x335_sum_1_io_b; // @[Math.scala 150:24:@27236.4]
  wire  x335_sum_1_io_flow; // @[Math.scala 150:24:@27236.4]
  wire [31:0] x335_sum_1_io_result; // @[Math.scala 150:24:@27236.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@27246.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@27246.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@27246.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@27246.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@27246.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@27255.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@27255.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@27255.4]
  wire [31:0] RetimeWrapper_26_io_in; // @[package.scala 93:22:@27255.4]
  wire [31:0] RetimeWrapper_26_io_out; // @[package.scala 93:22:@27255.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@27264.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@27264.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@27264.4]
  wire [31:0] RetimeWrapper_27_io_in; // @[package.scala 93:22:@27264.4]
  wire [31:0] RetimeWrapper_27_io_out; // @[package.scala 93:22:@27264.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@27276.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@27276.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@27276.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@27276.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@27276.4]
  wire  x340_rdcol_1_clock; // @[Math.scala 150:24:@27299.4]
  wire  x340_rdcol_1_reset; // @[Math.scala 150:24:@27299.4]
  wire [31:0] x340_rdcol_1_io_a; // @[Math.scala 150:24:@27299.4]
  wire [31:0] x340_rdcol_1_io_b; // @[Math.scala 150:24:@27299.4]
  wire  x340_rdcol_1_io_flow; // @[Math.scala 150:24:@27299.4]
  wire [31:0] x340_rdcol_1_io_result; // @[Math.scala 150:24:@27299.4]
  wire  x346_sum_1_clock; // @[Math.scala 150:24:@27342.4]
  wire  x346_sum_1_reset; // @[Math.scala 150:24:@27342.4]
  wire [31:0] x346_sum_1_io_a; // @[Math.scala 150:24:@27342.4]
  wire [31:0] x346_sum_1_io_b; // @[Math.scala 150:24:@27342.4]
  wire  x346_sum_1_io_flow; // @[Math.scala 150:24:@27342.4]
  wire [31:0] x346_sum_1_io_result; // @[Math.scala 150:24:@27342.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@27352.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@27352.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@27352.4]
  wire [31:0] RetimeWrapper_29_io_in; // @[package.scala 93:22:@27352.4]
  wire [31:0] RetimeWrapper_29_io_out; // @[package.scala 93:22:@27352.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@27361.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@27361.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@27361.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@27361.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@27361.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@27373.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@27373.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@27373.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@27373.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@27373.4]
  wire  x352_rdcol_1_clock; // @[Math.scala 150:24:@27396.4]
  wire  x352_rdcol_1_reset; // @[Math.scala 150:24:@27396.4]
  wire [31:0] x352_rdcol_1_io_a; // @[Math.scala 150:24:@27396.4]
  wire [31:0] x352_rdcol_1_io_b; // @[Math.scala 150:24:@27396.4]
  wire  x352_rdcol_1_io_flow; // @[Math.scala 150:24:@27396.4]
  wire [31:0] x352_rdcol_1_io_result; // @[Math.scala 150:24:@27396.4]
  wire  x358_sum_1_clock; // @[Math.scala 150:24:@27439.4]
  wire  x358_sum_1_reset; // @[Math.scala 150:24:@27439.4]
  wire [31:0] x358_sum_1_io_a; // @[Math.scala 150:24:@27439.4]
  wire [31:0] x358_sum_1_io_b; // @[Math.scala 150:24:@27439.4]
  wire  x358_sum_1_io_flow; // @[Math.scala 150:24:@27439.4]
  wire [31:0] x358_sum_1_io_result; // @[Math.scala 150:24:@27439.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@27449.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@27449.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@27449.4]
  wire [31:0] RetimeWrapper_32_io_in; // @[package.scala 93:22:@27449.4]
  wire [31:0] RetimeWrapper_32_io_out; // @[package.scala 93:22:@27449.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@27458.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@27458.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@27458.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@27458.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@27458.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@27470.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@27470.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@27470.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@27470.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@27470.4]
  wire  x364_rdrow_1_clock; // @[Math.scala 191:24:@27493.4]
  wire  x364_rdrow_1_reset; // @[Math.scala 191:24:@27493.4]
  wire [31:0] x364_rdrow_1_io_a; // @[Math.scala 191:24:@27493.4]
  wire [31:0] x364_rdrow_1_io_b; // @[Math.scala 191:24:@27493.4]
  wire  x364_rdrow_1_io_flow; // @[Math.scala 191:24:@27493.4]
  wire [31:0] x364_rdrow_1_io_result; // @[Math.scala 191:24:@27493.4]
  wire  x371_sum_1_clock; // @[Math.scala 150:24:@27547.4]
  wire  x371_sum_1_reset; // @[Math.scala 150:24:@27547.4]
  wire [31:0] x371_sum_1_io_a; // @[Math.scala 150:24:@27547.4]
  wire [31:0] x371_sum_1_io_b; // @[Math.scala 150:24:@27547.4]
  wire  x371_sum_1_io_flow; // @[Math.scala 150:24:@27547.4]
  wire [31:0] x371_sum_1_io_result; // @[Math.scala 150:24:@27547.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@27557.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@27557.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@27557.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@27557.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@27557.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@27566.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@27566.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@27566.4]
  wire [31:0] RetimeWrapper_36_io_in; // @[package.scala 93:22:@27566.4]
  wire [31:0] RetimeWrapper_36_io_out; // @[package.scala 93:22:@27566.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@27578.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@27578.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@27578.4]
  wire  RetimeWrapper_37_io_in; // @[package.scala 93:22:@27578.4]
  wire  RetimeWrapper_37_io_out; // @[package.scala 93:22:@27578.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@27599.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@27599.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@27599.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@27599.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@27599.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@27614.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@27614.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@27614.4]
  wire [31:0] RetimeWrapper_39_io_in; // @[package.scala 93:22:@27614.4]
  wire [31:0] RetimeWrapper_39_io_out; // @[package.scala 93:22:@27614.4]
  wire  x379_sum_1_clock; // @[Math.scala 150:24:@27625.4]
  wire  x379_sum_1_reset; // @[Math.scala 150:24:@27625.4]
  wire [31:0] x379_sum_1_io_a; // @[Math.scala 150:24:@27625.4]
  wire [31:0] x379_sum_1_io_b; // @[Math.scala 150:24:@27625.4]
  wire  x379_sum_1_io_flow; // @[Math.scala 150:24:@27625.4]
  wire [31:0] x379_sum_1_io_result; // @[Math.scala 150:24:@27625.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@27635.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@27635.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@27635.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@27635.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@27635.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@27647.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@27647.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@27647.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@27647.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@27647.4]
  wire  x386_sum_1_clock; // @[Math.scala 150:24:@27674.4]
  wire  x386_sum_1_reset; // @[Math.scala 150:24:@27674.4]
  wire [31:0] x386_sum_1_io_a; // @[Math.scala 150:24:@27674.4]
  wire [31:0] x386_sum_1_io_b; // @[Math.scala 150:24:@27674.4]
  wire  x386_sum_1_io_flow; // @[Math.scala 150:24:@27674.4]
  wire [31:0] x386_sum_1_io_result; // @[Math.scala 150:24:@27674.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@27684.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@27684.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@27684.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@27684.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@27684.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@27696.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@27696.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@27696.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@27696.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@27696.4]
  wire  x393_sum_1_clock; // @[Math.scala 150:24:@27723.4]
  wire  x393_sum_1_reset; // @[Math.scala 150:24:@27723.4]
  wire [31:0] x393_sum_1_io_a; // @[Math.scala 150:24:@27723.4]
  wire [31:0] x393_sum_1_io_b; // @[Math.scala 150:24:@27723.4]
  wire  x393_sum_1_io_flow; // @[Math.scala 150:24:@27723.4]
  wire [31:0] x393_sum_1_io_result; // @[Math.scala 150:24:@27723.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@27733.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@27733.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@27733.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@27733.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@27733.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@27745.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@27745.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@27745.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@27745.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@27745.4]
  wire  x398_rdrow_1_clock; // @[Math.scala 191:24:@27768.4]
  wire  x398_rdrow_1_reset; // @[Math.scala 191:24:@27768.4]
  wire [31:0] x398_rdrow_1_io_a; // @[Math.scala 191:24:@27768.4]
  wire [31:0] x398_rdrow_1_io_b; // @[Math.scala 191:24:@27768.4]
  wire  x398_rdrow_1_io_flow; // @[Math.scala 191:24:@27768.4]
  wire [31:0] x398_rdrow_1_io_result; // @[Math.scala 191:24:@27768.4]
  wire  x405_sum_1_clock; // @[Math.scala 150:24:@27822.4]
  wire  x405_sum_1_reset; // @[Math.scala 150:24:@27822.4]
  wire [31:0] x405_sum_1_io_a; // @[Math.scala 150:24:@27822.4]
  wire [31:0] x405_sum_1_io_b; // @[Math.scala 150:24:@27822.4]
  wire  x405_sum_1_io_flow; // @[Math.scala 150:24:@27822.4]
  wire [31:0] x405_sum_1_io_result; // @[Math.scala 150:24:@27822.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@27832.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@27832.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@27832.4]
  wire [31:0] RetimeWrapper_46_io_in; // @[package.scala 93:22:@27832.4]
  wire [31:0] RetimeWrapper_46_io_out; // @[package.scala 93:22:@27832.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@27841.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@27841.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@27841.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@27841.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@27841.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@27853.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@27853.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@27853.4]
  wire  RetimeWrapper_48_io_in; // @[package.scala 93:22:@27853.4]
  wire  RetimeWrapper_48_io_out; // @[package.scala 93:22:@27853.4]
  wire  x413_sum_1_clock; // @[Math.scala 150:24:@27880.4]
  wire  x413_sum_1_reset; // @[Math.scala 150:24:@27880.4]
  wire [31:0] x413_sum_1_io_a; // @[Math.scala 150:24:@27880.4]
  wire [31:0] x413_sum_1_io_b; // @[Math.scala 150:24:@27880.4]
  wire  x413_sum_1_io_flow; // @[Math.scala 150:24:@27880.4]
  wire [31:0] x413_sum_1_io_result; // @[Math.scala 150:24:@27880.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@27890.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@27890.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@27890.4]
  wire  RetimeWrapper_49_io_in; // @[package.scala 93:22:@27890.4]
  wire  RetimeWrapper_49_io_out; // @[package.scala 93:22:@27890.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@27902.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@27902.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@27902.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@27902.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@27902.4]
  wire  x420_sum_1_clock; // @[Math.scala 150:24:@27929.4]
  wire  x420_sum_1_reset; // @[Math.scala 150:24:@27929.4]
  wire [31:0] x420_sum_1_io_a; // @[Math.scala 150:24:@27929.4]
  wire [31:0] x420_sum_1_io_b; // @[Math.scala 150:24:@27929.4]
  wire  x420_sum_1_io_flow; // @[Math.scala 150:24:@27929.4]
  wire [31:0] x420_sum_1_io_result; // @[Math.scala 150:24:@27929.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@27939.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@27939.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@27939.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@27939.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@27939.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@27951.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@27951.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@27951.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@27951.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@27951.4]
  wire  x427_sum_1_clock; // @[Math.scala 150:24:@27978.4]
  wire  x427_sum_1_reset; // @[Math.scala 150:24:@27978.4]
  wire [31:0] x427_sum_1_io_a; // @[Math.scala 150:24:@27978.4]
  wire [31:0] x427_sum_1_io_b; // @[Math.scala 150:24:@27978.4]
  wire  x427_sum_1_io_flow; // @[Math.scala 150:24:@27978.4]
  wire [31:0] x427_sum_1_io_result; // @[Math.scala 150:24:@27978.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@27988.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@27988.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@27988.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@27988.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@27988.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@28000.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@28000.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@28000.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@28000.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@28000.4]
  wire  x437_x23_1_clock; // @[Math.scala 150:24:@28048.4]
  wire  x437_x23_1_reset; // @[Math.scala 150:24:@28048.4]
  wire [7:0] x437_x23_1_io_a; // @[Math.scala 150:24:@28048.4]
  wire [7:0] x437_x23_1_io_b; // @[Math.scala 150:24:@28048.4]
  wire  x437_x23_1_io_flow; // @[Math.scala 150:24:@28048.4]
  wire [7:0] x437_x23_1_io_result; // @[Math.scala 150:24:@28048.4]
  wire  x438_x24_1_clock; // @[Math.scala 150:24:@28058.4]
  wire  x438_x24_1_reset; // @[Math.scala 150:24:@28058.4]
  wire [7:0] x438_x24_1_io_a; // @[Math.scala 150:24:@28058.4]
  wire [7:0] x438_x24_1_io_b; // @[Math.scala 150:24:@28058.4]
  wire  x438_x24_1_io_flow; // @[Math.scala 150:24:@28058.4]
  wire [7:0] x438_x24_1_io_result; // @[Math.scala 150:24:@28058.4]
  wire  x439_x23_1_clock; // @[Math.scala 150:24:@28068.4]
  wire  x439_x23_1_reset; // @[Math.scala 150:24:@28068.4]
  wire [7:0] x439_x23_1_io_a; // @[Math.scala 150:24:@28068.4]
  wire [7:0] x439_x23_1_io_b; // @[Math.scala 150:24:@28068.4]
  wire  x439_x23_1_io_flow; // @[Math.scala 150:24:@28068.4]
  wire [7:0] x439_x23_1_io_result; // @[Math.scala 150:24:@28068.4]
  wire  x440_x24_1_clock; // @[Math.scala 150:24:@28078.4]
  wire  x440_x24_1_reset; // @[Math.scala 150:24:@28078.4]
  wire [7:0] x440_x24_1_io_a; // @[Math.scala 150:24:@28078.4]
  wire [7:0] x440_x24_1_io_b; // @[Math.scala 150:24:@28078.4]
  wire  x440_x24_1_io_flow; // @[Math.scala 150:24:@28078.4]
  wire [7:0] x440_x24_1_io_result; // @[Math.scala 150:24:@28078.4]
  wire [7:0] x441_x23_1_io_a; // @[Math.scala 150:24:@28088.4]
  wire [7:0] x441_x23_1_io_b; // @[Math.scala 150:24:@28088.4]
  wire [7:0] x441_x23_1_io_result; // @[Math.scala 150:24:@28088.4]
  wire [7:0] x442_x24_1_io_a; // @[Math.scala 150:24:@28098.4]
  wire [7:0] x442_x24_1_io_b; // @[Math.scala 150:24:@28098.4]
  wire [7:0] x442_x24_1_io_result; // @[Math.scala 150:24:@28098.4]
  wire [7:0] x443_x23_1_io_a; // @[Math.scala 150:24:@28108.4]
  wire [7:0] x443_x23_1_io_b; // @[Math.scala 150:24:@28108.4]
  wire [7:0] x443_x23_1_io_result; // @[Math.scala 150:24:@28108.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@28118.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@28118.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@28118.4]
  wire [7:0] RetimeWrapper_55_io_in; // @[package.scala 93:22:@28118.4]
  wire [7:0] RetimeWrapper_55_io_out; // @[package.scala 93:22:@28118.4]
  wire [7:0] x444_sum_1_io_a; // @[Math.scala 150:24:@28127.4]
  wire [7:0] x444_sum_1_io_b; // @[Math.scala 150:24:@28127.4]
  wire [7:0] x444_sum_1_io_result; // @[Math.scala 150:24:@28127.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@28141.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@28141.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@28141.4]
  wire [7:0] RetimeWrapper_56_io_in; // @[package.scala 93:22:@28141.4]
  wire [7:0] RetimeWrapper_56_io_out; // @[package.scala 93:22:@28141.4]
  wire  x451_x23_1_clock; // @[Math.scala 150:24:@28176.4]
  wire  x451_x23_1_reset; // @[Math.scala 150:24:@28176.4]
  wire [7:0] x451_x23_1_io_a; // @[Math.scala 150:24:@28176.4]
  wire [7:0] x451_x23_1_io_b; // @[Math.scala 150:24:@28176.4]
  wire  x451_x23_1_io_flow; // @[Math.scala 150:24:@28176.4]
  wire [7:0] x451_x23_1_io_result; // @[Math.scala 150:24:@28176.4]
  wire  x452_x24_1_clock; // @[Math.scala 150:24:@28186.4]
  wire  x452_x24_1_reset; // @[Math.scala 150:24:@28186.4]
  wire [7:0] x452_x24_1_io_a; // @[Math.scala 150:24:@28186.4]
  wire [7:0] x452_x24_1_io_b; // @[Math.scala 150:24:@28186.4]
  wire  x452_x24_1_io_flow; // @[Math.scala 150:24:@28186.4]
  wire [7:0] x452_x24_1_io_result; // @[Math.scala 150:24:@28186.4]
  wire  x453_x23_1_clock; // @[Math.scala 150:24:@28196.4]
  wire  x453_x23_1_reset; // @[Math.scala 150:24:@28196.4]
  wire [7:0] x453_x23_1_io_a; // @[Math.scala 150:24:@28196.4]
  wire [7:0] x453_x23_1_io_b; // @[Math.scala 150:24:@28196.4]
  wire  x453_x23_1_io_flow; // @[Math.scala 150:24:@28196.4]
  wire [7:0] x453_x23_1_io_result; // @[Math.scala 150:24:@28196.4]
  wire  x454_x24_1_clock; // @[Math.scala 150:24:@28206.4]
  wire  x454_x24_1_reset; // @[Math.scala 150:24:@28206.4]
  wire [7:0] x454_x24_1_io_a; // @[Math.scala 150:24:@28206.4]
  wire [7:0] x454_x24_1_io_b; // @[Math.scala 150:24:@28206.4]
  wire  x454_x24_1_io_flow; // @[Math.scala 150:24:@28206.4]
  wire [7:0] x454_x24_1_io_result; // @[Math.scala 150:24:@28206.4]
  wire [7:0] x455_x23_1_io_a; // @[Math.scala 150:24:@28216.4]
  wire [7:0] x455_x23_1_io_b; // @[Math.scala 150:24:@28216.4]
  wire [7:0] x455_x23_1_io_result; // @[Math.scala 150:24:@28216.4]
  wire [7:0] x456_x24_1_io_a; // @[Math.scala 150:24:@28226.4]
  wire [7:0] x456_x24_1_io_b; // @[Math.scala 150:24:@28226.4]
  wire [7:0] x456_x24_1_io_result; // @[Math.scala 150:24:@28226.4]
  wire [7:0] x457_x23_1_io_a; // @[Math.scala 150:24:@28236.4]
  wire [7:0] x457_x23_1_io_b; // @[Math.scala 150:24:@28236.4]
  wire [7:0] x457_x23_1_io_result; // @[Math.scala 150:24:@28236.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@28246.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@28246.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@28246.4]
  wire [7:0] RetimeWrapper_57_io_in; // @[package.scala 93:22:@28246.4]
  wire [7:0] RetimeWrapper_57_io_out; // @[package.scala 93:22:@28246.4]
  wire [7:0] x458_sum_1_io_a; // @[Math.scala 150:24:@28255.4]
  wire [7:0] x458_sum_1_io_b; // @[Math.scala 150:24:@28255.4]
  wire [7:0] x458_sum_1_io_result; // @[Math.scala 150:24:@28255.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@28269.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@28269.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@28269.4]
  wire [7:0] RetimeWrapper_58_io_in; // @[package.scala 93:22:@28269.4]
  wire [7:0] RetimeWrapper_58_io_out; // @[package.scala 93:22:@28269.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@28279.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@28279.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@28279.4]
  wire [31:0] RetimeWrapper_59_io_in; // @[package.scala 93:22:@28279.4]
  wire [31:0] RetimeWrapper_59_io_out; // @[package.scala 93:22:@28279.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@28288.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@28288.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@28288.4]
  wire  RetimeWrapper_60_io_in; // @[package.scala 93:22:@28288.4]
  wire  RetimeWrapper_60_io_out; // @[package.scala 93:22:@28288.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@28297.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@28297.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@28297.4]
  wire [31:0] RetimeWrapper_61_io_in; // @[package.scala 93:22:@28297.4]
  wire [31:0] RetimeWrapper_61_io_out; // @[package.scala 93:22:@28297.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@28306.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@28306.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@28306.4]
  wire  RetimeWrapper_62_io_in; // @[package.scala 93:22:@28306.4]
  wire  RetimeWrapper_62_io_out; // @[package.scala 93:22:@28306.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@28315.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@28315.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@28315.4]
  wire [31:0] RetimeWrapper_63_io_in; // @[package.scala 93:22:@28315.4]
  wire [31:0] RetimeWrapper_63_io_out; // @[package.scala 93:22:@28315.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@28326.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@28326.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@28326.4]
  wire  RetimeWrapper_64_io_in; // @[package.scala 93:22:@28326.4]
  wire  RetimeWrapper_64_io_out; // @[package.scala 93:22:@28326.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@28347.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@28347.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@28347.4]
  wire [31:0] RetimeWrapper_65_io_in; // @[package.scala 93:22:@28347.4]
  wire [31:0] RetimeWrapper_65_io_out; // @[package.scala 93:22:@28347.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@28356.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@28356.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@28356.4]
  wire [31:0] RetimeWrapper_66_io_in; // @[package.scala 93:22:@28356.4]
  wire [31:0] RetimeWrapper_66_io_out; // @[package.scala 93:22:@28356.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@28367.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@28367.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@28367.4]
  wire  RetimeWrapper_67_io_in; // @[package.scala 93:22:@28367.4]
  wire  RetimeWrapper_67_io_out; // @[package.scala 93:22:@28367.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@28388.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@28388.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@28388.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@28388.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@28388.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@28397.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@28397.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@28397.4]
  wire [31:0] RetimeWrapper_69_io_in; // @[package.scala 93:22:@28397.4]
  wire [31:0] RetimeWrapper_69_io_out; // @[package.scala 93:22:@28397.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@28406.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@28406.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@28406.4]
  wire [31:0] RetimeWrapper_70_io_in; // @[package.scala 93:22:@28406.4]
  wire [31:0] RetimeWrapper_70_io_out; // @[package.scala 93:22:@28406.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@28418.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@28418.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@28418.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@28418.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@28418.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@28439.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@28439.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@28439.4]
  wire  RetimeWrapper_72_io_in; // @[package.scala 93:22:@28439.4]
  wire  RetimeWrapper_72_io_out; // @[package.scala 93:22:@28439.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@28448.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@28448.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@28448.4]
  wire [31:0] RetimeWrapper_73_io_in; // @[package.scala 93:22:@28448.4]
  wire [31:0] RetimeWrapper_73_io_out; // @[package.scala 93:22:@28448.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@28460.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@28460.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@28460.4]
  wire  RetimeWrapper_74_io_in; // @[package.scala 93:22:@28460.4]
  wire  RetimeWrapper_74_io_out; // @[package.scala 93:22:@28460.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@28481.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@28481.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@28481.4]
  wire [31:0] RetimeWrapper_75_io_in; // @[package.scala 93:22:@28481.4]
  wire [31:0] RetimeWrapper_75_io_out; // @[package.scala 93:22:@28481.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@28490.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@28490.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@28490.4]
  wire  RetimeWrapper_76_io_in; // @[package.scala 93:22:@28490.4]
  wire  RetimeWrapper_76_io_out; // @[package.scala 93:22:@28490.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@28499.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@28499.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@28499.4]
  wire [31:0] RetimeWrapper_77_io_in; // @[package.scala 93:22:@28499.4]
  wire [31:0] RetimeWrapper_77_io_out; // @[package.scala 93:22:@28499.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@28511.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@28511.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@28511.4]
  wire  RetimeWrapper_78_io_in; // @[package.scala 93:22:@28511.4]
  wire  RetimeWrapper_78_io_out; // @[package.scala 93:22:@28511.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@28532.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@28532.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@28532.4]
  wire [31:0] RetimeWrapper_79_io_in; // @[package.scala 93:22:@28532.4]
  wire [31:0] RetimeWrapper_79_io_out; // @[package.scala 93:22:@28532.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@28541.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@28541.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@28541.4]
  wire  RetimeWrapper_80_io_in; // @[package.scala 93:22:@28541.4]
  wire  RetimeWrapper_80_io_out; // @[package.scala 93:22:@28541.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@28550.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@28550.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@28550.4]
  wire [31:0] RetimeWrapper_81_io_in; // @[package.scala 93:22:@28550.4]
  wire [31:0] RetimeWrapper_81_io_out; // @[package.scala 93:22:@28550.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@28562.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@28562.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@28562.4]
  wire  RetimeWrapper_82_io_in; // @[package.scala 93:22:@28562.4]
  wire  RetimeWrapper_82_io_out; // @[package.scala 93:22:@28562.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@28583.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@28583.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@28583.4]
  wire [31:0] RetimeWrapper_83_io_in; // @[package.scala 93:22:@28583.4]
  wire [31:0] RetimeWrapper_83_io_out; // @[package.scala 93:22:@28583.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@28592.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@28592.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@28592.4]
  wire  RetimeWrapper_84_io_in; // @[package.scala 93:22:@28592.4]
  wire  RetimeWrapper_84_io_out; // @[package.scala 93:22:@28592.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@28604.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@28604.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@28604.4]
  wire  RetimeWrapper_85_io_in; // @[package.scala 93:22:@28604.4]
  wire  RetimeWrapper_85_io_out; // @[package.scala 93:22:@28604.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@28625.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@28625.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@28625.4]
  wire  RetimeWrapper_86_io_in; // @[package.scala 93:22:@28625.4]
  wire  RetimeWrapper_86_io_out; // @[package.scala 93:22:@28625.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@28634.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@28634.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@28634.4]
  wire [31:0] RetimeWrapper_87_io_in; // @[package.scala 93:22:@28634.4]
  wire [31:0] RetimeWrapper_87_io_out; // @[package.scala 93:22:@28634.4]
  wire  RetimeWrapper_88_clock; // @[package.scala 93:22:@28646.4]
  wire  RetimeWrapper_88_reset; // @[package.scala 93:22:@28646.4]
  wire  RetimeWrapper_88_io_flow; // @[package.scala 93:22:@28646.4]
  wire  RetimeWrapper_88_io_in; // @[package.scala 93:22:@28646.4]
  wire  RetimeWrapper_88_io_out; // @[package.scala 93:22:@28646.4]
  wire [7:0] x478_x25_1_io_a; // @[Math.scala 150:24:@28679.4]
  wire [7:0] x478_x25_1_io_b; // @[Math.scala 150:24:@28679.4]
  wire [7:0] x478_x25_1_io_result; // @[Math.scala 150:24:@28679.4]
  wire [7:0] x479_x26_1_io_a; // @[Math.scala 150:24:@28689.4]
  wire [7:0] x479_x26_1_io_b; // @[Math.scala 150:24:@28689.4]
  wire [7:0] x479_x26_1_io_result; // @[Math.scala 150:24:@28689.4]
  wire [7:0] x480_sum_1_io_a; // @[Math.scala 150:24:@28699.4]
  wire [7:0] x480_sum_1_io_b; // @[Math.scala 150:24:@28699.4]
  wire [7:0] x480_sum_1_io_result; // @[Math.scala 150:24:@28699.4]
  wire  x481_div_1_clock; // @[Math.scala 327:24:@28711.4]
  wire  x481_div_1_reset; // @[Math.scala 327:24:@28711.4]
  wire [7:0] x481_div_1_io_a; // @[Math.scala 327:24:@28711.4]
  wire  x481_div_1_io_flow; // @[Math.scala 327:24:@28711.4]
  wire [7:0] x481_div_1_io_result; // @[Math.scala 327:24:@28711.4]
  wire [7:0] x484_x25_1_io_a; // @[Math.scala 150:24:@28731.4]
  wire [7:0] x484_x25_1_io_b; // @[Math.scala 150:24:@28731.4]
  wire [7:0] x484_x25_1_io_result; // @[Math.scala 150:24:@28731.4]
  wire [7:0] x485_x26_1_io_a; // @[Math.scala 150:24:@28741.4]
  wire [7:0] x485_x26_1_io_b; // @[Math.scala 150:24:@28741.4]
  wire [7:0] x485_x26_1_io_result; // @[Math.scala 150:24:@28741.4]
  wire [7:0] x486_sum_1_io_a; // @[Math.scala 150:24:@28751.4]
  wire [7:0] x486_sum_1_io_b; // @[Math.scala 150:24:@28751.4]
  wire [7:0] x486_sum_1_io_result; // @[Math.scala 150:24:@28751.4]
  wire  x487_div_1_clock; // @[Math.scala 327:24:@28763.4]
  wire  x487_div_1_reset; // @[Math.scala 327:24:@28763.4]
  wire [7:0] x487_div_1_io_a; // @[Math.scala 327:24:@28763.4]
  wire  x487_div_1_io_flow; // @[Math.scala 327:24:@28763.4]
  wire [7:0] x487_div_1_io_result; // @[Math.scala 327:24:@28763.4]
  wire  RetimeWrapper_89_clock; // @[package.scala 93:22:@28779.4]
  wire  RetimeWrapper_89_reset; // @[package.scala 93:22:@28779.4]
  wire  RetimeWrapper_89_io_flow; // @[package.scala 93:22:@28779.4]
  wire [15:0] RetimeWrapper_89_io_in; // @[package.scala 93:22:@28779.4]
  wire [15:0] RetimeWrapper_89_io_out; // @[package.scala 93:22:@28779.4]
  wire  RetimeWrapper_90_clock; // @[package.scala 93:22:@28788.4]
  wire  RetimeWrapper_90_reset; // @[package.scala 93:22:@28788.4]
  wire  RetimeWrapper_90_io_flow; // @[package.scala 93:22:@28788.4]
  wire  RetimeWrapper_90_io_in; // @[package.scala 93:22:@28788.4]
  wire  RetimeWrapper_90_io_out; // @[package.scala 93:22:@28788.4]
  wire  RetimeWrapper_91_clock; // @[package.scala 93:22:@28797.4]
  wire  RetimeWrapper_91_reset; // @[package.scala 93:22:@28797.4]
  wire  RetimeWrapper_91_io_flow; // @[package.scala 93:22:@28797.4]
  wire  RetimeWrapper_91_io_in; // @[package.scala 93:22:@28797.4]
  wire  RetimeWrapper_91_io_out; // @[package.scala 93:22:@28797.4]
  wire  RetimeWrapper_92_clock; // @[package.scala 93:22:@28806.4]
  wire  RetimeWrapper_92_reset; // @[package.scala 93:22:@28806.4]
  wire  RetimeWrapper_92_io_flow; // @[package.scala 93:22:@28806.4]
  wire  RetimeWrapper_92_io_in; // @[package.scala 93:22:@28806.4]
  wire  RetimeWrapper_92_io_out; // @[package.scala 93:22:@28806.4]
  wire  b286; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 62:18:@26575.4]
  wire  b287; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 63:18:@26576.4]
  wire  _T_207; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 69:30:@26728.4]
  wire  _T_208; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 69:37:@26729.4]
  wire  _T_212; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 71:76:@26734.4]
  wire  _T_213; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 71:62:@26735.4]
  wire  _T_215; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 71:101:@26736.4]
  wire [15:0] x571_x290_D1_0_number; // @[package.scala 96:25:@26745.4 package.scala 96:25:@26746.4]
  wire [31:0] b284_number; // @[Math.scala 712:22:@26560.4 Math.scala 713:14:@26561.4]
  wire [31:0] _T_243; // @[Math.scala 499:52:@26761.4]
  wire  x294; // @[Math.scala 499:44:@26769.4]
  wire  x295; // @[Math.scala 499:44:@26776.4]
  wire  x296; // @[Math.scala 499:44:@26783.4]
  wire [31:0] _T_290; // @[Mux.scala 19:72:@26795.4]
  wire [31:0] _T_292; // @[Mux.scala 19:72:@26796.4]
  wire [31:0] _T_294; // @[Mux.scala 19:72:@26797.4]
  wire [31:0] _T_296; // @[Mux.scala 19:72:@26799.4]
  wire [31:0] x297_number; // @[Mux.scala 19:72:@26800.4]
  wire [31:0] _T_308; // @[Math.scala 406:49:@26810.4]
  wire [31:0] _T_310; // @[Math.scala 406:56:@26812.4]
  wire [31:0] _T_311; // @[Math.scala 406:56:@26813.4]
  wire [31:0] b285_number; // @[Math.scala 712:22:@26572.4 Math.scala 713:14:@26573.4]
  wire [31:0] _T_320; // @[Math.scala 406:49:@26821.4]
  wire [31:0] _T_322; // @[Math.scala 406:56:@26823.4]
  wire [31:0] _T_323; // @[Math.scala 406:56:@26824.4]
  wire  _T_328; // @[FixedPoint.scala 50:25:@26830.4]
  wire [1:0] _T_332; // @[Bitwise.scala 72:12:@26832.4]
  wire [29:0] _T_333; // @[FixedPoint.scala 18:52:@26833.4]
  wire  _T_338; // @[FixedPoint.scala 50:25:@26839.4]
  wire [1:0] _T_342; // @[Bitwise.scala 72:12:@26841.4]
  wire [29:0] _T_343; // @[FixedPoint.scala 18:52:@26842.4]
  wire  _T_367; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 118:101:@26910.4]
  wire  _T_371; // @[package.scala 96:25:@26918.4 package.scala 96:25:@26919.4]
  wire  _T_373; // @[implicits.scala 55:10:@26920.4]
  wire  _T_374; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 118:118:@26921.4]
  wire  _T_376; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 118:205:@26923.4]
  wire  _T_377; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 118:224:@26924.4]
  wire  x574_b286_D2; // @[package.scala 96:25:@26880.4 package.scala 96:25:@26881.4]
  wire  _T_378; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 118:250:@26925.4]
  wire  x576_b287_D2; // @[package.scala 96:25:@26898.4 package.scala 96:25:@26899.4]
  wire [31:0] x309_rdcol_number; // @[Math.scala 154:22:@26942.4 Math.scala 155:14:@26943.4]
  wire [31:0] _T_395; // @[Math.scala 406:49:@26951.4]
  wire [31:0] _T_397; // @[Math.scala 406:56:@26953.4]
  wire [31:0] _T_398; // @[Math.scala 406:56:@26954.4]
  wire  _T_403; // @[FixedPoint.scala 50:25:@26960.4]
  wire [1:0] _T_407; // @[Bitwise.scala 72:12:@26962.4]
  wire [29:0] _T_408; // @[FixedPoint.scala 18:52:@26963.4]
  wire  _T_427; // @[package.scala 96:25:@27012.4 package.scala 96:25:@27013.4]
  wire  _T_429; // @[implicits.scala 55:10:@27014.4]
  wire  _T_430; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 139:118:@27015.4]
  wire  _T_432; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 139:205:@27017.4]
  wire  _T_433; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 139:224:@27018.4]
  wire  _T_434; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 139:250:@27019.4]
  wire [31:0] x581_b284_D4_number; // @[package.scala 96:25:@27033.4 package.scala 96:25:@27034.4]
  wire [31:0] _T_446; // @[Math.scala 406:49:@27040.4]
  wire [31:0] _T_448; // @[Math.scala 406:56:@27042.4]
  wire [31:0] _T_449; // @[Math.scala 406:56:@27043.4]
  wire [31:0] x563_number; // @[implicits.scala 133:21:@27044.4]
  wire  x320; // @[Math.scala 465:44:@27052.4]
  wire [31:0] x582_x309_rdcol_D4_number; // @[package.scala 96:25:@27060.4 package.scala 96:25:@27061.4]
  wire [31:0] _T_467; // @[Math.scala 465:37:@27066.4]
  wire  x321; // @[Math.scala 465:44:@27068.4]
  wire  x583_x320_D1; // @[package.scala 96:25:@27076.4 package.scala 96:25:@27077.4]
  wire  x322; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 154:24:@27080.4]
  wire [31:0] _T_484; // @[Math.scala 406:49:@27089.4]
  wire [31:0] _T_486; // @[Math.scala 406:56:@27091.4]
  wire [31:0] _T_487; // @[Math.scala 406:56:@27092.4]
  wire  _T_492; // @[FixedPoint.scala 50:25:@27098.4]
  wire [1:0] _T_496; // @[Bitwise.scala 72:12:@27100.4]
  wire [29:0] _T_497; // @[FixedPoint.scala 18:52:@27101.4]
  wire  _T_534; // @[package.scala 96:25:@27187.4 package.scala 96:25:@27188.4]
  wire  _T_536; // @[implicits.scala 55:10:@27189.4]
  wire  _T_537; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 187:194:@27190.4]
  wire  x588_x323_D1; // @[package.scala 96:25:@27157.4 package.scala 96:25:@27158.4]
  wire  _T_538; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 187:281:@27191.4]
  wire  x587_b286_D6; // @[package.scala 96:25:@27148.4 package.scala 96:25:@27149.4]
  wire  _T_539; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 187:289:@27192.4]
  wire  x589_b287_D6; // @[package.scala 96:25:@27166.4 package.scala 96:25:@27167.4]
  wire [31:0] x591_b285_D4_number; // @[package.scala 96:25:@27208.4 package.scala 96:25:@27209.4]
  wire [31:0] _T_552; // @[Math.scala 465:37:@27216.4]
  wire  x332; // @[Math.scala 465:44:@27218.4]
  wire  x333; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 197:59:@27221.4]
  wire  _T_585; // @[package.scala 96:25:@27281.4 package.scala 96:25:@27282.4]
  wire  _T_587; // @[implicits.scala 55:10:@27283.4]
  wire  _T_588; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 214:194:@27284.4]
  wire  x593_x334_D2; // @[package.scala 96:25:@27251.4 package.scala 96:25:@27252.4]
  wire  _T_589; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 214:281:@27285.4]
  wire  _T_590; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 214:289:@27286.4]
  wire [31:0] x340_rdcol_number; // @[Math.scala 154:22:@27305.4 Math.scala 155:14:@27306.4]
  wire [31:0] _T_605; // @[Math.scala 465:37:@27311.4]
  wire  x341; // @[Math.scala 465:44:@27313.4]
  wire  x342; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 222:59:@27316.4]
  wire [31:0] _T_621; // @[Math.scala 406:56:@27327.4]
  wire [31:0] _T_622; // @[Math.scala 406:56:@27328.4]
  wire  _T_627; // @[FixedPoint.scala 50:25:@27334.4]
  wire [1:0] _T_631; // @[Bitwise.scala 72:12:@27336.4]
  wire [29:0] _T_632; // @[FixedPoint.scala 18:52:@27337.4]
  wire  _T_654; // @[package.scala 96:25:@27378.4 package.scala 96:25:@27379.4]
  wire  _T_656; // @[implicits.scala 55:10:@27380.4]
  wire  _T_657; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 239:194:@27381.4]
  wire  x597_x343_D1; // @[package.scala 96:25:@27366.4 package.scala 96:25:@27367.4]
  wire  _T_658; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 239:281:@27382.4]
  wire  _T_659; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 239:289:@27383.4]
  wire [31:0] x352_rdcol_number; // @[Math.scala 154:22:@27402.4 Math.scala 155:14:@27403.4]
  wire [31:0] _T_674; // @[Math.scala 465:37:@27408.4]
  wire  x353; // @[Math.scala 465:44:@27410.4]
  wire  x354; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 247:59:@27413.4]
  wire [31:0] _T_690; // @[Math.scala 406:56:@27424.4]
  wire [31:0] _T_691; // @[Math.scala 406:56:@27425.4]
  wire  _T_696; // @[FixedPoint.scala 50:25:@27431.4]
  wire [1:0] _T_700; // @[Bitwise.scala 72:12:@27433.4]
  wire [29:0] _T_701; // @[FixedPoint.scala 18:52:@27434.4]
  wire  _T_723; // @[package.scala 96:25:@27475.4 package.scala 96:25:@27476.4]
  wire  _T_725; // @[implicits.scala 55:10:@27477.4]
  wire  _T_726; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 264:194:@27478.4]
  wire  x599_x355_D1; // @[package.scala 96:25:@27463.4 package.scala 96:25:@27464.4]
  wire  _T_727; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 264:281:@27479.4]
  wire  _T_728; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 264:289:@27480.4]
  wire [31:0] x364_rdrow_number; // @[Math.scala 195:22:@27499.4 Math.scala 196:14:@27500.4]
  wire [31:0] _T_745; // @[Math.scala 406:49:@27506.4]
  wire [31:0] _T_747; // @[Math.scala 406:56:@27508.4]
  wire [31:0] _T_748; // @[Math.scala 406:56:@27509.4]
  wire [31:0] x567_number; // @[implicits.scala 133:21:@27510.4]
  wire  x366; // @[Math.scala 465:44:@27518.4]
  wire  x367; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 274:24:@27521.4]
  wire [31:0] _T_769; // @[Math.scala 406:49:@27530.4]
  wire [31:0] _T_771; // @[Math.scala 406:56:@27532.4]
  wire [31:0] _T_772; // @[Math.scala 406:56:@27533.4]
  wire  _T_777; // @[FixedPoint.scala 50:25:@27539.4]
  wire [1:0] _T_781; // @[Bitwise.scala 72:12:@27541.4]
  wire [29:0] _T_782; // @[FixedPoint.scala 18:52:@27542.4]
  wire  _T_804; // @[package.scala 96:25:@27583.4 package.scala 96:25:@27584.4]
  wire  _T_806; // @[implicits.scala 55:10:@27585.4]
  wire  _T_807; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 291:194:@27586.4]
  wire  x600_x368_D1; // @[package.scala 96:25:@27562.4 package.scala 96:25:@27563.4]
  wire  _T_808; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 291:281:@27587.4]
  wire  _T_809; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 291:289:@27588.4]
  wire  x602_x332_D1; // @[package.scala 96:25:@27604.4 package.scala 96:25:@27605.4]
  wire  x377; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 303:59:@27608.4]
  wire  _T_841; // @[package.scala 96:25:@27652.4 package.scala 96:25:@27653.4]
  wire  _T_843; // @[implicits.scala 55:10:@27654.4]
  wire  _T_844; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 318:194:@27655.4]
  wire  x604_x378_D1; // @[package.scala 96:25:@27640.4 package.scala 96:25:@27641.4]
  wire  _T_845; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 318:281:@27656.4]
  wire  _T_846; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 318:289:@27657.4]
  wire  x384; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 322:59:@27668.4]
  wire  _T_870; // @[package.scala 96:25:@27701.4 package.scala 96:25:@27702.4]
  wire  _T_872; // @[implicits.scala 55:10:@27703.4]
  wire  _T_873; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 333:194:@27704.4]
  wire  x605_x385_D1; // @[package.scala 96:25:@27689.4 package.scala 96:25:@27690.4]
  wire  _T_874; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 333:281:@27705.4]
  wire  _T_875; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 333:289:@27706.4]
  wire  x391; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 337:59:@27717.4]
  wire  _T_899; // @[package.scala 96:25:@27750.4 package.scala 96:25:@27751.4]
  wire  _T_901; // @[implicits.scala 55:10:@27752.4]
  wire  _T_902; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 348:194:@27753.4]
  wire  x606_x392_D1; // @[package.scala 96:25:@27738.4 package.scala 96:25:@27739.4]
  wire  _T_903; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 348:281:@27754.4]
  wire  _T_904; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 348:289:@27755.4]
  wire [31:0] x398_rdrow_number; // @[Math.scala 195:22:@27774.4 Math.scala 196:14:@27775.4]
  wire [31:0] _T_921; // @[Math.scala 406:49:@27781.4]
  wire [31:0] _T_923; // @[Math.scala 406:56:@27783.4]
  wire [31:0] _T_924; // @[Math.scala 406:56:@27784.4]
  wire [31:0] x569_number; // @[implicits.scala 133:21:@27785.4]
  wire  x400; // @[Math.scala 465:44:@27793.4]
  wire  x401; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 358:24:@27796.4]
  wire [31:0] _T_945; // @[Math.scala 406:49:@27805.4]
  wire [31:0] _T_947; // @[Math.scala 406:56:@27807.4]
  wire [31:0] _T_948; // @[Math.scala 406:56:@27808.4]
  wire  _T_953; // @[FixedPoint.scala 50:25:@27814.4]
  wire [1:0] _T_957; // @[Bitwise.scala 72:12:@27816.4]
  wire [29:0] _T_958; // @[FixedPoint.scala 18:52:@27817.4]
  wire  _T_980; // @[package.scala 96:25:@27858.4 package.scala 96:25:@27859.4]
  wire  _T_982; // @[implicits.scala 55:10:@27860.4]
  wire  _T_983; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 375:194:@27861.4]
  wire  x608_x402_D1; // @[package.scala 96:25:@27846.4 package.scala 96:25:@27847.4]
  wire  _T_984; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 375:281:@27862.4]
  wire  _T_985; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 375:289:@27863.4]
  wire  x411; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 379:24:@27874.4]
  wire  _T_1009; // @[package.scala 96:25:@27907.4 package.scala 96:25:@27908.4]
  wire  _T_1011; // @[implicits.scala 55:10:@27909.4]
  wire  _T_1012; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 390:194:@27910.4]
  wire  x609_x412_D1; // @[package.scala 96:25:@27895.4 package.scala 96:25:@27896.4]
  wire  _T_1013; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 390:281:@27911.4]
  wire  _T_1014; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 390:289:@27912.4]
  wire  x418; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 394:24:@27923.4]
  wire  _T_1038; // @[package.scala 96:25:@27956.4 package.scala 96:25:@27957.4]
  wire  _T_1040; // @[implicits.scala 55:10:@27958.4]
  wire  _T_1041; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 405:194:@27959.4]
  wire  x610_x419_D1; // @[package.scala 96:25:@27944.4 package.scala 96:25:@27945.4]
  wire  _T_1042; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 405:281:@27960.4]
  wire  _T_1043; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 405:289:@27961.4]
  wire  x425; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 409:24:@27972.4]
  wire  _T_1067; // @[package.scala 96:25:@28005.4 package.scala 96:25:@28006.4]
  wire  _T_1069; // @[implicits.scala 55:10:@28007.4]
  wire  _T_1070; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 426:194:@28008.4]
  wire  x611_x426_D1; // @[package.scala 96:25:@27993.4 package.scala 96:25:@27994.4]
  wire  _T_1071; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 426:281:@28009.4]
  wire  _T_1072; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 426:324:@28010.4]
  wire [7:0] x338_rd_0_number; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 210:29:@27272.4 sm_x492_inr_Foreach_SAMPLER_BOX.scala 214:371:@27293.4]
  wire [8:0] _GEN_0; // @[Math.scala 450:32:@28024.4]
  wire [8:0] _T_1080; // @[Math.scala 450:32:@28024.4]
  wire [7:0] x375_rd_0_number; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 287:29:@27574.4 sm_x492_inr_Foreach_SAMPLER_BOX.scala 291:371:@27595.4]
  wire [8:0] _GEN_1; // @[Math.scala 450:32:@28029.4]
  wire [8:0] _T_1084; // @[Math.scala 450:32:@28029.4]
  wire [7:0] x382_rd_0_number; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 314:29:@27643.4 sm_x492_inr_Foreach_SAMPLER_BOX.scala 318:406:@27664.4]
  wire [9:0] _GEN_2; // @[Math.scala 450:32:@28034.4]
  wire [9:0] _T_1088; // @[Math.scala 450:32:@28034.4]
  wire [7:0] x389_rd_0_number; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 329:29:@27692.4 sm_x492_inr_Foreach_SAMPLER_BOX.scala 333:406:@27713.4]
  wire [8:0] _GEN_3; // @[Math.scala 450:32:@28039.4]
  wire [8:0] _T_1092; // @[Math.scala 450:32:@28039.4]
  wire [7:0] x416_rd_0_number; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 386:29:@27898.4 sm_x492_inr_Foreach_SAMPLER_BOX.scala 390:406:@27919.4]
  wire [8:0] _GEN_4; // @[Math.scala 450:32:@28044.4]
  wire [8:0] _T_1096; // @[Math.scala 450:32:@28044.4]
  wire [7:0] x444_sum_number; // @[Math.scala 154:22:@28133.4 Math.scala 155:14:@28134.4]
  wire [3:0] _T_1132; // @[FixedPoint.scala 18:52:@28139.4]
  wire [7:0] x350_rd_0_number; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 235:29:@27369.4 sm_x492_inr_Foreach_SAMPLER_BOX.scala 239:371:@27390.4]
  wire [8:0] _GEN_5; // @[Math.scala 450:32:@28152.4]
  wire [8:0] _T_1139; // @[Math.scala 450:32:@28152.4]
  wire [8:0] _GEN_6; // @[Math.scala 450:32:@28157.4]
  wire [8:0] _T_1143; // @[Math.scala 450:32:@28157.4]
  wire [9:0] _GEN_7; // @[Math.scala 450:32:@28162.4]
  wire [9:0] _T_1147; // @[Math.scala 450:32:@28162.4]
  wire [7:0] x396_rd_0_number; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 344:29:@27741.4 sm_x492_inr_Foreach_SAMPLER_BOX.scala 348:406:@27762.4]
  wire [8:0] _GEN_8; // @[Math.scala 450:32:@28167.4]
  wire [8:0] _T_1151; // @[Math.scala 450:32:@28167.4]
  wire [7:0] x423_rd_0_number; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 401:29:@27947.4 sm_x492_inr_Foreach_SAMPLER_BOX.scala 405:406:@27968.4]
  wire [8:0] _GEN_9; // @[Math.scala 450:32:@28172.4]
  wire [8:0] _T_1155; // @[Math.scala 450:32:@28172.4]
  wire [7:0] x458_sum_number; // @[Math.scala 154:22:@28261.4 Math.scala 155:14:@28262.4]
  wire [3:0] _T_1191; // @[FixedPoint.scala 18:52:@28267.4]
  wire  _T_1215; // @[package.scala 96:25:@28331.4 package.scala 96:25:@28332.4]
  wire  _T_1217; // @[implicits.scala 55:10:@28333.4]
  wire  _T_1218; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 506:167:@28334.4]
  wire  _T_1220; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 506:255:@28336.4]
  wire  _T_1221; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 506:274:@28337.4]
  wire  x615_b286_D10; // @[package.scala 96:25:@28293.4 package.scala 96:25:@28294.4]
  wire  _T_1222; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 506:300:@28338.4]
  wire  x617_b287_D10; // @[package.scala 96:25:@28311.4 package.scala 96:25:@28312.4]
  wire  _T_1235; // @[package.scala 96:25:@28372.4 package.scala 96:25:@28373.4]
  wire  _T_1237; // @[implicits.scala 55:10:@28374.4]
  wire  _T_1238; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 515:167:@28375.4]
  wire  _T_1240; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 515:255:@28377.4]
  wire  _T_1241; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 515:274:@28378.4]
  wire  _T_1242; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 515:300:@28379.4]
  wire  _T_1264; // @[package.scala 96:25:@28423.4 package.scala 96:25:@28424.4]
  wire  _T_1266; // @[implicits.scala 55:10:@28425.4]
  wire  _T_1267; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 527:195:@28426.4]
  wire  x621_x323_D5; // @[package.scala 96:25:@28393.4 package.scala 96:25:@28394.4]
  wire  _T_1268; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 527:283:@28427.4]
  wire  _T_1269; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 527:291:@28428.4]
  wire  _T_1289; // @[package.scala 96:25:@28465.4 package.scala 96:25:@28466.4]
  wire  _T_1291; // @[implicits.scala 55:10:@28467.4]
  wire  _T_1292; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 544:195:@28468.4]
  wire  x624_x334_D6; // @[package.scala 96:25:@28444.4 package.scala 96:25:@28445.4]
  wire  _T_1293; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 544:283:@28469.4]
  wire  _T_1294; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 544:326:@28470.4]
  wire  _T_1317; // @[package.scala 96:25:@28516.4 package.scala 96:25:@28517.4]
  wire  _T_1319; // @[implicits.scala 55:10:@28518.4]
  wire  _T_1320; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 557:195:@28519.4]
  wire  x627_x343_D5; // @[package.scala 96:25:@28495.4 package.scala 96:25:@28496.4]
  wire  _T_1321; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 557:283:@28520.4]
  wire  _T_1322; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 557:291:@28521.4]
  wire  _T_1345; // @[package.scala 96:25:@28567.4 package.scala 96:25:@28568.4]
  wire  _T_1347; // @[implicits.scala 55:10:@28569.4]
  wire  _T_1348; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 570:195:@28570.4]
  wire  x630_x368_D5; // @[package.scala 96:25:@28546.4 package.scala 96:25:@28547.4]
  wire  _T_1349; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 570:283:@28571.4]
  wire  _T_1350; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 570:291:@28572.4]
  wire  _T_1370; // @[package.scala 96:25:@28609.4 package.scala 96:25:@28610.4]
  wire  _T_1372; // @[implicits.scala 55:10:@28611.4]
  wire  _T_1373; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 581:195:@28612.4]
  wire  x633_x378_D5; // @[package.scala 96:25:@28597.4 package.scala 96:25:@28598.4]
  wire  _T_1374; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 581:283:@28613.4]
  wire  _T_1375; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 581:291:@28614.4]
  wire  _T_1395; // @[package.scala 96:25:@28651.4 package.scala 96:25:@28652.4]
  wire  _T_1397; // @[implicits.scala 55:10:@28653.4]
  wire  _T_1398; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 592:195:@28654.4]
  wire  x634_x385_D5; // @[package.scala 96:25:@28630.4 package.scala 96:25:@28631.4]
  wire  _T_1399; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 592:283:@28655.4]
  wire  _T_1400; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 592:291:@28656.4]
  wire [7:0] x466_rd_0_number; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 540:29:@28456.4 sm_x492_inr_Foreach_SAMPLER_BOX.scala 544:443:@28477.4]
  wire [8:0] _GEN_10; // @[Math.scala 450:32:@28670.4]
  wire [8:0] _T_1408; // @[Math.scala 450:32:@28670.4]
  wire [7:0] x470_rd_0_number; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 566:29:@28558.4 sm_x492_inr_Foreach_SAMPLER_BOX.scala 570:408:@28579.4]
  wire [8:0] _GEN_11; // @[Math.scala 450:32:@28675.4]
  wire [8:0] _T_1412; // @[Math.scala 450:32:@28675.4]
  wire [7:0] x468_rd_0_number; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 553:29:@28507.4 sm_x492_inr_Foreach_SAMPLER_BOX.scala 557:408:@28528.4]
  wire [8:0] _GEN_12; // @[Math.scala 450:32:@28722.4]
  wire [8:0] _T_1432; // @[Math.scala 450:32:@28722.4]
  wire [7:0] x472_rd_0_number; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 577:29:@28600.4 sm_x492_inr_Foreach_SAMPLER_BOX.scala 581:408:@28621.4]
  wire [8:0] _GEN_13; // @[Math.scala 450:32:@28727.4]
  wire [8:0] _T_1436; // @[Math.scala 450:32:@28727.4]
  wire [7:0] x481_div_number; // @[Math.scala 331:22:@28717.4 Math.scala 332:14:@28718.4]
  wire [7:0] x487_div_number; // @[Math.scala 331:22:@28769.4 Math.scala 332:14:@28770.4]
  wire  _T_1474; // @[package.scala 96:25:@28811.4 package.scala 96:25:@28812.4]
  wire  _T_1476; // @[implicits.scala 55:10:@28813.4]
  wire  x637_b286_D20; // @[package.scala 96:25:@28802.4 package.scala 96:25:@28803.4]
  wire  _T_1477; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 630:116:@28814.4]
  wire  x636_b287_D20; // @[package.scala 96:25:@28793.4 package.scala 96:25:@28794.4]
  wire  _T_1478; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 630:122:@28815.4]
  wire [31:0] x572_x561_D2_number; // @[package.scala 96:25:@26862.4 package.scala 96:25:@26863.4]
  wire [31:0] x575_x303_sum_D1_number; // @[package.scala 96:25:@26889.4 package.scala 96:25:@26890.4]
  wire [31:0] x577_x560_D2_number; // @[package.scala 96:25:@26907.4 package.scala 96:25:@26908.4]
  wire [31:0] x313_sum_number; // @[Math.scala 154:22:@26983.4 Math.scala 155:14:@26984.4]
  wire [31:0] x579_x562_D1_number; // @[package.scala 96:25:@26992.4 package.scala 96:25:@26993.4]
  wire [31:0] x326_sum_number; // @[Math.scala 154:22:@27130.4 Math.scala 155:14:@27131.4]
  wire [31:0] x586_x562_D5_number; // @[package.scala 96:25:@27139.4 package.scala 96:25:@27140.4]
  wire [31:0] x590_x564_D2_number; // @[package.scala 96:25:@27175.4 package.scala 96:25:@27176.4]
  wire [31:0] x594_x561_D6_number; // @[package.scala 96:25:@27260.4 package.scala 96:25:@27261.4]
  wire [31:0] x595_x335_sum_D1_number; // @[package.scala 96:25:@27269.4 package.scala 96:25:@27270.4]
  wire [31:0] x346_sum_number; // @[Math.scala 154:22:@27348.4 Math.scala 155:14:@27349.4]
  wire [31:0] x596_x565_D1_number; // @[package.scala 96:25:@27357.4 package.scala 96:25:@27358.4]
  wire [31:0] x358_sum_number; // @[Math.scala 154:22:@27445.4 Math.scala 155:14:@27446.4]
  wire [31:0] x598_x566_D1_number; // @[package.scala 96:25:@27454.4 package.scala 96:25:@27455.4]
  wire [31:0] x371_sum_number; // @[Math.scala 154:22:@27553.4 Math.scala 155:14:@27554.4]
  wire [31:0] x601_x568_D1_number; // @[package.scala 96:25:@27571.4 package.scala 96:25:@27572.4]
  wire [31:0] x379_sum_number; // @[Math.scala 154:22:@27631.4 Math.scala 155:14:@27632.4]
  wire [31:0] x386_sum_number; // @[Math.scala 154:22:@27680.4 Math.scala 155:14:@27681.4]
  wire [31:0] x393_sum_number; // @[Math.scala 154:22:@27729.4 Math.scala 155:14:@27730.4]
  wire [31:0] x405_sum_number; // @[Math.scala 154:22:@27828.4 Math.scala 155:14:@27829.4]
  wire [31:0] x607_x570_D1_number; // @[package.scala 96:25:@27837.4 package.scala 96:25:@27838.4]
  wire [31:0] x413_sum_number; // @[Math.scala 154:22:@27886.4 Math.scala 155:14:@27887.4]
  wire [31:0] x420_sum_number; // @[Math.scala 154:22:@27935.4 Math.scala 155:14:@27936.4]
  wire [31:0] x427_sum_number; // @[Math.scala 154:22:@27984.4 Math.scala 155:14:@27985.4]
  wire [31:0] x614_x561_D10_number; // @[package.scala 96:25:@28284.4 package.scala 96:25:@28285.4]
  wire [31:0] x616_x303_sum_D9_number; // @[package.scala 96:25:@28302.4 package.scala 96:25:@28303.4]
  wire [31:0] x618_x560_D10_number; // @[package.scala 96:25:@28320.4 package.scala 96:25:@28321.4]
  wire [31:0] x619_x562_D9_number; // @[package.scala 96:25:@28352.4 package.scala 96:25:@28353.4]
  wire [31:0] x620_x313_sum_D8_number; // @[package.scala 96:25:@28361.4 package.scala 96:25:@28362.4]
  wire [31:0] x622_x564_D6_number; // @[package.scala 96:25:@28402.4 package.scala 96:25:@28403.4]
  wire [31:0] x623_x326_sum_D4_number; // @[package.scala 96:25:@28411.4 package.scala 96:25:@28412.4]
  wire [31:0] x625_x335_sum_D5_number; // @[package.scala 96:25:@28453.4 package.scala 96:25:@28454.4]
  wire [31:0] x626_x565_D5_number; // @[package.scala 96:25:@28486.4 package.scala 96:25:@28487.4]
  wire [31:0] x628_x346_sum_D4_number; // @[package.scala 96:25:@28504.4 package.scala 96:25:@28505.4]
  wire [31:0] x629_x371_sum_D4_number; // @[package.scala 96:25:@28537.4 package.scala 96:25:@28538.4]
  wire [31:0] x631_x568_D5_number; // @[package.scala 96:25:@28555.4 package.scala 96:25:@28556.4]
  wire [31:0] x632_x379_sum_D4_number; // @[package.scala 96:25:@28588.4 package.scala 96:25:@28589.4]
  wire [31:0] x635_x386_sum_D4_number; // @[package.scala 96:25:@28639.4 package.scala 96:25:@28640.4]
  _ _ ( // @[Math.scala 709:24:@26555.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 709:24:@26567.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  x288_lb_0 x288_lb_0 ( // @[m_x288_lb_0.scala 39:17:@26577.4]
    .clock(x288_lb_0_clock),
    .reset(x288_lb_0_reset),
    .io_rPort_11_banks_1(x288_lb_0_io_rPort_11_banks_1),
    .io_rPort_11_banks_0(x288_lb_0_io_rPort_11_banks_0),
    .io_rPort_11_ofs_0(x288_lb_0_io_rPort_11_ofs_0),
    .io_rPort_11_en_0(x288_lb_0_io_rPort_11_en_0),
    .io_rPort_11_backpressure(x288_lb_0_io_rPort_11_backpressure),
    .io_rPort_11_output_0(x288_lb_0_io_rPort_11_output_0),
    .io_rPort_10_banks_1(x288_lb_0_io_rPort_10_banks_1),
    .io_rPort_10_banks_0(x288_lb_0_io_rPort_10_banks_0),
    .io_rPort_10_ofs_0(x288_lb_0_io_rPort_10_ofs_0),
    .io_rPort_10_en_0(x288_lb_0_io_rPort_10_en_0),
    .io_rPort_10_backpressure(x288_lb_0_io_rPort_10_backpressure),
    .io_rPort_10_output_0(x288_lb_0_io_rPort_10_output_0),
    .io_rPort_9_banks_1(x288_lb_0_io_rPort_9_banks_1),
    .io_rPort_9_banks_0(x288_lb_0_io_rPort_9_banks_0),
    .io_rPort_9_ofs_0(x288_lb_0_io_rPort_9_ofs_0),
    .io_rPort_9_en_0(x288_lb_0_io_rPort_9_en_0),
    .io_rPort_9_backpressure(x288_lb_0_io_rPort_9_backpressure),
    .io_rPort_9_output_0(x288_lb_0_io_rPort_9_output_0),
    .io_rPort_8_banks_1(x288_lb_0_io_rPort_8_banks_1),
    .io_rPort_8_banks_0(x288_lb_0_io_rPort_8_banks_0),
    .io_rPort_8_ofs_0(x288_lb_0_io_rPort_8_ofs_0),
    .io_rPort_8_en_0(x288_lb_0_io_rPort_8_en_0),
    .io_rPort_8_backpressure(x288_lb_0_io_rPort_8_backpressure),
    .io_rPort_8_output_0(x288_lb_0_io_rPort_8_output_0),
    .io_rPort_7_banks_1(x288_lb_0_io_rPort_7_banks_1),
    .io_rPort_7_banks_0(x288_lb_0_io_rPort_7_banks_0),
    .io_rPort_7_ofs_0(x288_lb_0_io_rPort_7_ofs_0),
    .io_rPort_7_en_0(x288_lb_0_io_rPort_7_en_0),
    .io_rPort_7_backpressure(x288_lb_0_io_rPort_7_backpressure),
    .io_rPort_7_output_0(x288_lb_0_io_rPort_7_output_0),
    .io_rPort_6_banks_1(x288_lb_0_io_rPort_6_banks_1),
    .io_rPort_6_banks_0(x288_lb_0_io_rPort_6_banks_0),
    .io_rPort_6_ofs_0(x288_lb_0_io_rPort_6_ofs_0),
    .io_rPort_6_en_0(x288_lb_0_io_rPort_6_en_0),
    .io_rPort_6_backpressure(x288_lb_0_io_rPort_6_backpressure),
    .io_rPort_6_output_0(x288_lb_0_io_rPort_6_output_0),
    .io_rPort_5_banks_1(x288_lb_0_io_rPort_5_banks_1),
    .io_rPort_5_banks_0(x288_lb_0_io_rPort_5_banks_0),
    .io_rPort_5_ofs_0(x288_lb_0_io_rPort_5_ofs_0),
    .io_rPort_5_en_0(x288_lb_0_io_rPort_5_en_0),
    .io_rPort_5_backpressure(x288_lb_0_io_rPort_5_backpressure),
    .io_rPort_5_output_0(x288_lb_0_io_rPort_5_output_0),
    .io_rPort_4_banks_1(x288_lb_0_io_rPort_4_banks_1),
    .io_rPort_4_banks_0(x288_lb_0_io_rPort_4_banks_0),
    .io_rPort_4_ofs_0(x288_lb_0_io_rPort_4_ofs_0),
    .io_rPort_4_en_0(x288_lb_0_io_rPort_4_en_0),
    .io_rPort_4_backpressure(x288_lb_0_io_rPort_4_backpressure),
    .io_rPort_4_output_0(x288_lb_0_io_rPort_4_output_0),
    .io_rPort_3_banks_1(x288_lb_0_io_rPort_3_banks_1),
    .io_rPort_3_banks_0(x288_lb_0_io_rPort_3_banks_0),
    .io_rPort_3_ofs_0(x288_lb_0_io_rPort_3_ofs_0),
    .io_rPort_3_en_0(x288_lb_0_io_rPort_3_en_0),
    .io_rPort_3_backpressure(x288_lb_0_io_rPort_3_backpressure),
    .io_rPort_3_output_0(x288_lb_0_io_rPort_3_output_0),
    .io_rPort_2_banks_1(x288_lb_0_io_rPort_2_banks_1),
    .io_rPort_2_banks_0(x288_lb_0_io_rPort_2_banks_0),
    .io_rPort_2_ofs_0(x288_lb_0_io_rPort_2_ofs_0),
    .io_rPort_2_en_0(x288_lb_0_io_rPort_2_en_0),
    .io_rPort_2_backpressure(x288_lb_0_io_rPort_2_backpressure),
    .io_rPort_2_output_0(x288_lb_0_io_rPort_2_output_0),
    .io_rPort_1_banks_1(x288_lb_0_io_rPort_1_banks_1),
    .io_rPort_1_banks_0(x288_lb_0_io_rPort_1_banks_0),
    .io_rPort_1_ofs_0(x288_lb_0_io_rPort_1_ofs_0),
    .io_rPort_1_en_0(x288_lb_0_io_rPort_1_en_0),
    .io_rPort_1_backpressure(x288_lb_0_io_rPort_1_backpressure),
    .io_rPort_1_output_0(x288_lb_0_io_rPort_1_output_0),
    .io_rPort_0_banks_1(x288_lb_0_io_rPort_0_banks_1),
    .io_rPort_0_banks_0(x288_lb_0_io_rPort_0_banks_0),
    .io_rPort_0_ofs_0(x288_lb_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x288_lb_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x288_lb_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x288_lb_0_io_rPort_0_output_0),
    .io_wPort_1_banks_1(x288_lb_0_io_wPort_1_banks_1),
    .io_wPort_1_banks_0(x288_lb_0_io_wPort_1_banks_0),
    .io_wPort_1_ofs_0(x288_lb_0_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(x288_lb_0_io_wPort_1_data_0),
    .io_wPort_1_en_0(x288_lb_0_io_wPort_1_en_0),
    .io_wPort_0_banks_1(x288_lb_0_io_wPort_0_banks_1),
    .io_wPort_0_banks_0(x288_lb_0_io_wPort_0_banks_0),
    .io_wPort_0_ofs_0(x288_lb_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x288_lb_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x288_lb_0_io_wPort_0_en_0)
  );
  x289_lb2_0 x289_lb2_0 ( // @[m_x289_lb2_0.scala 33:17:@26670.4]
    .clock(x289_lb2_0_clock),
    .reset(x289_lb2_0_reset),
    .io_rPort_5_banks_1(x289_lb2_0_io_rPort_5_banks_1),
    .io_rPort_5_banks_0(x289_lb2_0_io_rPort_5_banks_0),
    .io_rPort_5_ofs_0(x289_lb2_0_io_rPort_5_ofs_0),
    .io_rPort_5_en_0(x289_lb2_0_io_rPort_5_en_0),
    .io_rPort_5_backpressure(x289_lb2_0_io_rPort_5_backpressure),
    .io_rPort_5_output_0(x289_lb2_0_io_rPort_5_output_0),
    .io_rPort_4_banks_1(x289_lb2_0_io_rPort_4_banks_1),
    .io_rPort_4_banks_0(x289_lb2_0_io_rPort_4_banks_0),
    .io_rPort_4_ofs_0(x289_lb2_0_io_rPort_4_ofs_0),
    .io_rPort_4_en_0(x289_lb2_0_io_rPort_4_en_0),
    .io_rPort_4_backpressure(x289_lb2_0_io_rPort_4_backpressure),
    .io_rPort_4_output_0(x289_lb2_0_io_rPort_4_output_0),
    .io_rPort_3_banks_1(x289_lb2_0_io_rPort_3_banks_1),
    .io_rPort_3_banks_0(x289_lb2_0_io_rPort_3_banks_0),
    .io_rPort_3_ofs_0(x289_lb2_0_io_rPort_3_ofs_0),
    .io_rPort_3_en_0(x289_lb2_0_io_rPort_3_en_0),
    .io_rPort_3_backpressure(x289_lb2_0_io_rPort_3_backpressure),
    .io_rPort_3_output_0(x289_lb2_0_io_rPort_3_output_0),
    .io_rPort_2_banks_1(x289_lb2_0_io_rPort_2_banks_1),
    .io_rPort_2_banks_0(x289_lb2_0_io_rPort_2_banks_0),
    .io_rPort_2_ofs_0(x289_lb2_0_io_rPort_2_ofs_0),
    .io_rPort_2_en_0(x289_lb2_0_io_rPort_2_en_0),
    .io_rPort_2_backpressure(x289_lb2_0_io_rPort_2_backpressure),
    .io_rPort_2_output_0(x289_lb2_0_io_rPort_2_output_0),
    .io_rPort_1_banks_1(x289_lb2_0_io_rPort_1_banks_1),
    .io_rPort_1_banks_0(x289_lb2_0_io_rPort_1_banks_0),
    .io_rPort_1_ofs_0(x289_lb2_0_io_rPort_1_ofs_0),
    .io_rPort_1_en_0(x289_lb2_0_io_rPort_1_en_0),
    .io_rPort_1_backpressure(x289_lb2_0_io_rPort_1_backpressure),
    .io_rPort_1_output_0(x289_lb2_0_io_rPort_1_output_0),
    .io_rPort_0_banks_1(x289_lb2_0_io_rPort_0_banks_1),
    .io_rPort_0_banks_0(x289_lb2_0_io_rPort_0_banks_0),
    .io_rPort_0_ofs_0(x289_lb2_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x289_lb2_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x289_lb2_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x289_lb2_0_io_rPort_0_output_0),
    .io_wPort_1_banks_1(x289_lb2_0_io_wPort_1_banks_1),
    .io_wPort_1_banks_0(x289_lb2_0_io_wPort_1_banks_0),
    .io_wPort_1_ofs_0(x289_lb2_0_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(x289_lb2_0_io_wPort_1_data_0),
    .io_wPort_1_en_0(x289_lb2_0_io_wPort_1_en_0),
    .io_wPort_0_banks_1(x289_lb2_0_io_wPort_0_banks_1),
    .io_wPort_0_banks_0(x289_lb2_0_io_wPort_0_banks_0),
    .io_wPort_0_ofs_0(x289_lb2_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x289_lb2_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x289_lb2_0_io_wPort_0_en_0)
  );
  RetimeWrapper_228 RetimeWrapper ( // @[package.scala 93:22:@26740.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x303_sum x303_sum_1 ( // @[Math.scala 150:24:@26847.4]
    .clock(x303_sum_1_clock),
    .reset(x303_sum_1_reset),
    .io_a(x303_sum_1_io_a),
    .io_b(x303_sum_1_io_b),
    .io_flow(x303_sum_1_io_flow),
    .io_result(x303_sum_1_io_result)
  );
  RetimeWrapper_230 RetimeWrapper_1 ( // @[package.scala 93:22:@26857.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_2 ( // @[package.scala 93:22:@26866.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_3 ( // @[package.scala 93:22:@26875.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_229 RetimeWrapper_4 ( // @[package.scala 93:22:@26884.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_5 ( // @[package.scala 93:22:@26893.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_230 RetimeWrapper_6 ( // @[package.scala 93:22:@26902.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_7 ( // @[package.scala 93:22:@26913.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  x303_sum x309_rdcol_1 ( // @[Math.scala 150:24:@26936.4]
    .clock(x309_rdcol_1_clock),
    .reset(x309_rdcol_1_reset),
    .io_a(x309_rdcol_1_io_a),
    .io_b(x309_rdcol_1_io_b),
    .io_flow(x309_rdcol_1_io_flow),
    .io_result(x309_rdcol_1_io_result)
  );
  RetimeWrapper_229 RetimeWrapper_8 ( // @[package.scala 93:22:@26968.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  x303_sum x313_sum_1 ( // @[Math.scala 150:24:@26977.4]
    .clock(x313_sum_1_clock),
    .reset(x313_sum_1_reset),
    .io_a(x313_sum_1_io_a),
    .io_b(x313_sum_1_io_b),
    .io_flow(x313_sum_1_io_flow),
    .io_result(x313_sum_1_io_result)
  );
  RetimeWrapper_229 RetimeWrapper_9 ( // @[package.scala 93:22:@26987.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_10 ( // @[package.scala 93:22:@26996.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_11 ( // @[package.scala 93:22:@27007.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_243 RetimeWrapper_12 ( // @[package.scala 93:22:@27028.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_243 RetimeWrapper_13 ( // @[package.scala 93:22:@27055.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper RetimeWrapper_14 ( // @[package.scala 93:22:@27071.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_243 RetimeWrapper_15 ( // @[package.scala 93:22:@27106.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_229 RetimeWrapper_16 ( // @[package.scala 93:22:@27115.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  x303_sum x326_sum_1 ( // @[Math.scala 150:24:@27124.4]
    .clock(x326_sum_1_clock),
    .reset(x326_sum_1_reset),
    .io_a(x326_sum_1_io_a),
    .io_b(x326_sum_1_io_b),
    .io_flow(x326_sum_1_io_flow),
    .io_result(x326_sum_1_io_result)
  );
  RetimeWrapper_249 RetimeWrapper_17 ( // @[package.scala 93:22:@27134.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_250 RetimeWrapper_18 ( // @[package.scala 93:22:@27143.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper RetimeWrapper_19 ( // @[package.scala 93:22:@27152.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_250 RetimeWrapper_20 ( // @[package.scala 93:22:@27161.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_230 RetimeWrapper_21 ( // @[package.scala 93:22:@27170.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_250 RetimeWrapper_22 ( // @[package.scala 93:22:@27182.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_243 RetimeWrapper_23 ( // @[package.scala 93:22:@27203.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_243 RetimeWrapper_24 ( // @[package.scala 93:22:@27227.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  x303_sum x335_sum_1 ( // @[Math.scala 150:24:@27236.4]
    .clock(x335_sum_1_clock),
    .reset(x335_sum_1_reset),
    .io_a(x335_sum_1_io_a),
    .io_b(x335_sum_1_io_b),
    .io_flow(x335_sum_1_io_flow),
    .io_result(x335_sum_1_io_result)
  );
  RetimeWrapper_52 RetimeWrapper_25 ( // @[package.scala 93:22:@27246.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_259 RetimeWrapper_26 ( // @[package.scala 93:22:@27255.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_229 RetimeWrapper_27 ( // @[package.scala 93:22:@27264.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_250 RetimeWrapper_28 ( // @[package.scala 93:22:@27276.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  x303_sum x340_rdcol_1 ( // @[Math.scala 150:24:@27299.4]
    .clock(x340_rdcol_1_clock),
    .reset(x340_rdcol_1_reset),
    .io_a(x340_rdcol_1_io_a),
    .io_b(x340_rdcol_1_io_b),
    .io_flow(x340_rdcol_1_io_flow),
    .io_result(x340_rdcol_1_io_result)
  );
  x303_sum x346_sum_1 ( // @[Math.scala 150:24:@27342.4]
    .clock(x346_sum_1_clock),
    .reset(x346_sum_1_reset),
    .io_a(x346_sum_1_io_a),
    .io_b(x346_sum_1_io_b),
    .io_flow(x346_sum_1_io_flow),
    .io_result(x346_sum_1_io_result)
  );
  RetimeWrapper_229 RetimeWrapper_29 ( // @[package.scala 93:22:@27352.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper RetimeWrapper_30 ( // @[package.scala 93:22:@27361.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_250 RetimeWrapper_31 ( // @[package.scala 93:22:@27373.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  x303_sum x352_rdcol_1 ( // @[Math.scala 150:24:@27396.4]
    .clock(x352_rdcol_1_clock),
    .reset(x352_rdcol_1_reset),
    .io_a(x352_rdcol_1_io_a),
    .io_b(x352_rdcol_1_io_b),
    .io_flow(x352_rdcol_1_io_flow),
    .io_result(x352_rdcol_1_io_result)
  );
  x303_sum x358_sum_1 ( // @[Math.scala 150:24:@27439.4]
    .clock(x358_sum_1_clock),
    .reset(x358_sum_1_reset),
    .io_a(x358_sum_1_io_a),
    .io_b(x358_sum_1_io_b),
    .io_flow(x358_sum_1_io_flow),
    .io_result(x358_sum_1_io_result)
  );
  RetimeWrapper_229 RetimeWrapper_32 ( // @[package.scala 93:22:@27449.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper RetimeWrapper_33 ( // @[package.scala 93:22:@27458.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_250 RetimeWrapper_34 ( // @[package.scala 93:22:@27470.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  x364_rdrow x364_rdrow_1 ( // @[Math.scala 191:24:@27493.4]
    .clock(x364_rdrow_1_clock),
    .reset(x364_rdrow_1_reset),
    .io_a(x364_rdrow_1_io_a),
    .io_b(x364_rdrow_1_io_b),
    .io_flow(x364_rdrow_1_io_flow),
    .io_result(x364_rdrow_1_io_result)
  );
  x303_sum x371_sum_1 ( // @[Math.scala 150:24:@27547.4]
    .clock(x371_sum_1_clock),
    .reset(x371_sum_1_reset),
    .io_a(x371_sum_1_io_a),
    .io_b(x371_sum_1_io_b),
    .io_flow(x371_sum_1_io_flow),
    .io_result(x371_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_35 ( // @[package.scala 93:22:@27557.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_229 RetimeWrapper_36 ( // @[package.scala 93:22:@27566.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_250 RetimeWrapper_37 ( // @[package.scala 93:22:@27578.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper RetimeWrapper_38 ( // @[package.scala 93:22:@27599.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_249 RetimeWrapper_39 ( // @[package.scala 93:22:@27614.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  x303_sum x379_sum_1 ( // @[Math.scala 150:24:@27625.4]
    .clock(x379_sum_1_clock),
    .reset(x379_sum_1_reset),
    .io_a(x379_sum_1_io_a),
    .io_b(x379_sum_1_io_b),
    .io_flow(x379_sum_1_io_flow),
    .io_result(x379_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_40 ( // @[package.scala 93:22:@27635.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper_250 RetimeWrapper_41 ( // @[package.scala 93:22:@27647.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  x303_sum x386_sum_1 ( // @[Math.scala 150:24:@27674.4]
    .clock(x386_sum_1_clock),
    .reset(x386_sum_1_reset),
    .io_a(x386_sum_1_io_a),
    .io_b(x386_sum_1_io_b),
    .io_flow(x386_sum_1_io_flow),
    .io_result(x386_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_42 ( // @[package.scala 93:22:@27684.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_250 RetimeWrapper_43 ( // @[package.scala 93:22:@27696.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  x303_sum x393_sum_1 ( // @[Math.scala 150:24:@27723.4]
    .clock(x393_sum_1_clock),
    .reset(x393_sum_1_reset),
    .io_a(x393_sum_1_io_a),
    .io_b(x393_sum_1_io_b),
    .io_flow(x393_sum_1_io_flow),
    .io_result(x393_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_44 ( // @[package.scala 93:22:@27733.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_250 RetimeWrapper_45 ( // @[package.scala 93:22:@27745.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  x364_rdrow x398_rdrow_1 ( // @[Math.scala 191:24:@27768.4]
    .clock(x398_rdrow_1_clock),
    .reset(x398_rdrow_1_reset),
    .io_a(x398_rdrow_1_io_a),
    .io_b(x398_rdrow_1_io_b),
    .io_flow(x398_rdrow_1_io_flow),
    .io_result(x398_rdrow_1_io_result)
  );
  x303_sum x405_sum_1 ( // @[Math.scala 150:24:@27822.4]
    .clock(x405_sum_1_clock),
    .reset(x405_sum_1_reset),
    .io_a(x405_sum_1_io_a),
    .io_b(x405_sum_1_io_b),
    .io_flow(x405_sum_1_io_flow),
    .io_result(x405_sum_1_io_result)
  );
  RetimeWrapper_229 RetimeWrapper_46 ( // @[package.scala 93:22:@27832.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper RetimeWrapper_47 ( // @[package.scala 93:22:@27841.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_250 RetimeWrapper_48 ( // @[package.scala 93:22:@27853.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  x303_sum x413_sum_1 ( // @[Math.scala 150:24:@27880.4]
    .clock(x413_sum_1_clock),
    .reset(x413_sum_1_reset),
    .io_a(x413_sum_1_io_a),
    .io_b(x413_sum_1_io_b),
    .io_flow(x413_sum_1_io_flow),
    .io_result(x413_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_49 ( // @[package.scala 93:22:@27890.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_250 RetimeWrapper_50 ( // @[package.scala 93:22:@27902.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  x303_sum x420_sum_1 ( // @[Math.scala 150:24:@27929.4]
    .clock(x420_sum_1_clock),
    .reset(x420_sum_1_reset),
    .io_a(x420_sum_1_io_a),
    .io_b(x420_sum_1_io_b),
    .io_flow(x420_sum_1_io_flow),
    .io_result(x420_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_51 ( // @[package.scala 93:22:@27939.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_250 RetimeWrapper_52 ( // @[package.scala 93:22:@27951.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  x303_sum x427_sum_1 ( // @[Math.scala 150:24:@27978.4]
    .clock(x427_sum_1_clock),
    .reset(x427_sum_1_reset),
    .io_a(x427_sum_1_io_a),
    .io_b(x427_sum_1_io_b),
    .io_flow(x427_sum_1_io_flow),
    .io_result(x427_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_53 ( // @[package.scala 93:22:@27988.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper_250 RetimeWrapper_54 ( // @[package.scala 93:22:@28000.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  x437_x23 x437_x23_1 ( // @[Math.scala 150:24:@28048.4]
    .clock(x437_x23_1_clock),
    .reset(x437_x23_1_reset),
    .io_a(x437_x23_1_io_a),
    .io_b(x437_x23_1_io_b),
    .io_flow(x437_x23_1_io_flow),
    .io_result(x437_x23_1_io_result)
  );
  x437_x23 x438_x24_1 ( // @[Math.scala 150:24:@28058.4]
    .clock(x438_x24_1_clock),
    .reset(x438_x24_1_reset),
    .io_a(x438_x24_1_io_a),
    .io_b(x438_x24_1_io_b),
    .io_flow(x438_x24_1_io_flow),
    .io_result(x438_x24_1_io_result)
  );
  x437_x23 x439_x23_1 ( // @[Math.scala 150:24:@28068.4]
    .clock(x439_x23_1_clock),
    .reset(x439_x23_1_reset),
    .io_a(x439_x23_1_io_a),
    .io_b(x439_x23_1_io_b),
    .io_flow(x439_x23_1_io_flow),
    .io_result(x439_x23_1_io_result)
  );
  x437_x23 x440_x24_1 ( // @[Math.scala 150:24:@28078.4]
    .clock(x440_x24_1_clock),
    .reset(x440_x24_1_reset),
    .io_a(x440_x24_1_io_a),
    .io_b(x440_x24_1_io_b),
    .io_flow(x440_x24_1_io_flow),
    .io_result(x440_x24_1_io_result)
  );
  x441_x23 x441_x23_1 ( // @[Math.scala 150:24:@28088.4]
    .io_a(x441_x23_1_io_a),
    .io_b(x441_x23_1_io_b),
    .io_result(x441_x23_1_io_result)
  );
  x441_x23 x442_x24_1 ( // @[Math.scala 150:24:@28098.4]
    .io_a(x442_x24_1_io_a),
    .io_b(x442_x24_1_io_b),
    .io_result(x442_x24_1_io_result)
  );
  x441_x23 x443_x23_1 ( // @[Math.scala 150:24:@28108.4]
    .io_a(x443_x23_1_io_a),
    .io_b(x443_x23_1_io_b),
    .io_result(x443_x23_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_55 ( // @[package.scala 93:22:@28118.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  x441_x23 x444_sum_1 ( // @[Math.scala 150:24:@28127.4]
    .io_a(x444_sum_1_io_a),
    .io_b(x444_sum_1_io_b),
    .io_result(x444_sum_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_56 ( // @[package.scala 93:22:@28141.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  x437_x23 x451_x23_1 ( // @[Math.scala 150:24:@28176.4]
    .clock(x451_x23_1_clock),
    .reset(x451_x23_1_reset),
    .io_a(x451_x23_1_io_a),
    .io_b(x451_x23_1_io_b),
    .io_flow(x451_x23_1_io_flow),
    .io_result(x451_x23_1_io_result)
  );
  x437_x23 x452_x24_1 ( // @[Math.scala 150:24:@28186.4]
    .clock(x452_x24_1_clock),
    .reset(x452_x24_1_reset),
    .io_a(x452_x24_1_io_a),
    .io_b(x452_x24_1_io_b),
    .io_flow(x452_x24_1_io_flow),
    .io_result(x452_x24_1_io_result)
  );
  x437_x23 x453_x23_1 ( // @[Math.scala 150:24:@28196.4]
    .clock(x453_x23_1_clock),
    .reset(x453_x23_1_reset),
    .io_a(x453_x23_1_io_a),
    .io_b(x453_x23_1_io_b),
    .io_flow(x453_x23_1_io_flow),
    .io_result(x453_x23_1_io_result)
  );
  x437_x23 x454_x24_1 ( // @[Math.scala 150:24:@28206.4]
    .clock(x454_x24_1_clock),
    .reset(x454_x24_1_reset),
    .io_a(x454_x24_1_io_a),
    .io_b(x454_x24_1_io_b),
    .io_flow(x454_x24_1_io_flow),
    .io_result(x454_x24_1_io_result)
  );
  x441_x23 x455_x23_1 ( // @[Math.scala 150:24:@28216.4]
    .io_a(x455_x23_1_io_a),
    .io_b(x455_x23_1_io_b),
    .io_result(x455_x23_1_io_result)
  );
  x441_x23 x456_x24_1 ( // @[Math.scala 150:24:@28226.4]
    .io_a(x456_x24_1_io_a),
    .io_b(x456_x24_1_io_b),
    .io_result(x456_x24_1_io_result)
  );
  x441_x23 x457_x23_1 ( // @[Math.scala 150:24:@28236.4]
    .io_a(x457_x23_1_io_a),
    .io_b(x457_x23_1_io_b),
    .io_result(x457_x23_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_57 ( // @[package.scala 93:22:@28246.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  x441_x23 x458_sum_1 ( // @[Math.scala 150:24:@28255.4]
    .io_a(x458_sum_1_io_a),
    .io_b(x458_sum_1_io_b),
    .io_result(x458_sum_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_58 ( // @[package.scala 93:22:@28269.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_314 RetimeWrapper_59 ( // @[package.scala 93:22:@28279.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_315 RetimeWrapper_60 ( // @[package.scala 93:22:@28288.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_316 RetimeWrapper_61 ( // @[package.scala 93:22:@28297.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  RetimeWrapper_315 RetimeWrapper_62 ( // @[package.scala 93:22:@28306.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_314 RetimeWrapper_63 ( // @[package.scala 93:22:@28315.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  RetimeWrapper_315 RetimeWrapper_64 ( // @[package.scala 93:22:@28326.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_316 RetimeWrapper_65 ( // @[package.scala 93:22:@28347.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper_321 RetimeWrapper_66 ( // @[package.scala 93:22:@28356.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper_315 RetimeWrapper_67 ( // @[package.scala 93:22:@28367.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  RetimeWrapper_323 RetimeWrapper_68 ( // @[package.scala 93:22:@28388.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_259 RetimeWrapper_69 ( // @[package.scala 93:22:@28397.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  RetimeWrapper_243 RetimeWrapper_70 ( // @[package.scala 93:22:@28406.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_315 RetimeWrapper_71 ( // @[package.scala 93:22:@28418.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  RetimeWrapper_250 RetimeWrapper_72 ( // @[package.scala 93:22:@28439.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  RetimeWrapper_249 RetimeWrapper_73 ( // @[package.scala 93:22:@28448.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  RetimeWrapper_315 RetimeWrapper_74 ( // @[package.scala 93:22:@28460.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  RetimeWrapper_249 RetimeWrapper_75 ( // @[package.scala 93:22:@28481.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_323 RetimeWrapper_76 ( // @[package.scala 93:22:@28490.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  RetimeWrapper_243 RetimeWrapper_77 ( // @[package.scala 93:22:@28499.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  RetimeWrapper_315 RetimeWrapper_78 ( // @[package.scala 93:22:@28511.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  RetimeWrapper_243 RetimeWrapper_79 ( // @[package.scala 93:22:@28532.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper_323 RetimeWrapper_80 ( // @[package.scala 93:22:@28541.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  RetimeWrapper_249 RetimeWrapper_81 ( // @[package.scala 93:22:@28550.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_315 RetimeWrapper_82 ( // @[package.scala 93:22:@28562.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  RetimeWrapper_243 RetimeWrapper_83 ( // @[package.scala 93:22:@28583.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  RetimeWrapper_323 RetimeWrapper_84 ( // @[package.scala 93:22:@28592.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  RetimeWrapper_315 RetimeWrapper_85 ( // @[package.scala 93:22:@28604.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  RetimeWrapper_323 RetimeWrapper_86 ( // @[package.scala 93:22:@28625.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  RetimeWrapper_243 RetimeWrapper_87 ( // @[package.scala 93:22:@28634.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  RetimeWrapper_315 RetimeWrapper_88 ( // @[package.scala 93:22:@28646.4]
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  x441_x23 x478_x25_1 ( // @[Math.scala 150:24:@28679.4]
    .io_a(x478_x25_1_io_a),
    .io_b(x478_x25_1_io_b),
    .io_result(x478_x25_1_io_result)
  );
  x441_x23 x479_x26_1 ( // @[Math.scala 150:24:@28689.4]
    .io_a(x479_x26_1_io_a),
    .io_b(x479_x26_1_io_b),
    .io_result(x479_x26_1_io_result)
  );
  x441_x23 x480_sum_1 ( // @[Math.scala 150:24:@28699.4]
    .io_a(x480_sum_1_io_a),
    .io_b(x480_sum_1_io_b),
    .io_result(x480_sum_1_io_result)
  );
  x481_div x481_div_1 ( // @[Math.scala 327:24:@28711.4]
    .clock(x481_div_1_clock),
    .reset(x481_div_1_reset),
    .io_a(x481_div_1_io_a),
    .io_flow(x481_div_1_io_flow),
    .io_result(x481_div_1_io_result)
  );
  x441_x23 x484_x25_1 ( // @[Math.scala 150:24:@28731.4]
    .io_a(x484_x25_1_io_a),
    .io_b(x484_x25_1_io_b),
    .io_result(x484_x25_1_io_result)
  );
  x441_x23 x485_x26_1 ( // @[Math.scala 150:24:@28741.4]
    .io_a(x485_x26_1_io_a),
    .io_b(x485_x26_1_io_b),
    .io_result(x485_x26_1_io_result)
  );
  x441_x23 x486_sum_1 ( // @[Math.scala 150:24:@28751.4]
    .io_a(x486_sum_1_io_a),
    .io_b(x486_sum_1_io_b),
    .io_result(x486_sum_1_io_result)
  );
  x481_div x487_div_1 ( // @[Math.scala 327:24:@28763.4]
    .clock(x487_div_1_clock),
    .reset(x487_div_1_reset),
    .io_a(x487_div_1_io_a),
    .io_flow(x487_div_1_io_flow),
    .io_result(x487_div_1_io_result)
  );
  RetimeWrapper_346 RetimeWrapper_89 ( // @[package.scala 93:22:@28779.4]
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  RetimeWrapper_347 RetimeWrapper_90 ( // @[package.scala 93:22:@28788.4]
    .clock(RetimeWrapper_90_clock),
    .reset(RetimeWrapper_90_reset),
    .io_flow(RetimeWrapper_90_io_flow),
    .io_in(RetimeWrapper_90_io_in),
    .io_out(RetimeWrapper_90_io_out)
  );
  RetimeWrapper_347 RetimeWrapper_91 ( // @[package.scala 93:22:@28797.4]
    .clock(RetimeWrapper_91_clock),
    .reset(RetimeWrapper_91_reset),
    .io_flow(RetimeWrapper_91_io_flow),
    .io_in(RetimeWrapper_91_io_in),
    .io_out(RetimeWrapper_91_io_out)
  );
  RetimeWrapper_347 RetimeWrapper_92 ( // @[package.scala 93:22:@28806.4]
    .clock(RetimeWrapper_92_clock),
    .reset(RetimeWrapper_92_reset),
    .io_flow(RetimeWrapper_92_io_flow),
    .io_in(RetimeWrapper_92_io_in),
    .io_out(RetimeWrapper_92_io_out)
  );
  assign b286 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 62:18:@26575.4]
  assign b287 = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 63:18:@26576.4]
  assign _T_207 = b286 & b287; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 69:30:@26728.4]
  assign _T_208 = _T_207 & io_sigsIn_datapathEn; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 69:37:@26729.4]
  assign _T_212 = io_in_x275_TID == 8'h0; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 71:76:@26734.4]
  assign _T_213 = _T_208 & _T_212; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 71:62:@26735.4]
  assign _T_215 = io_in_x275_TDEST == 8'h0; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 71:101:@26736.4]
  assign x571_x290_D1_0_number = RetimeWrapper_io_out; // @[package.scala 96:25:@26745.4 package.scala 96:25:@26746.4]
  assign b284_number = __io_result; // @[Math.scala 712:22:@26560.4 Math.scala 713:14:@26561.4]
  assign _T_243 = $signed(b284_number); // @[Math.scala 499:52:@26761.4]
  assign x294 = $signed(32'sh1) == $signed(_T_243); // @[Math.scala 499:44:@26769.4]
  assign x295 = $signed(32'sh2) == $signed(_T_243); // @[Math.scala 499:44:@26776.4]
  assign x296 = $signed(32'sh3) == $signed(_T_243); // @[Math.scala 499:44:@26783.4]
  assign _T_290 = x294 ? 32'h1 : 32'h0; // @[Mux.scala 19:72:@26795.4]
  assign _T_292 = x295 ? 32'h2 : 32'h0; // @[Mux.scala 19:72:@26796.4]
  assign _T_294 = x296 ? 32'h3 : 32'h0; // @[Mux.scala 19:72:@26797.4]
  assign _T_296 = _T_290 | _T_292; // @[Mux.scala 19:72:@26799.4]
  assign x297_number = _T_296 | _T_294; // @[Mux.scala 19:72:@26800.4]
  assign _T_308 = $signed(x297_number); // @[Math.scala 406:49:@26810.4]
  assign _T_310 = $signed(_T_308) & $signed(32'sh3); // @[Math.scala 406:56:@26812.4]
  assign _T_311 = $signed(_T_310); // @[Math.scala 406:56:@26813.4]
  assign b285_number = __1_io_result; // @[Math.scala 712:22:@26572.4 Math.scala 713:14:@26573.4]
  assign _T_320 = $signed(b285_number); // @[Math.scala 406:49:@26821.4]
  assign _T_322 = $signed(_T_320) & $signed(32'sh3); // @[Math.scala 406:56:@26823.4]
  assign _T_323 = $signed(_T_322); // @[Math.scala 406:56:@26824.4]
  assign _T_328 = x297_number[31]; // @[FixedPoint.scala 50:25:@26830.4]
  assign _T_332 = _T_328 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@26832.4]
  assign _T_333 = x297_number[31:2]; // @[FixedPoint.scala 18:52:@26833.4]
  assign _T_338 = b285_number[31]; // @[FixedPoint.scala 50:25:@26839.4]
  assign _T_342 = _T_338 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@26841.4]
  assign _T_343 = b285_number[31:2]; // @[FixedPoint.scala 18:52:@26842.4]
  assign _T_367 = ~ io_sigsIn_break; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 118:101:@26910.4]
  assign _T_371 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@26918.4 package.scala 96:25:@26919.4]
  assign _T_373 = io_rr ? _T_371 : 1'h0; // @[implicits.scala 55:10:@26920.4]
  assign _T_374 = _T_367 & _T_373; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 118:118:@26921.4]
  assign _T_376 = _T_374 & _T_367; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 118:205:@26923.4]
  assign _T_377 = _T_376 & io_sigsIn_backpressure; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 118:224:@26924.4]
  assign x574_b286_D2 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@26880.4 package.scala 96:25:@26881.4]
  assign _T_378 = _T_377 & x574_b286_D2; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 118:250:@26925.4]
  assign x576_b287_D2 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@26898.4 package.scala 96:25:@26899.4]
  assign x309_rdcol_number = x309_rdcol_1_io_result; // @[Math.scala 154:22:@26942.4 Math.scala 155:14:@26943.4]
  assign _T_395 = $signed(x309_rdcol_number); // @[Math.scala 406:49:@26951.4]
  assign _T_397 = $signed(_T_395) & $signed(32'sh3); // @[Math.scala 406:56:@26953.4]
  assign _T_398 = $signed(_T_397); // @[Math.scala 406:56:@26954.4]
  assign _T_403 = x309_rdcol_number[31]; // @[FixedPoint.scala 50:25:@26960.4]
  assign _T_407 = _T_403 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@26962.4]
  assign _T_408 = x309_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@26963.4]
  assign _T_427 = RetimeWrapper_11_io_out; // @[package.scala 96:25:@27012.4 package.scala 96:25:@27013.4]
  assign _T_429 = io_rr ? _T_427 : 1'h0; // @[implicits.scala 55:10:@27014.4]
  assign _T_430 = _T_367 & _T_429; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 139:118:@27015.4]
  assign _T_432 = _T_430 & _T_367; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 139:205:@27017.4]
  assign _T_433 = _T_432 & io_sigsIn_backpressure; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 139:224:@27018.4]
  assign _T_434 = _T_433 & x574_b286_D2; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 139:250:@27019.4]
  assign x581_b284_D4_number = RetimeWrapper_12_io_out; // @[package.scala 96:25:@27033.4 package.scala 96:25:@27034.4]
  assign _T_446 = $signed(x581_b284_D4_number); // @[Math.scala 406:49:@27040.4]
  assign _T_448 = $signed(_T_446) & $signed(32'sh3); // @[Math.scala 406:56:@27042.4]
  assign _T_449 = $signed(_T_448); // @[Math.scala 406:56:@27043.4]
  assign x563_number = $unsigned(_T_449); // @[implicits.scala 133:21:@27044.4]
  assign x320 = $signed(_T_446) < $signed(32'sh0); // @[Math.scala 465:44:@27052.4]
  assign x582_x309_rdcol_D4_number = RetimeWrapper_13_io_out; // @[package.scala 96:25:@27060.4 package.scala 96:25:@27061.4]
  assign _T_467 = $signed(x582_x309_rdcol_D4_number); // @[Math.scala 465:37:@27066.4]
  assign x321 = $signed(_T_467) < $signed(32'sh0); // @[Math.scala 465:44:@27068.4]
  assign x583_x320_D1 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@27076.4 package.scala 96:25:@27077.4]
  assign x322 = x583_x320_D1 | x321; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 154:24:@27080.4]
  assign _T_484 = $signed(x563_number); // @[Math.scala 406:49:@27089.4]
  assign _T_486 = $signed(_T_484) & $signed(32'sh3); // @[Math.scala 406:56:@27091.4]
  assign _T_487 = $signed(_T_486); // @[Math.scala 406:56:@27092.4]
  assign _T_492 = x563_number[31]; // @[FixedPoint.scala 50:25:@27098.4]
  assign _T_496 = _T_492 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@27100.4]
  assign _T_497 = x563_number[31:2]; // @[FixedPoint.scala 18:52:@27101.4]
  assign _T_534 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@27187.4 package.scala 96:25:@27188.4]
  assign _T_536 = io_rr ? _T_534 : 1'h0; // @[implicits.scala 55:10:@27189.4]
  assign _T_537 = _T_367 & _T_536; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 187:194:@27190.4]
  assign x588_x323_D1 = RetimeWrapper_19_io_out; // @[package.scala 96:25:@27157.4 package.scala 96:25:@27158.4]
  assign _T_538 = _T_537 & x588_x323_D1; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 187:281:@27191.4]
  assign x587_b286_D6 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@27148.4 package.scala 96:25:@27149.4]
  assign _T_539 = _T_538 & x587_b286_D6; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 187:289:@27192.4]
  assign x589_b287_D6 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@27166.4 package.scala 96:25:@27167.4]
  assign x591_b285_D4_number = RetimeWrapper_23_io_out; // @[package.scala 96:25:@27208.4 package.scala 96:25:@27209.4]
  assign _T_552 = $signed(x591_b285_D4_number); // @[Math.scala 465:37:@27216.4]
  assign x332 = $signed(_T_552) < $signed(32'sh0); // @[Math.scala 465:44:@27218.4]
  assign x333 = x320 | x332; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 197:59:@27221.4]
  assign _T_585 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@27281.4 package.scala 96:25:@27282.4]
  assign _T_587 = io_rr ? _T_585 : 1'h0; // @[implicits.scala 55:10:@27283.4]
  assign _T_588 = _T_367 & _T_587; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 214:194:@27284.4]
  assign x593_x334_D2 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@27251.4 package.scala 96:25:@27252.4]
  assign _T_589 = _T_588 & x593_x334_D2; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 214:281:@27285.4]
  assign _T_590 = _T_589 & x587_b286_D6; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 214:289:@27286.4]
  assign x340_rdcol_number = x340_rdcol_1_io_result; // @[Math.scala 154:22:@27305.4 Math.scala 155:14:@27306.4]
  assign _T_605 = $signed(x340_rdcol_number); // @[Math.scala 465:37:@27311.4]
  assign x341 = $signed(_T_605) < $signed(32'sh0); // @[Math.scala 465:44:@27313.4]
  assign x342 = x583_x320_D1 | x341; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 222:59:@27316.4]
  assign _T_621 = $signed(_T_605) & $signed(32'sh3); // @[Math.scala 406:56:@27327.4]
  assign _T_622 = $signed(_T_621); // @[Math.scala 406:56:@27328.4]
  assign _T_627 = x340_rdcol_number[31]; // @[FixedPoint.scala 50:25:@27334.4]
  assign _T_631 = _T_627 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@27336.4]
  assign _T_632 = x340_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@27337.4]
  assign _T_654 = RetimeWrapper_31_io_out; // @[package.scala 96:25:@27378.4 package.scala 96:25:@27379.4]
  assign _T_656 = io_rr ? _T_654 : 1'h0; // @[implicits.scala 55:10:@27380.4]
  assign _T_657 = _T_367 & _T_656; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 239:194:@27381.4]
  assign x597_x343_D1 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@27366.4 package.scala 96:25:@27367.4]
  assign _T_658 = _T_657 & x597_x343_D1; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 239:281:@27382.4]
  assign _T_659 = _T_658 & x587_b286_D6; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 239:289:@27383.4]
  assign x352_rdcol_number = x352_rdcol_1_io_result; // @[Math.scala 154:22:@27402.4 Math.scala 155:14:@27403.4]
  assign _T_674 = $signed(x352_rdcol_number); // @[Math.scala 465:37:@27408.4]
  assign x353 = $signed(_T_674) < $signed(32'sh0); // @[Math.scala 465:44:@27410.4]
  assign x354 = x583_x320_D1 | x353; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 247:59:@27413.4]
  assign _T_690 = $signed(_T_674) & $signed(32'sh3); // @[Math.scala 406:56:@27424.4]
  assign _T_691 = $signed(_T_690); // @[Math.scala 406:56:@27425.4]
  assign _T_696 = x352_rdcol_number[31]; // @[FixedPoint.scala 50:25:@27431.4]
  assign _T_700 = _T_696 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@27433.4]
  assign _T_701 = x352_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@27434.4]
  assign _T_723 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@27475.4 package.scala 96:25:@27476.4]
  assign _T_725 = io_rr ? _T_723 : 1'h0; // @[implicits.scala 55:10:@27477.4]
  assign _T_726 = _T_367 & _T_725; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 264:194:@27478.4]
  assign x599_x355_D1 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@27463.4 package.scala 96:25:@27464.4]
  assign _T_727 = _T_726 & x599_x355_D1; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 264:281:@27479.4]
  assign _T_728 = _T_727 & x587_b286_D6; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 264:289:@27480.4]
  assign x364_rdrow_number = x364_rdrow_1_io_result; // @[Math.scala 195:22:@27499.4 Math.scala 196:14:@27500.4]
  assign _T_745 = $signed(x364_rdrow_number); // @[Math.scala 406:49:@27506.4]
  assign _T_747 = $signed(_T_745) & $signed(32'sh3); // @[Math.scala 406:56:@27508.4]
  assign _T_748 = $signed(_T_747); // @[Math.scala 406:56:@27509.4]
  assign x567_number = $unsigned(_T_748); // @[implicits.scala 133:21:@27510.4]
  assign x366 = $signed(_T_745) < $signed(32'sh0); // @[Math.scala 465:44:@27518.4]
  assign x367 = x366 | x321; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 274:24:@27521.4]
  assign _T_769 = $signed(x567_number); // @[Math.scala 406:49:@27530.4]
  assign _T_771 = $signed(_T_769) & $signed(32'sh3); // @[Math.scala 406:56:@27532.4]
  assign _T_772 = $signed(_T_771); // @[Math.scala 406:56:@27533.4]
  assign _T_777 = x567_number[31]; // @[FixedPoint.scala 50:25:@27539.4]
  assign _T_781 = _T_777 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@27541.4]
  assign _T_782 = x567_number[31:2]; // @[FixedPoint.scala 18:52:@27542.4]
  assign _T_804 = RetimeWrapper_37_io_out; // @[package.scala 96:25:@27583.4 package.scala 96:25:@27584.4]
  assign _T_806 = io_rr ? _T_804 : 1'h0; // @[implicits.scala 55:10:@27585.4]
  assign _T_807 = _T_367 & _T_806; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 291:194:@27586.4]
  assign x600_x368_D1 = RetimeWrapper_35_io_out; // @[package.scala 96:25:@27562.4 package.scala 96:25:@27563.4]
  assign _T_808 = _T_807 & x600_x368_D1; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 291:281:@27587.4]
  assign _T_809 = _T_808 & x587_b286_D6; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 291:289:@27588.4]
  assign x602_x332_D1 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@27604.4 package.scala 96:25:@27605.4]
  assign x377 = x366 | x602_x332_D1; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 303:59:@27608.4]
  assign _T_841 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@27652.4 package.scala 96:25:@27653.4]
  assign _T_843 = io_rr ? _T_841 : 1'h0; // @[implicits.scala 55:10:@27654.4]
  assign _T_844 = _T_367 & _T_843; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 318:194:@27655.4]
  assign x604_x378_D1 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@27640.4 package.scala 96:25:@27641.4]
  assign _T_845 = _T_844 & x604_x378_D1; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 318:281:@27656.4]
  assign _T_846 = _T_845 & x587_b286_D6; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 318:289:@27657.4]
  assign x384 = x366 | x341; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 322:59:@27668.4]
  assign _T_870 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@27701.4 package.scala 96:25:@27702.4]
  assign _T_872 = io_rr ? _T_870 : 1'h0; // @[implicits.scala 55:10:@27703.4]
  assign _T_873 = _T_367 & _T_872; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 333:194:@27704.4]
  assign x605_x385_D1 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@27689.4 package.scala 96:25:@27690.4]
  assign _T_874 = _T_873 & x605_x385_D1; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 333:281:@27705.4]
  assign _T_875 = _T_874 & x587_b286_D6; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 333:289:@27706.4]
  assign x391 = x366 | x353; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 337:59:@27717.4]
  assign _T_899 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@27750.4 package.scala 96:25:@27751.4]
  assign _T_901 = io_rr ? _T_899 : 1'h0; // @[implicits.scala 55:10:@27752.4]
  assign _T_902 = _T_367 & _T_901; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 348:194:@27753.4]
  assign x606_x392_D1 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@27738.4 package.scala 96:25:@27739.4]
  assign _T_903 = _T_902 & x606_x392_D1; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 348:281:@27754.4]
  assign _T_904 = _T_903 & x587_b286_D6; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 348:289:@27755.4]
  assign x398_rdrow_number = x398_rdrow_1_io_result; // @[Math.scala 195:22:@27774.4 Math.scala 196:14:@27775.4]
  assign _T_921 = $signed(x398_rdrow_number); // @[Math.scala 406:49:@27781.4]
  assign _T_923 = $signed(_T_921) & $signed(32'sh3); // @[Math.scala 406:56:@27783.4]
  assign _T_924 = $signed(_T_923); // @[Math.scala 406:56:@27784.4]
  assign x569_number = $unsigned(_T_924); // @[implicits.scala 133:21:@27785.4]
  assign x400 = $signed(_T_921) < $signed(32'sh0); // @[Math.scala 465:44:@27793.4]
  assign x401 = x400 | x321; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 358:24:@27796.4]
  assign _T_945 = $signed(x569_number); // @[Math.scala 406:49:@27805.4]
  assign _T_947 = $signed(_T_945) & $signed(32'sh3); // @[Math.scala 406:56:@27807.4]
  assign _T_948 = $signed(_T_947); // @[Math.scala 406:56:@27808.4]
  assign _T_953 = x569_number[31]; // @[FixedPoint.scala 50:25:@27814.4]
  assign _T_957 = _T_953 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@27816.4]
  assign _T_958 = x569_number[31:2]; // @[FixedPoint.scala 18:52:@27817.4]
  assign _T_980 = RetimeWrapper_48_io_out; // @[package.scala 96:25:@27858.4 package.scala 96:25:@27859.4]
  assign _T_982 = io_rr ? _T_980 : 1'h0; // @[implicits.scala 55:10:@27860.4]
  assign _T_983 = _T_367 & _T_982; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 375:194:@27861.4]
  assign x608_x402_D1 = RetimeWrapper_47_io_out; // @[package.scala 96:25:@27846.4 package.scala 96:25:@27847.4]
  assign _T_984 = _T_983 & x608_x402_D1; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 375:281:@27862.4]
  assign _T_985 = _T_984 & x587_b286_D6; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 375:289:@27863.4]
  assign x411 = x400 | x602_x332_D1; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 379:24:@27874.4]
  assign _T_1009 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@27907.4 package.scala 96:25:@27908.4]
  assign _T_1011 = io_rr ? _T_1009 : 1'h0; // @[implicits.scala 55:10:@27909.4]
  assign _T_1012 = _T_367 & _T_1011; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 390:194:@27910.4]
  assign x609_x412_D1 = RetimeWrapper_49_io_out; // @[package.scala 96:25:@27895.4 package.scala 96:25:@27896.4]
  assign _T_1013 = _T_1012 & x609_x412_D1; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 390:281:@27911.4]
  assign _T_1014 = _T_1013 & x587_b286_D6; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 390:289:@27912.4]
  assign x418 = x400 | x341; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 394:24:@27923.4]
  assign _T_1038 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@27956.4 package.scala 96:25:@27957.4]
  assign _T_1040 = io_rr ? _T_1038 : 1'h0; // @[implicits.scala 55:10:@27958.4]
  assign _T_1041 = _T_367 & _T_1040; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 405:194:@27959.4]
  assign x610_x419_D1 = RetimeWrapper_51_io_out; // @[package.scala 96:25:@27944.4 package.scala 96:25:@27945.4]
  assign _T_1042 = _T_1041 & x610_x419_D1; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 405:281:@27960.4]
  assign _T_1043 = _T_1042 & x587_b286_D6; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 405:289:@27961.4]
  assign x425 = x400 | x353; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 409:24:@27972.4]
  assign _T_1067 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@28005.4 package.scala 96:25:@28006.4]
  assign _T_1069 = io_rr ? _T_1067 : 1'h0; // @[implicits.scala 55:10:@28007.4]
  assign _T_1070 = _T_367 & _T_1069; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 426:194:@28008.4]
  assign x611_x426_D1 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@27993.4 package.scala 96:25:@27994.4]
  assign _T_1071 = _T_1070 & x611_x426_D1; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 426:281:@28009.4]
  assign _T_1072 = _T_1071 & x587_b286_D6; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 426:324:@28010.4]
  assign x338_rd_0_number = x288_lb_0_io_rPort_11_output_0; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 210:29:@27272.4 sm_x492_inr_Foreach_SAMPLER_BOX.scala 214:371:@27293.4]
  assign _GEN_0 = {{1'd0}, x338_rd_0_number}; // @[Math.scala 450:32:@28024.4]
  assign _T_1080 = _GEN_0 << 1; // @[Math.scala 450:32:@28024.4]
  assign x375_rd_0_number = x288_lb_0_io_rPort_4_output_0; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 287:29:@27574.4 sm_x492_inr_Foreach_SAMPLER_BOX.scala 291:371:@27595.4]
  assign _GEN_1 = {{1'd0}, x375_rd_0_number}; // @[Math.scala 450:32:@28029.4]
  assign _T_1084 = _GEN_1 << 1; // @[Math.scala 450:32:@28029.4]
  assign x382_rd_0_number = x288_lb_0_io_rPort_6_output_0; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 314:29:@27643.4 sm_x492_inr_Foreach_SAMPLER_BOX.scala 318:406:@27664.4]
  assign _GEN_2 = {{2'd0}, x382_rd_0_number}; // @[Math.scala 450:32:@28034.4]
  assign _T_1088 = _GEN_2 << 2; // @[Math.scala 450:32:@28034.4]
  assign x389_rd_0_number = x288_lb_0_io_rPort_0_output_0; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 329:29:@27692.4 sm_x492_inr_Foreach_SAMPLER_BOX.scala 333:406:@27713.4]
  assign _GEN_3 = {{1'd0}, x389_rd_0_number}; // @[Math.scala 450:32:@28039.4]
  assign _T_1092 = _GEN_3 << 1; // @[Math.scala 450:32:@28039.4]
  assign x416_rd_0_number = x288_lb_0_io_rPort_1_output_0; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 386:29:@27898.4 sm_x492_inr_Foreach_SAMPLER_BOX.scala 390:406:@27919.4]
  assign _GEN_4 = {{1'd0}, x416_rd_0_number}; // @[Math.scala 450:32:@28044.4]
  assign _T_1096 = _GEN_4 << 1; // @[Math.scala 450:32:@28044.4]
  assign x444_sum_number = x444_sum_1_io_result; // @[Math.scala 154:22:@28133.4 Math.scala 155:14:@28134.4]
  assign _T_1132 = x444_sum_number[7:4]; // @[FixedPoint.scala 18:52:@28139.4]
  assign x350_rd_0_number = x288_lb_0_io_rPort_7_output_0; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 235:29:@27369.4 sm_x492_inr_Foreach_SAMPLER_BOX.scala 239:371:@27390.4]
  assign _GEN_5 = {{1'd0}, x350_rd_0_number}; // @[Math.scala 450:32:@28152.4]
  assign _T_1139 = _GEN_5 << 1; // @[Math.scala 450:32:@28152.4]
  assign _GEN_6 = {{1'd0}, x382_rd_0_number}; // @[Math.scala 450:32:@28157.4]
  assign _T_1143 = _GEN_6 << 1; // @[Math.scala 450:32:@28157.4]
  assign _GEN_7 = {{2'd0}, x389_rd_0_number}; // @[Math.scala 450:32:@28162.4]
  assign _T_1147 = _GEN_7 << 2; // @[Math.scala 450:32:@28162.4]
  assign x396_rd_0_number = x288_lb_0_io_rPort_2_output_0; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 344:29:@27741.4 sm_x492_inr_Foreach_SAMPLER_BOX.scala 348:406:@27762.4]
  assign _GEN_8 = {{1'd0}, x396_rd_0_number}; // @[Math.scala 450:32:@28167.4]
  assign _T_1151 = _GEN_8 << 1; // @[Math.scala 450:32:@28167.4]
  assign x423_rd_0_number = x288_lb_0_io_rPort_5_output_0; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 401:29:@27947.4 sm_x492_inr_Foreach_SAMPLER_BOX.scala 405:406:@27968.4]
  assign _GEN_9 = {{1'd0}, x423_rd_0_number}; // @[Math.scala 450:32:@28172.4]
  assign _T_1155 = _GEN_9 << 1; // @[Math.scala 450:32:@28172.4]
  assign x458_sum_number = x458_sum_1_io_result; // @[Math.scala 154:22:@28261.4 Math.scala 155:14:@28262.4]
  assign _T_1191 = x458_sum_number[7:4]; // @[FixedPoint.scala 18:52:@28267.4]
  assign _T_1215 = RetimeWrapper_64_io_out; // @[package.scala 96:25:@28331.4 package.scala 96:25:@28332.4]
  assign _T_1217 = io_rr ? _T_1215 : 1'h0; // @[implicits.scala 55:10:@28333.4]
  assign _T_1218 = _T_367 & _T_1217; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 506:167:@28334.4]
  assign _T_1220 = _T_1218 & _T_367; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 506:255:@28336.4]
  assign _T_1221 = _T_1220 & io_sigsIn_backpressure; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 506:274:@28337.4]
  assign x615_b286_D10 = RetimeWrapper_60_io_out; // @[package.scala 96:25:@28293.4 package.scala 96:25:@28294.4]
  assign _T_1222 = _T_1221 & x615_b286_D10; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 506:300:@28338.4]
  assign x617_b287_D10 = RetimeWrapper_62_io_out; // @[package.scala 96:25:@28311.4 package.scala 96:25:@28312.4]
  assign _T_1235 = RetimeWrapper_67_io_out; // @[package.scala 96:25:@28372.4 package.scala 96:25:@28373.4]
  assign _T_1237 = io_rr ? _T_1235 : 1'h0; // @[implicits.scala 55:10:@28374.4]
  assign _T_1238 = _T_367 & _T_1237; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 515:167:@28375.4]
  assign _T_1240 = _T_1238 & _T_367; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 515:255:@28377.4]
  assign _T_1241 = _T_1240 & io_sigsIn_backpressure; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 515:274:@28378.4]
  assign _T_1242 = _T_1241 & x615_b286_D10; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 515:300:@28379.4]
  assign _T_1264 = RetimeWrapper_71_io_out; // @[package.scala 96:25:@28423.4 package.scala 96:25:@28424.4]
  assign _T_1266 = io_rr ? _T_1264 : 1'h0; // @[implicits.scala 55:10:@28425.4]
  assign _T_1267 = _T_367 & _T_1266; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 527:195:@28426.4]
  assign x621_x323_D5 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@28393.4 package.scala 96:25:@28394.4]
  assign _T_1268 = _T_1267 & x621_x323_D5; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 527:283:@28427.4]
  assign _T_1269 = _T_1268 & x615_b286_D10; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 527:291:@28428.4]
  assign _T_1289 = RetimeWrapper_74_io_out; // @[package.scala 96:25:@28465.4 package.scala 96:25:@28466.4]
  assign _T_1291 = io_rr ? _T_1289 : 1'h0; // @[implicits.scala 55:10:@28467.4]
  assign _T_1292 = _T_367 & _T_1291; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 544:195:@28468.4]
  assign x624_x334_D6 = RetimeWrapper_72_io_out; // @[package.scala 96:25:@28444.4 package.scala 96:25:@28445.4]
  assign _T_1293 = _T_1292 & x624_x334_D6; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 544:283:@28469.4]
  assign _T_1294 = _T_1293 & x615_b286_D10; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 544:326:@28470.4]
  assign _T_1317 = RetimeWrapper_78_io_out; // @[package.scala 96:25:@28516.4 package.scala 96:25:@28517.4]
  assign _T_1319 = io_rr ? _T_1317 : 1'h0; // @[implicits.scala 55:10:@28518.4]
  assign _T_1320 = _T_367 & _T_1319; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 557:195:@28519.4]
  assign x627_x343_D5 = RetimeWrapper_76_io_out; // @[package.scala 96:25:@28495.4 package.scala 96:25:@28496.4]
  assign _T_1321 = _T_1320 & x627_x343_D5; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 557:283:@28520.4]
  assign _T_1322 = _T_1321 & x615_b286_D10; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 557:291:@28521.4]
  assign _T_1345 = RetimeWrapper_82_io_out; // @[package.scala 96:25:@28567.4 package.scala 96:25:@28568.4]
  assign _T_1347 = io_rr ? _T_1345 : 1'h0; // @[implicits.scala 55:10:@28569.4]
  assign _T_1348 = _T_367 & _T_1347; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 570:195:@28570.4]
  assign x630_x368_D5 = RetimeWrapper_80_io_out; // @[package.scala 96:25:@28546.4 package.scala 96:25:@28547.4]
  assign _T_1349 = _T_1348 & x630_x368_D5; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 570:283:@28571.4]
  assign _T_1350 = _T_1349 & x615_b286_D10; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 570:291:@28572.4]
  assign _T_1370 = RetimeWrapper_85_io_out; // @[package.scala 96:25:@28609.4 package.scala 96:25:@28610.4]
  assign _T_1372 = io_rr ? _T_1370 : 1'h0; // @[implicits.scala 55:10:@28611.4]
  assign _T_1373 = _T_367 & _T_1372; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 581:195:@28612.4]
  assign x633_x378_D5 = RetimeWrapper_84_io_out; // @[package.scala 96:25:@28597.4 package.scala 96:25:@28598.4]
  assign _T_1374 = _T_1373 & x633_x378_D5; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 581:283:@28613.4]
  assign _T_1375 = _T_1374 & x615_b286_D10; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 581:291:@28614.4]
  assign _T_1395 = RetimeWrapper_88_io_out; // @[package.scala 96:25:@28651.4 package.scala 96:25:@28652.4]
  assign _T_1397 = io_rr ? _T_1395 : 1'h0; // @[implicits.scala 55:10:@28653.4]
  assign _T_1398 = _T_367 & _T_1397; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 592:195:@28654.4]
  assign x634_x385_D5 = RetimeWrapper_86_io_out; // @[package.scala 96:25:@28630.4 package.scala 96:25:@28631.4]
  assign _T_1399 = _T_1398 & x634_x385_D5; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 592:283:@28655.4]
  assign _T_1400 = _T_1399 & x615_b286_D10; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 592:291:@28656.4]
  assign x466_rd_0_number = x289_lb2_0_io_rPort_2_output_0; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 540:29:@28456.4 sm_x492_inr_Foreach_SAMPLER_BOX.scala 544:443:@28477.4]
  assign _GEN_10 = {{1'd0}, x466_rd_0_number}; // @[Math.scala 450:32:@28670.4]
  assign _T_1408 = _GEN_10 << 1; // @[Math.scala 450:32:@28670.4]
  assign x470_rd_0_number = x289_lb2_0_io_rPort_3_output_0; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 566:29:@28558.4 sm_x492_inr_Foreach_SAMPLER_BOX.scala 570:408:@28579.4]
  assign _GEN_11 = {{1'd0}, x470_rd_0_number}; // @[Math.scala 450:32:@28675.4]
  assign _T_1412 = _GEN_11 << 1; // @[Math.scala 450:32:@28675.4]
  assign x468_rd_0_number = x289_lb2_0_io_rPort_0_output_0; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 553:29:@28507.4 sm_x492_inr_Foreach_SAMPLER_BOX.scala 557:408:@28528.4]
  assign _GEN_12 = {{1'd0}, x468_rd_0_number}; // @[Math.scala 450:32:@28722.4]
  assign _T_1432 = _GEN_12 << 1; // @[Math.scala 450:32:@28722.4]
  assign x472_rd_0_number = x289_lb2_0_io_rPort_1_output_0; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 577:29:@28600.4 sm_x492_inr_Foreach_SAMPLER_BOX.scala 581:408:@28621.4]
  assign _GEN_13 = {{1'd0}, x472_rd_0_number}; // @[Math.scala 450:32:@28727.4]
  assign _T_1436 = _GEN_13 << 1; // @[Math.scala 450:32:@28727.4]
  assign x481_div_number = x481_div_1_io_result; // @[Math.scala 331:22:@28717.4 Math.scala 332:14:@28718.4]
  assign x487_div_number = x487_div_1_io_result; // @[Math.scala 331:22:@28769.4 Math.scala 332:14:@28770.4]
  assign _T_1474 = RetimeWrapper_92_io_out; // @[package.scala 96:25:@28811.4 package.scala 96:25:@28812.4]
  assign _T_1476 = io_rr ? _T_1474 : 1'h0; // @[implicits.scala 55:10:@28813.4]
  assign x637_b286_D20 = RetimeWrapper_91_io_out; // @[package.scala 96:25:@28802.4 package.scala 96:25:@28803.4]
  assign _T_1477 = _T_1476 & x637_b286_D20; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 630:116:@28814.4]
  assign x636_b287_D20 = RetimeWrapper_90_io_out; // @[package.scala 96:25:@28793.4 package.scala 96:25:@28794.4]
  assign _T_1478 = _T_1477 & x636_b287_D20; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 630:122:@28815.4]
  assign x572_x561_D2_number = RetimeWrapper_1_io_out; // @[package.scala 96:25:@26862.4 package.scala 96:25:@26863.4]
  assign x575_x303_sum_D1_number = RetimeWrapper_4_io_out; // @[package.scala 96:25:@26889.4 package.scala 96:25:@26890.4]
  assign x577_x560_D2_number = RetimeWrapper_6_io_out; // @[package.scala 96:25:@26907.4 package.scala 96:25:@26908.4]
  assign x313_sum_number = x313_sum_1_io_result; // @[Math.scala 154:22:@26983.4 Math.scala 155:14:@26984.4]
  assign x579_x562_D1_number = RetimeWrapper_9_io_out; // @[package.scala 96:25:@26992.4 package.scala 96:25:@26993.4]
  assign x326_sum_number = x326_sum_1_io_result; // @[Math.scala 154:22:@27130.4 Math.scala 155:14:@27131.4]
  assign x586_x562_D5_number = RetimeWrapper_17_io_out; // @[package.scala 96:25:@27139.4 package.scala 96:25:@27140.4]
  assign x590_x564_D2_number = RetimeWrapper_21_io_out; // @[package.scala 96:25:@27175.4 package.scala 96:25:@27176.4]
  assign x594_x561_D6_number = RetimeWrapper_26_io_out; // @[package.scala 96:25:@27260.4 package.scala 96:25:@27261.4]
  assign x595_x335_sum_D1_number = RetimeWrapper_27_io_out; // @[package.scala 96:25:@27269.4 package.scala 96:25:@27270.4]
  assign x346_sum_number = x346_sum_1_io_result; // @[Math.scala 154:22:@27348.4 Math.scala 155:14:@27349.4]
  assign x596_x565_D1_number = RetimeWrapper_29_io_out; // @[package.scala 96:25:@27357.4 package.scala 96:25:@27358.4]
  assign x358_sum_number = x358_sum_1_io_result; // @[Math.scala 154:22:@27445.4 Math.scala 155:14:@27446.4]
  assign x598_x566_D1_number = RetimeWrapper_32_io_out; // @[package.scala 96:25:@27454.4 package.scala 96:25:@27455.4]
  assign x371_sum_number = x371_sum_1_io_result; // @[Math.scala 154:22:@27553.4 Math.scala 155:14:@27554.4]
  assign x601_x568_D1_number = RetimeWrapper_36_io_out; // @[package.scala 96:25:@27571.4 package.scala 96:25:@27572.4]
  assign x379_sum_number = x379_sum_1_io_result; // @[Math.scala 154:22:@27631.4 Math.scala 155:14:@27632.4]
  assign x386_sum_number = x386_sum_1_io_result; // @[Math.scala 154:22:@27680.4 Math.scala 155:14:@27681.4]
  assign x393_sum_number = x393_sum_1_io_result; // @[Math.scala 154:22:@27729.4 Math.scala 155:14:@27730.4]
  assign x405_sum_number = x405_sum_1_io_result; // @[Math.scala 154:22:@27828.4 Math.scala 155:14:@27829.4]
  assign x607_x570_D1_number = RetimeWrapper_46_io_out; // @[package.scala 96:25:@27837.4 package.scala 96:25:@27838.4]
  assign x413_sum_number = x413_sum_1_io_result; // @[Math.scala 154:22:@27886.4 Math.scala 155:14:@27887.4]
  assign x420_sum_number = x420_sum_1_io_result; // @[Math.scala 154:22:@27935.4 Math.scala 155:14:@27936.4]
  assign x427_sum_number = x427_sum_1_io_result; // @[Math.scala 154:22:@27984.4 Math.scala 155:14:@27985.4]
  assign x614_x561_D10_number = RetimeWrapper_59_io_out; // @[package.scala 96:25:@28284.4 package.scala 96:25:@28285.4]
  assign x616_x303_sum_D9_number = RetimeWrapper_61_io_out; // @[package.scala 96:25:@28302.4 package.scala 96:25:@28303.4]
  assign x618_x560_D10_number = RetimeWrapper_63_io_out; // @[package.scala 96:25:@28320.4 package.scala 96:25:@28321.4]
  assign x619_x562_D9_number = RetimeWrapper_65_io_out; // @[package.scala 96:25:@28352.4 package.scala 96:25:@28353.4]
  assign x620_x313_sum_D8_number = RetimeWrapper_66_io_out; // @[package.scala 96:25:@28361.4 package.scala 96:25:@28362.4]
  assign x622_x564_D6_number = RetimeWrapper_69_io_out; // @[package.scala 96:25:@28402.4 package.scala 96:25:@28403.4]
  assign x623_x326_sum_D4_number = RetimeWrapper_70_io_out; // @[package.scala 96:25:@28411.4 package.scala 96:25:@28412.4]
  assign x625_x335_sum_D5_number = RetimeWrapper_73_io_out; // @[package.scala 96:25:@28453.4 package.scala 96:25:@28454.4]
  assign x626_x565_D5_number = RetimeWrapper_75_io_out; // @[package.scala 96:25:@28486.4 package.scala 96:25:@28487.4]
  assign x628_x346_sum_D4_number = RetimeWrapper_77_io_out; // @[package.scala 96:25:@28504.4 package.scala 96:25:@28505.4]
  assign x629_x371_sum_D4_number = RetimeWrapper_79_io_out; // @[package.scala 96:25:@28537.4 package.scala 96:25:@28538.4]
  assign x631_x568_D5_number = RetimeWrapper_81_io_out; // @[package.scala 96:25:@28555.4 package.scala 96:25:@28556.4]
  assign x632_x379_sum_D4_number = RetimeWrapper_83_io_out; // @[package.scala 96:25:@28588.4 package.scala 96:25:@28589.4]
  assign x635_x386_sum_D4_number = RetimeWrapper_87_io_out; // @[package.scala 96:25:@28639.4 package.scala 96:25:@28640.4]
  assign io_in_x276_TVALID = _T_1478 & io_sigsIn_backpressure; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 630:22:@28817.4]
  assign io_in_x276_TDATA = {{240'd0}, RetimeWrapper_89_io_out}; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 631:24:@28818.4]
  assign io_in_x275_TREADY = _T_213 & _T_215; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 69:22:@26730.4 sm_x492_inr_Foreach_SAMPLER_BOX.scala 71:22:@26738.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 710:17:@26558.4]
  assign __1_io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_1); // @[Math.scala 710:17:@26570.4]
  assign x288_lb_0_clock = clock; // @[:@26578.4]
  assign x288_lb_0_reset = reset; // @[:@26579.4]
  assign x288_lb_0_io_rPort_11_banks_1 = x594_x561_D6_number[2:0]; // @[MemInterfaceType.scala 106:58:@27289.4]
  assign x288_lb_0_io_rPort_11_banks_0 = x590_x564_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@27288.4]
  assign x288_lb_0_io_rPort_11_ofs_0 = x595_x335_sum_D1_number[0]; // @[MemInterfaceType.scala 107:54:@27290.4]
  assign x288_lb_0_io_rPort_11_en_0 = _T_590 & x589_b287_D6; // @[MemInterfaceType.scala 110:79:@27292.4]
  assign x288_lb_0_io_rPort_11_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@27291.4]
  assign x288_lb_0_io_rPort_10_banks_1 = x586_x562_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@27866.4]
  assign x288_lb_0_io_rPort_10_banks_0 = x607_x570_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@27865.4]
  assign x288_lb_0_io_rPort_10_ofs_0 = x405_sum_number[0]; // @[MemInterfaceType.scala 107:54:@27867.4]
  assign x288_lb_0_io_rPort_10_en_0 = _T_985 & x589_b287_D6; // @[MemInterfaceType.scala 110:79:@27869.4]
  assign x288_lb_0_io_rPort_10_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@27868.4]
  assign x288_lb_0_io_rPort_9_banks_1 = x586_x562_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@27195.4]
  assign x288_lb_0_io_rPort_9_banks_0 = x590_x564_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@27194.4]
  assign x288_lb_0_io_rPort_9_ofs_0 = x326_sum_number[0]; // @[MemInterfaceType.scala 107:54:@27196.4]
  assign x288_lb_0_io_rPort_9_en_0 = _T_539 & x589_b287_D6; // @[MemInterfaceType.scala 110:79:@27198.4]
  assign x288_lb_0_io_rPort_9_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@27197.4]
  assign x288_lb_0_io_rPort_8_banks_1 = x598_x566_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@27483.4]
  assign x288_lb_0_io_rPort_8_banks_0 = x590_x564_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@27482.4]
  assign x288_lb_0_io_rPort_8_ofs_0 = x358_sum_number[0]; // @[MemInterfaceType.scala 107:54:@27484.4]
  assign x288_lb_0_io_rPort_8_en_0 = _T_728 & x589_b287_D6; // @[MemInterfaceType.scala 110:79:@27486.4]
  assign x288_lb_0_io_rPort_8_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@27485.4]
  assign x288_lb_0_io_rPort_7_banks_1 = x596_x565_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@27386.4]
  assign x288_lb_0_io_rPort_7_banks_0 = x590_x564_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@27385.4]
  assign x288_lb_0_io_rPort_7_ofs_0 = x346_sum_number[0]; // @[MemInterfaceType.scala 107:54:@27387.4]
  assign x288_lb_0_io_rPort_7_en_0 = _T_659 & x589_b287_D6; // @[MemInterfaceType.scala 110:79:@27389.4]
  assign x288_lb_0_io_rPort_7_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@27388.4]
  assign x288_lb_0_io_rPort_6_banks_1 = x594_x561_D6_number[2:0]; // @[MemInterfaceType.scala 106:58:@27660.4]
  assign x288_lb_0_io_rPort_6_banks_0 = x601_x568_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@27659.4]
  assign x288_lb_0_io_rPort_6_ofs_0 = x379_sum_number[0]; // @[MemInterfaceType.scala 107:54:@27661.4]
  assign x288_lb_0_io_rPort_6_en_0 = _T_846 & x589_b287_D6; // @[MemInterfaceType.scala 110:79:@27663.4]
  assign x288_lb_0_io_rPort_6_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@27662.4]
  assign x288_lb_0_io_rPort_5_banks_1 = x596_x565_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@27964.4]
  assign x288_lb_0_io_rPort_5_banks_0 = x607_x570_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@27963.4]
  assign x288_lb_0_io_rPort_5_ofs_0 = x420_sum_number[0]; // @[MemInterfaceType.scala 107:54:@27965.4]
  assign x288_lb_0_io_rPort_5_en_0 = _T_1043 & x589_b287_D6; // @[MemInterfaceType.scala 110:79:@27967.4]
  assign x288_lb_0_io_rPort_5_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@27966.4]
  assign x288_lb_0_io_rPort_4_banks_1 = x586_x562_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@27591.4]
  assign x288_lb_0_io_rPort_4_banks_0 = x601_x568_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@27590.4]
  assign x288_lb_0_io_rPort_4_ofs_0 = x371_sum_number[0]; // @[MemInterfaceType.scala 107:54:@27592.4]
  assign x288_lb_0_io_rPort_4_en_0 = _T_809 & x589_b287_D6; // @[MemInterfaceType.scala 110:79:@27594.4]
  assign x288_lb_0_io_rPort_4_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@27593.4]
  assign x288_lb_0_io_rPort_3_banks_1 = x598_x566_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@28013.4]
  assign x288_lb_0_io_rPort_3_banks_0 = x607_x570_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@28012.4]
  assign x288_lb_0_io_rPort_3_ofs_0 = x427_sum_number[0]; // @[MemInterfaceType.scala 107:54:@28014.4]
  assign x288_lb_0_io_rPort_3_en_0 = _T_1072 & x589_b287_D6; // @[MemInterfaceType.scala 110:79:@28016.4]
  assign x288_lb_0_io_rPort_3_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@28015.4]
  assign x288_lb_0_io_rPort_2_banks_1 = x598_x566_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@27758.4]
  assign x288_lb_0_io_rPort_2_banks_0 = x601_x568_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@27757.4]
  assign x288_lb_0_io_rPort_2_ofs_0 = x393_sum_number[0]; // @[MemInterfaceType.scala 107:54:@27759.4]
  assign x288_lb_0_io_rPort_2_en_0 = _T_904 & x589_b287_D6; // @[MemInterfaceType.scala 110:79:@27761.4]
  assign x288_lb_0_io_rPort_2_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@27760.4]
  assign x288_lb_0_io_rPort_1_banks_1 = x594_x561_D6_number[2:0]; // @[MemInterfaceType.scala 106:58:@27915.4]
  assign x288_lb_0_io_rPort_1_banks_0 = x607_x570_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@27914.4]
  assign x288_lb_0_io_rPort_1_ofs_0 = x413_sum_number[0]; // @[MemInterfaceType.scala 107:54:@27916.4]
  assign x288_lb_0_io_rPort_1_en_0 = _T_1014 & x589_b287_D6; // @[MemInterfaceType.scala 110:79:@27918.4]
  assign x288_lb_0_io_rPort_1_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@27917.4]
  assign x288_lb_0_io_rPort_0_banks_1 = x596_x565_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@27709.4]
  assign x288_lb_0_io_rPort_0_banks_0 = x601_x568_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@27708.4]
  assign x288_lb_0_io_rPort_0_ofs_0 = x386_sum_number[0]; // @[MemInterfaceType.scala 107:54:@27710.4]
  assign x288_lb_0_io_rPort_0_en_0 = _T_875 & x589_b287_D6; // @[MemInterfaceType.scala 110:79:@27712.4]
  assign x288_lb_0_io_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@27711.4]
  assign x288_lb_0_io_wPort_1_banks_1 = x579_x562_D1_number[2:0]; // @[MemInterfaceType.scala 88:58:@27022.4]
  assign x288_lb_0_io_wPort_1_banks_0 = x577_x560_D2_number[2:0]; // @[MemInterfaceType.scala 88:58:@27021.4]
  assign x288_lb_0_io_wPort_1_ofs_0 = x313_sum_number[0]; // @[MemInterfaceType.scala 89:54:@27023.4]
  assign x288_lb_0_io_wPort_1_data_0 = RetimeWrapper_10_io_out; // @[MemInterfaceType.scala 90:56:@27024.4]
  assign x288_lb_0_io_wPort_1_en_0 = _T_434 & x576_b287_D2; // @[MemInterfaceType.scala 93:57:@27026.4]
  assign x288_lb_0_io_wPort_0_banks_1 = x572_x561_D2_number[2:0]; // @[MemInterfaceType.scala 88:58:@26928.4]
  assign x288_lb_0_io_wPort_0_banks_0 = x577_x560_D2_number[2:0]; // @[MemInterfaceType.scala 88:58:@26927.4]
  assign x288_lb_0_io_wPort_0_ofs_0 = x575_x303_sum_D1_number[0]; // @[MemInterfaceType.scala 89:54:@26929.4]
  assign x288_lb_0_io_wPort_0_data_0 = RetimeWrapper_2_io_out; // @[MemInterfaceType.scala 90:56:@26930.4]
  assign x288_lb_0_io_wPort_0_en_0 = _T_378 & x576_b287_D2; // @[MemInterfaceType.scala 93:57:@26932.4]
  assign x289_lb2_0_clock = clock; // @[:@26671.4]
  assign x289_lb2_0_reset = reset; // @[:@26672.4]
  assign x289_lb2_0_io_rPort_5_banks_1 = x619_x562_D9_number[2:0]; // @[MemInterfaceType.scala 106:58:@28431.4]
  assign x289_lb2_0_io_rPort_5_banks_0 = x622_x564_D6_number[2:0]; // @[MemInterfaceType.scala 106:58:@28430.4]
  assign x289_lb2_0_io_rPort_5_ofs_0 = x623_x326_sum_D4_number[0]; // @[MemInterfaceType.scala 107:54:@28432.4]
  assign x289_lb2_0_io_rPort_5_en_0 = _T_1269 & x617_b287_D10; // @[MemInterfaceType.scala 110:79:@28434.4]
  assign x289_lb2_0_io_rPort_5_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@28433.4]
  assign x289_lb2_0_io_rPort_4_banks_1 = x626_x565_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@28659.4]
  assign x289_lb2_0_io_rPort_4_banks_0 = x631_x568_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@28658.4]
  assign x289_lb2_0_io_rPort_4_ofs_0 = x635_x386_sum_D4_number[0]; // @[MemInterfaceType.scala 107:54:@28660.4]
  assign x289_lb2_0_io_rPort_4_en_0 = _T_1400 & x617_b287_D10; // @[MemInterfaceType.scala 110:79:@28662.4]
  assign x289_lb2_0_io_rPort_4_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@28661.4]
  assign x289_lb2_0_io_rPort_3_banks_1 = x619_x562_D9_number[2:0]; // @[MemInterfaceType.scala 106:58:@28575.4]
  assign x289_lb2_0_io_rPort_3_banks_0 = x631_x568_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@28574.4]
  assign x289_lb2_0_io_rPort_3_ofs_0 = x629_x371_sum_D4_number[0]; // @[MemInterfaceType.scala 107:54:@28576.4]
  assign x289_lb2_0_io_rPort_3_en_0 = _T_1350 & x617_b287_D10; // @[MemInterfaceType.scala 110:79:@28578.4]
  assign x289_lb2_0_io_rPort_3_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@28577.4]
  assign x289_lb2_0_io_rPort_2_banks_1 = x614_x561_D10_number[2:0]; // @[MemInterfaceType.scala 106:58:@28473.4]
  assign x289_lb2_0_io_rPort_2_banks_0 = x622_x564_D6_number[2:0]; // @[MemInterfaceType.scala 106:58:@28472.4]
  assign x289_lb2_0_io_rPort_2_ofs_0 = x625_x335_sum_D5_number[0]; // @[MemInterfaceType.scala 107:54:@28474.4]
  assign x289_lb2_0_io_rPort_2_en_0 = _T_1294 & x617_b287_D10; // @[MemInterfaceType.scala 110:79:@28476.4]
  assign x289_lb2_0_io_rPort_2_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@28475.4]
  assign x289_lb2_0_io_rPort_1_banks_1 = x614_x561_D10_number[2:0]; // @[MemInterfaceType.scala 106:58:@28617.4]
  assign x289_lb2_0_io_rPort_1_banks_0 = x631_x568_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@28616.4]
  assign x289_lb2_0_io_rPort_1_ofs_0 = x632_x379_sum_D4_number[0]; // @[MemInterfaceType.scala 107:54:@28618.4]
  assign x289_lb2_0_io_rPort_1_en_0 = _T_1375 & x617_b287_D10; // @[MemInterfaceType.scala 110:79:@28620.4]
  assign x289_lb2_0_io_rPort_1_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@28619.4]
  assign x289_lb2_0_io_rPort_0_banks_1 = x626_x565_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@28524.4]
  assign x289_lb2_0_io_rPort_0_banks_0 = x622_x564_D6_number[2:0]; // @[MemInterfaceType.scala 106:58:@28523.4]
  assign x289_lb2_0_io_rPort_0_ofs_0 = x628_x346_sum_D4_number[0]; // @[MemInterfaceType.scala 107:54:@28525.4]
  assign x289_lb2_0_io_rPort_0_en_0 = _T_1322 & x617_b287_D10; // @[MemInterfaceType.scala 110:79:@28527.4]
  assign x289_lb2_0_io_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@28526.4]
  assign x289_lb2_0_io_wPort_1_banks_1 = x619_x562_D9_number[2:0]; // @[MemInterfaceType.scala 88:58:@28382.4]
  assign x289_lb2_0_io_wPort_1_banks_0 = x618_x560_D10_number[2:0]; // @[MemInterfaceType.scala 88:58:@28381.4]
  assign x289_lb2_0_io_wPort_1_ofs_0 = x620_x313_sum_D8_number[0]; // @[MemInterfaceType.scala 89:54:@28383.4]
  assign x289_lb2_0_io_wPort_1_data_0 = RetimeWrapper_56_io_out; // @[MemInterfaceType.scala 90:56:@28384.4]
  assign x289_lb2_0_io_wPort_1_en_0 = _T_1242 & x617_b287_D10; // @[MemInterfaceType.scala 93:57:@28386.4]
  assign x289_lb2_0_io_wPort_0_banks_1 = x614_x561_D10_number[2:0]; // @[MemInterfaceType.scala 88:58:@28341.4]
  assign x289_lb2_0_io_wPort_0_banks_0 = x618_x560_D10_number[2:0]; // @[MemInterfaceType.scala 88:58:@28340.4]
  assign x289_lb2_0_io_wPort_0_ofs_0 = x616_x303_sum_D9_number[0]; // @[MemInterfaceType.scala 89:54:@28342.4]
  assign x289_lb2_0_io_wPort_0_data_0 = RetimeWrapper_58_io_out; // @[MemInterfaceType.scala 90:56:@28343.4]
  assign x289_lb2_0_io_wPort_0_en_0 = _T_1222 & x617_b287_D10; // @[MemInterfaceType.scala 93:57:@28345.4]
  assign RetimeWrapper_clock = clock; // @[:@26741.4]
  assign RetimeWrapper_reset = reset; // @[:@26742.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26744.4]
  assign RetimeWrapper_io_in = io_in_x275_TDATA[15:0]; // @[package.scala 94:16:@26743.4]
  assign x303_sum_1_clock = clock; // @[:@26848.4]
  assign x303_sum_1_reset = reset; // @[:@26849.4]
  assign x303_sum_1_io_a = {_T_332,_T_333}; // @[Math.scala 151:17:@26850.4]
  assign x303_sum_1_io_b = {_T_342,_T_343}; // @[Math.scala 152:17:@26851.4]
  assign x303_sum_1_io_flow = io_in_x276_TREADY; // @[Math.scala 153:20:@26852.4]
  assign RetimeWrapper_1_clock = clock; // @[:@26858.4]
  assign RetimeWrapper_1_reset = reset; // @[:@26859.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26861.4]
  assign RetimeWrapper_1_io_in = $unsigned(_T_323); // @[package.scala 94:16:@26860.4]
  assign RetimeWrapper_2_clock = clock; // @[:@26867.4]
  assign RetimeWrapper_2_reset = reset; // @[:@26868.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26870.4]
  assign RetimeWrapper_2_io_in = x571_x290_D1_0_number[7:0]; // @[package.scala 94:16:@26869.4]
  assign RetimeWrapper_3_clock = clock; // @[:@26876.4]
  assign RetimeWrapper_3_reset = reset; // @[:@26877.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26879.4]
  assign RetimeWrapper_3_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@26878.4]
  assign RetimeWrapper_4_clock = clock; // @[:@26885.4]
  assign RetimeWrapper_4_reset = reset; // @[:@26886.4]
  assign RetimeWrapper_4_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26888.4]
  assign RetimeWrapper_4_io_in = x303_sum_1_io_result; // @[package.scala 94:16:@26887.4]
  assign RetimeWrapper_5_clock = clock; // @[:@26894.4]
  assign RetimeWrapper_5_reset = reset; // @[:@26895.4]
  assign RetimeWrapper_5_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26897.4]
  assign RetimeWrapper_5_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@26896.4]
  assign RetimeWrapper_6_clock = clock; // @[:@26903.4]
  assign RetimeWrapper_6_reset = reset; // @[:@26904.4]
  assign RetimeWrapper_6_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26906.4]
  assign RetimeWrapper_6_io_in = $unsigned(_T_311); // @[package.scala 94:16:@26905.4]
  assign RetimeWrapper_7_clock = clock; // @[:@26914.4]
  assign RetimeWrapper_7_reset = reset; // @[:@26915.4]
  assign RetimeWrapper_7_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26917.4]
  assign RetimeWrapper_7_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@26916.4]
  assign x309_rdcol_1_clock = clock; // @[:@26937.4]
  assign x309_rdcol_1_reset = reset; // @[:@26938.4]
  assign x309_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@26939.4]
  assign x309_rdcol_1_io_b = 32'h1; // @[Math.scala 152:17:@26940.4]
  assign x309_rdcol_1_io_flow = io_in_x276_TREADY; // @[Math.scala 153:20:@26941.4]
  assign RetimeWrapper_8_clock = clock; // @[:@26969.4]
  assign RetimeWrapper_8_reset = reset; // @[:@26970.4]
  assign RetimeWrapper_8_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26972.4]
  assign RetimeWrapper_8_io_in = {_T_332,_T_333}; // @[package.scala 94:16:@26971.4]
  assign x313_sum_1_clock = clock; // @[:@26978.4]
  assign x313_sum_1_reset = reset; // @[:@26979.4]
  assign x313_sum_1_io_a = RetimeWrapper_8_io_out; // @[Math.scala 151:17:@26980.4]
  assign x313_sum_1_io_b = {_T_407,_T_408}; // @[Math.scala 152:17:@26981.4]
  assign x313_sum_1_io_flow = io_in_x276_TREADY; // @[Math.scala 153:20:@26982.4]
  assign RetimeWrapper_9_clock = clock; // @[:@26988.4]
  assign RetimeWrapper_9_reset = reset; // @[:@26989.4]
  assign RetimeWrapper_9_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26991.4]
  assign RetimeWrapper_9_io_in = $unsigned(_T_398); // @[package.scala 94:16:@26990.4]
  assign RetimeWrapper_10_clock = clock; // @[:@26997.4]
  assign RetimeWrapper_10_reset = reset; // @[:@26998.4]
  assign RetimeWrapper_10_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27000.4]
  assign RetimeWrapper_10_io_in = x571_x290_D1_0_number[15:8]; // @[package.scala 94:16:@26999.4]
  assign RetimeWrapper_11_clock = clock; // @[:@27008.4]
  assign RetimeWrapper_11_reset = reset; // @[:@27009.4]
  assign RetimeWrapper_11_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27011.4]
  assign RetimeWrapper_11_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@27010.4]
  assign RetimeWrapper_12_clock = clock; // @[:@27029.4]
  assign RetimeWrapper_12_reset = reset; // @[:@27030.4]
  assign RetimeWrapper_12_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27032.4]
  assign RetimeWrapper_12_io_in = __io_result; // @[package.scala 94:16:@27031.4]
  assign RetimeWrapper_13_clock = clock; // @[:@27056.4]
  assign RetimeWrapper_13_reset = reset; // @[:@27057.4]
  assign RetimeWrapper_13_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27059.4]
  assign RetimeWrapper_13_io_in = x309_rdcol_1_io_result; // @[package.scala 94:16:@27058.4]
  assign RetimeWrapper_14_clock = clock; // @[:@27072.4]
  assign RetimeWrapper_14_reset = reset; // @[:@27073.4]
  assign RetimeWrapper_14_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27075.4]
  assign RetimeWrapper_14_io_in = $signed(_T_446) < $signed(32'sh0); // @[package.scala 94:16:@27074.4]
  assign RetimeWrapper_15_clock = clock; // @[:@27107.4]
  assign RetimeWrapper_15_reset = reset; // @[:@27108.4]
  assign RetimeWrapper_15_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27110.4]
  assign RetimeWrapper_15_io_in = {_T_407,_T_408}; // @[package.scala 94:16:@27109.4]
  assign RetimeWrapper_16_clock = clock; // @[:@27116.4]
  assign RetimeWrapper_16_reset = reset; // @[:@27117.4]
  assign RetimeWrapper_16_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27119.4]
  assign RetimeWrapper_16_io_in = {_T_496,_T_497}; // @[package.scala 94:16:@27118.4]
  assign x326_sum_1_clock = clock; // @[:@27125.4]
  assign x326_sum_1_reset = reset; // @[:@27126.4]
  assign x326_sum_1_io_a = RetimeWrapper_16_io_out; // @[Math.scala 151:17:@27127.4]
  assign x326_sum_1_io_b = RetimeWrapper_15_io_out; // @[Math.scala 152:17:@27128.4]
  assign x326_sum_1_io_flow = io_in_x276_TREADY; // @[Math.scala 153:20:@27129.4]
  assign RetimeWrapper_17_clock = clock; // @[:@27135.4]
  assign RetimeWrapper_17_reset = reset; // @[:@27136.4]
  assign RetimeWrapper_17_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27138.4]
  assign RetimeWrapper_17_io_in = $unsigned(_T_398); // @[package.scala 94:16:@27137.4]
  assign RetimeWrapper_18_clock = clock; // @[:@27144.4]
  assign RetimeWrapper_18_reset = reset; // @[:@27145.4]
  assign RetimeWrapper_18_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27147.4]
  assign RetimeWrapper_18_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@27146.4]
  assign RetimeWrapper_19_clock = clock; // @[:@27153.4]
  assign RetimeWrapper_19_reset = reset; // @[:@27154.4]
  assign RetimeWrapper_19_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27156.4]
  assign RetimeWrapper_19_io_in = ~ x322; // @[package.scala 94:16:@27155.4]
  assign RetimeWrapper_20_clock = clock; // @[:@27162.4]
  assign RetimeWrapper_20_reset = reset; // @[:@27163.4]
  assign RetimeWrapper_20_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27165.4]
  assign RetimeWrapper_20_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@27164.4]
  assign RetimeWrapper_21_clock = clock; // @[:@27171.4]
  assign RetimeWrapper_21_reset = reset; // @[:@27172.4]
  assign RetimeWrapper_21_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27174.4]
  assign RetimeWrapper_21_io_in = $unsigned(_T_487); // @[package.scala 94:16:@27173.4]
  assign RetimeWrapper_22_clock = clock; // @[:@27183.4]
  assign RetimeWrapper_22_reset = reset; // @[:@27184.4]
  assign RetimeWrapper_22_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27186.4]
  assign RetimeWrapper_22_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@27185.4]
  assign RetimeWrapper_23_clock = clock; // @[:@27204.4]
  assign RetimeWrapper_23_reset = reset; // @[:@27205.4]
  assign RetimeWrapper_23_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27207.4]
  assign RetimeWrapper_23_io_in = __1_io_result; // @[package.scala 94:16:@27206.4]
  assign RetimeWrapper_24_clock = clock; // @[:@27228.4]
  assign RetimeWrapper_24_reset = reset; // @[:@27229.4]
  assign RetimeWrapper_24_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27231.4]
  assign RetimeWrapper_24_io_in = {_T_342,_T_343}; // @[package.scala 94:16:@27230.4]
  assign x335_sum_1_clock = clock; // @[:@27237.4]
  assign x335_sum_1_reset = reset; // @[:@27238.4]
  assign x335_sum_1_io_a = {_T_496,_T_497}; // @[Math.scala 151:17:@27239.4]
  assign x335_sum_1_io_b = RetimeWrapper_24_io_out; // @[Math.scala 152:17:@27240.4]
  assign x335_sum_1_io_flow = io_in_x276_TREADY; // @[Math.scala 153:20:@27241.4]
  assign RetimeWrapper_25_clock = clock; // @[:@27247.4]
  assign RetimeWrapper_25_reset = reset; // @[:@27248.4]
  assign RetimeWrapper_25_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27250.4]
  assign RetimeWrapper_25_io_in = ~ x333; // @[package.scala 94:16:@27249.4]
  assign RetimeWrapper_26_clock = clock; // @[:@27256.4]
  assign RetimeWrapper_26_reset = reset; // @[:@27257.4]
  assign RetimeWrapper_26_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27259.4]
  assign RetimeWrapper_26_io_in = $unsigned(_T_323); // @[package.scala 94:16:@27258.4]
  assign RetimeWrapper_27_clock = clock; // @[:@27265.4]
  assign RetimeWrapper_27_reset = reset; // @[:@27266.4]
  assign RetimeWrapper_27_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27268.4]
  assign RetimeWrapper_27_io_in = x335_sum_1_io_result; // @[package.scala 94:16:@27267.4]
  assign RetimeWrapper_28_clock = clock; // @[:@27277.4]
  assign RetimeWrapper_28_reset = reset; // @[:@27278.4]
  assign RetimeWrapper_28_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27280.4]
  assign RetimeWrapper_28_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@27279.4]
  assign x340_rdcol_1_clock = clock; // @[:@27300.4]
  assign x340_rdcol_1_reset = reset; // @[:@27301.4]
  assign x340_rdcol_1_io_a = RetimeWrapper_23_io_out; // @[Math.scala 151:17:@27302.4]
  assign x340_rdcol_1_io_b = 32'hffffffff; // @[Math.scala 152:17:@27303.4]
  assign x340_rdcol_1_io_flow = io_in_x276_TREADY; // @[Math.scala 153:20:@27304.4]
  assign x346_sum_1_clock = clock; // @[:@27343.4]
  assign x346_sum_1_reset = reset; // @[:@27344.4]
  assign x346_sum_1_io_a = RetimeWrapper_16_io_out; // @[Math.scala 151:17:@27345.4]
  assign x346_sum_1_io_b = {_T_631,_T_632}; // @[Math.scala 152:17:@27346.4]
  assign x346_sum_1_io_flow = io_in_x276_TREADY; // @[Math.scala 153:20:@27347.4]
  assign RetimeWrapper_29_clock = clock; // @[:@27353.4]
  assign RetimeWrapper_29_reset = reset; // @[:@27354.4]
  assign RetimeWrapper_29_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27356.4]
  assign RetimeWrapper_29_io_in = $unsigned(_T_622); // @[package.scala 94:16:@27355.4]
  assign RetimeWrapper_30_clock = clock; // @[:@27362.4]
  assign RetimeWrapper_30_reset = reset; // @[:@27363.4]
  assign RetimeWrapper_30_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27365.4]
  assign RetimeWrapper_30_io_in = ~ x342; // @[package.scala 94:16:@27364.4]
  assign RetimeWrapper_31_clock = clock; // @[:@27374.4]
  assign RetimeWrapper_31_reset = reset; // @[:@27375.4]
  assign RetimeWrapper_31_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27377.4]
  assign RetimeWrapper_31_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@27376.4]
  assign x352_rdcol_1_clock = clock; // @[:@27397.4]
  assign x352_rdcol_1_reset = reset; // @[:@27398.4]
  assign x352_rdcol_1_io_a = RetimeWrapper_23_io_out; // @[Math.scala 151:17:@27399.4]
  assign x352_rdcol_1_io_b = 32'hfffffffe; // @[Math.scala 152:17:@27400.4]
  assign x352_rdcol_1_io_flow = io_in_x276_TREADY; // @[Math.scala 153:20:@27401.4]
  assign x358_sum_1_clock = clock; // @[:@27440.4]
  assign x358_sum_1_reset = reset; // @[:@27441.4]
  assign x358_sum_1_io_a = RetimeWrapper_16_io_out; // @[Math.scala 151:17:@27442.4]
  assign x358_sum_1_io_b = {_T_700,_T_701}; // @[Math.scala 152:17:@27443.4]
  assign x358_sum_1_io_flow = io_in_x276_TREADY; // @[Math.scala 153:20:@27444.4]
  assign RetimeWrapper_32_clock = clock; // @[:@27450.4]
  assign RetimeWrapper_32_reset = reset; // @[:@27451.4]
  assign RetimeWrapper_32_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27453.4]
  assign RetimeWrapper_32_io_in = $unsigned(_T_691); // @[package.scala 94:16:@27452.4]
  assign RetimeWrapper_33_clock = clock; // @[:@27459.4]
  assign RetimeWrapper_33_reset = reset; // @[:@27460.4]
  assign RetimeWrapper_33_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27462.4]
  assign RetimeWrapper_33_io_in = ~ x354; // @[package.scala 94:16:@27461.4]
  assign RetimeWrapper_34_clock = clock; // @[:@27471.4]
  assign RetimeWrapper_34_reset = reset; // @[:@27472.4]
  assign RetimeWrapper_34_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27474.4]
  assign RetimeWrapper_34_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@27473.4]
  assign x364_rdrow_1_clock = clock; // @[:@27494.4]
  assign x364_rdrow_1_reset = reset; // @[:@27495.4]
  assign x364_rdrow_1_io_a = RetimeWrapper_12_io_out; // @[Math.scala 192:17:@27496.4]
  assign x364_rdrow_1_io_b = 32'h1; // @[Math.scala 193:17:@27497.4]
  assign x364_rdrow_1_io_flow = io_in_x276_TREADY; // @[Math.scala 194:20:@27498.4]
  assign x371_sum_1_clock = clock; // @[:@27548.4]
  assign x371_sum_1_reset = reset; // @[:@27549.4]
  assign x371_sum_1_io_a = {_T_781,_T_782}; // @[Math.scala 151:17:@27550.4]
  assign x371_sum_1_io_b = RetimeWrapper_15_io_out; // @[Math.scala 152:17:@27551.4]
  assign x371_sum_1_io_flow = io_in_x276_TREADY; // @[Math.scala 153:20:@27552.4]
  assign RetimeWrapper_35_clock = clock; // @[:@27558.4]
  assign RetimeWrapper_35_reset = reset; // @[:@27559.4]
  assign RetimeWrapper_35_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27561.4]
  assign RetimeWrapper_35_io_in = ~ x367; // @[package.scala 94:16:@27560.4]
  assign RetimeWrapper_36_clock = clock; // @[:@27567.4]
  assign RetimeWrapper_36_reset = reset; // @[:@27568.4]
  assign RetimeWrapper_36_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27570.4]
  assign RetimeWrapper_36_io_in = $unsigned(_T_772); // @[package.scala 94:16:@27569.4]
  assign RetimeWrapper_37_clock = clock; // @[:@27579.4]
  assign RetimeWrapper_37_reset = reset; // @[:@27580.4]
  assign RetimeWrapper_37_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27582.4]
  assign RetimeWrapper_37_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@27581.4]
  assign RetimeWrapper_38_clock = clock; // @[:@27600.4]
  assign RetimeWrapper_38_reset = reset; // @[:@27601.4]
  assign RetimeWrapper_38_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27603.4]
  assign RetimeWrapper_38_io_in = $signed(_T_552) < $signed(32'sh0); // @[package.scala 94:16:@27602.4]
  assign RetimeWrapper_39_clock = clock; // @[:@27615.4]
  assign RetimeWrapper_39_reset = reset; // @[:@27616.4]
  assign RetimeWrapper_39_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27618.4]
  assign RetimeWrapper_39_io_in = {_T_342,_T_343}; // @[package.scala 94:16:@27617.4]
  assign x379_sum_1_clock = clock; // @[:@27626.4]
  assign x379_sum_1_reset = reset; // @[:@27627.4]
  assign x379_sum_1_io_a = {_T_781,_T_782}; // @[Math.scala 151:17:@27628.4]
  assign x379_sum_1_io_b = RetimeWrapper_39_io_out; // @[Math.scala 152:17:@27629.4]
  assign x379_sum_1_io_flow = io_in_x276_TREADY; // @[Math.scala 153:20:@27630.4]
  assign RetimeWrapper_40_clock = clock; // @[:@27636.4]
  assign RetimeWrapper_40_reset = reset; // @[:@27637.4]
  assign RetimeWrapper_40_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27639.4]
  assign RetimeWrapper_40_io_in = ~ x377; // @[package.scala 94:16:@27638.4]
  assign RetimeWrapper_41_clock = clock; // @[:@27648.4]
  assign RetimeWrapper_41_reset = reset; // @[:@27649.4]
  assign RetimeWrapper_41_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27651.4]
  assign RetimeWrapper_41_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@27650.4]
  assign x386_sum_1_clock = clock; // @[:@27675.4]
  assign x386_sum_1_reset = reset; // @[:@27676.4]
  assign x386_sum_1_io_a = {_T_781,_T_782}; // @[Math.scala 151:17:@27677.4]
  assign x386_sum_1_io_b = {_T_631,_T_632}; // @[Math.scala 152:17:@27678.4]
  assign x386_sum_1_io_flow = io_in_x276_TREADY; // @[Math.scala 153:20:@27679.4]
  assign RetimeWrapper_42_clock = clock; // @[:@27685.4]
  assign RetimeWrapper_42_reset = reset; // @[:@27686.4]
  assign RetimeWrapper_42_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27688.4]
  assign RetimeWrapper_42_io_in = ~ x384; // @[package.scala 94:16:@27687.4]
  assign RetimeWrapper_43_clock = clock; // @[:@27697.4]
  assign RetimeWrapper_43_reset = reset; // @[:@27698.4]
  assign RetimeWrapper_43_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27700.4]
  assign RetimeWrapper_43_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@27699.4]
  assign x393_sum_1_clock = clock; // @[:@27724.4]
  assign x393_sum_1_reset = reset; // @[:@27725.4]
  assign x393_sum_1_io_a = {_T_781,_T_782}; // @[Math.scala 151:17:@27726.4]
  assign x393_sum_1_io_b = {_T_700,_T_701}; // @[Math.scala 152:17:@27727.4]
  assign x393_sum_1_io_flow = io_in_x276_TREADY; // @[Math.scala 153:20:@27728.4]
  assign RetimeWrapper_44_clock = clock; // @[:@27734.4]
  assign RetimeWrapper_44_reset = reset; // @[:@27735.4]
  assign RetimeWrapper_44_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27737.4]
  assign RetimeWrapper_44_io_in = ~ x391; // @[package.scala 94:16:@27736.4]
  assign RetimeWrapper_45_clock = clock; // @[:@27746.4]
  assign RetimeWrapper_45_reset = reset; // @[:@27747.4]
  assign RetimeWrapper_45_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27749.4]
  assign RetimeWrapper_45_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@27748.4]
  assign x398_rdrow_1_clock = clock; // @[:@27769.4]
  assign x398_rdrow_1_reset = reset; // @[:@27770.4]
  assign x398_rdrow_1_io_a = RetimeWrapper_12_io_out; // @[Math.scala 192:17:@27771.4]
  assign x398_rdrow_1_io_b = 32'h2; // @[Math.scala 193:17:@27772.4]
  assign x398_rdrow_1_io_flow = io_in_x276_TREADY; // @[Math.scala 194:20:@27773.4]
  assign x405_sum_1_clock = clock; // @[:@27823.4]
  assign x405_sum_1_reset = reset; // @[:@27824.4]
  assign x405_sum_1_io_a = {_T_957,_T_958}; // @[Math.scala 151:17:@27825.4]
  assign x405_sum_1_io_b = RetimeWrapper_15_io_out; // @[Math.scala 152:17:@27826.4]
  assign x405_sum_1_io_flow = io_in_x276_TREADY; // @[Math.scala 153:20:@27827.4]
  assign RetimeWrapper_46_clock = clock; // @[:@27833.4]
  assign RetimeWrapper_46_reset = reset; // @[:@27834.4]
  assign RetimeWrapper_46_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27836.4]
  assign RetimeWrapper_46_io_in = $unsigned(_T_948); // @[package.scala 94:16:@27835.4]
  assign RetimeWrapper_47_clock = clock; // @[:@27842.4]
  assign RetimeWrapper_47_reset = reset; // @[:@27843.4]
  assign RetimeWrapper_47_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27845.4]
  assign RetimeWrapper_47_io_in = ~ x401; // @[package.scala 94:16:@27844.4]
  assign RetimeWrapper_48_clock = clock; // @[:@27854.4]
  assign RetimeWrapper_48_reset = reset; // @[:@27855.4]
  assign RetimeWrapper_48_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27857.4]
  assign RetimeWrapper_48_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@27856.4]
  assign x413_sum_1_clock = clock; // @[:@27881.4]
  assign x413_sum_1_reset = reset; // @[:@27882.4]
  assign x413_sum_1_io_a = {_T_957,_T_958}; // @[Math.scala 151:17:@27883.4]
  assign x413_sum_1_io_b = RetimeWrapper_39_io_out; // @[Math.scala 152:17:@27884.4]
  assign x413_sum_1_io_flow = io_in_x276_TREADY; // @[Math.scala 153:20:@27885.4]
  assign RetimeWrapper_49_clock = clock; // @[:@27891.4]
  assign RetimeWrapper_49_reset = reset; // @[:@27892.4]
  assign RetimeWrapper_49_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27894.4]
  assign RetimeWrapper_49_io_in = ~ x411; // @[package.scala 94:16:@27893.4]
  assign RetimeWrapper_50_clock = clock; // @[:@27903.4]
  assign RetimeWrapper_50_reset = reset; // @[:@27904.4]
  assign RetimeWrapper_50_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27906.4]
  assign RetimeWrapper_50_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@27905.4]
  assign x420_sum_1_clock = clock; // @[:@27930.4]
  assign x420_sum_1_reset = reset; // @[:@27931.4]
  assign x420_sum_1_io_a = {_T_957,_T_958}; // @[Math.scala 151:17:@27932.4]
  assign x420_sum_1_io_b = {_T_631,_T_632}; // @[Math.scala 152:17:@27933.4]
  assign x420_sum_1_io_flow = io_in_x276_TREADY; // @[Math.scala 153:20:@27934.4]
  assign RetimeWrapper_51_clock = clock; // @[:@27940.4]
  assign RetimeWrapper_51_reset = reset; // @[:@27941.4]
  assign RetimeWrapper_51_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27943.4]
  assign RetimeWrapper_51_io_in = ~ x418; // @[package.scala 94:16:@27942.4]
  assign RetimeWrapper_52_clock = clock; // @[:@27952.4]
  assign RetimeWrapper_52_reset = reset; // @[:@27953.4]
  assign RetimeWrapper_52_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27955.4]
  assign RetimeWrapper_52_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@27954.4]
  assign x427_sum_1_clock = clock; // @[:@27979.4]
  assign x427_sum_1_reset = reset; // @[:@27980.4]
  assign x427_sum_1_io_a = {_T_957,_T_958}; // @[Math.scala 151:17:@27981.4]
  assign x427_sum_1_io_b = {_T_700,_T_701}; // @[Math.scala 152:17:@27982.4]
  assign x427_sum_1_io_flow = io_in_x276_TREADY; // @[Math.scala 153:20:@27983.4]
  assign RetimeWrapper_53_clock = clock; // @[:@27989.4]
  assign RetimeWrapper_53_reset = reset; // @[:@27990.4]
  assign RetimeWrapper_53_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27992.4]
  assign RetimeWrapper_53_io_in = ~ x425; // @[package.scala 94:16:@27991.4]
  assign RetimeWrapper_54_clock = clock; // @[:@28001.4]
  assign RetimeWrapper_54_reset = reset; // @[:@28002.4]
  assign RetimeWrapper_54_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28004.4]
  assign RetimeWrapper_54_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@28003.4]
  assign x437_x23_1_clock = clock; // @[:@28049.4]
  assign x437_x23_1_reset = reset; // @[:@28050.4]
  assign x437_x23_1_io_a = x288_lb_0_io_rPort_9_output_0; // @[Math.scala 151:17:@28051.4]
  assign x437_x23_1_io_b = _T_1080[7:0]; // @[Math.scala 152:17:@28052.4]
  assign x437_x23_1_io_flow = io_in_x276_TREADY; // @[Math.scala 153:20:@28053.4]
  assign x438_x24_1_clock = clock; // @[:@28059.4]
  assign x438_x24_1_reset = reset; // @[:@28060.4]
  assign x438_x24_1_io_a = x288_lb_0_io_rPort_7_output_0; // @[Math.scala 151:17:@28061.4]
  assign x438_x24_1_io_b = _T_1084[7:0]; // @[Math.scala 152:17:@28062.4]
  assign x438_x24_1_io_flow = io_in_x276_TREADY; // @[Math.scala 153:20:@28063.4]
  assign x439_x23_1_clock = clock; // @[:@28069.4]
  assign x439_x23_1_reset = reset; // @[:@28070.4]
  assign x439_x23_1_io_a = _T_1088[7:0]; // @[Math.scala 151:17:@28071.4]
  assign x439_x23_1_io_b = _T_1092[7:0]; // @[Math.scala 152:17:@28072.4]
  assign x439_x23_1_io_flow = io_in_x276_TREADY; // @[Math.scala 153:20:@28073.4]
  assign x440_x24_1_clock = clock; // @[:@28079.4]
  assign x440_x24_1_reset = reset; // @[:@28080.4]
  assign x440_x24_1_io_a = x288_lb_0_io_rPort_10_output_0; // @[Math.scala 151:17:@28081.4]
  assign x440_x24_1_io_b = _T_1096[7:0]; // @[Math.scala 152:17:@28082.4]
  assign x440_x24_1_io_flow = io_in_x276_TREADY; // @[Math.scala 153:20:@28083.4]
  assign x441_x23_1_io_a = x437_x23_1_io_result; // @[Math.scala 151:17:@28091.4]
  assign x441_x23_1_io_b = x438_x24_1_io_result; // @[Math.scala 152:17:@28092.4]
  assign x442_x24_1_io_a = x439_x23_1_io_result; // @[Math.scala 151:17:@28101.4]
  assign x442_x24_1_io_b = x440_x24_1_io_result; // @[Math.scala 152:17:@28102.4]
  assign x443_x23_1_io_a = x441_x23_1_io_result; // @[Math.scala 151:17:@28111.4]
  assign x443_x23_1_io_b = x442_x24_1_io_result; // @[Math.scala 152:17:@28112.4]
  assign RetimeWrapper_55_clock = clock; // @[:@28119.4]
  assign RetimeWrapper_55_reset = reset; // @[:@28120.4]
  assign RetimeWrapper_55_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28122.4]
  assign RetimeWrapper_55_io_in = x288_lb_0_io_rPort_5_output_0; // @[package.scala 94:16:@28121.4]
  assign x444_sum_1_io_a = x443_x23_1_io_result; // @[Math.scala 151:17:@28130.4]
  assign x444_sum_1_io_b = RetimeWrapper_55_io_out; // @[Math.scala 152:17:@28131.4]
  assign RetimeWrapper_56_clock = clock; // @[:@28142.4]
  assign RetimeWrapper_56_reset = reset; // @[:@28143.4]
  assign RetimeWrapper_56_io_flow = io_in_x276_TREADY; // @[package.scala 95:18:@28145.4]
  assign RetimeWrapper_56_io_in = {4'h0,_T_1132}; // @[package.scala 94:16:@28144.4]
  assign x451_x23_1_clock = clock; // @[:@28177.4]
  assign x451_x23_1_reset = reset; // @[:@28178.4]
  assign x451_x23_1_io_a = x288_lb_0_io_rPort_11_output_0; // @[Math.scala 151:17:@28179.4]
  assign x451_x23_1_io_b = _T_1139[7:0]; // @[Math.scala 152:17:@28180.4]
  assign x451_x23_1_io_flow = io_in_x276_TREADY; // @[Math.scala 153:20:@28181.4]
  assign x452_x24_1_clock = clock; // @[:@28187.4]
  assign x452_x24_1_reset = reset; // @[:@28188.4]
  assign x452_x24_1_io_a = x288_lb_0_io_rPort_8_output_0; // @[Math.scala 151:17:@28189.4]
  assign x452_x24_1_io_b = _T_1143[7:0]; // @[Math.scala 152:17:@28190.4]
  assign x452_x24_1_io_flow = io_in_x276_TREADY; // @[Math.scala 153:20:@28191.4]
  assign x453_x23_1_clock = clock; // @[:@28197.4]
  assign x453_x23_1_reset = reset; // @[:@28198.4]
  assign x453_x23_1_io_a = _T_1147[7:0]; // @[Math.scala 151:17:@28199.4]
  assign x453_x23_1_io_b = _T_1151[7:0]; // @[Math.scala 152:17:@28200.4]
  assign x453_x23_1_io_flow = io_in_x276_TREADY; // @[Math.scala 153:20:@28201.4]
  assign x454_x24_1_clock = clock; // @[:@28207.4]
  assign x454_x24_1_reset = reset; // @[:@28208.4]
  assign x454_x24_1_io_a = x288_lb_0_io_rPort_1_output_0; // @[Math.scala 151:17:@28209.4]
  assign x454_x24_1_io_b = _T_1155[7:0]; // @[Math.scala 152:17:@28210.4]
  assign x454_x24_1_io_flow = io_in_x276_TREADY; // @[Math.scala 153:20:@28211.4]
  assign x455_x23_1_io_a = x451_x23_1_io_result; // @[Math.scala 151:17:@28219.4]
  assign x455_x23_1_io_b = x452_x24_1_io_result; // @[Math.scala 152:17:@28220.4]
  assign x456_x24_1_io_a = x453_x23_1_io_result; // @[Math.scala 151:17:@28229.4]
  assign x456_x24_1_io_b = x454_x24_1_io_result; // @[Math.scala 152:17:@28230.4]
  assign x457_x23_1_io_a = x455_x23_1_io_result; // @[Math.scala 151:17:@28239.4]
  assign x457_x23_1_io_b = x456_x24_1_io_result; // @[Math.scala 152:17:@28240.4]
  assign RetimeWrapper_57_clock = clock; // @[:@28247.4]
  assign RetimeWrapper_57_reset = reset; // @[:@28248.4]
  assign RetimeWrapper_57_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28250.4]
  assign RetimeWrapper_57_io_in = x288_lb_0_io_rPort_3_output_0; // @[package.scala 94:16:@28249.4]
  assign x458_sum_1_io_a = x457_x23_1_io_result; // @[Math.scala 151:17:@28258.4]
  assign x458_sum_1_io_b = RetimeWrapper_57_io_out; // @[Math.scala 152:17:@28259.4]
  assign RetimeWrapper_58_clock = clock; // @[:@28270.4]
  assign RetimeWrapper_58_reset = reset; // @[:@28271.4]
  assign RetimeWrapper_58_io_flow = io_in_x276_TREADY; // @[package.scala 95:18:@28273.4]
  assign RetimeWrapper_58_io_in = {4'h0,_T_1191}; // @[package.scala 94:16:@28272.4]
  assign RetimeWrapper_59_clock = clock; // @[:@28280.4]
  assign RetimeWrapper_59_reset = reset; // @[:@28281.4]
  assign RetimeWrapper_59_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28283.4]
  assign RetimeWrapper_59_io_in = $unsigned(_T_323); // @[package.scala 94:16:@28282.4]
  assign RetimeWrapper_60_clock = clock; // @[:@28289.4]
  assign RetimeWrapper_60_reset = reset; // @[:@28290.4]
  assign RetimeWrapper_60_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28292.4]
  assign RetimeWrapper_60_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@28291.4]
  assign RetimeWrapper_61_clock = clock; // @[:@28298.4]
  assign RetimeWrapper_61_reset = reset; // @[:@28299.4]
  assign RetimeWrapper_61_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28301.4]
  assign RetimeWrapper_61_io_in = x303_sum_1_io_result; // @[package.scala 94:16:@28300.4]
  assign RetimeWrapper_62_clock = clock; // @[:@28307.4]
  assign RetimeWrapper_62_reset = reset; // @[:@28308.4]
  assign RetimeWrapper_62_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28310.4]
  assign RetimeWrapper_62_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@28309.4]
  assign RetimeWrapper_63_clock = clock; // @[:@28316.4]
  assign RetimeWrapper_63_reset = reset; // @[:@28317.4]
  assign RetimeWrapper_63_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28319.4]
  assign RetimeWrapper_63_io_in = $unsigned(_T_311); // @[package.scala 94:16:@28318.4]
  assign RetimeWrapper_64_clock = clock; // @[:@28327.4]
  assign RetimeWrapper_64_reset = reset; // @[:@28328.4]
  assign RetimeWrapper_64_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28330.4]
  assign RetimeWrapper_64_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@28329.4]
  assign RetimeWrapper_65_clock = clock; // @[:@28348.4]
  assign RetimeWrapper_65_reset = reset; // @[:@28349.4]
  assign RetimeWrapper_65_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28351.4]
  assign RetimeWrapper_65_io_in = $unsigned(_T_398); // @[package.scala 94:16:@28350.4]
  assign RetimeWrapper_66_clock = clock; // @[:@28357.4]
  assign RetimeWrapper_66_reset = reset; // @[:@28358.4]
  assign RetimeWrapper_66_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28360.4]
  assign RetimeWrapper_66_io_in = x313_sum_1_io_result; // @[package.scala 94:16:@28359.4]
  assign RetimeWrapper_67_clock = clock; // @[:@28368.4]
  assign RetimeWrapper_67_reset = reset; // @[:@28369.4]
  assign RetimeWrapper_67_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28371.4]
  assign RetimeWrapper_67_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@28370.4]
  assign RetimeWrapper_68_clock = clock; // @[:@28389.4]
  assign RetimeWrapper_68_reset = reset; // @[:@28390.4]
  assign RetimeWrapper_68_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28392.4]
  assign RetimeWrapper_68_io_in = ~ x322; // @[package.scala 94:16:@28391.4]
  assign RetimeWrapper_69_clock = clock; // @[:@28398.4]
  assign RetimeWrapper_69_reset = reset; // @[:@28399.4]
  assign RetimeWrapper_69_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28401.4]
  assign RetimeWrapper_69_io_in = $unsigned(_T_487); // @[package.scala 94:16:@28400.4]
  assign RetimeWrapper_70_clock = clock; // @[:@28407.4]
  assign RetimeWrapper_70_reset = reset; // @[:@28408.4]
  assign RetimeWrapper_70_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28410.4]
  assign RetimeWrapper_70_io_in = x326_sum_1_io_result; // @[package.scala 94:16:@28409.4]
  assign RetimeWrapper_71_clock = clock; // @[:@28419.4]
  assign RetimeWrapper_71_reset = reset; // @[:@28420.4]
  assign RetimeWrapper_71_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28422.4]
  assign RetimeWrapper_71_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@28421.4]
  assign RetimeWrapper_72_clock = clock; // @[:@28440.4]
  assign RetimeWrapper_72_reset = reset; // @[:@28441.4]
  assign RetimeWrapper_72_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28443.4]
  assign RetimeWrapper_72_io_in = ~ x333; // @[package.scala 94:16:@28442.4]
  assign RetimeWrapper_73_clock = clock; // @[:@28449.4]
  assign RetimeWrapper_73_reset = reset; // @[:@28450.4]
  assign RetimeWrapper_73_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28452.4]
  assign RetimeWrapper_73_io_in = x335_sum_1_io_result; // @[package.scala 94:16:@28451.4]
  assign RetimeWrapper_74_clock = clock; // @[:@28461.4]
  assign RetimeWrapper_74_reset = reset; // @[:@28462.4]
  assign RetimeWrapper_74_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28464.4]
  assign RetimeWrapper_74_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@28463.4]
  assign RetimeWrapper_75_clock = clock; // @[:@28482.4]
  assign RetimeWrapper_75_reset = reset; // @[:@28483.4]
  assign RetimeWrapper_75_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28485.4]
  assign RetimeWrapper_75_io_in = $unsigned(_T_622); // @[package.scala 94:16:@28484.4]
  assign RetimeWrapper_76_clock = clock; // @[:@28491.4]
  assign RetimeWrapper_76_reset = reset; // @[:@28492.4]
  assign RetimeWrapper_76_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28494.4]
  assign RetimeWrapper_76_io_in = ~ x342; // @[package.scala 94:16:@28493.4]
  assign RetimeWrapper_77_clock = clock; // @[:@28500.4]
  assign RetimeWrapper_77_reset = reset; // @[:@28501.4]
  assign RetimeWrapper_77_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28503.4]
  assign RetimeWrapper_77_io_in = x346_sum_1_io_result; // @[package.scala 94:16:@28502.4]
  assign RetimeWrapper_78_clock = clock; // @[:@28512.4]
  assign RetimeWrapper_78_reset = reset; // @[:@28513.4]
  assign RetimeWrapper_78_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28515.4]
  assign RetimeWrapper_78_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@28514.4]
  assign RetimeWrapper_79_clock = clock; // @[:@28533.4]
  assign RetimeWrapper_79_reset = reset; // @[:@28534.4]
  assign RetimeWrapper_79_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28536.4]
  assign RetimeWrapper_79_io_in = x371_sum_1_io_result; // @[package.scala 94:16:@28535.4]
  assign RetimeWrapper_80_clock = clock; // @[:@28542.4]
  assign RetimeWrapper_80_reset = reset; // @[:@28543.4]
  assign RetimeWrapper_80_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28545.4]
  assign RetimeWrapper_80_io_in = ~ x367; // @[package.scala 94:16:@28544.4]
  assign RetimeWrapper_81_clock = clock; // @[:@28551.4]
  assign RetimeWrapper_81_reset = reset; // @[:@28552.4]
  assign RetimeWrapper_81_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28554.4]
  assign RetimeWrapper_81_io_in = $unsigned(_T_772); // @[package.scala 94:16:@28553.4]
  assign RetimeWrapper_82_clock = clock; // @[:@28563.4]
  assign RetimeWrapper_82_reset = reset; // @[:@28564.4]
  assign RetimeWrapper_82_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28566.4]
  assign RetimeWrapper_82_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@28565.4]
  assign RetimeWrapper_83_clock = clock; // @[:@28584.4]
  assign RetimeWrapper_83_reset = reset; // @[:@28585.4]
  assign RetimeWrapper_83_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28587.4]
  assign RetimeWrapper_83_io_in = x379_sum_1_io_result; // @[package.scala 94:16:@28586.4]
  assign RetimeWrapper_84_clock = clock; // @[:@28593.4]
  assign RetimeWrapper_84_reset = reset; // @[:@28594.4]
  assign RetimeWrapper_84_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28596.4]
  assign RetimeWrapper_84_io_in = ~ x377; // @[package.scala 94:16:@28595.4]
  assign RetimeWrapper_85_clock = clock; // @[:@28605.4]
  assign RetimeWrapper_85_reset = reset; // @[:@28606.4]
  assign RetimeWrapper_85_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28608.4]
  assign RetimeWrapper_85_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@28607.4]
  assign RetimeWrapper_86_clock = clock; // @[:@28626.4]
  assign RetimeWrapper_86_reset = reset; // @[:@28627.4]
  assign RetimeWrapper_86_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28629.4]
  assign RetimeWrapper_86_io_in = ~ x384; // @[package.scala 94:16:@28628.4]
  assign RetimeWrapper_87_clock = clock; // @[:@28635.4]
  assign RetimeWrapper_87_reset = reset; // @[:@28636.4]
  assign RetimeWrapper_87_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28638.4]
  assign RetimeWrapper_87_io_in = x386_sum_1_io_result; // @[package.scala 94:16:@28637.4]
  assign RetimeWrapper_88_clock = clock; // @[:@28647.4]
  assign RetimeWrapper_88_reset = reset; // @[:@28648.4]
  assign RetimeWrapper_88_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28650.4]
  assign RetimeWrapper_88_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@28649.4]
  assign x478_x25_1_io_a = x289_lb2_0_io_rPort_5_output_0; // @[Math.scala 151:17:@28682.4]
  assign x478_x25_1_io_b = _T_1408[7:0]; // @[Math.scala 152:17:@28683.4]
  assign x479_x26_1_io_a = _T_1412[7:0]; // @[Math.scala 151:17:@28692.4]
  assign x479_x26_1_io_b = x289_lb2_0_io_rPort_1_output_0; // @[Math.scala 152:17:@28693.4]
  assign x480_sum_1_io_a = x478_x25_1_io_result; // @[Math.scala 151:17:@28702.4]
  assign x480_sum_1_io_b = x479_x26_1_io_result; // @[Math.scala 152:17:@28703.4]
  assign x481_div_1_clock = clock; // @[:@28712.4]
  assign x481_div_1_reset = reset; // @[:@28713.4]
  assign x481_div_1_io_a = x480_sum_1_io_result; // @[Math.scala 328:17:@28714.4]
  assign x481_div_1_io_flow = io_in_x276_TREADY; // @[Math.scala 330:20:@28716.4]
  assign x484_x25_1_io_a = x289_lb2_0_io_rPort_2_output_0; // @[Math.scala 151:17:@28734.4]
  assign x484_x25_1_io_b = _T_1432[7:0]; // @[Math.scala 152:17:@28735.4]
  assign x485_x26_1_io_a = _T_1436[7:0]; // @[Math.scala 151:17:@28744.4]
  assign x485_x26_1_io_b = x289_lb2_0_io_rPort_4_output_0; // @[Math.scala 152:17:@28745.4]
  assign x486_sum_1_io_a = x484_x25_1_io_result; // @[Math.scala 151:17:@28754.4]
  assign x486_sum_1_io_b = x485_x26_1_io_result; // @[Math.scala 152:17:@28755.4]
  assign x487_div_1_clock = clock; // @[:@28764.4]
  assign x487_div_1_reset = reset; // @[:@28765.4]
  assign x487_div_1_io_a = x486_sum_1_io_result; // @[Math.scala 328:17:@28766.4]
  assign x487_div_1_io_flow = io_in_x276_TREADY; // @[Math.scala 330:20:@28768.4]
  assign RetimeWrapper_89_clock = clock; // @[:@28780.4]
  assign RetimeWrapper_89_reset = reset; // @[:@28781.4]
  assign RetimeWrapper_89_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28783.4]
  assign RetimeWrapper_89_io_in = {x481_div_number,x487_div_number}; // @[package.scala 94:16:@28782.4]
  assign RetimeWrapper_90_clock = clock; // @[:@28789.4]
  assign RetimeWrapper_90_reset = reset; // @[:@28790.4]
  assign RetimeWrapper_90_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28792.4]
  assign RetimeWrapper_90_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@28791.4]
  assign RetimeWrapper_91_clock = clock; // @[:@28798.4]
  assign RetimeWrapper_91_reset = reset; // @[:@28799.4]
  assign RetimeWrapper_91_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28801.4]
  assign RetimeWrapper_91_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@28800.4]
  assign RetimeWrapper_92_clock = clock; // @[:@28807.4]
  assign RetimeWrapper_92_reset = reset; // @[:@28808.4]
  assign RetimeWrapper_92_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28810.4]
  assign RetimeWrapper_92_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@28809.4]
endmodule
module x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1( // @[:@28828.2]
  input          clock, // @[:@28829.4]
  input          reset, // @[:@28830.4]
  output         io_in_x276_TVALID, // @[:@28831.4]
  input          io_in_x276_TREADY, // @[:@28831.4]
  output [255:0] io_in_x276_TDATA, // @[:@28831.4]
  input          io_in_x275_TVALID, // @[:@28831.4]
  output         io_in_x275_TREADY, // @[:@28831.4]
  input  [255:0] io_in_x275_TDATA, // @[:@28831.4]
  input  [7:0]   io_in_x275_TID, // @[:@28831.4]
  input  [7:0]   io_in_x275_TDEST, // @[:@28831.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@28831.4]
  input          io_sigsIn_smChildAcks_0, // @[:@28831.4]
  output         io_sigsOut_smDoneIn_0, // @[:@28831.4]
  output         io_sigsOut_smCtrCopyDone_0, // @[:@28831.4]
  input          io_rr // @[:@28831.4]
);
  wire  x283_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@28841.4]
  wire  x283_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@28841.4]
  wire  x283_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@28841.4]
  wire  x283_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@28841.4]
  wire [31:0] x283_ctrchain_io_output_counts_1; // @[SpatialBlocks.scala 37:22:@28841.4]
  wire [31:0] x283_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@28841.4]
  wire  x283_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@28841.4]
  wire  x283_ctrchain_io_output_oobs_1; // @[SpatialBlocks.scala 37:22:@28841.4]
  wire  x283_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@28841.4]
  wire  x492_inr_Foreach_SAMPLER_BOX_sm_clock; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 32:18:@28900.4]
  wire  x492_inr_Foreach_SAMPLER_BOX_sm_reset; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 32:18:@28900.4]
  wire  x492_inr_Foreach_SAMPLER_BOX_sm_io_enable; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 32:18:@28900.4]
  wire  x492_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 32:18:@28900.4]
  wire  x492_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 32:18:@28900.4]
  wire  x492_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 32:18:@28900.4]
  wire  x492_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 32:18:@28900.4]
  wire  x492_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 32:18:@28900.4]
  wire  x492_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 32:18:@28900.4]
  wire  x492_inr_Foreach_SAMPLER_BOX_sm_io_parentAck; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 32:18:@28900.4]
  wire  x492_inr_Foreach_SAMPLER_BOX_sm_io_backpressure; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 32:18:@28900.4]
  wire  x492_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 32:18:@28900.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@28928.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@28928.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@28928.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@28928.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@28928.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@28970.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@28970.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@28970.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@28970.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@28970.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@28978.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@28978.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@28978.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@28978.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@28978.4]
  wire  x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_clock; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 643:24:@29010.4]
  wire  x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_reset; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 643:24:@29010.4]
  wire  x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x276_TVALID; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 643:24:@29010.4]
  wire  x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x276_TREADY; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 643:24:@29010.4]
  wire [255:0] x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x276_TDATA; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 643:24:@29010.4]
  wire  x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x275_TREADY; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 643:24:@29010.4]
  wire [255:0] x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x275_TDATA; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 643:24:@29010.4]
  wire [7:0] x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x275_TID; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 643:24:@29010.4]
  wire [7:0] x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x275_TDEST; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 643:24:@29010.4]
  wire  x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 643:24:@29010.4]
  wire  x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 643:24:@29010.4]
  wire  x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 643:24:@29010.4]
  wire [31:0] x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 643:24:@29010.4]
  wire [31:0] x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 643:24:@29010.4]
  wire  x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 643:24:@29010.4]
  wire  x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 643:24:@29010.4]
  wire  x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_rr; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 643:24:@29010.4]
  wire  _T_239; // @[package.scala 96:25:@28933.4 package.scala 96:25:@28934.4]
  wire  x492_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[sm_x493_outr_UnitPipe.scala 68:66:@28939.4]
  wire  _T_252; // @[package.scala 96:25:@28975.4 package.scala 96:25:@28976.4]
  wire  _T_258; // @[package.scala 96:25:@28983.4 package.scala 96:25:@28984.4]
  wire  _T_261; // @[SpatialBlocks.scala 110:93:@28986.4]
  wire  x492_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn; // @[SpatialBlocks.scala 110:90:@28987.4]
  wire  _T_263; // @[SpatialBlocks.scala 128:36:@28995.4]
  wire  _T_264; // @[SpatialBlocks.scala 128:78:@28996.4]
  wire  _T_269; // @[SpatialBlocks.scala 130:61:@29005.4]
  x283_ctrchain x283_ctrchain ( // @[SpatialBlocks.scala 37:22:@28841.4]
    .clock(x283_ctrchain_clock),
    .reset(x283_ctrchain_reset),
    .io_input_reset(x283_ctrchain_io_input_reset),
    .io_input_enable(x283_ctrchain_io_input_enable),
    .io_output_counts_1(x283_ctrchain_io_output_counts_1),
    .io_output_counts_0(x283_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x283_ctrchain_io_output_oobs_0),
    .io_output_oobs_1(x283_ctrchain_io_output_oobs_1),
    .io_output_done(x283_ctrchain_io_output_done)
  );
  x492_inr_Foreach_SAMPLER_BOX_sm x492_inr_Foreach_SAMPLER_BOX_sm ( // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 32:18:@28900.4]
    .clock(x492_inr_Foreach_SAMPLER_BOX_sm_clock),
    .reset(x492_inr_Foreach_SAMPLER_BOX_sm_reset),
    .io_enable(x492_inr_Foreach_SAMPLER_BOX_sm_io_enable),
    .io_done(x492_inr_Foreach_SAMPLER_BOX_sm_io_done),
    .io_doneLatch(x492_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch),
    .io_ctrDone(x492_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone),
    .io_datapathEn(x492_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn),
    .io_ctrInc(x492_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc),
    .io_ctrRst(x492_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst),
    .io_parentAck(x492_inr_Foreach_SAMPLER_BOX_sm_io_parentAck),
    .io_backpressure(x492_inr_Foreach_SAMPLER_BOX_sm_io_backpressure),
    .io_break(x492_inr_Foreach_SAMPLER_BOX_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@28928.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@28970.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@28978.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1 x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1 ( // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 643:24:@29010.4]
    .clock(x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_clock),
    .reset(x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_reset),
    .io_in_x276_TVALID(x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x276_TVALID),
    .io_in_x276_TREADY(x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x276_TREADY),
    .io_in_x276_TDATA(x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x276_TDATA),
    .io_in_x275_TREADY(x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x275_TREADY),
    .io_in_x275_TDATA(x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x275_TDATA),
    .io_in_x275_TID(x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x275_TID),
    .io_in_x275_TDEST(x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x275_TDEST),
    .io_sigsIn_backpressure(x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_1(x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsIn_cchainOutputs_0_oobs_1(x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1),
    .io_rr(x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_rr)
  );
  assign _T_239 = RetimeWrapper_io_out; // @[package.scala 96:25:@28933.4 package.scala 96:25:@28934.4]
  assign x492_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure = io_in_x275_TVALID | x492_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x493_outr_UnitPipe.scala 68:66:@28939.4]
  assign _T_252 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@28975.4 package.scala 96:25:@28976.4]
  assign _T_258 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@28983.4 package.scala 96:25:@28984.4]
  assign _T_261 = ~ _T_258; // @[SpatialBlocks.scala 110:93:@28986.4]
  assign x492_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn = _T_252 & _T_261; // @[SpatialBlocks.scala 110:90:@28987.4]
  assign _T_263 = x492_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[SpatialBlocks.scala 128:36:@28995.4]
  assign _T_264 = ~ x492_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[SpatialBlocks.scala 128:78:@28996.4]
  assign _T_269 = x492_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[SpatialBlocks.scala 130:61:@29005.4]
  assign io_in_x276_TVALID = x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x276_TVALID; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 48:23:@29068.4]
  assign io_in_x276_TDATA = x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x276_TDATA; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 48:23:@29066.4]
  assign io_in_x275_TREADY = x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x275_TREADY; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 49:23:@29076.4]
  assign io_sigsOut_smDoneIn_0 = x492_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[SpatialBlocks.scala 127:53:@28993.4]
  assign io_sigsOut_smCtrCopyDone_0 = x492_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[SpatialBlocks.scala 139:125:@29009.4]
  assign x283_ctrchain_clock = clock; // @[:@28842.4]
  assign x283_ctrchain_reset = reset; // @[:@28843.4]
  assign x283_ctrchain_io_input_reset = x492_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[SpatialBlocks.scala 130:103:@29008.4]
  assign x283_ctrchain_io_input_enable = _T_269 & x492_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 104:75:@28963.4 SpatialBlocks.scala 130:45:@29007.4]
  assign x492_inr_Foreach_SAMPLER_BOX_sm_clock = clock; // @[:@28901.4]
  assign x492_inr_Foreach_SAMPLER_BOX_sm_reset = reset; // @[:@28902.4]
  assign x492_inr_Foreach_SAMPLER_BOX_sm_io_enable = x492_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn & x492_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 112:18:@28990.4]
  assign x492_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone = io_rr ? _T_239 : 1'h0; // @[sm_x493_outr_UnitPipe.scala 66:50:@28936.4]
  assign x492_inr_Foreach_SAMPLER_BOX_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 114:21:@28992.4]
  assign x492_inr_Foreach_SAMPLER_BOX_sm_io_backpressure = io_in_x276_TREADY | x492_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[SpatialBlocks.scala 105:24:@28964.4]
  assign x492_inr_Foreach_SAMPLER_BOX_sm_io_break = 1'h0; // @[sm_x493_outr_UnitPipe.scala 70:48:@28942.4]
  assign RetimeWrapper_clock = clock; // @[:@28929.4]
  assign RetimeWrapper_reset = reset; // @[:@28930.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@28932.4]
  assign RetimeWrapper_io_in = x283_ctrchain_io_output_done; // @[package.scala 94:16:@28931.4]
  assign RetimeWrapper_1_clock = clock; // @[:@28971.4]
  assign RetimeWrapper_1_reset = reset; // @[:@28972.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@28974.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@28973.4]
  assign RetimeWrapper_2_clock = clock; // @[:@28979.4]
  assign RetimeWrapper_2_reset = reset; // @[:@28980.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@28982.4]
  assign RetimeWrapper_2_io_in = x492_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[package.scala 94:16:@28981.4]
  assign x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_clock = clock; // @[:@29011.4]
  assign x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_reset = reset; // @[:@29012.4]
  assign x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x276_TREADY = io_in_x276_TREADY; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 48:23:@29067.4]
  assign x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x275_TDATA = io_in_x275_TDATA; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 49:23:@29075.4]
  assign x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x275_TID = io_in_x275_TID; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 49:23:@29071.4]
  assign x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x275_TDEST = io_in_x275_TDEST; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 49:23:@29070.4]
  assign x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure = io_in_x276_TREADY | x492_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 647:22:@29094.4]
  assign x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn = _T_263 & _T_264; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 647:22:@29092.4]
  assign x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break = x492_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 647:22:@29090.4]
  assign x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1 = x283_ctrchain_io_output_counts_1; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 647:22:@29085.4]
  assign x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = x283_ctrchain_io_output_counts_0; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 647:22:@29084.4]
  assign x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x283_ctrchain_io_output_oobs_0; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 647:22:@29082.4]
  assign x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1 = x283_ctrchain_io_output_oobs_1; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 647:22:@29083.4]
  assign x492_inr_Foreach_SAMPLER_BOX_kernelx492_inr_Foreach_SAMPLER_BOX_concrete1_io_rr = io_rr; // @[sm_x492_inr_Foreach_SAMPLER_BOX.scala 646:18:@29078.4]
endmodule
module RootController_kernelRootController_concrete1( // @[:@29107.2]
  input          clock, // @[:@29108.4]
  input          reset, // @[:@29109.4]
  output         io_in_x276_TVALID, // @[:@29110.4]
  input          io_in_x276_TREADY, // @[:@29110.4]
  output [255:0] io_in_x276_TDATA, // @[:@29110.4]
  input          io_in_x275_TVALID, // @[:@29110.4]
  output         io_in_x275_TREADY, // @[:@29110.4]
  input  [255:0] io_in_x275_TDATA, // @[:@29110.4]
  input  [7:0]   io_in_x275_TID, // @[:@29110.4]
  input  [7:0]   io_in_x275_TDEST, // @[:@29110.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@29110.4]
  input          io_sigsIn_smChildAcks_0, // @[:@29110.4]
  output         io_sigsOut_smDoneIn_0, // @[:@29110.4]
  input          io_rr // @[:@29110.4]
);
  wire  x493_outr_UnitPipe_sm_clock; // @[sm_x493_outr_UnitPipe.scala 32:18:@29251.4]
  wire  x493_outr_UnitPipe_sm_reset; // @[sm_x493_outr_UnitPipe.scala 32:18:@29251.4]
  wire  x493_outr_UnitPipe_sm_io_enable; // @[sm_x493_outr_UnitPipe.scala 32:18:@29251.4]
  wire  x493_outr_UnitPipe_sm_io_done; // @[sm_x493_outr_UnitPipe.scala 32:18:@29251.4]
  wire  x493_outr_UnitPipe_sm_io_parentAck; // @[sm_x493_outr_UnitPipe.scala 32:18:@29251.4]
  wire  x493_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x493_outr_UnitPipe.scala 32:18:@29251.4]
  wire  x493_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x493_outr_UnitPipe.scala 32:18:@29251.4]
  wire  x493_outr_UnitPipe_sm_io_childAck_0; // @[sm_x493_outr_UnitPipe.scala 32:18:@29251.4]
  wire  x493_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x493_outr_UnitPipe.scala 32:18:@29251.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@29303.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@29303.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@29303.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@29303.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@29303.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@29311.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@29311.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@29311.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@29311.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@29311.4]
  wire  x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_clock; // @[sm_x493_outr_UnitPipe.scala 75:24:@29338.4]
  wire  x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_reset; // @[sm_x493_outr_UnitPipe.scala 75:24:@29338.4]
  wire  x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x276_TVALID; // @[sm_x493_outr_UnitPipe.scala 75:24:@29338.4]
  wire  x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x276_TREADY; // @[sm_x493_outr_UnitPipe.scala 75:24:@29338.4]
  wire [255:0] x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x276_TDATA; // @[sm_x493_outr_UnitPipe.scala 75:24:@29338.4]
  wire  x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x275_TVALID; // @[sm_x493_outr_UnitPipe.scala 75:24:@29338.4]
  wire  x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x275_TREADY; // @[sm_x493_outr_UnitPipe.scala 75:24:@29338.4]
  wire [255:0] x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x275_TDATA; // @[sm_x493_outr_UnitPipe.scala 75:24:@29338.4]
  wire [7:0] x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x275_TID; // @[sm_x493_outr_UnitPipe.scala 75:24:@29338.4]
  wire [7:0] x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x275_TDEST; // @[sm_x493_outr_UnitPipe.scala 75:24:@29338.4]
  wire  x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x493_outr_UnitPipe.scala 75:24:@29338.4]
  wire  x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x493_outr_UnitPipe.scala 75:24:@29338.4]
  wire  x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x493_outr_UnitPipe.scala 75:24:@29338.4]
  wire  x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x493_outr_UnitPipe.scala 75:24:@29338.4]
  wire  x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_rr; // @[sm_x493_outr_UnitPipe.scala 75:24:@29338.4]
  wire  _T_246; // @[package.scala 96:25:@29308.4 package.scala 96:25:@29309.4]
  wire  _T_252; // @[package.scala 96:25:@29316.4 package.scala 96:25:@29317.4]
  wire  _T_255; // @[SpatialBlocks.scala 110:93:@29319.4]
  x493_outr_UnitPipe_sm x493_outr_UnitPipe_sm ( // @[sm_x493_outr_UnitPipe.scala 32:18:@29251.4]
    .clock(x493_outr_UnitPipe_sm_clock),
    .reset(x493_outr_UnitPipe_sm_reset),
    .io_enable(x493_outr_UnitPipe_sm_io_enable),
    .io_done(x493_outr_UnitPipe_sm_io_done),
    .io_parentAck(x493_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x493_outr_UnitPipe_sm_io_doneIn_0),
    .io_enableOut_0(x493_outr_UnitPipe_sm_io_enableOut_0),
    .io_childAck_0(x493_outr_UnitPipe_sm_io_childAck_0),
    .io_ctrCopyDone_0(x493_outr_UnitPipe_sm_io_ctrCopyDone_0)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@29303.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@29311.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1 x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1 ( // @[sm_x493_outr_UnitPipe.scala 75:24:@29338.4]
    .clock(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_clock),
    .reset(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_reset),
    .io_in_x276_TVALID(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x276_TVALID),
    .io_in_x276_TREADY(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x276_TREADY),
    .io_in_x276_TDATA(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x276_TDATA),
    .io_in_x275_TVALID(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x275_TVALID),
    .io_in_x275_TREADY(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x275_TREADY),
    .io_in_x275_TDATA(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x275_TDATA),
    .io_in_x275_TID(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x275_TID),
    .io_in_x275_TDEST(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x275_TDEST),
    .io_sigsIn_smEnableOuts_0(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smCtrCopyDone_0(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_rr(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_246 = RetimeWrapper_io_out; // @[package.scala 96:25:@29308.4 package.scala 96:25:@29309.4]
  assign _T_252 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@29316.4 package.scala 96:25:@29317.4]
  assign _T_255 = ~ _T_252; // @[SpatialBlocks.scala 110:93:@29319.4]
  assign io_in_x276_TVALID = x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x276_TVALID; // @[sm_x493_outr_UnitPipe.scala 48:23:@29394.4]
  assign io_in_x276_TDATA = x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x276_TDATA; // @[sm_x493_outr_UnitPipe.scala 48:23:@29392.4]
  assign io_in_x275_TREADY = x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x275_TREADY; // @[sm_x493_outr_UnitPipe.scala 49:23:@29402.4]
  assign io_sigsOut_smDoneIn_0 = x493_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 127:53:@29326.4]
  assign x493_outr_UnitPipe_sm_clock = clock; // @[:@29252.4]
  assign x493_outr_UnitPipe_sm_reset = reset; // @[:@29253.4]
  assign x493_outr_UnitPipe_sm_io_enable = _T_246 & _T_255; // @[SpatialBlocks.scala 112:18:@29323.4]
  assign x493_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 114:21:@29325.4]
  assign x493_outr_UnitPipe_sm_io_doneIn_0 = x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 102:67:@29295.4]
  assign x493_outr_UnitPipe_sm_io_ctrCopyDone_0 = x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 132:80:@29337.4]
  assign RetimeWrapper_clock = clock; // @[:@29304.4]
  assign RetimeWrapper_reset = reset; // @[:@29305.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@29307.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@29306.4]
  assign RetimeWrapper_1_clock = clock; // @[:@29312.4]
  assign RetimeWrapper_1_reset = reset; // @[:@29313.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@29315.4]
  assign RetimeWrapper_1_io_in = x493_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@29314.4]
  assign x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_clock = clock; // @[:@29339.4]
  assign x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_reset = reset; // @[:@29340.4]
  assign x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x276_TREADY = io_in_x276_TREADY; // @[sm_x493_outr_UnitPipe.scala 48:23:@29393.4]
  assign x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x275_TVALID = io_in_x275_TVALID; // @[sm_x493_outr_UnitPipe.scala 49:23:@29403.4]
  assign x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x275_TDATA = io_in_x275_TDATA; // @[sm_x493_outr_UnitPipe.scala 49:23:@29401.4]
  assign x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x275_TID = io_in_x275_TID; // @[sm_x493_outr_UnitPipe.scala 49:23:@29397.4]
  assign x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x275_TDEST = io_in_x275_TDEST; // @[sm_x493_outr_UnitPipe.scala 49:23:@29396.4]
  assign x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x493_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x493_outr_UnitPipe.scala 79:22:@29412.4]
  assign x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x493_outr_UnitPipe_sm_io_childAck_0; // @[sm_x493_outr_UnitPipe.scala 79:22:@29410.4]
  assign x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x493_outr_UnitPipe.scala 78:18:@29404.4]
endmodule
module AccelUnit( // @[:@29431.2]
  input          clock, // @[:@29432.4]
  input          reset, // @[:@29433.4]
  input          io_enable, // @[:@29434.4]
  output         io_done, // @[:@29434.4]
  input          io_reset, // @[:@29434.4]
  input          io_memStreams_loads_0_cmd_ready, // @[:@29434.4]
  output         io_memStreams_loads_0_cmd_valid, // @[:@29434.4]
  output [63:0]  io_memStreams_loads_0_cmd_bits_addr, // @[:@29434.4]
  output [31:0]  io_memStreams_loads_0_cmd_bits_size, // @[:@29434.4]
  output         io_memStreams_loads_0_data_ready, // @[:@29434.4]
  input          io_memStreams_loads_0_data_valid, // @[:@29434.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_0, // @[:@29434.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_1, // @[:@29434.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_2, // @[:@29434.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_3, // @[:@29434.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_4, // @[:@29434.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_5, // @[:@29434.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_6, // @[:@29434.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_7, // @[:@29434.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_8, // @[:@29434.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_9, // @[:@29434.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_10, // @[:@29434.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_11, // @[:@29434.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_12, // @[:@29434.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_13, // @[:@29434.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_14, // @[:@29434.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_15, // @[:@29434.4]
  input          io_memStreams_stores_0_cmd_ready, // @[:@29434.4]
  output         io_memStreams_stores_0_cmd_valid, // @[:@29434.4]
  output [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@29434.4]
  output [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@29434.4]
  input          io_memStreams_stores_0_data_ready, // @[:@29434.4]
  output         io_memStreams_stores_0_data_valid, // @[:@29434.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_0, // @[:@29434.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_1, // @[:@29434.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_2, // @[:@29434.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_3, // @[:@29434.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_4, // @[:@29434.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_5, // @[:@29434.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_6, // @[:@29434.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_7, // @[:@29434.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_8, // @[:@29434.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_9, // @[:@29434.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_10, // @[:@29434.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_11, // @[:@29434.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_12, // @[:@29434.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_13, // @[:@29434.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_14, // @[:@29434.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_15, // @[:@29434.4]
  output [15:0]  io_memStreams_stores_0_data_bits_wstrb, // @[:@29434.4]
  output         io_memStreams_stores_0_wresp_ready, // @[:@29434.4]
  input          io_memStreams_stores_0_wresp_valid, // @[:@29434.4]
  input          io_memStreams_stores_0_wresp_bits, // @[:@29434.4]
  input          io_memStreams_gathers_0_cmd_ready, // @[:@29434.4]
  output         io_memStreams_gathers_0_cmd_valid, // @[:@29434.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_0, // @[:@29434.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_1, // @[:@29434.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_2, // @[:@29434.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_3, // @[:@29434.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_4, // @[:@29434.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_5, // @[:@29434.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_6, // @[:@29434.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_7, // @[:@29434.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_8, // @[:@29434.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_9, // @[:@29434.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_10, // @[:@29434.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_11, // @[:@29434.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_12, // @[:@29434.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_13, // @[:@29434.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_14, // @[:@29434.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_15, // @[:@29434.4]
  output         io_memStreams_gathers_0_data_ready, // @[:@29434.4]
  input          io_memStreams_gathers_0_data_valid, // @[:@29434.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_0, // @[:@29434.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_1, // @[:@29434.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_2, // @[:@29434.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_3, // @[:@29434.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_4, // @[:@29434.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_5, // @[:@29434.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_6, // @[:@29434.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_7, // @[:@29434.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_8, // @[:@29434.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_9, // @[:@29434.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_10, // @[:@29434.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_11, // @[:@29434.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_12, // @[:@29434.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_13, // @[:@29434.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_14, // @[:@29434.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_15, // @[:@29434.4]
  input          io_memStreams_scatters_0_cmd_ready, // @[:@29434.4]
  output         io_memStreams_scatters_0_cmd_valid, // @[:@29434.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_0, // @[:@29434.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_1, // @[:@29434.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_2, // @[:@29434.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_3, // @[:@29434.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_4, // @[:@29434.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_5, // @[:@29434.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_6, // @[:@29434.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_7, // @[:@29434.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_8, // @[:@29434.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_9, // @[:@29434.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_10, // @[:@29434.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_11, // @[:@29434.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_12, // @[:@29434.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_13, // @[:@29434.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_14, // @[:@29434.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_15, // @[:@29434.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_0, // @[:@29434.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_1, // @[:@29434.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_2, // @[:@29434.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_3, // @[:@29434.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_4, // @[:@29434.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_5, // @[:@29434.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_6, // @[:@29434.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_7, // @[:@29434.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_8, // @[:@29434.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_9, // @[:@29434.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_10, // @[:@29434.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_11, // @[:@29434.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_12, // @[:@29434.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_13, // @[:@29434.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_14, // @[:@29434.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_15, // @[:@29434.4]
  output         io_memStreams_scatters_0_wresp_ready, // @[:@29434.4]
  input          io_memStreams_scatters_0_wresp_valid, // @[:@29434.4]
  input          io_memStreams_scatters_0_wresp_bits, // @[:@29434.4]
  input          io_axiStreamsIn_0_TVALID, // @[:@29434.4]
  output         io_axiStreamsIn_0_TREADY, // @[:@29434.4]
  input  [255:0] io_axiStreamsIn_0_TDATA, // @[:@29434.4]
  input  [31:0]  io_axiStreamsIn_0_TSTRB, // @[:@29434.4]
  input  [31:0]  io_axiStreamsIn_0_TKEEP, // @[:@29434.4]
  input          io_axiStreamsIn_0_TLAST, // @[:@29434.4]
  input  [7:0]   io_axiStreamsIn_0_TID, // @[:@29434.4]
  input  [7:0]   io_axiStreamsIn_0_TDEST, // @[:@29434.4]
  input  [31:0]  io_axiStreamsIn_0_TUSER, // @[:@29434.4]
  output         io_axiStreamsOut_0_TVALID, // @[:@29434.4]
  input          io_axiStreamsOut_0_TREADY, // @[:@29434.4]
  output [255:0] io_axiStreamsOut_0_TDATA, // @[:@29434.4]
  output [31:0]  io_axiStreamsOut_0_TSTRB, // @[:@29434.4]
  output [31:0]  io_axiStreamsOut_0_TKEEP, // @[:@29434.4]
  output         io_axiStreamsOut_0_TLAST, // @[:@29434.4]
  output [7:0]   io_axiStreamsOut_0_TID, // @[:@29434.4]
  output [7:0]   io_axiStreamsOut_0_TDEST, // @[:@29434.4]
  output [31:0]  io_axiStreamsOut_0_TUSER, // @[:@29434.4]
  output         io_heap_0_req_valid, // @[:@29434.4]
  output         io_heap_0_req_bits_allocDealloc, // @[:@29434.4]
  output [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@29434.4]
  input          io_heap_0_resp_valid, // @[:@29434.4]
  input          io_heap_0_resp_bits_allocDealloc, // @[:@29434.4]
  input  [63:0]  io_heap_0_resp_bits_sizeAddr, // @[:@29434.4]
  input  [63:0]  io_argIns_0, // @[:@29434.4]
  input  [63:0]  io_argIns_1, // @[:@29434.4]
  input          io_argOuts_0_port_ready, // @[:@29434.4]
  output         io_argOuts_0_port_valid, // @[:@29434.4]
  output [63:0]  io_argOuts_0_port_bits, // @[:@29434.4]
  input  [63:0]  io_argOuts_0_echo // @[:@29434.4]
);
  wire  SingleCounter_clock; // @[Main.scala 35:32:@29597.4]
  wire  SingleCounter_reset; // @[Main.scala 35:32:@29597.4]
  wire  SingleCounter_io_input_reset; // @[Main.scala 35:32:@29597.4]
  wire  SingleCounter_io_output_done; // @[Main.scala 35:32:@29597.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@29615.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@29615.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@29615.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@29615.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@29615.4]
  wire  SRFF_clock; // @[Main.scala 39:28:@29624.4]
  wire  SRFF_reset; // @[Main.scala 39:28:@29624.4]
  wire  SRFF_io_input_set; // @[Main.scala 39:28:@29624.4]
  wire  SRFF_io_input_reset; // @[Main.scala 39:28:@29624.4]
  wire  SRFF_io_input_asyn_reset; // @[Main.scala 39:28:@29624.4]
  wire  SRFF_io_output; // @[Main.scala 39:28:@29624.4]
  wire  RootController_sm_clock; // @[sm_RootController.scala 32:18:@29662.4]
  wire  RootController_sm_reset; // @[sm_RootController.scala 32:18:@29662.4]
  wire  RootController_sm_io_enable; // @[sm_RootController.scala 32:18:@29662.4]
  wire  RootController_sm_io_done; // @[sm_RootController.scala 32:18:@29662.4]
  wire  RootController_sm_io_rst; // @[sm_RootController.scala 32:18:@29662.4]
  wire  RootController_sm_io_ctrDone; // @[sm_RootController.scala 32:18:@29662.4]
  wire  RootController_sm_io_ctrInc; // @[sm_RootController.scala 32:18:@29662.4]
  wire  RootController_sm_io_doneIn_0; // @[sm_RootController.scala 32:18:@29662.4]
  wire  RootController_sm_io_enableOut_0; // @[sm_RootController.scala 32:18:@29662.4]
  wire  RootController_sm_io_childAck_0; // @[sm_RootController.scala 32:18:@29662.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@29694.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@29694.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@29694.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@29694.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@29694.4]
  wire  RootController_kernelRootController_concrete1_clock; // @[sm_RootController.scala 73:24:@29753.4]
  wire  RootController_kernelRootController_concrete1_reset; // @[sm_RootController.scala 73:24:@29753.4]
  wire  RootController_kernelRootController_concrete1_io_in_x276_TVALID; // @[sm_RootController.scala 73:24:@29753.4]
  wire  RootController_kernelRootController_concrete1_io_in_x276_TREADY; // @[sm_RootController.scala 73:24:@29753.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x276_TDATA; // @[sm_RootController.scala 73:24:@29753.4]
  wire  RootController_kernelRootController_concrete1_io_in_x275_TVALID; // @[sm_RootController.scala 73:24:@29753.4]
  wire  RootController_kernelRootController_concrete1_io_in_x275_TREADY; // @[sm_RootController.scala 73:24:@29753.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x275_TDATA; // @[sm_RootController.scala 73:24:@29753.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x275_TID; // @[sm_RootController.scala 73:24:@29753.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x275_TDEST; // @[sm_RootController.scala 73:24:@29753.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_RootController.scala 73:24:@29753.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0; // @[sm_RootController.scala 73:24:@29753.4]
  wire  RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[sm_RootController.scala 73:24:@29753.4]
  wire  RootController_kernelRootController_concrete1_io_rr; // @[sm_RootController.scala 73:24:@29753.4]
  wire  _T_599; // @[package.scala 96:25:@29620.4 package.scala 96:25:@29621.4]
  wire  _T_664; // @[Main.scala 41:50:@29690.4]
  wire  _T_665; // @[Main.scala 41:59:@29691.4]
  wire  _T_677; // @[package.scala 100:49:@29711.4]
  reg  _T_680; // @[package.scala 48:56:@29712.4]
  reg [31:0] _RAND_0;
  SingleCounter SingleCounter ( // @[Main.scala 35:32:@29597.4]
    .clock(SingleCounter_clock),
    .reset(SingleCounter_reset),
    .io_input_reset(SingleCounter_io_input_reset),
    .io_output_done(SingleCounter_io_output_done)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@29615.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  SRFF SRFF ( // @[Main.scala 39:28:@29624.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  RootController_sm RootController_sm ( // @[sm_RootController.scala 32:18:@29662.4]
    .clock(RootController_sm_clock),
    .reset(RootController_sm_reset),
    .io_enable(RootController_sm_io_enable),
    .io_done(RootController_sm_io_done),
    .io_rst(RootController_sm_io_rst),
    .io_ctrDone(RootController_sm_io_ctrDone),
    .io_ctrInc(RootController_sm_io_ctrInc),
    .io_doneIn_0(RootController_sm_io_doneIn_0),
    .io_enableOut_0(RootController_sm_io_enableOut_0),
    .io_childAck_0(RootController_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@29694.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RootController_kernelRootController_concrete1 RootController_kernelRootController_concrete1 ( // @[sm_RootController.scala 73:24:@29753.4]
    .clock(RootController_kernelRootController_concrete1_clock),
    .reset(RootController_kernelRootController_concrete1_reset),
    .io_in_x276_TVALID(RootController_kernelRootController_concrete1_io_in_x276_TVALID),
    .io_in_x276_TREADY(RootController_kernelRootController_concrete1_io_in_x276_TREADY),
    .io_in_x276_TDATA(RootController_kernelRootController_concrete1_io_in_x276_TDATA),
    .io_in_x275_TVALID(RootController_kernelRootController_concrete1_io_in_x275_TVALID),
    .io_in_x275_TREADY(RootController_kernelRootController_concrete1_io_in_x275_TREADY),
    .io_in_x275_TDATA(RootController_kernelRootController_concrete1_io_in_x275_TDATA),
    .io_in_x275_TID(RootController_kernelRootController_concrete1_io_in_x275_TID),
    .io_in_x275_TDEST(RootController_kernelRootController_concrete1_io_in_x275_TDEST),
    .io_sigsIn_smEnableOuts_0(RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(RootController_kernelRootController_concrete1_io_rr)
  );
  assign _T_599 = RetimeWrapper_io_out; // @[package.scala 96:25:@29620.4 package.scala 96:25:@29621.4]
  assign _T_664 = io_enable & _T_599; // @[Main.scala 41:50:@29690.4]
  assign _T_665 = ~ SRFF_io_output; // @[Main.scala 41:59:@29691.4]
  assign _T_677 = RootController_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@29711.4]
  assign io_done = SRFF_io_output; // @[Main.scala 48:23:@29710.4]
  assign io_memStreams_loads_0_cmd_valid = 1'h0;
  assign io_memStreams_loads_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_loads_0_cmd_bits_size = 32'h0;
  assign io_memStreams_loads_0_data_ready = 1'h0;
  assign io_memStreams_stores_0_cmd_valid = 1'h0;
  assign io_memStreams_stores_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_stores_0_cmd_bits_size = 32'h0;
  assign io_memStreams_stores_0_data_valid = 1'h0;
  assign io_memStreams_stores_0_data_bits_wdata_0 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_1 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_2 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_3 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_4 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_5 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_6 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_7 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_8 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_9 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_10 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_11 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_12 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_13 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_14 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_15 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wstrb = 16'h0;
  assign io_memStreams_stores_0_wresp_ready = 1'h0;
  assign io_memStreams_gathers_0_cmd_valid = 1'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_0 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_1 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_2 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_3 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_4 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_5 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_6 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_7 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_8 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_9 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_10 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_11 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_12 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_13 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_14 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_15 = 64'h0;
  assign io_memStreams_gathers_0_data_ready = 1'h0;
  assign io_memStreams_scatters_0_cmd_valid = 1'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_0 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_1 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_2 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_3 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_4 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_5 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_6 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_7 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_8 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_9 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_10 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_11 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_12 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_13 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_14 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_15 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_0 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_1 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_2 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_3 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_4 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_5 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_6 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_7 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_8 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_9 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_10 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_11 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_12 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_13 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_14 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_15 = 32'h0;
  assign io_memStreams_scatters_0_wresp_ready = 1'h0;
  assign io_axiStreamsIn_0_TREADY = RootController_kernelRootController_concrete1_io_in_x275_TREADY; // @[sm_RootController.scala 49:23:@29817.4]
  assign io_axiStreamsOut_0_TVALID = RootController_kernelRootController_concrete1_io_in_x276_TVALID; // @[sm_RootController.scala 48:23:@29809.4]
  assign io_axiStreamsOut_0_TDATA = RootController_kernelRootController_concrete1_io_in_x276_TDATA; // @[sm_RootController.scala 48:23:@29807.4]
  assign io_axiStreamsOut_0_TSTRB = 32'hffffffff; // @[sm_RootController.scala 48:23:@29806.4]
  assign io_axiStreamsOut_0_TKEEP = 32'hffffffff; // @[sm_RootController.scala 48:23:@29805.4]
  assign io_axiStreamsOut_0_TLAST = 1'h0; // @[sm_RootController.scala 48:23:@29804.4]
  assign io_axiStreamsOut_0_TID = 8'h0; // @[sm_RootController.scala 48:23:@29803.4]
  assign io_axiStreamsOut_0_TDEST = 8'h0; // @[sm_RootController.scala 48:23:@29802.4]
  assign io_axiStreamsOut_0_TUSER = 32'h4; // @[sm_RootController.scala 48:23:@29801.4]
  assign io_heap_0_req_valid = 1'h0;
  assign io_heap_0_req_bits_allocDealloc = 1'h0;
  assign io_heap_0_req_bits_sizeAddr = 64'h0;
  assign io_argOuts_0_port_valid = 1'h0;
  assign io_argOuts_0_port_bits = 64'h0;
  assign SingleCounter_clock = clock; // @[:@29598.4]
  assign SingleCounter_reset = reset; // @[:@29599.4]
  assign SingleCounter_io_input_reset = reset; // @[Main.scala 36:79:@29613.4]
  assign RetimeWrapper_clock = clock; // @[:@29616.4]
  assign RetimeWrapper_reset = reset; // @[:@29617.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@29619.4]
  assign RetimeWrapper_io_in = SingleCounter_io_output_done; // @[package.scala 94:16:@29618.4]
  assign SRFF_clock = clock; // @[:@29625.4]
  assign SRFF_reset = reset; // @[:@29626.4]
  assign SRFF_io_input_set = RootController_sm_io_done; // @[Main.scala 57:29:@29845.4]
  assign SRFF_io_input_reset = RetimeWrapper_1_io_out; // @[Main.scala 46:31:@29708.4]
  assign SRFF_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[Main.scala 47:36:@29709.4]
  assign RootController_sm_clock = clock; // @[:@29663.4]
  assign RootController_sm_reset = reset; // @[:@29664.4]
  assign RootController_sm_io_enable = _T_664 & _T_665; // @[Main.scala 45:33:@29707.4 SpatialBlocks.scala 112:18:@29741.4]
  assign RootController_sm_io_rst = RetimeWrapper_1_io_out; // @[SpatialBlocks.scala 106:15:@29735.4]
  assign RootController_sm_io_ctrDone = RootController_sm_io_ctrInc & _T_680; // @[Main.scala 49:34:@29715.4]
  assign RootController_sm_io_doneIn_0 = RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 102:67:@29732.4]
  assign RetimeWrapper_1_clock = clock; // @[:@29695.4]
  assign RetimeWrapper_1_reset = reset; // @[:@29696.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@29698.4]
  assign RetimeWrapper_1_io_in = reset | io_reset; // @[package.scala 94:16:@29697.4]
  assign RootController_kernelRootController_concrete1_clock = clock; // @[:@29754.4]
  assign RootController_kernelRootController_concrete1_reset = reset; // @[:@29755.4]
  assign RootController_kernelRootController_concrete1_io_in_x276_TREADY = io_axiStreamsOut_0_TREADY; // @[sm_RootController.scala 48:23:@29808.4]
  assign RootController_kernelRootController_concrete1_io_in_x275_TVALID = io_axiStreamsIn_0_TVALID; // @[sm_RootController.scala 49:23:@29818.4]
  assign RootController_kernelRootController_concrete1_io_in_x275_TDATA = io_axiStreamsIn_0_TDATA; // @[sm_RootController.scala 49:23:@29816.4]
  assign RootController_kernelRootController_concrete1_io_in_x275_TID = io_axiStreamsIn_0_TID; // @[sm_RootController.scala 49:23:@29812.4]
  assign RootController_kernelRootController_concrete1_io_in_x275_TDEST = io_axiStreamsIn_0_TDEST; // @[sm_RootController.scala 49:23:@29811.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0 = RootController_sm_io_enableOut_0; // @[sm_RootController.scala 77:22:@29827.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0 = RootController_sm_io_childAck_0; // @[sm_RootController.scala 77:22:@29825.4]
  assign RootController_kernelRootController_concrete1_io_rr = RetimeWrapper_io_out; // @[sm_RootController.scala 76:18:@29819.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_680 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_680 <= 1'h0;
    end else begin
      _T_680 <= _T_677;
    end
  end
endmodule
module SpatialIP( // @[:@29847.2]
  input         clock, // @[:@29848.4]
  input         reset, // @[:@29849.4]
  input  [31:0] io_raddr, // @[:@29850.4]
  input         io_wen, // @[:@29850.4]
  input  [31:0] io_waddr, // @[:@29850.4]
  input  [63:0] io_wdata, // @[:@29850.4]
  output [63:0] io_rdata // @[:@29850.4]
);
  wire  accel_clock; // @[Instantiator.scala 53:44:@29852.4]
  wire  accel_reset; // @[Instantiator.scala 53:44:@29852.4]
  wire  accel_io_enable; // @[Instantiator.scala 53:44:@29852.4]
  wire  accel_io_done; // @[Instantiator.scala 53:44:@29852.4]
  wire  accel_io_reset; // @[Instantiator.scala 53:44:@29852.4]
  wire  accel_io_memStreams_loads_0_cmd_ready; // @[Instantiator.scala 53:44:@29852.4]
  wire  accel_io_memStreams_loads_0_cmd_valid; // @[Instantiator.scala 53:44:@29852.4]
  wire [63:0] accel_io_memStreams_loads_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_loads_0_cmd_bits_size; // @[Instantiator.scala 53:44:@29852.4]
  wire  accel_io_memStreams_loads_0_data_ready; // @[Instantiator.scala 53:44:@29852.4]
  wire  accel_io_memStreams_loads_0_data_valid; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_0; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_1; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_2; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_3; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_4; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_5; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_6; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_7; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_8; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_9; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_10; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_11; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_12; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_13; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_14; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_15; // @[Instantiator.scala 53:44:@29852.4]
  wire  accel_io_memStreams_stores_0_cmd_ready; // @[Instantiator.scala 53:44:@29852.4]
  wire  accel_io_memStreams_stores_0_cmd_valid; // @[Instantiator.scala 53:44:@29852.4]
  wire [63:0] accel_io_memStreams_stores_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_stores_0_cmd_bits_size; // @[Instantiator.scala 53:44:@29852.4]
  wire  accel_io_memStreams_stores_0_data_ready; // @[Instantiator.scala 53:44:@29852.4]
  wire  accel_io_memStreams_stores_0_data_valid; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_1; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_2; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_3; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_4; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_5; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_6; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_7; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_8; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_9; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_10; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_11; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_12; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_13; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_14; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_15; // @[Instantiator.scala 53:44:@29852.4]
  wire [15:0] accel_io_memStreams_stores_0_data_bits_wstrb; // @[Instantiator.scala 53:44:@29852.4]
  wire  accel_io_memStreams_stores_0_wresp_ready; // @[Instantiator.scala 53:44:@29852.4]
  wire  accel_io_memStreams_stores_0_wresp_valid; // @[Instantiator.scala 53:44:@29852.4]
  wire  accel_io_memStreams_stores_0_wresp_bits; // @[Instantiator.scala 53:44:@29852.4]
  wire  accel_io_memStreams_gathers_0_cmd_ready; // @[Instantiator.scala 53:44:@29852.4]
  wire  accel_io_memStreams_gathers_0_cmd_valid; // @[Instantiator.scala 53:44:@29852.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_0; // @[Instantiator.scala 53:44:@29852.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_1; // @[Instantiator.scala 53:44:@29852.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_2; // @[Instantiator.scala 53:44:@29852.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_3; // @[Instantiator.scala 53:44:@29852.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_4; // @[Instantiator.scala 53:44:@29852.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_5; // @[Instantiator.scala 53:44:@29852.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_6; // @[Instantiator.scala 53:44:@29852.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_7; // @[Instantiator.scala 53:44:@29852.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_8; // @[Instantiator.scala 53:44:@29852.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_9; // @[Instantiator.scala 53:44:@29852.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_10; // @[Instantiator.scala 53:44:@29852.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_11; // @[Instantiator.scala 53:44:@29852.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_12; // @[Instantiator.scala 53:44:@29852.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_13; // @[Instantiator.scala 53:44:@29852.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_14; // @[Instantiator.scala 53:44:@29852.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_15; // @[Instantiator.scala 53:44:@29852.4]
  wire  accel_io_memStreams_gathers_0_data_ready; // @[Instantiator.scala 53:44:@29852.4]
  wire  accel_io_memStreams_gathers_0_data_valid; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_0; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_1; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_2; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_3; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_4; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_5; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_6; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_7; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_8; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_9; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_10; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_11; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_12; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_13; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_14; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_15; // @[Instantiator.scala 53:44:@29852.4]
  wire  accel_io_memStreams_scatters_0_cmd_ready; // @[Instantiator.scala 53:44:@29852.4]
  wire  accel_io_memStreams_scatters_0_cmd_valid; // @[Instantiator.scala 53:44:@29852.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0; // @[Instantiator.scala 53:44:@29852.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1; // @[Instantiator.scala 53:44:@29852.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2; // @[Instantiator.scala 53:44:@29852.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3; // @[Instantiator.scala 53:44:@29852.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4; // @[Instantiator.scala 53:44:@29852.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5; // @[Instantiator.scala 53:44:@29852.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6; // @[Instantiator.scala 53:44:@29852.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7; // @[Instantiator.scala 53:44:@29852.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8; // @[Instantiator.scala 53:44:@29852.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9; // @[Instantiator.scala 53:44:@29852.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10; // @[Instantiator.scala 53:44:@29852.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11; // @[Instantiator.scala 53:44:@29852.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12; // @[Instantiator.scala 53:44:@29852.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13; // @[Instantiator.scala 53:44:@29852.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14; // @[Instantiator.scala 53:44:@29852.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_0; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_1; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_2; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_3; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_4; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_5; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_6; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_7; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_8; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_9; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_10; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_11; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_12; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_13; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_14; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_15; // @[Instantiator.scala 53:44:@29852.4]
  wire  accel_io_memStreams_scatters_0_wresp_ready; // @[Instantiator.scala 53:44:@29852.4]
  wire  accel_io_memStreams_scatters_0_wresp_valid; // @[Instantiator.scala 53:44:@29852.4]
  wire  accel_io_memStreams_scatters_0_wresp_bits; // @[Instantiator.scala 53:44:@29852.4]
  wire  accel_io_axiStreamsIn_0_TVALID; // @[Instantiator.scala 53:44:@29852.4]
  wire  accel_io_axiStreamsIn_0_TREADY; // @[Instantiator.scala 53:44:@29852.4]
  wire [255:0] accel_io_axiStreamsIn_0_TDATA; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_axiStreamsIn_0_TSTRB; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_axiStreamsIn_0_TKEEP; // @[Instantiator.scala 53:44:@29852.4]
  wire  accel_io_axiStreamsIn_0_TLAST; // @[Instantiator.scala 53:44:@29852.4]
  wire [7:0] accel_io_axiStreamsIn_0_TID; // @[Instantiator.scala 53:44:@29852.4]
  wire [7:0] accel_io_axiStreamsIn_0_TDEST; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_axiStreamsIn_0_TUSER; // @[Instantiator.scala 53:44:@29852.4]
  wire  accel_io_axiStreamsOut_0_TVALID; // @[Instantiator.scala 53:44:@29852.4]
  wire  accel_io_axiStreamsOut_0_TREADY; // @[Instantiator.scala 53:44:@29852.4]
  wire [255:0] accel_io_axiStreamsOut_0_TDATA; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_axiStreamsOut_0_TSTRB; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_axiStreamsOut_0_TKEEP; // @[Instantiator.scala 53:44:@29852.4]
  wire  accel_io_axiStreamsOut_0_TLAST; // @[Instantiator.scala 53:44:@29852.4]
  wire [7:0] accel_io_axiStreamsOut_0_TID; // @[Instantiator.scala 53:44:@29852.4]
  wire [7:0] accel_io_axiStreamsOut_0_TDEST; // @[Instantiator.scala 53:44:@29852.4]
  wire [31:0] accel_io_axiStreamsOut_0_TUSER; // @[Instantiator.scala 53:44:@29852.4]
  wire  accel_io_heap_0_req_valid; // @[Instantiator.scala 53:44:@29852.4]
  wire  accel_io_heap_0_req_bits_allocDealloc; // @[Instantiator.scala 53:44:@29852.4]
  wire [63:0] accel_io_heap_0_req_bits_sizeAddr; // @[Instantiator.scala 53:44:@29852.4]
  wire  accel_io_heap_0_resp_valid; // @[Instantiator.scala 53:44:@29852.4]
  wire  accel_io_heap_0_resp_bits_allocDealloc; // @[Instantiator.scala 53:44:@29852.4]
  wire [63:0] accel_io_heap_0_resp_bits_sizeAddr; // @[Instantiator.scala 53:44:@29852.4]
  wire [63:0] accel_io_argIns_0; // @[Instantiator.scala 53:44:@29852.4]
  wire [63:0] accel_io_argIns_1; // @[Instantiator.scala 53:44:@29852.4]
  wire  accel_io_argOuts_0_port_ready; // @[Instantiator.scala 53:44:@29852.4]
  wire  accel_io_argOuts_0_port_valid; // @[Instantiator.scala 53:44:@29852.4]
  wire [63:0] accel_io_argOuts_0_port_bits; // @[Instantiator.scala 53:44:@29852.4]
  wire [63:0] accel_io_argOuts_0_echo; // @[Instantiator.scala 53:44:@29852.4]
  AccelUnit accel ( // @[Instantiator.scala 53:44:@29852.4]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_enable(accel_io_enable),
    .io_done(accel_io_done),
    .io_reset(accel_io_reset),
    .io_memStreams_loads_0_cmd_ready(accel_io_memStreams_loads_0_cmd_ready),
    .io_memStreams_loads_0_cmd_valid(accel_io_memStreams_loads_0_cmd_valid),
    .io_memStreams_loads_0_cmd_bits_addr(accel_io_memStreams_loads_0_cmd_bits_addr),
    .io_memStreams_loads_0_cmd_bits_size(accel_io_memStreams_loads_0_cmd_bits_size),
    .io_memStreams_loads_0_data_ready(accel_io_memStreams_loads_0_data_ready),
    .io_memStreams_loads_0_data_valid(accel_io_memStreams_loads_0_data_valid),
    .io_memStreams_loads_0_data_bits_rdata_0(accel_io_memStreams_loads_0_data_bits_rdata_0),
    .io_memStreams_loads_0_data_bits_rdata_1(accel_io_memStreams_loads_0_data_bits_rdata_1),
    .io_memStreams_loads_0_data_bits_rdata_2(accel_io_memStreams_loads_0_data_bits_rdata_2),
    .io_memStreams_loads_0_data_bits_rdata_3(accel_io_memStreams_loads_0_data_bits_rdata_3),
    .io_memStreams_loads_0_data_bits_rdata_4(accel_io_memStreams_loads_0_data_bits_rdata_4),
    .io_memStreams_loads_0_data_bits_rdata_5(accel_io_memStreams_loads_0_data_bits_rdata_5),
    .io_memStreams_loads_0_data_bits_rdata_6(accel_io_memStreams_loads_0_data_bits_rdata_6),
    .io_memStreams_loads_0_data_bits_rdata_7(accel_io_memStreams_loads_0_data_bits_rdata_7),
    .io_memStreams_loads_0_data_bits_rdata_8(accel_io_memStreams_loads_0_data_bits_rdata_8),
    .io_memStreams_loads_0_data_bits_rdata_9(accel_io_memStreams_loads_0_data_bits_rdata_9),
    .io_memStreams_loads_0_data_bits_rdata_10(accel_io_memStreams_loads_0_data_bits_rdata_10),
    .io_memStreams_loads_0_data_bits_rdata_11(accel_io_memStreams_loads_0_data_bits_rdata_11),
    .io_memStreams_loads_0_data_bits_rdata_12(accel_io_memStreams_loads_0_data_bits_rdata_12),
    .io_memStreams_loads_0_data_bits_rdata_13(accel_io_memStreams_loads_0_data_bits_rdata_13),
    .io_memStreams_loads_0_data_bits_rdata_14(accel_io_memStreams_loads_0_data_bits_rdata_14),
    .io_memStreams_loads_0_data_bits_rdata_15(accel_io_memStreams_loads_0_data_bits_rdata_15),
    .io_memStreams_stores_0_cmd_ready(accel_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(accel_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(accel_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(accel_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(accel_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(accel_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(accel_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wdata_1(accel_io_memStreams_stores_0_data_bits_wdata_1),
    .io_memStreams_stores_0_data_bits_wdata_2(accel_io_memStreams_stores_0_data_bits_wdata_2),
    .io_memStreams_stores_0_data_bits_wdata_3(accel_io_memStreams_stores_0_data_bits_wdata_3),
    .io_memStreams_stores_0_data_bits_wdata_4(accel_io_memStreams_stores_0_data_bits_wdata_4),
    .io_memStreams_stores_0_data_bits_wdata_5(accel_io_memStreams_stores_0_data_bits_wdata_5),
    .io_memStreams_stores_0_data_bits_wdata_6(accel_io_memStreams_stores_0_data_bits_wdata_6),
    .io_memStreams_stores_0_data_bits_wdata_7(accel_io_memStreams_stores_0_data_bits_wdata_7),
    .io_memStreams_stores_0_data_bits_wdata_8(accel_io_memStreams_stores_0_data_bits_wdata_8),
    .io_memStreams_stores_0_data_bits_wdata_9(accel_io_memStreams_stores_0_data_bits_wdata_9),
    .io_memStreams_stores_0_data_bits_wdata_10(accel_io_memStreams_stores_0_data_bits_wdata_10),
    .io_memStreams_stores_0_data_bits_wdata_11(accel_io_memStreams_stores_0_data_bits_wdata_11),
    .io_memStreams_stores_0_data_bits_wdata_12(accel_io_memStreams_stores_0_data_bits_wdata_12),
    .io_memStreams_stores_0_data_bits_wdata_13(accel_io_memStreams_stores_0_data_bits_wdata_13),
    .io_memStreams_stores_0_data_bits_wdata_14(accel_io_memStreams_stores_0_data_bits_wdata_14),
    .io_memStreams_stores_0_data_bits_wdata_15(accel_io_memStreams_stores_0_data_bits_wdata_15),
    .io_memStreams_stores_0_data_bits_wstrb(accel_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(accel_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(accel_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(accel_io_memStreams_stores_0_wresp_bits),
    .io_memStreams_gathers_0_cmd_ready(accel_io_memStreams_gathers_0_cmd_ready),
    .io_memStreams_gathers_0_cmd_valid(accel_io_memStreams_gathers_0_cmd_valid),
    .io_memStreams_gathers_0_cmd_bits_addr_0(accel_io_memStreams_gathers_0_cmd_bits_addr_0),
    .io_memStreams_gathers_0_cmd_bits_addr_1(accel_io_memStreams_gathers_0_cmd_bits_addr_1),
    .io_memStreams_gathers_0_cmd_bits_addr_2(accel_io_memStreams_gathers_0_cmd_bits_addr_2),
    .io_memStreams_gathers_0_cmd_bits_addr_3(accel_io_memStreams_gathers_0_cmd_bits_addr_3),
    .io_memStreams_gathers_0_cmd_bits_addr_4(accel_io_memStreams_gathers_0_cmd_bits_addr_4),
    .io_memStreams_gathers_0_cmd_bits_addr_5(accel_io_memStreams_gathers_0_cmd_bits_addr_5),
    .io_memStreams_gathers_0_cmd_bits_addr_6(accel_io_memStreams_gathers_0_cmd_bits_addr_6),
    .io_memStreams_gathers_0_cmd_bits_addr_7(accel_io_memStreams_gathers_0_cmd_bits_addr_7),
    .io_memStreams_gathers_0_cmd_bits_addr_8(accel_io_memStreams_gathers_0_cmd_bits_addr_8),
    .io_memStreams_gathers_0_cmd_bits_addr_9(accel_io_memStreams_gathers_0_cmd_bits_addr_9),
    .io_memStreams_gathers_0_cmd_bits_addr_10(accel_io_memStreams_gathers_0_cmd_bits_addr_10),
    .io_memStreams_gathers_0_cmd_bits_addr_11(accel_io_memStreams_gathers_0_cmd_bits_addr_11),
    .io_memStreams_gathers_0_cmd_bits_addr_12(accel_io_memStreams_gathers_0_cmd_bits_addr_12),
    .io_memStreams_gathers_0_cmd_bits_addr_13(accel_io_memStreams_gathers_0_cmd_bits_addr_13),
    .io_memStreams_gathers_0_cmd_bits_addr_14(accel_io_memStreams_gathers_0_cmd_bits_addr_14),
    .io_memStreams_gathers_0_cmd_bits_addr_15(accel_io_memStreams_gathers_0_cmd_bits_addr_15),
    .io_memStreams_gathers_0_data_ready(accel_io_memStreams_gathers_0_data_ready),
    .io_memStreams_gathers_0_data_valid(accel_io_memStreams_gathers_0_data_valid),
    .io_memStreams_gathers_0_data_bits_0(accel_io_memStreams_gathers_0_data_bits_0),
    .io_memStreams_gathers_0_data_bits_1(accel_io_memStreams_gathers_0_data_bits_1),
    .io_memStreams_gathers_0_data_bits_2(accel_io_memStreams_gathers_0_data_bits_2),
    .io_memStreams_gathers_0_data_bits_3(accel_io_memStreams_gathers_0_data_bits_3),
    .io_memStreams_gathers_0_data_bits_4(accel_io_memStreams_gathers_0_data_bits_4),
    .io_memStreams_gathers_0_data_bits_5(accel_io_memStreams_gathers_0_data_bits_5),
    .io_memStreams_gathers_0_data_bits_6(accel_io_memStreams_gathers_0_data_bits_6),
    .io_memStreams_gathers_0_data_bits_7(accel_io_memStreams_gathers_0_data_bits_7),
    .io_memStreams_gathers_0_data_bits_8(accel_io_memStreams_gathers_0_data_bits_8),
    .io_memStreams_gathers_0_data_bits_9(accel_io_memStreams_gathers_0_data_bits_9),
    .io_memStreams_gathers_0_data_bits_10(accel_io_memStreams_gathers_0_data_bits_10),
    .io_memStreams_gathers_0_data_bits_11(accel_io_memStreams_gathers_0_data_bits_11),
    .io_memStreams_gathers_0_data_bits_12(accel_io_memStreams_gathers_0_data_bits_12),
    .io_memStreams_gathers_0_data_bits_13(accel_io_memStreams_gathers_0_data_bits_13),
    .io_memStreams_gathers_0_data_bits_14(accel_io_memStreams_gathers_0_data_bits_14),
    .io_memStreams_gathers_0_data_bits_15(accel_io_memStreams_gathers_0_data_bits_15),
    .io_memStreams_scatters_0_cmd_ready(accel_io_memStreams_scatters_0_cmd_ready),
    .io_memStreams_scatters_0_cmd_valid(accel_io_memStreams_scatters_0_cmd_valid),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_0(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_1(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_2(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_3(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_4(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_5(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_6(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_7(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_8(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_9(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_10(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_11(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_12(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_13(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_14(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_15(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15),
    .io_memStreams_scatters_0_cmd_bits_wdata_0(accel_io_memStreams_scatters_0_cmd_bits_wdata_0),
    .io_memStreams_scatters_0_cmd_bits_wdata_1(accel_io_memStreams_scatters_0_cmd_bits_wdata_1),
    .io_memStreams_scatters_0_cmd_bits_wdata_2(accel_io_memStreams_scatters_0_cmd_bits_wdata_2),
    .io_memStreams_scatters_0_cmd_bits_wdata_3(accel_io_memStreams_scatters_0_cmd_bits_wdata_3),
    .io_memStreams_scatters_0_cmd_bits_wdata_4(accel_io_memStreams_scatters_0_cmd_bits_wdata_4),
    .io_memStreams_scatters_0_cmd_bits_wdata_5(accel_io_memStreams_scatters_0_cmd_bits_wdata_5),
    .io_memStreams_scatters_0_cmd_bits_wdata_6(accel_io_memStreams_scatters_0_cmd_bits_wdata_6),
    .io_memStreams_scatters_0_cmd_bits_wdata_7(accel_io_memStreams_scatters_0_cmd_bits_wdata_7),
    .io_memStreams_scatters_0_cmd_bits_wdata_8(accel_io_memStreams_scatters_0_cmd_bits_wdata_8),
    .io_memStreams_scatters_0_cmd_bits_wdata_9(accel_io_memStreams_scatters_0_cmd_bits_wdata_9),
    .io_memStreams_scatters_0_cmd_bits_wdata_10(accel_io_memStreams_scatters_0_cmd_bits_wdata_10),
    .io_memStreams_scatters_0_cmd_bits_wdata_11(accel_io_memStreams_scatters_0_cmd_bits_wdata_11),
    .io_memStreams_scatters_0_cmd_bits_wdata_12(accel_io_memStreams_scatters_0_cmd_bits_wdata_12),
    .io_memStreams_scatters_0_cmd_bits_wdata_13(accel_io_memStreams_scatters_0_cmd_bits_wdata_13),
    .io_memStreams_scatters_0_cmd_bits_wdata_14(accel_io_memStreams_scatters_0_cmd_bits_wdata_14),
    .io_memStreams_scatters_0_cmd_bits_wdata_15(accel_io_memStreams_scatters_0_cmd_bits_wdata_15),
    .io_memStreams_scatters_0_wresp_ready(accel_io_memStreams_scatters_0_wresp_ready),
    .io_memStreams_scatters_0_wresp_valid(accel_io_memStreams_scatters_0_wresp_valid),
    .io_memStreams_scatters_0_wresp_bits(accel_io_memStreams_scatters_0_wresp_bits),
    .io_axiStreamsIn_0_TVALID(accel_io_axiStreamsIn_0_TVALID),
    .io_axiStreamsIn_0_TREADY(accel_io_axiStreamsIn_0_TREADY),
    .io_axiStreamsIn_0_TDATA(accel_io_axiStreamsIn_0_TDATA),
    .io_axiStreamsIn_0_TSTRB(accel_io_axiStreamsIn_0_TSTRB),
    .io_axiStreamsIn_0_TKEEP(accel_io_axiStreamsIn_0_TKEEP),
    .io_axiStreamsIn_0_TLAST(accel_io_axiStreamsIn_0_TLAST),
    .io_axiStreamsIn_0_TID(accel_io_axiStreamsIn_0_TID),
    .io_axiStreamsIn_0_TDEST(accel_io_axiStreamsIn_0_TDEST),
    .io_axiStreamsIn_0_TUSER(accel_io_axiStreamsIn_0_TUSER),
    .io_axiStreamsOut_0_TVALID(accel_io_axiStreamsOut_0_TVALID),
    .io_axiStreamsOut_0_TREADY(accel_io_axiStreamsOut_0_TREADY),
    .io_axiStreamsOut_0_TDATA(accel_io_axiStreamsOut_0_TDATA),
    .io_axiStreamsOut_0_TSTRB(accel_io_axiStreamsOut_0_TSTRB),
    .io_axiStreamsOut_0_TKEEP(accel_io_axiStreamsOut_0_TKEEP),
    .io_axiStreamsOut_0_TLAST(accel_io_axiStreamsOut_0_TLAST),
    .io_axiStreamsOut_0_TID(accel_io_axiStreamsOut_0_TID),
    .io_axiStreamsOut_0_TDEST(accel_io_axiStreamsOut_0_TDEST),
    .io_axiStreamsOut_0_TUSER(accel_io_axiStreamsOut_0_TUSER),
    .io_heap_0_req_valid(accel_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(accel_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(accel_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(accel_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(accel_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(accel_io_heap_0_resp_bits_sizeAddr),
    .io_argIns_0(accel_io_argIns_0),
    .io_argIns_1(accel_io_argIns_1),
    .io_argOuts_0_port_ready(accel_io_argOuts_0_port_ready),
    .io_argOuts_0_port_valid(accel_io_argOuts_0_port_valid),
    .io_argOuts_0_port_bits(accel_io_argOuts_0_port_bits),
    .io_argOuts_0_echo(accel_io_argOuts_0_echo)
  );
  assign io_rdata = 64'h0;
  assign accel_clock = clock; // @[:@29853.4]
  assign accel_reset = reset; // @[:@29854.4]
  assign accel_io_enable = 1'h0;
  assign accel_io_reset = 1'h0;
  assign accel_io_memStreams_loads_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_loads_0_data_valid = 1'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_0 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_1 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_2 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_3 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_4 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_5 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_6 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_7 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_8 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_9 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_10 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_11 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_12 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_13 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_14 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_15 = 32'h0;
  assign accel_io_memStreams_stores_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_stores_0_data_ready = 1'h0;
  assign accel_io_memStreams_stores_0_wresp_valid = 1'h0;
  assign accel_io_memStreams_stores_0_wresp_bits = 1'h0;
  assign accel_io_memStreams_gathers_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_gathers_0_data_valid = 1'h0;
  assign accel_io_memStreams_gathers_0_data_bits_0 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_1 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_2 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_3 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_4 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_5 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_6 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_7 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_8 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_9 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_10 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_11 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_12 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_13 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_14 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_15 = 32'h0;
  assign accel_io_memStreams_scatters_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_scatters_0_wresp_valid = 1'h0;
  assign accel_io_memStreams_scatters_0_wresp_bits = 1'h0;
  assign accel_io_axiStreamsIn_0_TVALID = 1'h0;
  assign accel_io_axiStreamsIn_0_TDATA = 256'h0;
  assign accel_io_axiStreamsIn_0_TSTRB = 32'h0;
  assign accel_io_axiStreamsIn_0_TKEEP = 32'h0;
  assign accel_io_axiStreamsIn_0_TLAST = 1'h0;
  assign accel_io_axiStreamsIn_0_TID = 8'h0;
  assign accel_io_axiStreamsIn_0_TDEST = 8'h0;
  assign accel_io_axiStreamsIn_0_TUSER = 32'h0;
  assign accel_io_axiStreamsOut_0_TREADY = 1'h0;
  assign accel_io_heap_0_resp_valid = 1'h0;
  assign accel_io_heap_0_resp_bits_allocDealloc = 1'h0;
  assign accel_io_heap_0_resp_bits_sizeAddr = 64'h0;
  assign accel_io_argIns_0 = 64'h0;
  assign accel_io_argIns_1 = 64'h0;
  assign accel_io_argOuts_0_port_ready = 1'h0;
  assign accel_io_argOuts_0_echo = 64'h0;
endmodule
