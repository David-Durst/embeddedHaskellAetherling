module coreir_ugt #(parameter width = 1) (input [width-1:0] in0/*verilator public*/, input [width-1:0] in1/*verilator public*/, output out/*verilator public*/);
  assign out = in0 > in1;
endmodule

module coreir_reg #(parameter width = 1, parameter clk_posedge = 1, parameter init = 1) (input clk/*verilator public*/, input [width-1:0] in/*verilator public*/, output [width-1:0] out/*verilator public*/);
  reg [width-1:0] outReg/*verilator public*/=init;
  wire real_clk;
  assign real_clk = clk_posedge ? clk : ~clk;
  always @(posedge real_clk) begin
    outReg <= in;
  end
  assign out = outReg;
endmodule

module coreir_neg #(parameter width = 1) (input [width-1:0] in/*verilator public*/, output [width-1:0] out/*verilator public*/);
  assign out = -in;
endmodule

module coreir_mux #(parameter width = 1) (input [width-1:0] in0/*verilator public*/, input [width-1:0] in1/*verilator public*/, input sel/*verilator public*/, output [width-1:0] out/*verilator public*/);
  assign out = sel ? in1 : in0;
endmodule

module corebit_and (input in0/*verilator public*/, input in1/*verilator public*/, output out/*verilator public*/);
  assign out = in0 & in1;
endmodule

module top (input CLK/*verilator public*/, output [7:0] O_0/*verilator public*/, output [7:0] O_1/*verilator public*/, output [7:0] O_2/*verilator public*/, output [7:0] O_3/*verilator public*/, input [7:0] hi_0/*verilator public*/, input [7:0] hi_1/*verilator public*/, input [7:0] hi_2/*verilator public*/, input [7:0] hi_3/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst10$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst11$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst12$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst13$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst14$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst15$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst16$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst17$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst18$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst19$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst20$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst21$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst22$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst23$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst24$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst25$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst26$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst27$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst28$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst29$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst30$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst31$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst8$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst9$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Bitt_0init_FalseCE_FalseRESET_inst0$Register1_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst10$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst11$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst12$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst13$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst14$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst15$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst16$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst17$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst18$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst19$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst20$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst21$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst22$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst23$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst24$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst25$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst26$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst27$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst28$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst29$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst30$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst31$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst8$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst9$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Bitt_0init_FalseCE_FalseRESET_inst0$Register1_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst10$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst11$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst12$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst13$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst14$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst15$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst16$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst17$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst18$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst19$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst20$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst21$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst22$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst23$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst24$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst25$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst26$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst27$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst28$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst29$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst30$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst31$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst8$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst9$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Bitt_0init_FalseCE_FalseRESET_inst0$Register1_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst10$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst11$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst12$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst13$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst14$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst15$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst16$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst17$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst18$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst19$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst20$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst21$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst22$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst23$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst24$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst25$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst26$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst27$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst28$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst29$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst30$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst31$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst8$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst9$reg_P_inst0_out;
wire [0:0] FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Bitt_0init_FalseCE_FalseRESET_inst0$Register1_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out;
wire [7:0] NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst0$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out;
wire [7:0] NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst0$Negate8_inst0$coreir_neg_inst0_out;
wire NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst0$coreir_ugt8_inst0_out;
wire [7:0] NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst1$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out;
wire [7:0] NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst1$Negate8_inst0$coreir_neg_inst0_out;
wire NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst1$coreir_ugt8_inst0_out;
wire [7:0] NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst2$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out;
wire [7:0] NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst2$Negate8_inst0$coreir_neg_inst0_out;
wire NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst2$coreir_ugt8_inst0_out;
wire [7:0] NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst3$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out;
wire [7:0] NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst3$Negate8_inst0$coreir_neg_inst0_out;
wire NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst3$coreir_ugt8_inst0_out;
wire NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$and_inst0_out;
wire NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$and_inst1_out;
wire NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$and_inst2_out;
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(.clk(CLK), .in(hi_0[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0(.clk(CLK), .in(hi_0[1]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst10$reg_P_inst0(.clk(CLK), .in(hi_1[2]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst10$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst11$reg_P_inst0(.clk(CLK), .in(hi_1[3]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst11$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst12$reg_P_inst0(.clk(CLK), .in(hi_1[4]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst12$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst13$reg_P_inst0(.clk(CLK), .in(hi_1[5]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst13$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst14$reg_P_inst0(.clk(CLK), .in(hi_1[6]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst14$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst15$reg_P_inst0(.clk(CLK), .in(hi_1[7]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst15$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst16$reg_P_inst0(.clk(CLK), .in(hi_2[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst16$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst17$reg_P_inst0(.clk(CLK), .in(hi_2[1]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst17$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst18$reg_P_inst0(.clk(CLK), .in(hi_2[2]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst18$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst19$reg_P_inst0(.clk(CLK), .in(hi_2[3]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst19$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2$reg_P_inst0(.clk(CLK), .in(hi_0[2]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst20$reg_P_inst0(.clk(CLK), .in(hi_2[4]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst20$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst21$reg_P_inst0(.clk(CLK), .in(hi_2[5]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst21$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst22$reg_P_inst0(.clk(CLK), .in(hi_2[6]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst22$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst23$reg_P_inst0(.clk(CLK), .in(hi_2[7]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst23$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst24$reg_P_inst0(.clk(CLK), .in(hi_3[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst24$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst25$reg_P_inst0(.clk(CLK), .in(hi_3[1]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst25$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst26$reg_P_inst0(.clk(CLK), .in(hi_3[2]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst26$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst27$reg_P_inst0(.clk(CLK), .in(hi_3[3]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst27$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst28$reg_P_inst0(.clk(CLK), .in(hi_3[4]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst28$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst29$reg_P_inst0(.clk(CLK), .in(hi_3[5]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst29$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3$reg_P_inst0(.clk(CLK), .in(hi_0[3]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst30$reg_P_inst0(.clk(CLK), .in(hi_3[6]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst30$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst31$reg_P_inst0(.clk(CLK), .in(hi_3[7]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst31$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4$reg_P_inst0(.clk(CLK), .in(hi_0[4]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5$reg_P_inst0(.clk(CLK), .in(hi_0[5]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6$reg_P_inst0(.clk(CLK), .in(hi_0[6]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7$reg_P_inst0(.clk(CLK), .in(hi_0[7]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst8$reg_P_inst0(.clk(CLK), .in(hi_1[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst8$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst9$reg_P_inst0(.clk(CLK), .in(hi_1[1]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst9$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Bitt_0init_FalseCE_FalseRESET_inst0$Register1_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(.clk(CLK), .in(valid_up), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Bitt_0init_FalseCE_FalseRESET_inst0$Register1_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(.clk(CLK), .in(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst0$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0(.clk(CLK), .in(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst0$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out[1]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst10$reg_P_inst0(.clk(CLK), .in(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst1$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out[2]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst10$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst11$reg_P_inst0(.clk(CLK), .in(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst1$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out[3]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst11$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst12$reg_P_inst0(.clk(CLK), .in(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst1$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out[4]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst12$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst13$reg_P_inst0(.clk(CLK), .in(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst1$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out[5]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst13$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst14$reg_P_inst0(.clk(CLK), .in(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst1$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out[6]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst14$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst15$reg_P_inst0(.clk(CLK), .in(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst1$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out[7]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst15$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst16$reg_P_inst0(.clk(CLK), .in(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst2$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst16$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst17$reg_P_inst0(.clk(CLK), .in(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst2$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out[1]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst17$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst18$reg_P_inst0(.clk(CLK), .in(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst2$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out[2]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst18$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst19$reg_P_inst0(.clk(CLK), .in(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst2$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out[3]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst19$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2$reg_P_inst0(.clk(CLK), .in(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst0$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out[2]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst20$reg_P_inst0(.clk(CLK), .in(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst2$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out[4]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst20$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst21$reg_P_inst0(.clk(CLK), .in(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst2$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out[5]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst21$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst22$reg_P_inst0(.clk(CLK), .in(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst2$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out[6]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst22$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst23$reg_P_inst0(.clk(CLK), .in(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst2$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out[7]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst23$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst24$reg_P_inst0(.clk(CLK), .in(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst3$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst24$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst25$reg_P_inst0(.clk(CLK), .in(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst3$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out[1]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst25$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst26$reg_P_inst0(.clk(CLK), .in(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst3$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out[2]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst26$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst27$reg_P_inst0(.clk(CLK), .in(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst3$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out[3]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst27$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst28$reg_P_inst0(.clk(CLK), .in(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst3$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out[4]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst28$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst29$reg_P_inst0(.clk(CLK), .in(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst3$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out[5]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst29$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3$reg_P_inst0(.clk(CLK), .in(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst0$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out[3]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst30$reg_P_inst0(.clk(CLK), .in(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst3$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out[6]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst30$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst31$reg_P_inst0(.clk(CLK), .in(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst3$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out[7]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst31$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4$reg_P_inst0(.clk(CLK), .in(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst0$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out[4]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5$reg_P_inst0(.clk(CLK), .in(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst0$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out[5]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6$reg_P_inst0(.clk(CLK), .in(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst0$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out[6]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7$reg_P_inst0(.clk(CLK), .in(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst0$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out[7]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst8$reg_P_inst0(.clk(CLK), .in(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst1$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst8$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst9$reg_P_inst0(.clk(CLK), .in(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst1$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out[1]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst9$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Bitt_0init_FalseCE_FalseRESET_inst0$Register1_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(.clk(CLK), .in(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$and_inst2_out), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Bitt_0init_FalseCE_FalseRESET_inst0$Register1_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst10$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst10$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst10$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst11$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst11$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst11$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst12$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst12$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst12$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst13$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst13$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst13$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst14$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst14$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst14$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst15$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst15$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst15$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst16$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst16$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst16$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst17$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst17$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst17$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst18$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst18$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst18$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst19$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst19$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst19$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst20$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst20$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst20$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst21$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst21$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst21$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst22$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst22$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst22$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst23$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst23$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst23$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst24$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst24$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst24$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst25$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst25$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst25$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst26$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst26$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst26$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst27$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst27$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst27$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst28$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst28$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst28$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst29$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst29$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst29$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst30$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst30$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst30$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst31$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst31$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst31$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst8$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst8$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst8$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst9$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst9$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst9$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Bitt_0init_FalseCE_FalseRESET_inst0$Register1_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1$Register_Bitt_0init_FalseCE_FalseRESET_inst0$Register1_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Bitt_0init_FalseCE_FalseRESET_inst0$Register1_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst10$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst10$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst10$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst11$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst11$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst11$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst12$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst12$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst12$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst13$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst13$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst13$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst14$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst14$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst14$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst15$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst15$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst15$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst16$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst16$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst16$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst17$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst17$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst17$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst18$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst18$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst18$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst19$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst19$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst19$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst20$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst20$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst20$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst21$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst21$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst21$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst22$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst22$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst22$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst23$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst23$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst23$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst24$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst24$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst24$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst25$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst25$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst25$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst26$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst26$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst26$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst27$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst27$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst27$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst28$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst28$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst28$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst29$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst29$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst29$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst30$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst30$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst30$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst31$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst31$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst31$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst8$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst8$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst8$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst9$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst9$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst9$reg_P_inst0_out));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Bitt_0init_FalseCE_FalseRESET_inst0$Register1_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(.clk(CLK), .in(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2$Register_Bitt_0init_FalseCE_FalseRESET_inst0$Register1_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out[0]), .out(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Bitt_0init_FalseCE_FalseRESET_inst0$Register1_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out));
coreir_mux #(.width(8)) NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst0$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join(.in0({FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out[0]}), .in1({NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst0$Negate8_inst0$coreir_neg_inst0_out[7],NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst0$Negate8_inst0$coreir_neg_inst0_out[6],NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst0$Negate8_inst0$coreir_neg_inst0_out[5],NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst0$Negate8_inst0$coreir_neg_inst0_out[4],NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst0$Negate8_inst0$coreir_neg_inst0_out[3],NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst0$Negate8_inst0$coreir_neg_inst0_out[2],NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst0$Negate8_inst0$coreir_neg_inst0_out[1],NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst0$Negate8_inst0$coreir_neg_inst0_out[0]}), .out(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst0$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out), .sel(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst0$coreir_ugt8_inst0_out));
coreir_neg #(.width(8)) NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst0$Negate8_inst0$coreir_neg_inst0(.in({FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out[0]}), .out(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst0$Negate8_inst0$coreir_neg_inst0_out));
coreir_ugt #(.width(8)) NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst0$coreir_ugt8_inst0(.in0({FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out[0]}), .in1(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst0$Negate8_inst0$coreir_neg_inst0_out), .out(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst0$coreir_ugt8_inst0_out));
coreir_mux #(.width(8)) NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst1$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join(.in0({FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst15$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst14$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst13$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst12$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst11$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst10$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst9$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst8$reg_P_inst0_out[0]}), .in1({NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst1$Negate8_inst0$coreir_neg_inst0_out[7],NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst1$Negate8_inst0$coreir_neg_inst0_out[6],NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst1$Negate8_inst0$coreir_neg_inst0_out[5],NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst1$Negate8_inst0$coreir_neg_inst0_out[4],NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst1$Negate8_inst0$coreir_neg_inst0_out[3],NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst1$Negate8_inst0$coreir_neg_inst0_out[2],NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst1$Negate8_inst0$coreir_neg_inst0_out[1],NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst1$Negate8_inst0$coreir_neg_inst0_out[0]}), .out(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst1$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out), .sel(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst1$coreir_ugt8_inst0_out));
coreir_neg #(.width(8)) NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst1$Negate8_inst0$coreir_neg_inst0(.in({FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst15$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst14$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst13$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst12$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst11$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst10$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst9$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst8$reg_P_inst0_out[0]}), .out(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst1$Negate8_inst0$coreir_neg_inst0_out));
coreir_ugt #(.width(8)) NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst1$coreir_ugt8_inst0(.in0({FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst15$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst14$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst13$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst12$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst11$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst10$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst9$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst8$reg_P_inst0_out[0]}), .in1(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst1$Negate8_inst0$coreir_neg_inst0_out), .out(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst1$coreir_ugt8_inst0_out));
coreir_mux #(.width(8)) NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst2$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join(.in0({FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst23$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst22$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst21$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst20$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst19$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst18$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst17$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst16$reg_P_inst0_out[0]}), .in1({NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst2$Negate8_inst0$coreir_neg_inst0_out[7],NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst2$Negate8_inst0$coreir_neg_inst0_out[6],NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst2$Negate8_inst0$coreir_neg_inst0_out[5],NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst2$Negate8_inst0$coreir_neg_inst0_out[4],NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst2$Negate8_inst0$coreir_neg_inst0_out[3],NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst2$Negate8_inst0$coreir_neg_inst0_out[2],NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst2$Negate8_inst0$coreir_neg_inst0_out[1],NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst2$Negate8_inst0$coreir_neg_inst0_out[0]}), .out(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst2$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out), .sel(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst2$coreir_ugt8_inst0_out));
coreir_neg #(.width(8)) NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst2$Negate8_inst0$coreir_neg_inst0(.in({FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst23$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst22$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst21$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst20$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst19$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst18$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst17$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst16$reg_P_inst0_out[0]}), .out(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst2$Negate8_inst0$coreir_neg_inst0_out));
coreir_ugt #(.width(8)) NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst2$coreir_ugt8_inst0(.in0({FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst23$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst22$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst21$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst20$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst19$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst18$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst17$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst16$reg_P_inst0_out[0]}), .in1(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst2$Negate8_inst0$coreir_neg_inst0_out), .out(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst2$coreir_ugt8_inst0_out));
coreir_mux #(.width(8)) NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst3$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join(.in0({FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst31$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst30$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst29$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst28$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst27$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst26$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst25$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst24$reg_P_inst0_out[0]}), .in1({NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst3$Negate8_inst0$coreir_neg_inst0_out[7],NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst3$Negate8_inst0$coreir_neg_inst0_out[6],NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst3$Negate8_inst0$coreir_neg_inst0_out[5],NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst3$Negate8_inst0$coreir_neg_inst0_out[4],NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst3$Negate8_inst0$coreir_neg_inst0_out[3],NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst3$Negate8_inst0$coreir_neg_inst0_out[2],NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst3$Negate8_inst0$coreir_neg_inst0_out[1],NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst3$Negate8_inst0$coreir_neg_inst0_out[0]}), .out(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst3$Mux_Array_8_Bit_t_2n_inst0$CommonlibMuxN_n2_w8_inst0$_join_out), .sel(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst3$coreir_ugt8_inst0_out));
coreir_neg #(.width(8)) NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst3$Negate8_inst0$coreir_neg_inst0(.in({FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst31$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst30$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst29$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst28$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst27$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst26$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst25$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst24$reg_P_inst0_out[0]}), .out(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst3$Negate8_inst0$coreir_neg_inst0_out));
coreir_ugt #(.width(8)) NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst3$coreir_ugt8_inst0(.in0({FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst31$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst30$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst29$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst28$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst27$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst26$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst25$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst24$reg_P_inst0_out[0]}), .in1(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst3$Negate8_inst0$coreir_neg_inst0_out), .out(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$Abs_Atom_inst3$coreir_ugt8_inst0_out));
corebit_and NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$and_inst0(.in0(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Bitt_0init_FalseCE_FalseRESET_inst0$Register1_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out[0]), .in1(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Bitt_0init_FalseCE_FalseRESET_inst0$Register1_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out[0]), .out(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$and_inst0_out));
corebit_and NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$and_inst1(.in0(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$and_inst0_out), .in1(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Bitt_0init_FalseCE_FalseRESET_inst0$Register1_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out[0]), .out(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$and_inst1_out));
corebit_and NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$and_inst2(.in0(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$and_inst1_out), .in1(FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0$Register_Bitt_0init_FalseCE_FalseRESET_inst0$Register1_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out[0]), .out(NativeMapParallel_n4_opAbs_Atom_I_Array_8_In_Bit___O_Array_8_Out_Bit___valid_up_In_Bit__valid_down_Out_Bit___inst0$and_inst2_out));
assign O_0 = {FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out[0]};
assign O_1 = {FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst15$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst14$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst13$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst12$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst11$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst10$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst9$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst8$reg_P_inst0_out[0]};
assign O_2 = {FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst23$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst22$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst21$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst20$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst19$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst18$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst17$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst16$reg_P_inst0_out[0]};
assign O_3 = {FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst31$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst30$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst29$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst28$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst27$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst26$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst25$reg_P_inst0_out[0],FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Array_4_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0$Register32_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst24$reg_P_inst0_out[0]};
assign valid_down = FIFO_tSSeq_4_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3$Register_Bitt_0init_FalseCE_FalseRESET_inst0$Register1_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0_out[0];
endmodule

