// Latency = 4
module Top(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  input  [7:0] I_2,
  input  [7:0] I_3,
  output [7:0] O_0_0_0,
  output [7:0] O_1_0_0,
  output [7:0] O_2_0_0,
  output [7:0] O_3_0_0
);
  wire dontcare;
  wire [31:0] io_output_counts_1;
  wire [31:0] io_output_counts_0;

  x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1 sampler_box ( // @[m_x55_ctr_0.scala 26:17:@1721.4]
    .clock(clock), // @[:@1296.4]
    .reset('b0), // @[:@1297.4]
    .io_in_x480_TREADY(dontcare), // @[:@1298.4]
    .io_in_x480_TDATA({I_0,I_1,I_2,I_3}), // @[:@1298.4]
    .io_in_x480_TID(8'h0),
    .io_in_x480_TDEST(8'h0),
    .io_in_x481_TVALID(valid_down), // @[:@1298.4]
    .io_in_x481_TDATA({O_0_0_0,O_1_0_0,O_2_0_0,O_3_0_0}), // @[:@1298.4]
    .io_in_x481_TREADY(1'b1), // @[:@1298.4]
    .io_sigsIn_datapathEn(valid_up), // @[:@1298.4]
    .io_sigsIn_backpressure(1'b1), // @[:@20563.4]
    .io_sigsIn_break(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_1(io_output_counts_1), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_0(io_output_counts_0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_0(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_1(1'b0), // @[:@20563.4]
    .io_rr('b1) // @[:@1298.4]
  );

  wire dontcare2;

  wire io_output_oobs_0;
  wire io_output_oobs_1;
  x488_ctrchain cchain ( // @[:@2879.2]
    .clock(clock), // @[:@2880.4]
    .reset(1'b0), // @[:@2881.4]
    .io_input_reset(1'b0), // @[:@2882.4]
    .io_input_enable(valid_up), // @[:@2882.4]
    .io_output_counts_1(io_output_counts_1), // @[:@2882.4]
    .io_output_counts_0(io_output_counts_0), // @[:@2882.4]
    .io_output_oobs_0(io_output_oobs_0), // @[:@2882.4]
    .io_output_oobs_1(io_output_oobs_1), // @[:@2882.4]
    .io_output_done(dontcare2) // @[:@2882.4]
  );

endmodule

module SRAMVerilogSim
#(
    parameter WORDS = 1024,
    parameter AWIDTH = 10,
    parameter DWIDTH = 32)
(
    input clk,
    input [AWIDTH-1:0] raddr,
    input [AWIDTH-1:0] waddr,
    input raddrEn,
    input waddrEn,
    input wen,
    input [DWIDTH-1:0] wdata,
    input backpressure,
    output reg [DWIDTH-1:0] rdata
);

    reg [DWIDTH-1:0] mem [0:WORDS-1];

    always @(posedge clk) begin
      if (wen) mem[waddr] <= wdata;
      if (backpressure) rdata <= mem[raddr];
    end

endmodule
module RetimeShiftRegister
#(
    parameter WIDTH = 1,
    parameter STAGES = 1)
(
    input clock,
    input reset,
    input flow,
    input [WIDTH-1:0] init,
    input [WIDTH-1:0] in,
    output reg [WIDTH-1:0] out
);
  integer i;
  reg [WIDTH-1:0] sr[STAGES:0]; // Create 'STAGES' number of register, each 'WIDTH' bits wide

   /* synopsys dc_tcl_script_begin
    set_ungroup [current_design] true
    set_flatten true -effort high -phase true -design [current_design]
    set_dont_retime [current_design] false
    set_optimize_registers true -design [current_design]
    */
  always @(posedge clock) begin
    if (reset) begin
      for(i=0; i<STAGES; i=i+1) begin
        sr[i] <= init;
      end
    end else begin
      if (flow) begin 
        sr[0] <= in;
        for(i=1; i<STAGES; i=i+1) begin
          sr[i] <= sr[i-1];
        end
      end
    end
  end

  always @(*) begin
    out = sr[STAGES-1];
  end
endmodule
module FF( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  output [31:0] io_rPort_0_output_0, // @[:@6.4]
  input  [31:0] io_wPort_0_data_0, // @[:@6.4]
  input         io_wPort_0_reset // @[:@6.4]
);
  reg [31:0] ff; // @[MemPrimitives.scala 311:19:@21.4]
  reg [31:0] _RAND_0;
  wire [31:0] _T_69; // @[MemPrimitives.scala 315:12:@24.4]
  assign _T_69 = io_wPort_0_reset ? 32'h0 : io_wPort_0_data_0; // @[MemPrimitives.scala 315:12:@24.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 316:34:@26.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 32'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 32'h0;
      end else begin
        ff <= io_wPort_0_data_0;
      end
    end
  end
endmodule
module SRFF( // @[:@28.2]
  input   clock, // @[:@29.4]
  input   reset, // @[:@30.4]
  input   io_input_set, // @[:@31.4]
  input   io_input_reset, // @[:@31.4]
  input   io_input_asyn_reset, // @[:@31.4]
  output  io_output // @[:@31.4]
);
  reg  _T_15; // @[SRFF.scala 20:21:@33.4]
  reg [31:0] _RAND_0;
  wire  _T_19; // @[SRFF.scala 21:74:@34.4]
  wire  _T_20; // @[SRFF.scala 21:48:@35.4]
  wire  _T_21; // @[SRFF.scala 21:14:@36.4]
  assign _T_19 = io_input_reset ? 1'h0 : _T_15; // @[SRFF.scala 21:74:@34.4]
  assign _T_20 = io_input_set ? 1'h1 : _T_19; // @[SRFF.scala 21:48:@35.4]
  assign _T_21 = io_input_asyn_reset ? 1'h0 : _T_20; // @[SRFF.scala 21:14:@36.4]
  assign io_output = io_input_asyn_reset ? 1'h0 : _T_15; // @[SRFF.scala 22:15:@39.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_15 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_15 <= 1'h0;
    end else begin
      if (io_input_asyn_reset) begin
        _T_15 <= 1'h0;
      end else begin
        if (io_input_set) begin
          _T_15 <= 1'h1;
        end else begin
          if (io_input_reset) begin
            _T_15 <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module SingleCounter( // @[:@41.2]
  input   clock, // @[:@42.4]
  input   reset, // @[:@43.4]
  input   io_input_reset, // @[:@44.4]
  output  io_output_done // @[:@44.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@57.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@57.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@57.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@57.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@57.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@73.4]
  wire [31:0] _T_48; // @[Counter.scala 287:52:@101.4]
  wire [32:0] _T_50; // @[Counter.scala 291:33:@102.4]
  wire [31:0] _T_51; // @[Counter.scala 291:33:@103.4]
  wire [31:0] _T_52; // @[Counter.scala 291:33:@104.4]
  wire  _T_57; // @[Counter.scala 293:18:@106.4]
  wire [31:0] _T_68; // @[Counter.scala 299:115:@114.4]
  wire [31:0] _T_71; // @[Counter.scala 299:152:@117.4]
  wire [31:0] _T_72; // @[Counter.scala 299:74:@118.4]
  FF bases_0 ( // @[Counter.scala 261:53:@57.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@73.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@101.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@102.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@103.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@104.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh37); // @[Counter.scala 293:18:@106.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@114.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@117.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 299:74:@118.4]
  assign io_output_done = $signed(_T_52) >= $signed(32'sh37); // @[Counter.scala 333:20:@127.4]
  assign bases_0_clock = clock; // @[:@58.4]
  assign bases_0_reset = reset; // @[:@59.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 299:31:@120.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@99.4]
  assign SRFF_clock = clock; // @[:@74.4]
  assign SRFF_reset = reset; // @[:@75.4]
  assign SRFF_io_input_set = io_input_reset == 1'h0; // @[Counter.scala 264:23:@78.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@80.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@81.4]
endmodule
module RetimeWrapper( // @[:@144.2]
  input   clock, // @[:@145.4]
  input   reset, // @[:@146.4]
  input   io_flow, // @[:@147.4]
  input   io_in, // @[:@147.4]
  output  io_out // @[:@147.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@149.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@149.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@162.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@161.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@160.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@159.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@158.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@156.4]
endmodule
module RootController_sm( // @[:@312.2]
  input   clock, // @[:@313.4]
  input   reset, // @[:@314.4]
  input   io_enable, // @[:@315.4]
  output  io_done, // @[:@315.4]
  input   io_rst, // @[:@315.4]
  input   io_ctrDone, // @[:@315.4]
  output  io_ctrInc, // @[:@315.4]
  input   io_parentAck, // @[:@315.4]
  input   io_doneIn_0, // @[:@315.4]
  output  io_enableOut_0, // @[:@315.4]
  output  io_childAck_0 // @[:@315.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@318.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@321.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@338.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@433.4]
  wire  finished; // @[Controllers.scala 81:26:@324.4]
  wire  _T_81; // @[Controllers.scala 86:43:@328.4]
  wire  synchronize; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  wire  _T_93; // @[Controllers.scala 92:52:@342.4]
  wire  _T_122; // @[Controllers.scala 128:33:@371.4]
  wire  _T_124; // @[Controllers.scala 128:54:@372.4]
  wire  _T_125; // @[Controllers.scala 128:52:@373.4]
  wire  _T_126; // @[Controllers.scala 128:66:@374.4]
  wire  _T_128; // @[Controllers.scala 128:98:@376.4]
  wire  _T_129; // @[Controllers.scala 128:96:@377.4]
  wire  _T_131; // @[Controllers.scala 128:123:@378.4]
  wire  _T_133; // @[Controllers.scala 129:48:@381.4]
  wire  _T_134; // @[Controllers.scala 129:57:@382.4]
  wire  _T_138; // @[Controllers.scala 130:52:@386.4]
  wire  _T_139; // @[Controllers.scala 130:50:@387.4]
  wire  _T_147; // @[Controllers.scala 130:129:@393.4]
  wire  _T_150; // @[Controllers.scala 131:45:@396.4]
  wire  _T_154; // @[Controllers.scala 213:68:@402.4]
  wire  _T_156; // @[Controllers.scala 213:90:@404.4]
  wire  _T_158; // @[Controllers.scala 213:132:@406.4]
  wire  _T_159; // @[Controllers.scala 213:130:@407.4]
  wire  _T_160; // @[Controllers.scala 213:156:@408.4]
  reg  _T_166; // @[package.scala 48:56:@412.4]
  reg [31:0] _RAND_0;
  wire  _T_167; // @[package.scala 100:41:@414.4]
  reg  _T_180; // @[package.scala 48:56:@430.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@318.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@321.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@338.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@357.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@416.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@433.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  assign finished = done_0_io_output | io_done; // @[Controllers.scala 81:26:@324.4]
  assign _T_81 = io_rst | done_0_io_output; // @[Controllers.scala 86:43:@328.4]
  assign synchronize = RetimeWrapper_io_out; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  assign _T_93 = synchronize | io_rst; // @[Controllers.scala 92:52:@342.4]
  assign _T_122 = done_0_io_output == 1'h0; // @[Controllers.scala 128:33:@371.4]
  assign _T_124 = io_ctrDone == 1'h0; // @[Controllers.scala 128:54:@372.4]
  assign _T_125 = _T_122 & _T_124; // @[Controllers.scala 128:52:@373.4]
  assign _T_126 = _T_125 & io_enable; // @[Controllers.scala 128:66:@374.4]
  assign _T_128 = ~ iterDone_0_io_output; // @[Controllers.scala 128:98:@376.4]
  assign _T_129 = _T_126 & _T_128; // @[Controllers.scala 128:96:@377.4]
  assign _T_131 = io_doneIn_0 == 1'h0; // @[Controllers.scala 128:123:@378.4]
  assign _T_133 = io_doneIn_0 | io_rst; // @[Controllers.scala 129:48:@381.4]
  assign _T_134 = _T_133 | io_parentAck; // @[Controllers.scala 129:57:@382.4]
  assign _T_138 = synchronize == 1'h0; // @[Controllers.scala 130:52:@386.4]
  assign _T_139 = io_doneIn_0 & _T_138; // @[Controllers.scala 130:50:@387.4]
  assign _T_147 = finished == 1'h0; // @[Controllers.scala 130:129:@393.4]
  assign _T_150 = io_rst == 1'h0; // @[Controllers.scala 131:45:@396.4]
  assign _T_154 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@402.4]
  assign _T_156 = _T_154 & _T_128; // @[Controllers.scala 213:90:@404.4]
  assign _T_158 = ~ done_0_io_output; // @[Controllers.scala 213:132:@406.4]
  assign _T_159 = _T_156 & _T_158; // @[Controllers.scala 213:130:@407.4]
  assign _T_160 = ~ io_ctrDone; // @[Controllers.scala 213:156:@408.4]
  assign _T_167 = done_0_io_output & _T_166; // @[package.scala 100:41:@414.4]
  assign io_done = RetimeWrapper_2_io_out; // @[Controllers.scala 245:13:@440.4]
  assign io_ctrInc = io_doneIn_0; // @[Controllers.scala 122:17:@356.4]
  assign io_enableOut_0 = _T_159 & _T_160; // @[Controllers.scala 213:55:@410.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@401.4]
  assign active_0_clock = clock; // @[:@319.4]
  assign active_0_reset = reset; // @[:@320.4]
  assign active_0_io_input_set = _T_129 & _T_131; // @[Controllers.scala 128:30:@380.4]
  assign active_0_io_input_reset = _T_134 | done_0_io_output; // @[Controllers.scala 129:32:@385.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@326.4]
  assign done_0_clock = clock; // @[:@322.4]
  assign done_0_reset = reset; // @[:@323.4]
  assign done_0_io_input_set = io_ctrDone & _T_150; // @[Controllers.scala 131:28:@399.4]
  assign done_0_io_input_reset = _T_81 | io_parentAck; // @[Controllers.scala 86:33:@336.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@327.4]
  assign iterDone_0_clock = clock; // @[:@339.4]
  assign iterDone_0_reset = reset; // @[:@340.4]
  assign iterDone_0_io_input_set = _T_139 & _T_147; // @[Controllers.scala 130:32:@395.4]
  assign iterDone_0_io_input_reset = _T_93 | io_parentAck; // @[Controllers.scala 92:37:@350.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@341.4]
  assign RetimeWrapper_clock = clock; // @[:@358.4]
  assign RetimeWrapper_reset = reset; // @[:@359.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@361.4]
  assign RetimeWrapper_io_in = io_doneIn_0; // @[package.scala 94:16:@360.4]
  assign RetimeWrapper_1_clock = clock; // @[:@417.4]
  assign RetimeWrapper_1_reset = reset; // @[:@418.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@420.4]
  assign RetimeWrapper_1_io_in = _T_167 | io_parentAck; // @[package.scala 94:16:@419.4]
  assign RetimeWrapper_2_clock = clock; // @[:@434.4]
  assign RetimeWrapper_2_reset = reset; // @[:@435.4]
  assign RetimeWrapper_2_io_flow = io_enable; // @[package.scala 95:18:@437.4]
  assign RetimeWrapper_2_io_in = done_0_io_output & _T_180; // @[package.scala 94:16:@436.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_166 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_180 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_166 <= 1'h0;
    end else begin
      _T_166 <= _T_122;
    end
    if (reset) begin
      _T_180 <= 1'h0;
    end else begin
      _T_180 <= _T_122;
    end
  end
endmodule
module SRAM( // @[:@507.2]
  input         clock, // @[:@508.4]
  input  [20:0] io_raddr, // @[:@510.4]
  output [7:0]  io_rdata, // @[:@510.4]
  input         io_backpressure // @[:@510.4]
);
  wire [7:0] SRAMVerilogSim_rdata; // @[SRAM.scala 185:23:@512.4]
  wire [7:0] SRAMVerilogSim_wdata; // @[SRAM.scala 185:23:@512.4]
  wire  SRAMVerilogSim_backpressure; // @[SRAM.scala 185:23:@512.4]
  wire  SRAMVerilogSim_wen; // @[SRAM.scala 185:23:@512.4]
  wire  SRAMVerilogSim_waddrEn; // @[SRAM.scala 185:23:@512.4]
  wire  SRAMVerilogSim_raddrEn; // @[SRAM.scala 185:23:@512.4]
  wire [20:0] SRAMVerilogSim_waddr; // @[SRAM.scala 185:23:@512.4]
  wire [20:0] SRAMVerilogSim_raddr; // @[SRAM.scala 185:23:@512.4]
  wire  SRAMVerilogSim_clk; // @[SRAM.scala 185:23:@512.4]
  SRAMVerilogSim #(.DWIDTH(8), .WORDS(2073600), .AWIDTH(21)) SRAMVerilogSim ( // @[SRAM.scala 185:23:@512.4]
    .rdata(SRAMVerilogSim_rdata),
    .wdata(SRAMVerilogSim_wdata),
    .backpressure(SRAMVerilogSim_backpressure),
    .wen(SRAMVerilogSim_wen),
    .waddrEn(SRAMVerilogSim_waddrEn),
    .raddrEn(SRAMVerilogSim_raddrEn),
    .waddr(SRAMVerilogSim_waddr),
    .raddr(SRAMVerilogSim_raddr),
    .clk(SRAMVerilogSim_clk)
  );
  assign io_rdata = SRAMVerilogSim_rdata; // @[SRAM.scala 195:16:@532.4]
  assign SRAMVerilogSim_wdata = 8'h0; // @[SRAM.scala 190:20:@526.4]
  assign SRAMVerilogSim_backpressure = io_backpressure; // @[SRAM.scala 191:27:@527.4]
  assign SRAMVerilogSim_wen = 1'h0; // @[SRAM.scala 188:18:@524.4]
  assign SRAMVerilogSim_waddrEn = 1'h1; // @[SRAM.scala 193:22:@529.4]
  assign SRAMVerilogSim_raddrEn = 1'h1; // @[SRAM.scala 192:22:@528.4]
  assign SRAMVerilogSim_waddr = 21'h0; // @[SRAM.scala 189:20:@525.4]
  assign SRAMVerilogSim_raddr = io_raddr; // @[SRAM.scala 187:20:@523.4]
  assign SRAMVerilogSim_clk = clock; // @[SRAM.scala 186:18:@522.4]
endmodule
module RetimeWrapper_5( // @[:@546.2]
  input         clock, // @[:@547.4]
  input         reset, // @[:@548.4]
  input         io_flow, // @[:@549.4]
  input  [20:0] io_in, // @[:@549.4]
  output [20:0] io_out // @[:@549.4]
);
  wire [20:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@551.4]
  wire [20:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@551.4]
  wire [20:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@551.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@551.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@551.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@551.4]
  RetimeShiftRegister #(.WIDTH(21), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@551.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@564.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@563.4]
  assign sr_init = 21'h0; // @[RetimeShiftRegister.scala 19:16:@562.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@561.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@560.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@558.4]
endmodule
module Mem1D( // @[:@566.2]
  input         clock, // @[:@567.4]
  input         reset, // @[:@568.4]
  input  [20:0] io_r_ofs_0, // @[:@569.4]
  input         io_r_backpressure, // @[:@569.4]
  output [7:0]  io_output // @[:@569.4]
);
  wire  SRAM_clock; // @[MemPrimitives.scala 705:21:@573.4]
  wire [20:0] SRAM_io_raddr; // @[MemPrimitives.scala 705:21:@573.4]
  wire [7:0] SRAM_io_rdata; // @[MemPrimitives.scala 705:21:@573.4]
  wire  SRAM_io_backpressure; // @[MemPrimitives.scala 705:21:@573.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@576.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@576.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@576.4]
  wire [20:0] RetimeWrapper_io_in; // @[package.scala 93:22:@576.4]
  wire [20:0] RetimeWrapper_io_out; // @[package.scala 93:22:@576.4]
  SRAM SRAM ( // @[MemPrimitives.scala 705:21:@573.4]
    .clock(SRAM_clock),
    .io_raddr(SRAM_io_raddr),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  RetimeWrapper_5 RetimeWrapper ( // @[package.scala 93:22:@576.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_output = SRAM_io_rdata; // @[MemPrimitives.scala 712:17:@589.4]
  assign SRAM_clock = clock; // @[:@574.4]
  assign SRAM_io_raddr = RetimeWrapper_io_out; // @[MemPrimitives.scala 706:37:@583.4]
  assign SRAM_io_backpressure = io_r_backpressure; // @[MemPrimitives.scala 711:30:@588.4]
  assign RetimeWrapper_clock = clock; // @[:@577.4]
  assign RetimeWrapper_reset = reset; // @[:@578.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@580.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@579.4]
endmodule
module StickySelects( // @[:@591.2]
  input   io_ins_0, // @[:@594.4]
  output  io_outs_0 // @[:@594.4]
);
  assign io_outs_0 = io_ins_0; // @[StickySelects.scala 34:26:@596.4]
endmodule
module RetimeWrapper_6( // @[:@610.2]
  input   clock, // @[:@611.4]
  input   reset, // @[:@612.4]
  input   io_flow, // @[:@613.4]
  input   io_in, // @[:@613.4]
  output  io_out // @[:@613.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@615.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@615.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@615.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@615.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@615.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@615.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@615.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@628.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@627.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@626.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@625.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@624.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@622.4]
endmodule
module x482_outbuf_0( // @[:@630.2]
  input         clock, // @[:@631.4]
  input         reset, // @[:@632.4]
  input  [20:0] io_rPort_0_ofs_0, // @[:@633.4]
  input         io_rPort_0_en_0, // @[:@633.4]
  input         io_rPort_0_backpressure, // @[:@633.4]
  output [7:0]  io_rPort_0_output_0 // @[:@633.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@648.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@648.4]
  wire [20:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@648.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@648.4]
  wire [7:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@648.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 121:29:@674.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 121:29:@674.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@688.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@688.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@688.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@688.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@688.4]
  wire  _T_76; // @[MemPrimitives.scala 123:41:@678.4]
  wire [22:0] _T_78; // @[Cat.scala 30:58:@680.4]
  Mem1D Mem1D ( // @[MemPrimitives.scala 64:21:@648.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_output(Mem1D_io_output)
  );
  StickySelects StickySelects ( // @[MemPrimitives.scala 121:29:@674.4]
    .io_ins_0(StickySelects_io_ins_0),
    .io_outs_0(StickySelects_io_outs_0)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@688.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_76 = StickySelects_io_outs_0; // @[MemPrimitives.scala 123:41:@678.4]
  assign _T_78 = {_T_76,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@680.4]
  assign io_rPort_0_output_0 = Mem1D_io_output; // @[MemPrimitives.scala 148:13:@695.4]
  assign Mem1D_clock = clock; // @[:@649.4]
  assign Mem1D_reset = reset; // @[:@650.4]
  assign Mem1D_io_r_ofs_0 = _T_78[20:0]; // @[MemPrimitives.scala 127:28:@684.4]
  assign Mem1D_io_r_backpressure = _T_78[21]; // @[MemPrimitives.scala 128:32:@685.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0; // @[MemPrimitives.scala 122:60:@677.4]
  assign RetimeWrapper_clock = clock; // @[:@689.4]
  assign RetimeWrapper_reset = reset; // @[:@690.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@692.4]
  assign RetimeWrapper_io_in = io_rPort_0_en_0; // @[package.scala 94:16:@691.4]
endmodule
module x819_sm( // @[:@839.2]
  input   clock, // @[:@840.4]
  input   reset, // @[:@841.4]
  input   io_enable, // @[:@842.4]
  output  io_done, // @[:@842.4]
  input   io_ctrDone, // @[:@842.4]
  output  io_ctrInc, // @[:@842.4]
  input   io_parentAck, // @[:@842.4]
  input   io_doneIn_0, // @[:@842.4]
  input   io_doneIn_1, // @[:@842.4]
  output  io_enableOut_0, // @[:@842.4]
  output  io_enableOut_1, // @[:@842.4]
  output  io_childAck_0, // @[:@842.4]
  output  io_childAck_1 // @[:@842.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@845.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@845.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@845.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@845.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@845.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@845.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@848.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@848.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@848.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@848.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@848.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@848.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@851.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@851.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@851.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@851.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@851.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@851.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@854.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@854.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@854.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@854.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@854.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@854.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@883.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@883.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@883.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@883.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@883.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@883.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@886.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@886.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@886.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@886.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@886.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@886.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@987.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@987.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@987.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@987.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@987.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@1004.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@1004.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@1004.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@1004.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@1004.4]
  wire  allDone; // @[Controllers.scala 80:47:@857.4]
  wire  synchronize; // @[Controllers.scala 146:56:@911.4]
  wire  _T_127; // @[Controllers.scala 150:35:@913.4]
  wire  _T_129; // @[Controllers.scala 150:60:@914.4]
  wire  _T_130; // @[Controllers.scala 150:58:@915.4]
  wire  _T_132; // @[Controllers.scala 150:76:@916.4]
  wire  _T_133; // @[Controllers.scala 150:74:@917.4]
  wire  _T_135; // @[Controllers.scala 150:97:@918.4]
  wire  _T_136; // @[Controllers.scala 150:95:@919.4]
  wire  _T_152; // @[Controllers.scala 150:35:@937.4]
  wire  _T_154; // @[Controllers.scala 150:60:@938.4]
  wire  _T_155; // @[Controllers.scala 150:58:@939.4]
  wire  _T_157; // @[Controllers.scala 150:76:@940.4]
  wire  _T_158; // @[Controllers.scala 150:74:@941.4]
  wire  _T_161; // @[Controllers.scala 150:95:@943.4]
  wire  _T_179; // @[Controllers.scala 213:68:@965.4]
  wire  _T_181; // @[Controllers.scala 213:90:@967.4]
  wire  _T_183; // @[Controllers.scala 213:132:@969.4]
  wire  _T_184; // @[Controllers.scala 213:130:@970.4]
  wire  _T_185; // @[Controllers.scala 213:156:@971.4]
  wire  _T_187; // @[Controllers.scala 213:68:@974.4]
  wire  _T_189; // @[Controllers.scala 213:90:@976.4]
  wire  _T_196; // @[package.scala 100:49:@982.4]
  reg  _T_199; // @[package.scala 48:56:@983.4]
  reg [31:0] _RAND_0;
  wire  _T_200; // @[package.scala 100:41:@985.4]
  reg  _T_213; // @[package.scala 48:56:@1001.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@845.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@848.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@851.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@854.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@883.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@886.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@987.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@1004.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign allDone = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@857.4]
  assign synchronize = iterDone_0_io_output & iterDone_1_io_output; // @[Controllers.scala 146:56:@911.4]
  assign _T_127 = ~ iterDone_0_io_output; // @[Controllers.scala 150:35:@913.4]
  assign _T_129 = io_doneIn_0 == 1'h0; // @[Controllers.scala 150:60:@914.4]
  assign _T_130 = _T_127 & _T_129; // @[Controllers.scala 150:58:@915.4]
  assign _T_132 = done_0_io_output == 1'h0; // @[Controllers.scala 150:76:@916.4]
  assign _T_133 = _T_130 & _T_132; // @[Controllers.scala 150:74:@917.4]
  assign _T_135 = io_ctrDone == 1'h0; // @[Controllers.scala 150:97:@918.4]
  assign _T_136 = _T_133 & _T_135; // @[Controllers.scala 150:95:@919.4]
  assign _T_152 = ~ iterDone_1_io_output; // @[Controllers.scala 150:35:@937.4]
  assign _T_154 = io_doneIn_1 == 1'h0; // @[Controllers.scala 150:60:@938.4]
  assign _T_155 = _T_152 & _T_154; // @[Controllers.scala 150:58:@939.4]
  assign _T_157 = done_1_io_output == 1'h0; // @[Controllers.scala 150:76:@940.4]
  assign _T_158 = _T_155 & _T_157; // @[Controllers.scala 150:74:@941.4]
  assign _T_161 = _T_158 & _T_135; // @[Controllers.scala 150:95:@943.4]
  assign _T_179 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@965.4]
  assign _T_181 = _T_179 & _T_127; // @[Controllers.scala 213:90:@967.4]
  assign _T_183 = ~ allDone; // @[Controllers.scala 213:132:@969.4]
  assign _T_184 = _T_181 & _T_183; // @[Controllers.scala 213:130:@970.4]
  assign _T_185 = ~ io_ctrDone; // @[Controllers.scala 213:156:@971.4]
  assign _T_187 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@974.4]
  assign _T_189 = _T_187 & _T_152; // @[Controllers.scala 213:90:@976.4]
  assign _T_196 = allDone == 1'h0; // @[package.scala 100:49:@982.4]
  assign _T_200 = allDone & _T_199; // @[package.scala 100:41:@985.4]
  assign io_done = RetimeWrapper_1_io_out; // @[Controllers.scala 245:13:@1011.4]
  assign io_ctrInc = iterDone_0_io_output & iterDone_1_io_output; // @[Controllers.scala 143:17:@910.4]
  assign io_enableOut_0 = _T_184 & _T_185; // @[Controllers.scala 213:55:@973.4]
  assign io_enableOut_1 = _T_189 & _T_183; // @[Controllers.scala 213:55:@981.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@962.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@964.4]
  assign active_0_clock = clock; // @[:@846.4]
  assign active_0_reset = reset; // @[:@847.4]
  assign active_0_io_input_set = _T_136 & io_enable; // @[Controllers.scala 150:32:@922.4]
  assign active_0_io_input_reset = io_doneIn_0 | io_parentAck; // @[Controllers.scala 151:34:@926.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@860.4]
  assign active_1_clock = clock; // @[:@849.4]
  assign active_1_reset = reset; // @[:@850.4]
  assign active_1_io_input_set = _T_161 & io_enable; // @[Controllers.scala 150:32:@946.4]
  assign active_1_io_input_reset = io_doneIn_1 | io_parentAck; // @[Controllers.scala 151:34:@950.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@861.4]
  assign done_0_clock = clock; // @[:@852.4]
  assign done_0_reset = reset; // @[:@853.4]
  assign done_0_io_input_set = io_ctrDone; // @[Controllers.scala 153:30:@936.4]
  assign done_0_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@872.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@862.4]
  assign done_1_clock = clock; // @[:@855.4]
  assign done_1_reset = reset; // @[:@856.4]
  assign done_1_io_input_set = io_ctrDone; // @[Controllers.scala 153:30:@960.4]
  assign done_1_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@881.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@863.4]
  assign iterDone_0_clock = clock; // @[:@884.4]
  assign iterDone_0_reset = reset; // @[:@885.4]
  assign iterDone_0_io_input_set = io_doneIn_0; // @[Controllers.scala 152:34:@932.4]
  assign iterDone_0_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@899.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@889.4]
  assign iterDone_1_clock = clock; // @[:@887.4]
  assign iterDone_1_reset = reset; // @[:@888.4]
  assign iterDone_1_io_input_set = io_doneIn_1; // @[Controllers.scala 152:34:@956.4]
  assign iterDone_1_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@908.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@890.4]
  assign RetimeWrapper_clock = clock; // @[:@988.4]
  assign RetimeWrapper_reset = reset; // @[:@989.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@991.4]
  assign RetimeWrapper_io_in = _T_200 | io_parentAck; // @[package.scala 94:16:@990.4]
  assign RetimeWrapper_1_clock = clock; // @[:@1005.4]
  assign RetimeWrapper_1_reset = reset; // @[:@1006.4]
  assign RetimeWrapper_1_io_flow = io_enable; // @[package.scala 95:18:@1008.4]
  assign RetimeWrapper_1_io_in = allDone & _T_213; // @[package.scala 94:16:@1007.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_199 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_213 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_199 <= 1'h0;
    end else begin
      _T_199 <= _T_196;
    end
    if (reset) begin
      _T_213 <= 1'h0;
    end else begin
      _T_213 <= _T_196;
    end
  end
endmodule
module x738_outr_UnitPipe_sm( // @[:@1428.2]
  input   clock, // @[:@1429.4]
  input   reset, // @[:@1430.4]
  input   io_enable, // @[:@1431.4]
  output  io_done, // @[:@1431.4]
  input   io_parentAck, // @[:@1431.4]
  input   io_doneIn_0, // @[:@1431.4]
  input   io_doneIn_1, // @[:@1431.4]
  output  io_enableOut_0, // @[:@1431.4]
  output  io_enableOut_1, // @[:@1431.4]
  output  io_childAck_0, // @[:@1431.4]
  output  io_childAck_1, // @[:@1431.4]
  input   io_ctrCopyDone_0, // @[:@1431.4]
  input   io_ctrCopyDone_1 // @[:@1431.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@1434.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@1434.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@1434.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@1434.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@1434.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@1434.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@1437.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@1437.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@1437.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@1437.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@1437.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@1437.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@1440.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@1440.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@1440.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@1440.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@1440.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@1440.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@1443.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@1443.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@1443.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@1443.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@1443.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@1443.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@1472.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@1472.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@1472.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@1472.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@1472.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@1472.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@1475.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@1475.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@1475.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@1475.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@1475.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@1475.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@1516.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@1516.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@1516.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@1516.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@1516.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@1530.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@1530.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@1530.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@1530.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@1530.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@1548.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@1548.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@1548.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@1548.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@1548.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@1585.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@1585.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@1585.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@1585.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@1585.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@1599.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@1599.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@1599.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@1599.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@1599.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@1617.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@1617.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@1617.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@1617.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@1617.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@1664.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@1664.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@1664.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@1664.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@1664.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@1681.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@1681.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@1681.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@1681.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@1681.4]
  wire  allDone; // @[Controllers.scala 80:47:@1446.4]
  wire  _T_127; // @[Controllers.scala 165:35:@1500.4]
  wire  _T_129; // @[Controllers.scala 165:60:@1501.4]
  wire  _T_130; // @[Controllers.scala 165:58:@1502.4]
  wire  _T_132; // @[Controllers.scala 165:76:@1503.4]
  wire  _T_133; // @[Controllers.scala 165:74:@1504.4]
  wire  _T_137; // @[Controllers.scala 165:109:@1507.4]
  wire  _T_140; // @[Controllers.scala 165:141:@1509.4]
  wire  _T_148; // @[package.scala 96:25:@1521.4 package.scala 96:25:@1522.4]
  wire  _T_152; // @[Controllers.scala 167:54:@1524.4]
  wire  _T_153; // @[Controllers.scala 167:52:@1525.4]
  wire  _T_160; // @[package.scala 96:25:@1535.4 package.scala 96:25:@1536.4]
  wire  _T_178; // @[package.scala 96:25:@1553.4 package.scala 96:25:@1554.4]
  wire  _T_182; // @[Controllers.scala 169:67:@1556.4]
  wire  _T_183; // @[Controllers.scala 169:86:@1557.4]
  wire  _T_195; // @[Controllers.scala 165:35:@1569.4]
  wire  _T_197; // @[Controllers.scala 165:60:@1570.4]
  wire  _T_198; // @[Controllers.scala 165:58:@1571.4]
  wire  _T_200; // @[Controllers.scala 165:76:@1572.4]
  wire  _T_201; // @[Controllers.scala 165:74:@1573.4]
  wire  _T_205; // @[Controllers.scala 165:109:@1576.4]
  wire  _T_208; // @[Controllers.scala 165:141:@1578.4]
  wire  _T_216; // @[package.scala 96:25:@1590.4 package.scala 96:25:@1591.4]
  wire  _T_220; // @[Controllers.scala 167:54:@1593.4]
  wire  _T_221; // @[Controllers.scala 167:52:@1594.4]
  wire  _T_228; // @[package.scala 96:25:@1604.4 package.scala 96:25:@1605.4]
  wire  _T_246; // @[package.scala 96:25:@1622.4 package.scala 96:25:@1623.4]
  wire  _T_250; // @[Controllers.scala 169:67:@1625.4]
  wire  _T_251; // @[Controllers.scala 169:86:@1626.4]
  wire  _T_265; // @[Controllers.scala 213:68:@1642.4]
  wire  _T_267; // @[Controllers.scala 213:90:@1644.4]
  wire  _T_269; // @[Controllers.scala 213:132:@1646.4]
  wire  _T_273; // @[Controllers.scala 213:68:@1651.4]
  wire  _T_275; // @[Controllers.scala 213:90:@1653.4]
  wire  _T_282; // @[package.scala 100:49:@1659.4]
  reg  _T_285; // @[package.scala 48:56:@1660.4]
  reg [31:0] _RAND_0;
  wire  _T_286; // @[package.scala 100:41:@1662.4]
  reg  _T_299; // @[package.scala 48:56:@1678.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@1434.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@1437.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@1440.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@1443.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@1472.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@1475.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@1516.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@1530.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@1548.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@1585.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@1599.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@1617.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@1664.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@1681.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  assign allDone = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@1446.4]
  assign _T_127 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@1500.4]
  assign _T_129 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@1501.4]
  assign _T_130 = _T_127 & _T_129; // @[Controllers.scala 165:58:@1502.4]
  assign _T_132 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@1503.4]
  assign _T_133 = _T_130 & _T_132; // @[Controllers.scala 165:74:@1504.4]
  assign _T_137 = _T_133 & io_enable; // @[Controllers.scala 165:109:@1507.4]
  assign _T_140 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@1509.4]
  assign _T_148 = RetimeWrapper_io_out; // @[package.scala 96:25:@1521.4 package.scala 96:25:@1522.4]
  assign _T_152 = _T_148 == 1'h0; // @[Controllers.scala 167:54:@1524.4]
  assign _T_153 = io_doneIn_0 | _T_152; // @[Controllers.scala 167:52:@1525.4]
  assign _T_160 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@1535.4 package.scala 96:25:@1536.4]
  assign _T_178 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@1553.4 package.scala 96:25:@1554.4]
  assign _T_182 = _T_178 == 1'h0; // @[Controllers.scala 169:67:@1556.4]
  assign _T_183 = _T_182 & io_enable; // @[Controllers.scala 169:86:@1557.4]
  assign _T_195 = ~ iterDone_1_io_output; // @[Controllers.scala 165:35:@1569.4]
  assign _T_197 = io_doneIn_1 == 1'h0; // @[Controllers.scala 165:60:@1570.4]
  assign _T_198 = _T_195 & _T_197; // @[Controllers.scala 165:58:@1571.4]
  assign _T_200 = done_1_io_output == 1'h0; // @[Controllers.scala 165:76:@1572.4]
  assign _T_201 = _T_198 & _T_200; // @[Controllers.scala 165:74:@1573.4]
  assign _T_205 = _T_201 & io_enable; // @[Controllers.scala 165:109:@1576.4]
  assign _T_208 = io_ctrCopyDone_1 == 1'h0; // @[Controllers.scala 165:141:@1578.4]
  assign _T_216 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@1590.4 package.scala 96:25:@1591.4]
  assign _T_220 = _T_216 == 1'h0; // @[Controllers.scala 167:54:@1593.4]
  assign _T_221 = io_doneIn_1 | _T_220; // @[Controllers.scala 167:52:@1594.4]
  assign _T_228 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@1604.4 package.scala 96:25:@1605.4]
  assign _T_246 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@1622.4 package.scala 96:25:@1623.4]
  assign _T_250 = _T_246 == 1'h0; // @[Controllers.scala 169:67:@1625.4]
  assign _T_251 = _T_250 & io_enable; // @[Controllers.scala 169:86:@1626.4]
  assign _T_265 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@1642.4]
  assign _T_267 = _T_265 & _T_127; // @[Controllers.scala 213:90:@1644.4]
  assign _T_269 = ~ allDone; // @[Controllers.scala 213:132:@1646.4]
  assign _T_273 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@1651.4]
  assign _T_275 = _T_273 & _T_195; // @[Controllers.scala 213:90:@1653.4]
  assign _T_282 = allDone == 1'h0; // @[package.scala 100:49:@1659.4]
  assign _T_286 = allDone & _T_285; // @[package.scala 100:41:@1662.4]
  assign io_done = RetimeWrapper_7_io_out; // @[Controllers.scala 245:13:@1688.4]
  assign io_enableOut_0 = _T_267 & _T_269; // @[Controllers.scala 213:55:@1650.4]
  assign io_enableOut_1 = _T_275 & _T_269; // @[Controllers.scala 213:55:@1658.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@1639.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@1641.4]
  assign active_0_clock = clock; // @[:@1435.4]
  assign active_0_reset = reset; // @[:@1436.4]
  assign active_0_io_input_set = _T_137 & _T_140; // @[Controllers.scala 165:32:@1511.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@1515.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@1449.4]
  assign active_1_clock = clock; // @[:@1438.4]
  assign active_1_reset = reset; // @[:@1439.4]
  assign active_1_io_input_set = _T_205 & _T_208; // @[Controllers.scala 165:32:@1580.4]
  assign active_1_io_input_reset = io_ctrCopyDone_1 | io_parentAck; // @[Controllers.scala 166:34:@1584.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@1450.4]
  assign done_0_clock = clock; // @[:@1441.4]
  assign done_0_reset = reset; // @[:@1442.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_183; // @[Controllers.scala 169:30:@1561.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@1461.4 Controllers.scala 170:32:@1568.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@1451.4]
  assign done_1_clock = clock; // @[:@1444.4]
  assign done_1_reset = reset; // @[:@1445.4]
  assign done_1_io_input_set = io_ctrCopyDone_1 | _T_251; // @[Controllers.scala 169:30:@1630.4]
  assign done_1_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@1470.4 Controllers.scala 170:32:@1637.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@1452.4]
  assign iterDone_0_clock = clock; // @[:@1473.4]
  assign iterDone_0_reset = reset; // @[:@1474.4]
  assign iterDone_0_io_input_set = _T_153 & io_enable; // @[Controllers.scala 167:34:@1529.4]
  assign iterDone_0_io_input_reset = _T_160 | io_parentAck; // @[Controllers.scala 92:37:@1488.4 Controllers.scala 168:36:@1545.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@1478.4]
  assign iterDone_1_clock = clock; // @[:@1476.4]
  assign iterDone_1_reset = reset; // @[:@1477.4]
  assign iterDone_1_io_input_set = _T_221 & io_enable; // @[Controllers.scala 167:34:@1598.4]
  assign iterDone_1_io_input_reset = _T_228 | io_parentAck; // @[Controllers.scala 92:37:@1497.4 Controllers.scala 168:36:@1614.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@1479.4]
  assign RetimeWrapper_clock = clock; // @[:@1517.4]
  assign RetimeWrapper_reset = reset; // @[:@1518.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@1520.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@1519.4]
  assign RetimeWrapper_1_clock = clock; // @[:@1531.4]
  assign RetimeWrapper_1_reset = reset; // @[:@1532.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@1534.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@1533.4]
  assign RetimeWrapper_2_clock = clock; // @[:@1549.4]
  assign RetimeWrapper_2_reset = reset; // @[:@1550.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@1552.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@1551.4]
  assign RetimeWrapper_3_clock = clock; // @[:@1586.4]
  assign RetimeWrapper_3_reset = reset; // @[:@1587.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@1589.4]
  assign RetimeWrapper_3_io_in = 1'h1; // @[package.scala 94:16:@1588.4]
  assign RetimeWrapper_4_clock = clock; // @[:@1600.4]
  assign RetimeWrapper_4_reset = reset; // @[:@1601.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@1603.4]
  assign RetimeWrapper_4_io_in = io_doneIn_1; // @[package.scala 94:16:@1602.4]
  assign RetimeWrapper_5_clock = clock; // @[:@1618.4]
  assign RetimeWrapper_5_reset = reset; // @[:@1619.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@1621.4]
  assign RetimeWrapper_5_io_in = 1'h1; // @[package.scala 94:16:@1620.4]
  assign RetimeWrapper_6_clock = clock; // @[:@1665.4]
  assign RetimeWrapper_6_reset = reset; // @[:@1666.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@1668.4]
  assign RetimeWrapper_6_io_in = _T_286 | io_parentAck; // @[package.scala 94:16:@1667.4]
  assign RetimeWrapper_7_clock = clock; // @[:@1682.4]
  assign RetimeWrapper_7_reset = reset; // @[:@1683.4]
  assign RetimeWrapper_7_io_flow = io_enable; // @[package.scala 95:18:@1685.4]
  assign RetimeWrapper_7_io_in = allDone & _T_299; // @[package.scala 94:16:@1684.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_285 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_299 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_285 <= 1'h0;
    end else begin
      _T_285 <= _T_282;
    end
    if (reset) begin
      _T_299 <= 1'h0;
    end else begin
      _T_299 <= _T_282;
    end
  end
endmodule
module CompactingIncDincCtr( // @[:@1917.2]
  input   clock, // @[:@1918.4]
  input   reset, // @[:@1919.4]
  input   io_input_inc_en_0, // @[:@1920.4]
  input   io_input_dinc_en_0, // @[:@1920.4]
  output  io_output_full // @[:@1920.4]
);
  reg [31:0] cnt; // @[Counter.scala 170:20:@1922.4]
  reg [31:0] _RAND_0;
  wire [14:0] numPushed; // @[Counter.scala 172:47:@1923.4]
  wire [14:0] numPopped; // @[Counter.scala 173:48:@1924.4]
  wire [31:0] _GEN_0; // @[Counter.scala 174:14:@1925.4]
  wire [32:0] _T_37; // @[Counter.scala 174:14:@1925.4]
  wire [31:0] _T_38; // @[Counter.scala 174:14:@1926.4]
  wire [31:0] _T_39; // @[Counter.scala 174:14:@1927.4]
  wire [31:0] _GEN_1; // @[Counter.scala 174:26:@1928.4]
  wire [32:0] _T_40; // @[Counter.scala 174:26:@1928.4]
  wire [31:0] _T_41; // @[Counter.scala 174:26:@1929.4]
  wire [31:0] _T_42; // @[Counter.scala 174:26:@1930.4]
  assign numPushed = io_input_inc_en_0 ? $signed(15'sh1) : $signed(15'sh0); // @[Counter.scala 172:47:@1923.4]
  assign numPopped = io_input_dinc_en_0 ? $signed(15'sh1) : $signed(15'sh0); // @[Counter.scala 173:48:@1924.4]
  assign _GEN_0 = {{17{numPushed[14]}},numPushed}; // @[Counter.scala 174:14:@1925.4]
  assign _T_37 = $signed(cnt) + $signed(_GEN_0); // @[Counter.scala 174:14:@1925.4]
  assign _T_38 = $signed(cnt) + $signed(_GEN_0); // @[Counter.scala 174:14:@1926.4]
  assign _T_39 = $signed(_T_38); // @[Counter.scala 174:14:@1927.4]
  assign _GEN_1 = {{17{numPopped[14]}},numPopped}; // @[Counter.scala 174:26:@1928.4]
  assign _T_40 = $signed(_T_39) - $signed(_GEN_1); // @[Counter.scala 174:26:@1928.4]
  assign _T_41 = $signed(_T_39) - $signed(_GEN_1); // @[Counter.scala 174:26:@1929.4]
  assign _T_42 = $signed(_T_41); // @[Counter.scala 174:26:@1930.4]
  assign io_output_full = $signed(cnt) > $signed(32'sh1dff); // @[Counter.scala 180:18:@1944.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 32'sh0;
    end else begin
      cnt <= _T_42;
    end
  end
endmodule
module x483_fifoinraw_0( // @[:@2067.2]
  input   clock, // @[:@2068.4]
  input   reset // @[:@2069.4]
);
  wire  elements_clock; // @[MemPrimitives.scala 382:24:@2114.4]
  wire  elements_reset; // @[MemPrimitives.scala 382:24:@2114.4]
  wire  elements_io_input_inc_en_0; // @[MemPrimitives.scala 382:24:@2114.4]
  wire  elements_io_input_dinc_en_0; // @[MemPrimitives.scala 382:24:@2114.4]
  wire  elements_io_output_full; // @[MemPrimitives.scala 382:24:@2114.4]
  CompactingIncDincCtr elements ( // @[MemPrimitives.scala 382:24:@2114.4]
    .clock(elements_clock),
    .reset(elements_reset),
    .io_input_inc_en_0(elements_io_input_inc_en_0),
    .io_input_dinc_en_0(elements_io_input_dinc_en_0),
    .io_output_full(elements_io_output_full)
  );
  assign elements_clock = clock; // @[:@2115.4]
  assign elements_reset = reset; // @[:@2116.4]
  assign elements_io_input_inc_en_0 = 1'h0; // @[MemPrimitives.scala 384:79:@2126.4]
  assign elements_io_input_dinc_en_0 = 1'h0; // @[MemPrimitives.scala 385:80:@2127.4]
endmodule
module x484_fifoinpacked_0( // @[:@2490.2]
  input   clock, // @[:@2491.4]
  input   reset, // @[:@2492.4]
  input   io_wPort_0_en_0, // @[:@2493.4]
  output  io_full, // @[:@2493.4]
  input   io_active_0_in, // @[:@2493.4]
  output  io_active_0_out // @[:@2493.4]
);
  wire  elements_clock; // @[MemPrimitives.scala 382:24:@2537.4]
  wire  elements_reset; // @[MemPrimitives.scala 382:24:@2537.4]
  wire  elements_io_input_inc_en_0; // @[MemPrimitives.scala 382:24:@2537.4]
  wire  elements_io_input_dinc_en_0; // @[MemPrimitives.scala 382:24:@2537.4]
  wire  elements_io_output_full; // @[MemPrimitives.scala 382:24:@2537.4]
  CompactingIncDincCtr elements ( // @[MemPrimitives.scala 382:24:@2537.4]
    .clock(elements_clock),
    .reset(elements_reset),
    .io_input_inc_en_0(elements_io_input_inc_en_0),
    .io_input_dinc_en_0(elements_io_input_dinc_en_0),
    .io_output_full(elements_io_output_full)
  );
  assign io_full = elements_io_output_full; // @[MemPrimitives.scala 429:39:@2611.4]
  assign io_active_0_out = io_active_0_in; // @[MemPrimitives.scala 427:129:@2609.4]
  assign elements_clock = clock; // @[:@2538.4]
  assign elements_reset = reset; // @[:@2539.4]
  assign elements_io_input_inc_en_0 = io_wPort_0_en_0; // @[MemPrimitives.scala 384:79:@2549.4]
  assign elements_io_input_dinc_en_0 = 1'h0; // @[MemPrimitives.scala 385:80:@2550.4]
endmodule
module FF_7( // @[:@3040.2]
  input         clock, // @[:@3041.4]
  input         reset, // @[:@3042.4]
  output [12:0] io_rPort_0_output_0, // @[:@3043.4]
  input  [12:0] io_wPort_0_data_0, // @[:@3043.4]
  input         io_wPort_0_reset, // @[:@3043.4]
  input         io_wPort_0_en_0 // @[:@3043.4]
);
  reg [12:0] ff; // @[MemPrimitives.scala 311:19:@3058.4]
  reg [31:0] _RAND_0;
  wire [12:0] _T_68; // @[MemPrimitives.scala 315:32:@3060.4]
  wire [12:0] _T_69; // @[MemPrimitives.scala 315:12:@3061.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 315:32:@3060.4]
  assign _T_69 = io_wPort_0_reset ? 13'h0 : _T_68; // @[MemPrimitives.scala 315:12:@3061.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 316:34:@3063.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[12:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 13'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 13'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SingleCounter_1( // @[:@3078.2]
  input         clock, // @[:@3079.4]
  input         reset, // @[:@3080.4]
  input         io_setup_saturate, // @[:@3081.4]
  input         io_input_reset, // @[:@3081.4]
  input         io_input_enable, // @[:@3081.4]
  output [12:0] io_output_count_0, // @[:@3081.4]
  output        io_output_oobs_0, // @[:@3081.4]
  output        io_output_done, // @[:@3081.4]
  output        io_output_saturated // @[:@3081.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@3094.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@3094.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@3094.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@3094.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@3094.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@3094.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@3110.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@3110.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@3110.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@3110.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@3110.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@3110.4]
  wire  _T_36; // @[Counter.scala 264:45:@3113.4]
  wire [12:0] _T_48; // @[Counter.scala 287:52:@3138.4]
  wire [13:0] _T_50; // @[Counter.scala 291:33:@3139.4]
  wire [12:0] _T_51; // @[Counter.scala 291:33:@3140.4]
  wire [12:0] _T_52; // @[Counter.scala 291:33:@3141.4]
  wire  _T_57; // @[Counter.scala 293:18:@3143.4]
  wire [12:0] _T_68; // @[Counter.scala 299:115:@3151.4]
  wire [12:0] _T_70; // @[Counter.scala 299:85:@3153.4]
  wire [12:0] _T_71; // @[Counter.scala 299:152:@3154.4]
  wire [12:0] _T_72; // @[Counter.scala 299:74:@3155.4]
  wire  _T_75; // @[Counter.scala 322:102:@3159.4]
  wire  _T_77; // @[Counter.scala 322:130:@3160.4]
  FF_7 bases_0 ( // @[Counter.scala 261:53:@3094.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@3110.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@3113.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@3138.4]
  assign _T_50 = $signed(_T_48) + $signed(13'sh1); // @[Counter.scala 291:33:@3139.4]
  assign _T_51 = $signed(_T_48) + $signed(13'sh1); // @[Counter.scala 291:33:@3140.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@3141.4]
  assign _T_57 = $signed(_T_52) >= $signed(13'sh438); // @[Counter.scala 293:18:@3143.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@3151.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 13'h0; // @[Counter.scala 299:85:@3153.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@3154.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 299:74:@3155.4]
  assign _T_75 = $signed(_T_48) < $signed(13'sh0); // @[Counter.scala 322:102:@3159.4]
  assign _T_77 = $signed(_T_48) >= $signed(13'sh438); // @[Counter.scala 322:130:@3160.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@3158.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@3162.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@3164.4]
  assign io_output_saturated = io_setup_saturate & _T_57; // @[Counter.scala 340:25:@3167.4]
  assign bases_0_clock = clock; // @[:@3095.4]
  assign bases_0_reset = reset; // @[:@3096.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 13'h0 : _T_72; // @[Counter.scala 299:31:@3157.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@3136.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@3137.4]
  assign SRFF_clock = clock; // @[:@3111.4]
  assign SRFF_reset = reset; // @[:@3112.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@3115.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@3117.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@3118.4]
endmodule
module SingleCounter_2( // @[:@3207.2]
  input         clock, // @[:@3208.4]
  input         reset, // @[:@3209.4]
  input         io_setup_saturate, // @[:@3210.4]
  input         io_input_reset, // @[:@3210.4]
  input         io_input_enable, // @[:@3210.4]
  output [12:0] io_output_count_0, // @[:@3210.4]
  output        io_output_oobs_0, // @[:@3210.4]
  output        io_output_done // @[:@3210.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@3223.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@3223.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@3223.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@3223.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@3223.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@3223.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@3239.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@3239.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@3239.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@3239.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@3239.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@3239.4]
  wire  _T_36; // @[Counter.scala 264:45:@3242.4]
  wire [12:0] _T_48; // @[Counter.scala 287:52:@3267.4]
  wire [13:0] _T_50; // @[Counter.scala 291:33:@3268.4]
  wire [12:0] _T_51; // @[Counter.scala 291:33:@3269.4]
  wire [12:0] _T_52; // @[Counter.scala 291:33:@3270.4]
  wire  _T_57; // @[Counter.scala 293:18:@3272.4]
  wire [12:0] _T_68; // @[Counter.scala 299:115:@3280.4]
  wire [12:0] _T_70; // @[Counter.scala 299:85:@3282.4]
  wire [12:0] _T_71; // @[Counter.scala 299:152:@3283.4]
  wire [12:0] _T_72; // @[Counter.scala 299:74:@3284.4]
  wire  _T_75; // @[Counter.scala 322:102:@3288.4]
  wire  _T_77; // @[Counter.scala 322:130:@3289.4]
  FF_7 bases_0 ( // @[Counter.scala 261:53:@3223.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@3239.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@3242.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@3267.4]
  assign _T_50 = $signed(_T_48) + $signed(13'sh4); // @[Counter.scala 291:33:@3268.4]
  assign _T_51 = $signed(_T_48) + $signed(13'sh4); // @[Counter.scala 291:33:@3269.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@3270.4]
  assign _T_57 = $signed(_T_52) >= $signed(13'sh780); // @[Counter.scala 293:18:@3272.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@3280.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 13'h0; // @[Counter.scala 299:85:@3282.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@3283.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 299:74:@3284.4]
  assign _T_75 = $signed(_T_48) < $signed(13'sh0); // @[Counter.scala 322:102:@3288.4]
  assign _T_77 = $signed(_T_48) >= $signed(13'sh780); // @[Counter.scala 322:130:@3289.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@3287.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@3291.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@3293.4]
  assign bases_0_clock = clock; // @[:@3224.4]
  assign bases_0_reset = reset; // @[:@3225.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 13'h0 : _T_72; // @[Counter.scala 299:31:@3286.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@3265.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@3266.4]
  assign SRFF_clock = clock; // @[:@3240.4]
  assign SRFF_reset = reset; // @[:@3241.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@3244.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@3246.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@3247.4]
endmodule
module x488_ctrchain( // @[:@3298.2]
  input         clock, // @[:@3299.4]
  input         reset, // @[:@3300.4]
  input         io_input_reset, // @[:@3301.4]
  input         io_input_enable, // @[:@3301.4]
  output [12:0] io_output_counts_1, // @[:@3301.4]
  output [12:0] io_output_counts_0, // @[:@3301.4]
  output        io_output_oobs_0, // @[:@3301.4]
  output        io_output_oobs_1, // @[:@3301.4]
  output        io_output_done // @[:@3301.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 513:46:@3303.4]
  wire  ctrs_0_reset; // @[Counter.scala 513:46:@3303.4]
  wire  ctrs_0_io_setup_saturate; // @[Counter.scala 513:46:@3303.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 513:46:@3303.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 513:46:@3303.4]
  wire [12:0] ctrs_0_io_output_count_0; // @[Counter.scala 513:46:@3303.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 513:46:@3303.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 513:46:@3303.4]
  wire  ctrs_0_io_output_saturated; // @[Counter.scala 513:46:@3303.4]
  wire  ctrs_1_clock; // @[Counter.scala 513:46:@3306.4]
  wire  ctrs_1_reset; // @[Counter.scala 513:46:@3306.4]
  wire  ctrs_1_io_setup_saturate; // @[Counter.scala 513:46:@3306.4]
  wire  ctrs_1_io_input_reset; // @[Counter.scala 513:46:@3306.4]
  wire  ctrs_1_io_input_enable; // @[Counter.scala 513:46:@3306.4]
  wire [12:0] ctrs_1_io_output_count_0; // @[Counter.scala 513:46:@3306.4]
  wire  ctrs_1_io_output_oobs_0; // @[Counter.scala 513:46:@3306.4]
  wire  ctrs_1_io_output_done; // @[Counter.scala 513:46:@3306.4]
  wire  isDone; // @[Counter.scala 541:51:@3323.4]
  reg  wasDone; // @[Counter.scala 542:24:@3324.4]
  reg [31:0] _RAND_0;
  wire  _T_64; // @[Counter.scala 546:69:@3332.4]
  wire  _T_66; // @[Counter.scala 546:80:@3333.4]
  reg  doneLatch; // @[Counter.scala 550:26:@3338.4]
  reg [31:0] _RAND_1;
  wire  _T_73; // @[Counter.scala 551:48:@3339.4]
  wire  _T_74; // @[Counter.scala 551:19:@3340.4]
  SingleCounter_1 ctrs_0 ( // @[Counter.scala 513:46:@3303.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_setup_saturate(ctrs_0_io_setup_saturate),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done),
    .io_output_saturated(ctrs_0_io_output_saturated)
  );
  SingleCounter_2 ctrs_1 ( // @[Counter.scala 513:46:@3306.4]
    .clock(ctrs_1_clock),
    .reset(ctrs_1_reset),
    .io_setup_saturate(ctrs_1_io_setup_saturate),
    .io_input_reset(ctrs_1_io_input_reset),
    .io_input_enable(ctrs_1_io_input_enable),
    .io_output_count_0(ctrs_1_io_output_count_0),
    .io_output_oobs_0(ctrs_1_io_output_oobs_0),
    .io_output_done(ctrs_1_io_output_done)
  );
  assign isDone = ctrs_0_io_output_done & ctrs_1_io_output_done; // @[Counter.scala 541:51:@3323.4]
  assign _T_64 = io_input_enable & isDone; // @[Counter.scala 546:69:@3332.4]
  assign _T_66 = wasDone == 1'h0; // @[Counter.scala 546:80:@3333.4]
  assign _T_73 = isDone ? 1'h1 : doneLatch; // @[Counter.scala 551:48:@3339.4]
  assign _T_74 = io_input_reset ? 1'h0 : _T_73; // @[Counter.scala 551:19:@3340.4]
  assign io_output_counts_1 = ctrs_1_io_output_count_0; // @[Counter.scala 557:32:@3345.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 557:32:@3342.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@3344.4]
  assign io_output_oobs_1 = ctrs_1_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@3347.4]
  assign io_output_done = _T_64 & _T_66; // @[Counter.scala 546:18:@3335.4]
  assign ctrs_0_clock = clock; // @[:@3304.4]
  assign ctrs_0_reset = reset; // @[:@3305.4]
  assign ctrs_0_io_setup_saturate = 1'h1; // @[Counter.scala 530:29:@3320.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@3312.4]
  assign ctrs_0_io_input_enable = ctrs_1_io_output_done & io_input_enable; // @[Counter.scala 526:29:@3319.4]
  assign ctrs_1_clock = clock; // @[:@3307.4]
  assign ctrs_1_reset = reset; // @[:@3308.4]
  assign ctrs_1_io_setup_saturate = ctrs_0_io_output_saturated; // @[Counter.scala 532:31:@3322.4]
  assign ctrs_1_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@3316.4]
  assign ctrs_1_io_input_enable = io_input_enable; // @[Counter.scala 524:33:@3317.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= isDone;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (isDone) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module RetimeWrapper_21( // @[:@3387.2]
  input   clock, // @[:@3388.4]
  input   reset, // @[:@3389.4]
  input   io_flow, // @[:@3390.4]
  input   io_in, // @[:@3390.4]
  output  io_out // @[:@3390.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3392.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3392.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3392.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3392.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3392.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3392.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(5)) sr ( // @[RetimeShiftRegister.scala 15:20:@3392.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3405.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3404.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3403.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3402.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3401.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3399.4]
endmodule
module RetimeWrapper_25( // @[:@3515.2]
  input   clock, // @[:@3516.4]
  input   reset, // @[:@3517.4]
  input   io_flow, // @[:@3518.4]
  input   io_in, // @[:@3518.4]
  output  io_out // @[:@3518.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3520.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3520.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3520.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3520.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3520.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3520.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(4)) sr ( // @[RetimeShiftRegister.scala 15:20:@3520.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3533.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3532.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3531.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3530.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3529.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3527.4]
endmodule
module x514_inr_Foreach_sm( // @[:@3535.2]
  input   clock, // @[:@3536.4]
  input   reset, // @[:@3537.4]
  input   io_enable, // @[:@3538.4]
  output  io_done, // @[:@3538.4]
  output  io_doneLatch, // @[:@3538.4]
  input   io_ctrDone, // @[:@3538.4]
  output  io_datapathEn, // @[:@3538.4]
  output  io_ctrInc, // @[:@3538.4]
  output  io_ctrRst, // @[:@3538.4]
  input   io_parentAck, // @[:@3538.4]
  input   io_backpressure, // @[:@3538.4]
  input   io_break // @[:@3538.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@3540.4]
  wire  active_reset; // @[Controllers.scala 261:22:@3540.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@3540.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@3540.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@3540.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@3540.4]
  wire  done_clock; // @[Controllers.scala 262:20:@3543.4]
  wire  done_reset; // @[Controllers.scala 262:20:@3543.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@3543.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@3543.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@3543.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@3543.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3577.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3577.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3577.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@3577.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@3577.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@3599.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@3599.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@3599.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@3599.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@3599.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@3611.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@3611.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@3611.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@3611.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@3611.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@3619.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@3619.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@3619.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@3619.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@3619.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@3635.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@3635.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@3635.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@3635.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@3635.4]
  wire  _T_80; // @[Controllers.scala 264:48:@3548.4]
  wire  _T_81; // @[Controllers.scala 264:46:@3549.4]
  wire  _T_82; // @[Controllers.scala 264:62:@3550.4]
  wire  _T_83; // @[Controllers.scala 264:60:@3551.4]
  wire  _T_100; // @[package.scala 100:49:@3568.4]
  reg  _T_103; // @[package.scala 48:56:@3569.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@3582.4 package.scala 96:25:@3583.4]
  wire  _T_110; // @[package.scala 100:49:@3584.4]
  reg  _T_113; // @[package.scala 48:56:@3585.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@3587.4]
  wire  _T_118; // @[Controllers.scala 283:41:@3592.4]
  wire  _T_119; // @[Controllers.scala 283:59:@3593.4]
  wire  _T_121; // @[Controllers.scala 284:37:@3596.4]
  wire  _T_124; // @[package.scala 96:25:@3604.4 package.scala 96:25:@3605.4]
  wire  _T_126; // @[package.scala 100:49:@3606.4]
  reg  _T_129; // @[package.scala 48:56:@3607.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@3629.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@3631.4]
  reg  _T_153; // @[package.scala 48:56:@3632.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@3640.4 package.scala 96:25:@3641.4]
  wire  _T_158; // @[Controllers.scala 292:61:@3642.4]
  wire  _T_159; // @[Controllers.scala 292:24:@3643.4]
  SRFF active ( // @[Controllers.scala 261:22:@3540.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@3543.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_21 RetimeWrapper ( // @[package.scala 93:22:@3577.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_1 ( // @[package.scala 93:22:@3599.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@3611.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@3619.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_4 ( // @[package.scala 93:22:@3635.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@3548.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@3549.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@3550.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@3551.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@3568.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@3582.4 package.scala 96:25:@3583.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@3584.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@3587.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@3592.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@3593.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@3596.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@3604.4 package.scala 96:25:@3605.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@3606.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@3631.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@3640.4 package.scala 96:25:@3641.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@3642.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@3643.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@3610.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@3645.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@3595.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@3598.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@3590.4]
  assign active_clock = clock; // @[:@3541.4]
  assign active_reset = reset; // @[:@3542.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@3553.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@3557.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@3558.4]
  assign done_clock = clock; // @[:@3544.4]
  assign done_reset = reset; // @[:@3545.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@3573.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@3566.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@3567.4]
  assign RetimeWrapper_clock = clock; // @[:@3578.4]
  assign RetimeWrapper_reset = reset; // @[:@3579.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@3581.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@3580.4]
  assign RetimeWrapper_1_clock = clock; // @[:@3600.4]
  assign RetimeWrapper_1_reset = reset; // @[:@3601.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@3603.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@3602.4]
  assign RetimeWrapper_2_clock = clock; // @[:@3612.4]
  assign RetimeWrapper_2_reset = reset; // @[:@3613.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@3615.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@3614.4]
  assign RetimeWrapper_3_clock = clock; // @[:@3620.4]
  assign RetimeWrapper_3_reset = reset; // @[:@3621.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@3623.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@3622.4]
  assign RetimeWrapper_4_clock = clock; // @[:@3636.4]
  assign RetimeWrapper_4_reset = reset; // @[:@3637.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@3639.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@3638.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module SimBlackBoxesfix2fixBox( // @[:@3752.2]
  input  [31:0] io_a, // @[:@3755.4]
  output [31:0] io_b // @[:@3755.4]
);
  assign io_b = io_a; // @[SimBlackBoxes.scala 99:40:@3768.4]
endmodule
module _( // @[:@3770.2]
  input  [31:0] io_b, // @[:@3773.4]
  output [31:0] io_result // @[:@3773.4]
);
  wire [31:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@3778.4]
  wire [31:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@3778.4]
  SimBlackBoxesfix2fixBox SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@3778.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@3791.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@3786.4]
endmodule
module SimBlackBoxesfix2fixBox_2( // @[:@3834.2]
  input  [31:0] io_a, // @[:@3837.4]
  output [32:0] io_b // @[:@3837.4]
);
  wire  _T_20; // @[implicits.scala 69:16:@3847.4]
  assign _T_20 = io_a[31]; // @[implicits.scala 69:16:@3847.4]
  assign io_b = {_T_20,io_a}; // @[SimBlackBoxes.scala 99:40:@3852.4]
endmodule
module __2( // @[:@3854.2]
  input  [31:0] io_b, // @[:@3857.4]
  output [32:0] io_result // @[:@3857.4]
);
  wire [31:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@3862.4]
  wire [32:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@3862.4]
  SimBlackBoxesfix2fixBox_2 SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@3862.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@3875.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@3870.4]
endmodule
module RetimeWrapper_29( // @[:@3932.2]
  input         clock, // @[:@3933.4]
  input         reset, // @[:@3934.4]
  input         io_flow, // @[:@3935.4]
  input  [31:0] io_in, // @[:@3935.4]
  output [31:0] io_out // @[:@3935.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@3937.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@3937.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@3937.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3937.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3937.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3937.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@3937.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3950.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3949.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@3948.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3947.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3946.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3944.4]
endmodule
module fix2fixBox( // @[:@3952.2]
  input         clock, // @[:@3953.4]
  input         reset, // @[:@3954.4]
  input  [32:0] io_a, // @[:@3955.4]
  input         io_flow, // @[:@3955.4]
  output [31:0] io_b // @[:@3955.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3968.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3968.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3968.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@3968.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@3968.4]
  RetimeWrapper_29 RetimeWrapper ( // @[package.scala 93:22:@3968.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@3975.4]
  assign RetimeWrapper_clock = clock; // @[:@3969.4]
  assign RetimeWrapper_reset = reset; // @[:@3970.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@3972.4]
  assign RetimeWrapper_io_in = io_a[31:0]; // @[package.scala 94:16:@3971.4]
endmodule
module x787_sub( // @[:@3977.2]
  input         clock, // @[:@3978.4]
  input         reset, // @[:@3979.4]
  input  [31:0] io_a, // @[:@3980.4]
  input  [31:0] io_b, // @[:@3980.4]
  input         io_flow, // @[:@3980.4]
  output [31:0] io_result // @[:@3980.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@3988.4]
  wire [32:0] __io_result; // @[Math.scala 709:24:@3988.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@3995.4]
  wire [32:0] __1_io_result; // @[Math.scala 709:24:@3995.4]
  wire  fix2fixBox_clock; // @[Math.scala 182:30:@4014.4]
  wire  fix2fixBox_reset; // @[Math.scala 182:30:@4014.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 182:30:@4014.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 182:30:@4014.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 182:30:@4014.4]
  wire [32:0] a_upcast_number; // @[Math.scala 712:22:@3993.4 Math.scala 713:14:@3994.4]
  wire [32:0] b_upcast_number; // @[Math.scala 712:22:@4000.4 Math.scala 713:14:@4001.4]
  wire [33:0] _T_21; // @[Math.scala 177:37:@4002.4]
  wire [33:0] _T_22; // @[Math.scala 177:37:@4003.4]
  __2 _ ( // @[Math.scala 709:24:@3988.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 709:24:@3995.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox fix2fixBox ( // @[Math.scala 182:30:@4014.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@3993.4 Math.scala 713:14:@3994.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@4000.4 Math.scala 713:14:@4001.4]
  assign _T_21 = a_upcast_number - b_upcast_number; // @[Math.scala 177:37:@4002.4]
  assign _T_22 = $unsigned(_T_21); // @[Math.scala 177:37:@4003.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 188:17:@4022.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@3991.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@3998.4]
  assign fix2fixBox_clock = clock; // @[:@4015.4]
  assign fix2fixBox_reset = reset; // @[:@4016.4]
  assign fix2fixBox_io_a = _T_22[32:0]; // @[Math.scala 183:23:@4017.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 186:26:@4020.4]
endmodule
module x494_sum( // @[:@4199.2]
  input         clock, // @[:@4200.4]
  input         reset, // @[:@4201.4]
  input  [31:0] io_a, // @[:@4202.4]
  input  [31:0] io_b, // @[:@4202.4]
  input         io_flow, // @[:@4202.4]
  output [31:0] io_result // @[:@4202.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@4210.4]
  wire [32:0] __io_result; // @[Math.scala 709:24:@4210.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@4217.4]
  wire [32:0] __1_io_result; // @[Math.scala 709:24:@4217.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@4235.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@4235.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@4235.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@4235.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@4235.4]
  wire [32:0] a_upcast_number; // @[Math.scala 712:22:@4215.4 Math.scala 713:14:@4216.4]
  wire [32:0] b_upcast_number; // @[Math.scala 712:22:@4222.4 Math.scala 713:14:@4223.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@4224.4]
  __2 _ ( // @[Math.scala 709:24:@4210.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 709:24:@4217.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox fix2fixBox ( // @[Math.scala 141:30:@4235.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@4215.4 Math.scala 713:14:@4216.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@4222.4 Math.scala 713:14:@4223.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@4224.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@4243.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@4213.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@4220.4]
  assign fix2fixBox_clock = clock; // @[:@4236.4]
  assign fix2fixBox_reset = reset; // @[:@4237.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@4238.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@4241.4]
endmodule
module x514_inr_Foreach_kernelx514_inr_Foreach_concrete1( // @[:@6017.2]
  input         clock, // @[:@6018.4]
  input         reset, // @[:@6019.4]
  output        io_in_x484_fifoinpacked_0_wPort_0_en_0, // @[:@6020.4]
  input         io_in_x484_fifoinpacked_0_full, // @[:@6020.4]
  output        io_in_x484_fifoinpacked_0_active_0_in, // @[:@6020.4]
  input         io_in_x484_fifoinpacked_0_active_0_out, // @[:@6020.4]
  input         io_sigsIn_backpressure, // @[:@6020.4]
  input         io_sigsIn_datapathEn, // @[:@6020.4]
  input         io_sigsIn_break, // @[:@6020.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_1, // @[:@6020.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@6020.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@6020.4]
  input         io_sigsIn_cchainOutputs_0_oobs_1, // @[:@6020.4]
  input         io_rr // @[:@6020.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@6054.4]
  wire [31:0] __io_result; // @[Math.scala 709:24:@6054.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@6066.4]
  wire [31:0] __1_io_result; // @[Math.scala 709:24:@6066.4]
  wire  x787_sub_1_clock; // @[Math.scala 191:24:@6093.4]
  wire  x787_sub_1_reset; // @[Math.scala 191:24:@6093.4]
  wire [31:0] x787_sub_1_io_a; // @[Math.scala 191:24:@6093.4]
  wire [31:0] x787_sub_1_io_b; // @[Math.scala 191:24:@6093.4]
  wire  x787_sub_1_io_flow; // @[Math.scala 191:24:@6093.4]
  wire [31:0] x787_sub_1_io_result; // @[Math.scala 191:24:@6093.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@6103.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@6103.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@6103.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@6103.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@6103.4]
  wire  x494_sum_1_clock; // @[Math.scala 150:24:@6112.4]
  wire  x494_sum_1_reset; // @[Math.scala 150:24:@6112.4]
  wire [31:0] x494_sum_1_io_a; // @[Math.scala 150:24:@6112.4]
  wire [31:0] x494_sum_1_io_b; // @[Math.scala 150:24:@6112.4]
  wire  x494_sum_1_io_flow; // @[Math.scala 150:24:@6112.4]
  wire [31:0] x494_sum_1_io_result; // @[Math.scala 150:24:@6112.4]
  wire  x495_sum_1_clock; // @[Math.scala 150:24:@6124.4]
  wire  x495_sum_1_reset; // @[Math.scala 150:24:@6124.4]
  wire [31:0] x495_sum_1_io_a; // @[Math.scala 150:24:@6124.4]
  wire [31:0] x495_sum_1_io_b; // @[Math.scala 150:24:@6124.4]
  wire  x495_sum_1_io_flow; // @[Math.scala 150:24:@6124.4]
  wire [31:0] x495_sum_1_io_result; // @[Math.scala 150:24:@6124.4]
  wire  x789_sum_1_clock; // @[Math.scala 150:24:@6139.4]
  wire  x789_sum_1_reset; // @[Math.scala 150:24:@6139.4]
  wire [31:0] x789_sum_1_io_a; // @[Math.scala 150:24:@6139.4]
  wire [31:0] x789_sum_1_io_b; // @[Math.scala 150:24:@6139.4]
  wire  x789_sum_1_io_flow; // @[Math.scala 150:24:@6139.4]
  wire [31:0] x789_sum_1_io_result; // @[Math.scala 150:24:@6139.4]
  wire  x499_sum_1_clock; // @[Math.scala 150:24:@6171.4]
  wire  x499_sum_1_reset; // @[Math.scala 150:24:@6171.4]
  wire [31:0] x499_sum_1_io_a; // @[Math.scala 150:24:@6171.4]
  wire [31:0] x499_sum_1_io_b; // @[Math.scala 150:24:@6171.4]
  wire  x499_sum_1_io_flow; // @[Math.scala 150:24:@6171.4]
  wire [31:0] x499_sum_1_io_result; // @[Math.scala 150:24:@6171.4]
  wire  x792_sum_1_clock; // @[Math.scala 150:24:@6186.4]
  wire  x792_sum_1_reset; // @[Math.scala 150:24:@6186.4]
  wire [31:0] x792_sum_1_io_a; // @[Math.scala 150:24:@6186.4]
  wire [31:0] x792_sum_1_io_b; // @[Math.scala 150:24:@6186.4]
  wire  x792_sum_1_io_flow; // @[Math.scala 150:24:@6186.4]
  wire [31:0] x792_sum_1_io_result; // @[Math.scala 150:24:@6186.4]
  wire  x503_sum_1_clock; // @[Math.scala 150:24:@6218.4]
  wire  x503_sum_1_reset; // @[Math.scala 150:24:@6218.4]
  wire [31:0] x503_sum_1_io_a; // @[Math.scala 150:24:@6218.4]
  wire [31:0] x503_sum_1_io_b; // @[Math.scala 150:24:@6218.4]
  wire  x503_sum_1_io_flow; // @[Math.scala 150:24:@6218.4]
  wire [31:0] x503_sum_1_io_result; // @[Math.scala 150:24:@6218.4]
  wire  x795_sum_1_clock; // @[Math.scala 150:24:@6233.4]
  wire  x795_sum_1_reset; // @[Math.scala 150:24:@6233.4]
  wire [31:0] x795_sum_1_io_a; // @[Math.scala 150:24:@6233.4]
  wire [31:0] x795_sum_1_io_b; // @[Math.scala 150:24:@6233.4]
  wire  x795_sum_1_io_flow; // @[Math.scala 150:24:@6233.4]
  wire [31:0] x795_sum_1_io_result; // @[Math.scala 150:24:@6233.4]
  wire  x507_sum_1_clock; // @[Math.scala 150:24:@6265.4]
  wire  x507_sum_1_reset; // @[Math.scala 150:24:@6265.4]
  wire [31:0] x507_sum_1_io_a; // @[Math.scala 150:24:@6265.4]
  wire [31:0] x507_sum_1_io_b; // @[Math.scala 150:24:@6265.4]
  wire  x507_sum_1_io_flow; // @[Math.scala 150:24:@6265.4]
  wire [31:0] x507_sum_1_io_result; // @[Math.scala 150:24:@6265.4]
  wire  x798_sum_1_clock; // @[Math.scala 150:24:@6280.4]
  wire  x798_sum_1_reset; // @[Math.scala 150:24:@6280.4]
  wire [31:0] x798_sum_1_io_a; // @[Math.scala 150:24:@6280.4]
  wire [31:0] x798_sum_1_io_b; // @[Math.scala 150:24:@6280.4]
  wire  x798_sum_1_io_flow; // @[Math.scala 150:24:@6280.4]
  wire [31:0] x798_sum_1_io_result; // @[Math.scala 150:24:@6280.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@6320.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@6320.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@6320.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@6320.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@6320.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@6329.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@6329.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@6329.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@6329.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@6329.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@6340.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@6340.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@6340.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@6340.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@6340.4]
  wire  _T_327; // @[sm_x514_inr_Foreach.scala 62:18:@6079.4]
  wire  _T_328; // @[sm_x514_inr_Foreach.scala 62:55:@6080.4]
  wire [31:0] b489_number; // @[Math.scala 712:22:@6059.4 Math.scala 713:14:@6060.4]
  wire [42:0] _GEN_0; // @[Math.scala 450:32:@6084.4]
  wire [42:0] _T_332; // @[Math.scala 450:32:@6084.4]
  wire [38:0] _GEN_1; // @[Math.scala 450:32:@6089.4]
  wire [38:0] _T_336; // @[Math.scala 450:32:@6089.4]
  wire [31:0] x495_sum_number; // @[Math.scala 154:22:@6130.4 Math.scala 155:14:@6131.4]
  wire [33:0] _GEN_2; // @[Math.scala 450:32:@6135.4]
  wire [33:0] _T_356; // @[Math.scala 450:32:@6135.4]
  wire [31:0] x499_sum_number; // @[Math.scala 154:22:@6177.4 Math.scala 155:14:@6178.4]
  wire [33:0] _GEN_3; // @[Math.scala 450:32:@6182.4]
  wire [33:0] _T_385; // @[Math.scala 450:32:@6182.4]
  wire [31:0] x503_sum_number; // @[Math.scala 154:22:@6224.4 Math.scala 155:14:@6225.4]
  wire [33:0] _GEN_4; // @[Math.scala 450:32:@6229.4]
  wire [33:0] _T_414; // @[Math.scala 450:32:@6229.4]
  wire [31:0] x507_sum_number; // @[Math.scala 154:22:@6271.4 Math.scala 155:14:@6272.4]
  wire [33:0] _GEN_5; // @[Math.scala 450:32:@6276.4]
  wire [33:0] _T_443; // @[Math.scala 450:32:@6276.4]
  wire  _T_481; // @[sm_x514_inr_Foreach.scala 123:131:@6337.4]
  wire  _T_485; // @[package.scala 96:25:@6345.4 package.scala 96:25:@6346.4]
  wire  _T_487; // @[implicits.scala 55:10:@6347.4]
  wire  _T_488; // @[sm_x514_inr_Foreach.scala 123:148:@6348.4]
  wire  _T_490; // @[sm_x514_inr_Foreach.scala 123:236:@6350.4]
  wire  _T_491; // @[sm_x514_inr_Foreach.scala 123:255:@6351.4]
  wire  x822_b491_D4; // @[package.scala 96:25:@6325.4 package.scala 96:25:@6326.4]
  wire  _T_494; // @[sm_x514_inr_Foreach.scala 123:291:@6353.4]
  wire  x823_b492_D4; // @[package.scala 96:25:@6334.4 package.scala 96:25:@6335.4]
  _ _ ( // @[Math.scala 709:24:@6054.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 709:24:@6066.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  x787_sub x787_sub_1 ( // @[Math.scala 191:24:@6093.4]
    .clock(x787_sub_1_clock),
    .reset(x787_sub_1_reset),
    .io_a(x787_sub_1_io_a),
    .io_b(x787_sub_1_io_b),
    .io_flow(x787_sub_1_io_flow),
    .io_result(x787_sub_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper ( // @[package.scala 93:22:@6103.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x494_sum x494_sum_1 ( // @[Math.scala 150:24:@6112.4]
    .clock(x494_sum_1_clock),
    .reset(x494_sum_1_reset),
    .io_a(x494_sum_1_io_a),
    .io_b(x494_sum_1_io_b),
    .io_flow(x494_sum_1_io_flow),
    .io_result(x494_sum_1_io_result)
  );
  x494_sum x495_sum_1 ( // @[Math.scala 150:24:@6124.4]
    .clock(x495_sum_1_clock),
    .reset(x495_sum_1_reset),
    .io_a(x495_sum_1_io_a),
    .io_b(x495_sum_1_io_b),
    .io_flow(x495_sum_1_io_flow),
    .io_result(x495_sum_1_io_result)
  );
  x494_sum x789_sum_1 ( // @[Math.scala 150:24:@6139.4]
    .clock(x789_sum_1_clock),
    .reset(x789_sum_1_reset),
    .io_a(x789_sum_1_io_a),
    .io_b(x789_sum_1_io_b),
    .io_flow(x789_sum_1_io_flow),
    .io_result(x789_sum_1_io_result)
  );
  x494_sum x499_sum_1 ( // @[Math.scala 150:24:@6171.4]
    .clock(x499_sum_1_clock),
    .reset(x499_sum_1_reset),
    .io_a(x499_sum_1_io_a),
    .io_b(x499_sum_1_io_b),
    .io_flow(x499_sum_1_io_flow),
    .io_result(x499_sum_1_io_result)
  );
  x494_sum x792_sum_1 ( // @[Math.scala 150:24:@6186.4]
    .clock(x792_sum_1_clock),
    .reset(x792_sum_1_reset),
    .io_a(x792_sum_1_io_a),
    .io_b(x792_sum_1_io_b),
    .io_flow(x792_sum_1_io_flow),
    .io_result(x792_sum_1_io_result)
  );
  x494_sum x503_sum_1 ( // @[Math.scala 150:24:@6218.4]
    .clock(x503_sum_1_clock),
    .reset(x503_sum_1_reset),
    .io_a(x503_sum_1_io_a),
    .io_b(x503_sum_1_io_b),
    .io_flow(x503_sum_1_io_flow),
    .io_result(x503_sum_1_io_result)
  );
  x494_sum x795_sum_1 ( // @[Math.scala 150:24:@6233.4]
    .clock(x795_sum_1_clock),
    .reset(x795_sum_1_reset),
    .io_a(x795_sum_1_io_a),
    .io_b(x795_sum_1_io_b),
    .io_flow(x795_sum_1_io_flow),
    .io_result(x795_sum_1_io_result)
  );
  x494_sum x507_sum_1 ( // @[Math.scala 150:24:@6265.4]
    .clock(x507_sum_1_clock),
    .reset(x507_sum_1_reset),
    .io_a(x507_sum_1_io_a),
    .io_b(x507_sum_1_io_b),
    .io_flow(x507_sum_1_io_flow),
    .io_result(x507_sum_1_io_result)
  );
  x494_sum x798_sum_1 ( // @[Math.scala 150:24:@6280.4]
    .clock(x798_sum_1_clock),
    .reset(x798_sum_1_reset),
    .io_a(x798_sum_1_io_a),
    .io_b(x798_sum_1_io_b),
    .io_flow(x798_sum_1_io_flow),
    .io_result(x798_sum_1_io_result)
  );
  RetimeWrapper_25 RetimeWrapper_1 ( // @[package.scala 93:22:@6320.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_2 ( // @[package.scala 93:22:@6329.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_3 ( // @[package.scala 93:22:@6340.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  assign _T_327 = ~ io_in_x484_fifoinpacked_0_full; // @[sm_x514_inr_Foreach.scala 62:18:@6079.4]
  assign _T_328 = ~ io_in_x484_fifoinpacked_0_active_0_out; // @[sm_x514_inr_Foreach.scala 62:55:@6080.4]
  assign b489_number = __io_result; // @[Math.scala 712:22:@6059.4 Math.scala 713:14:@6060.4]
  assign _GEN_0 = {{11'd0}, b489_number}; // @[Math.scala 450:32:@6084.4]
  assign _T_332 = _GEN_0 << 11; // @[Math.scala 450:32:@6084.4]
  assign _GEN_1 = {{7'd0}, b489_number}; // @[Math.scala 450:32:@6089.4]
  assign _T_336 = _GEN_1 << 7; // @[Math.scala 450:32:@6089.4]
  assign x495_sum_number = x495_sum_1_io_result; // @[Math.scala 154:22:@6130.4 Math.scala 155:14:@6131.4]
  assign _GEN_2 = {{2'd0}, x495_sum_number}; // @[Math.scala 450:32:@6135.4]
  assign _T_356 = _GEN_2 << 2; // @[Math.scala 450:32:@6135.4]
  assign x499_sum_number = x499_sum_1_io_result; // @[Math.scala 154:22:@6177.4 Math.scala 155:14:@6178.4]
  assign _GEN_3 = {{2'd0}, x499_sum_number}; // @[Math.scala 450:32:@6182.4]
  assign _T_385 = _GEN_3 << 2; // @[Math.scala 450:32:@6182.4]
  assign x503_sum_number = x503_sum_1_io_result; // @[Math.scala 154:22:@6224.4 Math.scala 155:14:@6225.4]
  assign _GEN_4 = {{2'd0}, x503_sum_number}; // @[Math.scala 450:32:@6229.4]
  assign _T_414 = _GEN_4 << 2; // @[Math.scala 450:32:@6229.4]
  assign x507_sum_number = x507_sum_1_io_result; // @[Math.scala 154:22:@6271.4 Math.scala 155:14:@6272.4]
  assign _GEN_5 = {{2'd0}, x507_sum_number}; // @[Math.scala 450:32:@6276.4]
  assign _T_443 = _GEN_5 << 2; // @[Math.scala 450:32:@6276.4]
  assign _T_481 = ~ io_sigsIn_break; // @[sm_x514_inr_Foreach.scala 123:131:@6337.4]
  assign _T_485 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@6345.4 package.scala 96:25:@6346.4]
  assign _T_487 = io_rr ? _T_485 : 1'h0; // @[implicits.scala 55:10:@6347.4]
  assign _T_488 = _T_481 & _T_487; // @[sm_x514_inr_Foreach.scala 123:148:@6348.4]
  assign _T_490 = _T_488 & _T_481; // @[sm_x514_inr_Foreach.scala 123:236:@6350.4]
  assign _T_491 = _T_490 & io_sigsIn_backpressure; // @[sm_x514_inr_Foreach.scala 123:255:@6351.4]
  assign x822_b491_D4 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@6325.4 package.scala 96:25:@6326.4]
  assign _T_494 = _T_491 & x822_b491_D4; // @[sm_x514_inr_Foreach.scala 123:291:@6353.4]
  assign x823_b492_D4 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@6334.4 package.scala 96:25:@6335.4]
  assign io_in_x484_fifoinpacked_0_wPort_0_en_0 = _T_494 & x823_b492_D4; // @[MemInterfaceType.scala 93:57:@6357.4]
  assign io_in_x484_fifoinpacked_0_active_0_in = x822_b491_D4 & x823_b492_D4; // @[MemInterfaceType.scala 147:18:@6360.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 710:17:@6057.4]
  assign __1_io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_1); // @[Math.scala 710:17:@6069.4]
  assign x787_sub_1_clock = clock; // @[:@6094.4]
  assign x787_sub_1_reset = reset; // @[:@6095.4]
  assign x787_sub_1_io_a = _T_332[31:0]; // @[Math.scala 192:17:@6096.4]
  assign x787_sub_1_io_b = _T_336[31:0]; // @[Math.scala 193:17:@6097.4]
  assign x787_sub_1_io_flow = _T_327 | _T_328; // @[Math.scala 194:20:@6098.4]
  assign RetimeWrapper_clock = clock; // @[:@6104.4]
  assign RetimeWrapper_reset = reset; // @[:@6105.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@6107.4]
  assign RetimeWrapper_io_in = __1_io_result; // @[package.scala 94:16:@6106.4]
  assign x494_sum_1_clock = clock; // @[:@6113.4]
  assign x494_sum_1_reset = reset; // @[:@6114.4]
  assign x494_sum_1_io_a = x787_sub_1_io_result; // @[Math.scala 151:17:@6115.4]
  assign x494_sum_1_io_b = RetimeWrapper_io_out; // @[Math.scala 152:17:@6116.4]
  assign x494_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@6117.4]
  assign x495_sum_1_clock = clock; // @[:@6125.4]
  assign x495_sum_1_reset = reset; // @[:@6126.4]
  assign x495_sum_1_io_a = x494_sum_1_io_result; // @[Math.scala 151:17:@6127.4]
  assign x495_sum_1_io_b = 32'h1; // @[Math.scala 152:17:@6128.4]
  assign x495_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@6129.4]
  assign x789_sum_1_clock = clock; // @[:@6140.4]
  assign x789_sum_1_reset = reset; // @[:@6141.4]
  assign x789_sum_1_io_a = _T_356[31:0]; // @[Math.scala 151:17:@6142.4]
  assign x789_sum_1_io_b = x495_sum_1_io_result; // @[Math.scala 152:17:@6143.4]
  assign x789_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@6144.4]
  assign x499_sum_1_clock = clock; // @[:@6172.4]
  assign x499_sum_1_reset = reset; // @[:@6173.4]
  assign x499_sum_1_io_a = x494_sum_1_io_result; // @[Math.scala 151:17:@6174.4]
  assign x499_sum_1_io_b = 32'h2; // @[Math.scala 152:17:@6175.4]
  assign x499_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@6176.4]
  assign x792_sum_1_clock = clock; // @[:@6187.4]
  assign x792_sum_1_reset = reset; // @[:@6188.4]
  assign x792_sum_1_io_a = _T_385[31:0]; // @[Math.scala 151:17:@6189.4]
  assign x792_sum_1_io_b = x499_sum_1_io_result; // @[Math.scala 152:17:@6190.4]
  assign x792_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@6191.4]
  assign x503_sum_1_clock = clock; // @[:@6219.4]
  assign x503_sum_1_reset = reset; // @[:@6220.4]
  assign x503_sum_1_io_a = x494_sum_1_io_result; // @[Math.scala 151:17:@6221.4]
  assign x503_sum_1_io_b = 32'h3; // @[Math.scala 152:17:@6222.4]
  assign x503_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@6223.4]
  assign x795_sum_1_clock = clock; // @[:@6234.4]
  assign x795_sum_1_reset = reset; // @[:@6235.4]
  assign x795_sum_1_io_a = _T_414[31:0]; // @[Math.scala 151:17:@6236.4]
  assign x795_sum_1_io_b = x503_sum_1_io_result; // @[Math.scala 152:17:@6237.4]
  assign x795_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@6238.4]
  assign x507_sum_1_clock = clock; // @[:@6266.4]
  assign x507_sum_1_reset = reset; // @[:@6267.4]
  assign x507_sum_1_io_a = x494_sum_1_io_result; // @[Math.scala 151:17:@6268.4]
  assign x507_sum_1_io_b = 32'h4; // @[Math.scala 152:17:@6269.4]
  assign x507_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@6270.4]
  assign x798_sum_1_clock = clock; // @[:@6281.4]
  assign x798_sum_1_reset = reset; // @[:@6282.4]
  assign x798_sum_1_io_a = _T_443[31:0]; // @[Math.scala 151:17:@6283.4]
  assign x798_sum_1_io_b = x507_sum_1_io_result; // @[Math.scala 152:17:@6284.4]
  assign x798_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@6285.4]
  assign RetimeWrapper_1_clock = clock; // @[:@6321.4]
  assign RetimeWrapper_1_reset = reset; // @[:@6322.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@6324.4]
  assign RetimeWrapper_1_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@6323.4]
  assign RetimeWrapper_2_clock = clock; // @[:@6330.4]
  assign RetimeWrapper_2_reset = reset; // @[:@6331.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@6333.4]
  assign RetimeWrapper_2_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@6332.4]
  assign RetimeWrapper_3_clock = clock; // @[:@6341.4]
  assign RetimeWrapper_3_reset = reset; // @[:@6342.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@6344.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@6343.4]
endmodule
module RetimeWrapper_48( // @[:@7478.2]
  input   clock, // @[:@7479.4]
  input   reset, // @[:@7480.4]
  input   io_flow, // @[:@7481.4]
  input   io_in, // @[:@7481.4]
  output  io_out // @[:@7481.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@7483.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@7483.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@7483.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@7483.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@7483.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@7483.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(55)) sr ( // @[RetimeShiftRegister.scala 15:20:@7483.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@7496.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@7495.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@7494.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@7493.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@7492.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@7490.4]
endmodule
module RetimeWrapper_52( // @[:@7606.2]
  input   clock, // @[:@7607.4]
  input   reset, // @[:@7608.4]
  input   io_flow, // @[:@7609.4]
  input   io_in, // @[:@7609.4]
  output  io_out // @[:@7609.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@7611.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@7611.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@7611.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@7611.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@7611.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@7611.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(54)) sr ( // @[RetimeShiftRegister.scala 15:20:@7611.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@7624.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@7623.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@7622.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@7621.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@7620.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@7618.4]
endmodule
module x736_inr_Foreach_SAMPLER_BOX_sm( // @[:@7626.2]
  input   clock, // @[:@7627.4]
  input   reset, // @[:@7628.4]
  input   io_enable, // @[:@7629.4]
  output  io_done, // @[:@7629.4]
  output  io_doneLatch, // @[:@7629.4]
  input   io_ctrDone, // @[:@7629.4]
  output  io_datapathEn, // @[:@7629.4]
  output  io_ctrInc, // @[:@7629.4]
  output  io_ctrRst, // @[:@7629.4]
  input   io_parentAck, // @[:@7629.4]
  input   io_backpressure, // @[:@7629.4]
  input   io_break // @[:@7629.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@7631.4]
  wire  active_reset; // @[Controllers.scala 261:22:@7631.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@7631.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@7631.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@7631.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@7631.4]
  wire  done_clock; // @[Controllers.scala 262:20:@7634.4]
  wire  done_reset; // @[Controllers.scala 262:20:@7634.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@7634.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@7634.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@7634.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@7634.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@7668.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@7668.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@7668.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@7668.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@7668.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@7690.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@7690.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@7690.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@7690.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@7690.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@7702.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@7702.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@7702.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@7702.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@7702.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@7710.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@7710.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@7710.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@7710.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@7710.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@7726.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@7726.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@7726.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@7726.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@7726.4]
  wire  _T_80; // @[Controllers.scala 264:48:@7639.4]
  wire  _T_81; // @[Controllers.scala 264:46:@7640.4]
  wire  _T_82; // @[Controllers.scala 264:62:@7641.4]
  wire  _T_83; // @[Controllers.scala 264:60:@7642.4]
  wire  _T_100; // @[package.scala 100:49:@7659.4]
  reg  _T_103; // @[package.scala 48:56:@7660.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@7673.4 package.scala 96:25:@7674.4]
  wire  _T_110; // @[package.scala 100:49:@7675.4]
  reg  _T_113; // @[package.scala 48:56:@7676.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@7678.4]
  wire  _T_118; // @[Controllers.scala 283:41:@7683.4]
  wire  _T_119; // @[Controllers.scala 283:59:@7684.4]
  wire  _T_121; // @[Controllers.scala 284:37:@7687.4]
  wire  _T_124; // @[package.scala 96:25:@7695.4 package.scala 96:25:@7696.4]
  wire  _T_126; // @[package.scala 100:49:@7697.4]
  reg  _T_129; // @[package.scala 48:56:@7698.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@7720.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@7722.4]
  reg  _T_153; // @[package.scala 48:56:@7723.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@7731.4 package.scala 96:25:@7732.4]
  wire  _T_158; // @[Controllers.scala 292:61:@7733.4]
  wire  _T_159; // @[Controllers.scala 292:24:@7734.4]
  SRFF active ( // @[Controllers.scala 261:22:@7631.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@7634.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_48 RetimeWrapper ( // @[package.scala 93:22:@7668.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_48 RetimeWrapper_1 ( // @[package.scala 93:22:@7690.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@7702.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@7710.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_4 ( // @[package.scala 93:22:@7726.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@7639.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@7640.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@7641.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@7642.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@7659.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@7673.4 package.scala 96:25:@7674.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@7675.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@7678.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@7683.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@7684.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@7687.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@7695.4 package.scala 96:25:@7696.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@7697.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@7722.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@7731.4 package.scala 96:25:@7732.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@7733.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@7734.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@7701.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@7736.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@7686.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@7689.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@7681.4]
  assign active_clock = clock; // @[:@7632.4]
  assign active_reset = reset; // @[:@7633.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@7644.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@7648.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@7649.4]
  assign done_clock = clock; // @[:@7635.4]
  assign done_reset = reset; // @[:@7636.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@7664.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@7657.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@7658.4]
  assign RetimeWrapper_clock = clock; // @[:@7669.4]
  assign RetimeWrapper_reset = reset; // @[:@7670.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@7672.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@7671.4]
  assign RetimeWrapper_1_clock = clock; // @[:@7691.4]
  assign RetimeWrapper_1_reset = reset; // @[:@7692.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@7694.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@7693.4]
  assign RetimeWrapper_2_clock = clock; // @[:@7703.4]
  assign RetimeWrapper_2_reset = reset; // @[:@7704.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@7706.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@7705.4]
  assign RetimeWrapper_3_clock = clock; // @[:@7711.4]
  assign RetimeWrapper_3_reset = reset; // @[:@7712.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@7714.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@7713.4]
  assign RetimeWrapper_4_clock = clock; // @[:@7727.4]
  assign RetimeWrapper_4_reset = reset; // @[:@7728.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@7730.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@7729.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module SRAM_1( // @[:@7973.2]
  input        clock, // @[:@7974.4]
  input  [8:0] io_raddr, // @[:@7976.4]
  input        io_wen, // @[:@7976.4]
  input  [8:0] io_waddr, // @[:@7976.4]
  input  [7:0] io_wdata, // @[:@7976.4]
  output [7:0] io_rdata, // @[:@7976.4]
  input        io_backpressure // @[:@7976.4]
);
  wire [7:0] SRAMVerilogSim_rdata; // @[SRAM.scala 185:23:@7978.4]
  wire [7:0] SRAMVerilogSim_wdata; // @[SRAM.scala 185:23:@7978.4]
  wire  SRAMVerilogSim_backpressure; // @[SRAM.scala 185:23:@7978.4]
  wire  SRAMVerilogSim_wen; // @[SRAM.scala 185:23:@7978.4]
  wire  SRAMVerilogSim_waddrEn; // @[SRAM.scala 185:23:@7978.4]
  wire  SRAMVerilogSim_raddrEn; // @[SRAM.scala 185:23:@7978.4]
  wire [8:0] SRAMVerilogSim_waddr; // @[SRAM.scala 185:23:@7978.4]
  wire [8:0] SRAMVerilogSim_raddr; // @[SRAM.scala 185:23:@7978.4]
  wire  SRAMVerilogSim_clk; // @[SRAM.scala 185:23:@7978.4]
  SRAMVerilogSim #(.DWIDTH(8), .WORDS(320), .AWIDTH(9)) SRAMVerilogSim ( // @[SRAM.scala 185:23:@7978.4]
    .rdata(SRAMVerilogSim_rdata),
    .wdata(SRAMVerilogSim_wdata),
    .backpressure(SRAMVerilogSim_backpressure),
    .wen(SRAMVerilogSim_wen),
    .waddrEn(SRAMVerilogSim_waddrEn),
    .raddrEn(SRAMVerilogSim_raddrEn),
    .waddr(SRAMVerilogSim_waddr),
    .raddr(SRAMVerilogSim_raddr),
    .clk(SRAMVerilogSim_clk)
  );
  assign io_rdata = SRAMVerilogSim_rdata; // @[SRAM.scala 195:16:@7998.4]
  assign SRAMVerilogSim_wdata = io_wdata; // @[SRAM.scala 190:20:@7992.4]
  assign SRAMVerilogSim_backpressure = io_backpressure; // @[SRAM.scala 191:27:@7993.4]
  assign SRAMVerilogSim_wen = io_wen; // @[SRAM.scala 188:18:@7990.4]
  assign SRAMVerilogSim_waddrEn = 1'h1; // @[SRAM.scala 193:22:@7995.4]
  assign SRAMVerilogSim_raddrEn = 1'h1; // @[SRAM.scala 192:22:@7994.4]
  assign SRAMVerilogSim_waddr = io_waddr; // @[SRAM.scala 189:20:@7991.4]
  assign SRAMVerilogSim_raddr = io_raddr; // @[SRAM.scala 187:20:@7989.4]
  assign SRAMVerilogSim_clk = clock; // @[SRAM.scala 186:18:@7988.4]
endmodule
module RetimeWrapper_57( // @[:@8012.2]
  input        clock, // @[:@8013.4]
  input        reset, // @[:@8014.4]
  input        io_flow, // @[:@8015.4]
  input  [8:0] io_in, // @[:@8015.4]
  output [8:0] io_out // @[:@8015.4]
);
  wire [8:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@8017.4]
  wire [8:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@8017.4]
  wire [8:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@8017.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@8017.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@8017.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@8017.4]
  RetimeShiftRegister #(.WIDTH(9), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@8017.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@8030.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@8029.4]
  assign sr_init = 9'h0; // @[RetimeShiftRegister.scala 19:16:@8028.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@8027.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@8026.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@8024.4]
endmodule
module Mem1D_5( // @[:@8032.2]
  input        clock, // @[:@8033.4]
  input        reset, // @[:@8034.4]
  input  [8:0] io_r_ofs_0, // @[:@8035.4]
  input        io_r_backpressure, // @[:@8035.4]
  input  [8:0] io_w_ofs_0, // @[:@8035.4]
  input  [7:0] io_w_data_0, // @[:@8035.4]
  input        io_w_en_0, // @[:@8035.4]
  output [7:0] io_output // @[:@8035.4]
);
  wire  SRAM_clock; // @[MemPrimitives.scala 705:21:@8039.4]
  wire [8:0] SRAM_io_raddr; // @[MemPrimitives.scala 705:21:@8039.4]
  wire  SRAM_io_wen; // @[MemPrimitives.scala 705:21:@8039.4]
  wire [8:0] SRAM_io_waddr; // @[MemPrimitives.scala 705:21:@8039.4]
  wire [7:0] SRAM_io_wdata; // @[MemPrimitives.scala 705:21:@8039.4]
  wire [7:0] SRAM_io_rdata; // @[MemPrimitives.scala 705:21:@8039.4]
  wire  SRAM_io_backpressure; // @[MemPrimitives.scala 705:21:@8039.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@8042.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@8042.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@8042.4]
  wire [8:0] RetimeWrapper_io_in; // @[package.scala 93:22:@8042.4]
  wire [8:0] RetimeWrapper_io_out; // @[package.scala 93:22:@8042.4]
  wire  wInBound; // @[MemPrimitives.scala 692:32:@8037.4]
  SRAM_1 SRAM ( // @[MemPrimitives.scala 705:21:@8039.4]
    .clock(SRAM_clock),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata(SRAM_io_wdata),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  RetimeWrapper_57 RetimeWrapper ( // @[package.scala 93:22:@8042.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign wInBound = io_w_ofs_0 <= 9'h140; // @[MemPrimitives.scala 692:32:@8037.4]
  assign io_output = SRAM_io_rdata; // @[MemPrimitives.scala 712:17:@8055.4]
  assign SRAM_clock = clock; // @[:@8040.4]
  assign SRAM_io_raddr = RetimeWrapper_io_out; // @[MemPrimitives.scala 706:37:@8049.4]
  assign SRAM_io_wen = io_w_en_0 & wInBound; // @[MemPrimitives.scala 709:22:@8052.4]
  assign SRAM_io_waddr = io_w_ofs_0; // @[MemPrimitives.scala 708:22:@8050.4]
  assign SRAM_io_wdata = io_w_data_0; // @[MemPrimitives.scala 710:22:@8053.4]
  assign SRAM_io_backpressure = io_r_backpressure; // @[MemPrimitives.scala 711:30:@8054.4]
  assign RetimeWrapper_clock = clock; // @[:@8043.4]
  assign RetimeWrapper_reset = reset; // @[:@8044.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@8046.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@8045.4]
endmodule
module StickySelects_1( // @[:@10357.2]
  input   clock, // @[:@10358.4]
  input   reset, // @[:@10359.4]
  input   io_ins_0, // @[:@10360.4]
  input   io_ins_1, // @[:@10360.4]
  input   io_ins_2, // @[:@10360.4]
  input   io_ins_3, // @[:@10360.4]
  input   io_ins_4, // @[:@10360.4]
  input   io_ins_5, // @[:@10360.4]
  input   io_ins_6, // @[:@10360.4]
  input   io_ins_7, // @[:@10360.4]
  input   io_ins_8, // @[:@10360.4]
  output  io_outs_0, // @[:@10360.4]
  output  io_outs_1, // @[:@10360.4]
  output  io_outs_2, // @[:@10360.4]
  output  io_outs_3, // @[:@10360.4]
  output  io_outs_4, // @[:@10360.4]
  output  io_outs_5, // @[:@10360.4]
  output  io_outs_6, // @[:@10360.4]
  output  io_outs_7, // @[:@10360.4]
  output  io_outs_8 // @[:@10360.4]
);
  reg  _T_19; // @[StickySelects.scala 37:46:@10362.4]
  reg [31:0] _RAND_0;
  reg  _T_22; // @[StickySelects.scala 37:46:@10363.4]
  reg [31:0] _RAND_1;
  reg  _T_25; // @[StickySelects.scala 37:46:@10364.4]
  reg [31:0] _RAND_2;
  reg  _T_28; // @[StickySelects.scala 37:46:@10365.4]
  reg [31:0] _RAND_3;
  reg  _T_31; // @[StickySelects.scala 37:46:@10366.4]
  reg [31:0] _RAND_4;
  reg  _T_34; // @[StickySelects.scala 37:46:@10367.4]
  reg [31:0] _RAND_5;
  reg  _T_37; // @[StickySelects.scala 37:46:@10368.4]
  reg [31:0] _RAND_6;
  reg  _T_40; // @[StickySelects.scala 37:46:@10369.4]
  reg [31:0] _RAND_7;
  reg  _T_43; // @[StickySelects.scala 37:46:@10370.4]
  reg [31:0] _RAND_8;
  wire  _T_44; // @[StickySelects.scala 47:46:@10371.4]
  wire  _T_45; // @[StickySelects.scala 47:46:@10372.4]
  wire  _T_46; // @[StickySelects.scala 47:46:@10373.4]
  wire  _T_47; // @[StickySelects.scala 47:46:@10374.4]
  wire  _T_48; // @[StickySelects.scala 47:46:@10375.4]
  wire  _T_49; // @[StickySelects.scala 47:46:@10376.4]
  wire  _T_50; // @[StickySelects.scala 47:46:@10377.4]
  wire  _T_51; // @[StickySelects.scala 49:53:@10378.4]
  wire  _T_52; // @[StickySelects.scala 49:21:@10379.4]
  wire  _T_53; // @[StickySelects.scala 47:46:@10381.4]
  wire  _T_54; // @[StickySelects.scala 47:46:@10382.4]
  wire  _T_55; // @[StickySelects.scala 47:46:@10383.4]
  wire  _T_56; // @[StickySelects.scala 47:46:@10384.4]
  wire  _T_57; // @[StickySelects.scala 47:46:@10385.4]
  wire  _T_58; // @[StickySelects.scala 47:46:@10386.4]
  wire  _T_59; // @[StickySelects.scala 47:46:@10387.4]
  wire  _T_60; // @[StickySelects.scala 49:53:@10388.4]
  wire  _T_61; // @[StickySelects.scala 49:21:@10389.4]
  wire  _T_62; // @[StickySelects.scala 47:46:@10391.4]
  wire  _T_63; // @[StickySelects.scala 47:46:@10392.4]
  wire  _T_64; // @[StickySelects.scala 47:46:@10393.4]
  wire  _T_65; // @[StickySelects.scala 47:46:@10394.4]
  wire  _T_66; // @[StickySelects.scala 47:46:@10395.4]
  wire  _T_67; // @[StickySelects.scala 47:46:@10396.4]
  wire  _T_68; // @[StickySelects.scala 47:46:@10397.4]
  wire  _T_69; // @[StickySelects.scala 49:53:@10398.4]
  wire  _T_70; // @[StickySelects.scala 49:21:@10399.4]
  wire  _T_72; // @[StickySelects.scala 47:46:@10402.4]
  wire  _T_73; // @[StickySelects.scala 47:46:@10403.4]
  wire  _T_74; // @[StickySelects.scala 47:46:@10404.4]
  wire  _T_75; // @[StickySelects.scala 47:46:@10405.4]
  wire  _T_76; // @[StickySelects.scala 47:46:@10406.4]
  wire  _T_77; // @[StickySelects.scala 47:46:@10407.4]
  wire  _T_78; // @[StickySelects.scala 49:53:@10408.4]
  wire  _T_79; // @[StickySelects.scala 49:21:@10409.4]
  wire  _T_82; // @[StickySelects.scala 47:46:@10413.4]
  wire  _T_83; // @[StickySelects.scala 47:46:@10414.4]
  wire  _T_84; // @[StickySelects.scala 47:46:@10415.4]
  wire  _T_85; // @[StickySelects.scala 47:46:@10416.4]
  wire  _T_86; // @[StickySelects.scala 47:46:@10417.4]
  wire  _T_87; // @[StickySelects.scala 49:53:@10418.4]
  wire  _T_88; // @[StickySelects.scala 49:21:@10419.4]
  wire  _T_92; // @[StickySelects.scala 47:46:@10424.4]
  wire  _T_93; // @[StickySelects.scala 47:46:@10425.4]
  wire  _T_94; // @[StickySelects.scala 47:46:@10426.4]
  wire  _T_95; // @[StickySelects.scala 47:46:@10427.4]
  wire  _T_96; // @[StickySelects.scala 49:53:@10428.4]
  wire  _T_97; // @[StickySelects.scala 49:21:@10429.4]
  wire  _T_102; // @[StickySelects.scala 47:46:@10435.4]
  wire  _T_103; // @[StickySelects.scala 47:46:@10436.4]
  wire  _T_104; // @[StickySelects.scala 47:46:@10437.4]
  wire  _T_105; // @[StickySelects.scala 49:53:@10438.4]
  wire  _T_106; // @[StickySelects.scala 49:21:@10439.4]
  wire  _T_112; // @[StickySelects.scala 47:46:@10446.4]
  wire  _T_113; // @[StickySelects.scala 47:46:@10447.4]
  wire  _T_114; // @[StickySelects.scala 49:53:@10448.4]
  wire  _T_115; // @[StickySelects.scala 49:21:@10449.4]
  wire  _T_122; // @[StickySelects.scala 47:46:@10457.4]
  wire  _T_123; // @[StickySelects.scala 49:53:@10458.4]
  wire  _T_124; // @[StickySelects.scala 49:21:@10459.4]
  assign _T_44 = io_ins_1 | io_ins_2; // @[StickySelects.scala 47:46:@10371.4]
  assign _T_45 = _T_44 | io_ins_3; // @[StickySelects.scala 47:46:@10372.4]
  assign _T_46 = _T_45 | io_ins_4; // @[StickySelects.scala 47:46:@10373.4]
  assign _T_47 = _T_46 | io_ins_5; // @[StickySelects.scala 47:46:@10374.4]
  assign _T_48 = _T_47 | io_ins_6; // @[StickySelects.scala 47:46:@10375.4]
  assign _T_49 = _T_48 | io_ins_7; // @[StickySelects.scala 47:46:@10376.4]
  assign _T_50 = _T_49 | io_ins_8; // @[StickySelects.scala 47:46:@10377.4]
  assign _T_51 = io_ins_0 | _T_19; // @[StickySelects.scala 49:53:@10378.4]
  assign _T_52 = _T_50 ? io_ins_0 : _T_51; // @[StickySelects.scala 49:21:@10379.4]
  assign _T_53 = io_ins_0 | io_ins_2; // @[StickySelects.scala 47:46:@10381.4]
  assign _T_54 = _T_53 | io_ins_3; // @[StickySelects.scala 47:46:@10382.4]
  assign _T_55 = _T_54 | io_ins_4; // @[StickySelects.scala 47:46:@10383.4]
  assign _T_56 = _T_55 | io_ins_5; // @[StickySelects.scala 47:46:@10384.4]
  assign _T_57 = _T_56 | io_ins_6; // @[StickySelects.scala 47:46:@10385.4]
  assign _T_58 = _T_57 | io_ins_7; // @[StickySelects.scala 47:46:@10386.4]
  assign _T_59 = _T_58 | io_ins_8; // @[StickySelects.scala 47:46:@10387.4]
  assign _T_60 = io_ins_1 | _T_22; // @[StickySelects.scala 49:53:@10388.4]
  assign _T_61 = _T_59 ? io_ins_1 : _T_60; // @[StickySelects.scala 49:21:@10389.4]
  assign _T_62 = io_ins_0 | io_ins_1; // @[StickySelects.scala 47:46:@10391.4]
  assign _T_63 = _T_62 | io_ins_3; // @[StickySelects.scala 47:46:@10392.4]
  assign _T_64 = _T_63 | io_ins_4; // @[StickySelects.scala 47:46:@10393.4]
  assign _T_65 = _T_64 | io_ins_5; // @[StickySelects.scala 47:46:@10394.4]
  assign _T_66 = _T_65 | io_ins_6; // @[StickySelects.scala 47:46:@10395.4]
  assign _T_67 = _T_66 | io_ins_7; // @[StickySelects.scala 47:46:@10396.4]
  assign _T_68 = _T_67 | io_ins_8; // @[StickySelects.scala 47:46:@10397.4]
  assign _T_69 = io_ins_2 | _T_25; // @[StickySelects.scala 49:53:@10398.4]
  assign _T_70 = _T_68 ? io_ins_2 : _T_69; // @[StickySelects.scala 49:21:@10399.4]
  assign _T_72 = _T_62 | io_ins_2; // @[StickySelects.scala 47:46:@10402.4]
  assign _T_73 = _T_72 | io_ins_4; // @[StickySelects.scala 47:46:@10403.4]
  assign _T_74 = _T_73 | io_ins_5; // @[StickySelects.scala 47:46:@10404.4]
  assign _T_75 = _T_74 | io_ins_6; // @[StickySelects.scala 47:46:@10405.4]
  assign _T_76 = _T_75 | io_ins_7; // @[StickySelects.scala 47:46:@10406.4]
  assign _T_77 = _T_76 | io_ins_8; // @[StickySelects.scala 47:46:@10407.4]
  assign _T_78 = io_ins_3 | _T_28; // @[StickySelects.scala 49:53:@10408.4]
  assign _T_79 = _T_77 ? io_ins_3 : _T_78; // @[StickySelects.scala 49:21:@10409.4]
  assign _T_82 = _T_72 | io_ins_3; // @[StickySelects.scala 47:46:@10413.4]
  assign _T_83 = _T_82 | io_ins_5; // @[StickySelects.scala 47:46:@10414.4]
  assign _T_84 = _T_83 | io_ins_6; // @[StickySelects.scala 47:46:@10415.4]
  assign _T_85 = _T_84 | io_ins_7; // @[StickySelects.scala 47:46:@10416.4]
  assign _T_86 = _T_85 | io_ins_8; // @[StickySelects.scala 47:46:@10417.4]
  assign _T_87 = io_ins_4 | _T_31; // @[StickySelects.scala 49:53:@10418.4]
  assign _T_88 = _T_86 ? io_ins_4 : _T_87; // @[StickySelects.scala 49:21:@10419.4]
  assign _T_92 = _T_82 | io_ins_4; // @[StickySelects.scala 47:46:@10424.4]
  assign _T_93 = _T_92 | io_ins_6; // @[StickySelects.scala 47:46:@10425.4]
  assign _T_94 = _T_93 | io_ins_7; // @[StickySelects.scala 47:46:@10426.4]
  assign _T_95 = _T_94 | io_ins_8; // @[StickySelects.scala 47:46:@10427.4]
  assign _T_96 = io_ins_5 | _T_34; // @[StickySelects.scala 49:53:@10428.4]
  assign _T_97 = _T_95 ? io_ins_5 : _T_96; // @[StickySelects.scala 49:21:@10429.4]
  assign _T_102 = _T_92 | io_ins_5; // @[StickySelects.scala 47:46:@10435.4]
  assign _T_103 = _T_102 | io_ins_7; // @[StickySelects.scala 47:46:@10436.4]
  assign _T_104 = _T_103 | io_ins_8; // @[StickySelects.scala 47:46:@10437.4]
  assign _T_105 = io_ins_6 | _T_37; // @[StickySelects.scala 49:53:@10438.4]
  assign _T_106 = _T_104 ? io_ins_6 : _T_105; // @[StickySelects.scala 49:21:@10439.4]
  assign _T_112 = _T_102 | io_ins_6; // @[StickySelects.scala 47:46:@10446.4]
  assign _T_113 = _T_112 | io_ins_8; // @[StickySelects.scala 47:46:@10447.4]
  assign _T_114 = io_ins_7 | _T_40; // @[StickySelects.scala 49:53:@10448.4]
  assign _T_115 = _T_113 ? io_ins_7 : _T_114; // @[StickySelects.scala 49:21:@10449.4]
  assign _T_122 = _T_112 | io_ins_7; // @[StickySelects.scala 47:46:@10457.4]
  assign _T_123 = io_ins_8 | _T_43; // @[StickySelects.scala 49:53:@10458.4]
  assign _T_124 = _T_122 ? io_ins_8 : _T_123; // @[StickySelects.scala 49:21:@10459.4]
  assign io_outs_0 = _T_50 ? io_ins_0 : _T_51; // @[StickySelects.scala 53:57:@10461.4]
  assign io_outs_1 = _T_59 ? io_ins_1 : _T_60; // @[StickySelects.scala 53:57:@10462.4]
  assign io_outs_2 = _T_68 ? io_ins_2 : _T_69; // @[StickySelects.scala 53:57:@10463.4]
  assign io_outs_3 = _T_77 ? io_ins_3 : _T_78; // @[StickySelects.scala 53:57:@10464.4]
  assign io_outs_4 = _T_86 ? io_ins_4 : _T_87; // @[StickySelects.scala 53:57:@10465.4]
  assign io_outs_5 = _T_95 ? io_ins_5 : _T_96; // @[StickySelects.scala 53:57:@10466.4]
  assign io_outs_6 = _T_104 ? io_ins_6 : _T_105; // @[StickySelects.scala 53:57:@10467.4]
  assign io_outs_7 = _T_113 ? io_ins_7 : _T_114; // @[StickySelects.scala 53:57:@10468.4]
  assign io_outs_8 = _T_122 ? io_ins_8 : _T_123; // @[StickySelects.scala 53:57:@10469.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_22 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_25 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_28 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_31 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_34 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_37 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_40 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_43 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (_T_50) begin
        _T_19 <= io_ins_0;
      end else begin
        _T_19 <= _T_51;
      end
    end
    if (reset) begin
      _T_22 <= 1'h0;
    end else begin
      if (_T_59) begin
        _T_22 <= io_ins_1;
      end else begin
        _T_22 <= _T_60;
      end
    end
    if (reset) begin
      _T_25 <= 1'h0;
    end else begin
      if (_T_68) begin
        _T_25 <= io_ins_2;
      end else begin
        _T_25 <= _T_69;
      end
    end
    if (reset) begin
      _T_28 <= 1'h0;
    end else begin
      if (_T_77) begin
        _T_28 <= io_ins_3;
      end else begin
        _T_28 <= _T_78;
      end
    end
    if (reset) begin
      _T_31 <= 1'h0;
    end else begin
      if (_T_86) begin
        _T_31 <= io_ins_4;
      end else begin
        _T_31 <= _T_87;
      end
    end
    if (reset) begin
      _T_34 <= 1'h0;
    end else begin
      if (_T_95) begin
        _T_34 <= io_ins_5;
      end else begin
        _T_34 <= _T_96;
      end
    end
    if (reset) begin
      _T_37 <= 1'h0;
    end else begin
      if (_T_104) begin
        _T_37 <= io_ins_6;
      end else begin
        _T_37 <= _T_105;
      end
    end
    if (reset) begin
      _T_40 <= 1'h0;
    end else begin
      if (_T_113) begin
        _T_40 <= io_ins_7;
      end else begin
        _T_40 <= _T_114;
      end
    end
    if (reset) begin
      _T_43 <= 1'h0;
    end else begin
      if (_T_122) begin
        _T_43 <= io_ins_8;
      end else begin
        _T_43 <= _T_123;
      end
    end
  end
endmodule
module x525_lb_0( // @[:@20005.2]
  input        clock, // @[:@20006.4]
  input        reset, // @[:@20007.4]
  input  [2:0] io_rPort_17_banks_1, // @[:@20008.4]
  input  [2:0] io_rPort_17_banks_0, // @[:@20008.4]
  input  [8:0] io_rPort_17_ofs_0, // @[:@20008.4]
  input        io_rPort_17_en_0, // @[:@20008.4]
  input        io_rPort_17_backpressure, // @[:@20008.4]
  output [7:0] io_rPort_17_output_0, // @[:@20008.4]
  input  [2:0] io_rPort_16_banks_1, // @[:@20008.4]
  input  [2:0] io_rPort_16_banks_0, // @[:@20008.4]
  input  [8:0] io_rPort_16_ofs_0, // @[:@20008.4]
  input        io_rPort_16_en_0, // @[:@20008.4]
  input        io_rPort_16_backpressure, // @[:@20008.4]
  output [7:0] io_rPort_16_output_0, // @[:@20008.4]
  input  [2:0] io_rPort_15_banks_1, // @[:@20008.4]
  input  [2:0] io_rPort_15_banks_0, // @[:@20008.4]
  input  [8:0] io_rPort_15_ofs_0, // @[:@20008.4]
  input        io_rPort_15_en_0, // @[:@20008.4]
  input        io_rPort_15_backpressure, // @[:@20008.4]
  output [7:0] io_rPort_15_output_0, // @[:@20008.4]
  input  [2:0] io_rPort_14_banks_1, // @[:@20008.4]
  input  [2:0] io_rPort_14_banks_0, // @[:@20008.4]
  input  [8:0] io_rPort_14_ofs_0, // @[:@20008.4]
  input        io_rPort_14_en_0, // @[:@20008.4]
  input        io_rPort_14_backpressure, // @[:@20008.4]
  output [7:0] io_rPort_14_output_0, // @[:@20008.4]
  input  [2:0] io_rPort_13_banks_1, // @[:@20008.4]
  input  [2:0] io_rPort_13_banks_0, // @[:@20008.4]
  input  [8:0] io_rPort_13_ofs_0, // @[:@20008.4]
  input        io_rPort_13_en_0, // @[:@20008.4]
  input        io_rPort_13_backpressure, // @[:@20008.4]
  output [7:0] io_rPort_13_output_0, // @[:@20008.4]
  input  [2:0] io_rPort_12_banks_1, // @[:@20008.4]
  input  [2:0] io_rPort_12_banks_0, // @[:@20008.4]
  input  [8:0] io_rPort_12_ofs_0, // @[:@20008.4]
  input        io_rPort_12_en_0, // @[:@20008.4]
  input        io_rPort_12_backpressure, // @[:@20008.4]
  output [7:0] io_rPort_12_output_0, // @[:@20008.4]
  input  [2:0] io_rPort_11_banks_1, // @[:@20008.4]
  input  [2:0] io_rPort_11_banks_0, // @[:@20008.4]
  input  [8:0] io_rPort_11_ofs_0, // @[:@20008.4]
  input        io_rPort_11_en_0, // @[:@20008.4]
  input        io_rPort_11_backpressure, // @[:@20008.4]
  output [7:0] io_rPort_11_output_0, // @[:@20008.4]
  input  [2:0] io_rPort_10_banks_1, // @[:@20008.4]
  input  [2:0] io_rPort_10_banks_0, // @[:@20008.4]
  input  [8:0] io_rPort_10_ofs_0, // @[:@20008.4]
  input        io_rPort_10_en_0, // @[:@20008.4]
  input        io_rPort_10_backpressure, // @[:@20008.4]
  output [7:0] io_rPort_10_output_0, // @[:@20008.4]
  input  [2:0] io_rPort_9_banks_1, // @[:@20008.4]
  input  [2:0] io_rPort_9_banks_0, // @[:@20008.4]
  input  [8:0] io_rPort_9_ofs_0, // @[:@20008.4]
  input        io_rPort_9_en_0, // @[:@20008.4]
  input        io_rPort_9_backpressure, // @[:@20008.4]
  output [7:0] io_rPort_9_output_0, // @[:@20008.4]
  input  [2:0] io_rPort_8_banks_1, // @[:@20008.4]
  input  [2:0] io_rPort_8_banks_0, // @[:@20008.4]
  input  [8:0] io_rPort_8_ofs_0, // @[:@20008.4]
  input        io_rPort_8_en_0, // @[:@20008.4]
  input        io_rPort_8_backpressure, // @[:@20008.4]
  output [7:0] io_rPort_8_output_0, // @[:@20008.4]
  input  [2:0] io_rPort_7_banks_1, // @[:@20008.4]
  input  [2:0] io_rPort_7_banks_0, // @[:@20008.4]
  input  [8:0] io_rPort_7_ofs_0, // @[:@20008.4]
  input        io_rPort_7_en_0, // @[:@20008.4]
  input        io_rPort_7_backpressure, // @[:@20008.4]
  output [7:0] io_rPort_7_output_0, // @[:@20008.4]
  input  [2:0] io_rPort_6_banks_1, // @[:@20008.4]
  input  [2:0] io_rPort_6_banks_0, // @[:@20008.4]
  input  [8:0] io_rPort_6_ofs_0, // @[:@20008.4]
  input        io_rPort_6_en_0, // @[:@20008.4]
  input        io_rPort_6_backpressure, // @[:@20008.4]
  output [7:0] io_rPort_6_output_0, // @[:@20008.4]
  input  [2:0] io_rPort_5_banks_1, // @[:@20008.4]
  input  [2:0] io_rPort_5_banks_0, // @[:@20008.4]
  input  [8:0] io_rPort_5_ofs_0, // @[:@20008.4]
  input        io_rPort_5_en_0, // @[:@20008.4]
  input        io_rPort_5_backpressure, // @[:@20008.4]
  output [7:0] io_rPort_5_output_0, // @[:@20008.4]
  input  [2:0] io_rPort_4_banks_1, // @[:@20008.4]
  input  [2:0] io_rPort_4_banks_0, // @[:@20008.4]
  input  [8:0] io_rPort_4_ofs_0, // @[:@20008.4]
  input        io_rPort_4_en_0, // @[:@20008.4]
  input        io_rPort_4_backpressure, // @[:@20008.4]
  output [7:0] io_rPort_4_output_0, // @[:@20008.4]
  input  [2:0] io_rPort_3_banks_1, // @[:@20008.4]
  input  [2:0] io_rPort_3_banks_0, // @[:@20008.4]
  input  [8:0] io_rPort_3_ofs_0, // @[:@20008.4]
  input        io_rPort_3_en_0, // @[:@20008.4]
  input        io_rPort_3_backpressure, // @[:@20008.4]
  output [7:0] io_rPort_3_output_0, // @[:@20008.4]
  input  [2:0] io_rPort_2_banks_1, // @[:@20008.4]
  input  [2:0] io_rPort_2_banks_0, // @[:@20008.4]
  input  [8:0] io_rPort_2_ofs_0, // @[:@20008.4]
  input        io_rPort_2_en_0, // @[:@20008.4]
  input        io_rPort_2_backpressure, // @[:@20008.4]
  output [7:0] io_rPort_2_output_0, // @[:@20008.4]
  input  [2:0] io_rPort_1_banks_1, // @[:@20008.4]
  input  [2:0] io_rPort_1_banks_0, // @[:@20008.4]
  input  [8:0] io_rPort_1_ofs_0, // @[:@20008.4]
  input        io_rPort_1_en_0, // @[:@20008.4]
  input        io_rPort_1_backpressure, // @[:@20008.4]
  output [7:0] io_rPort_1_output_0, // @[:@20008.4]
  input  [2:0] io_rPort_0_banks_1, // @[:@20008.4]
  input  [2:0] io_rPort_0_banks_0, // @[:@20008.4]
  input  [8:0] io_rPort_0_ofs_0, // @[:@20008.4]
  input        io_rPort_0_en_0, // @[:@20008.4]
  input        io_rPort_0_backpressure, // @[:@20008.4]
  output [7:0] io_rPort_0_output_0, // @[:@20008.4]
  input  [2:0] io_wPort_3_banks_1, // @[:@20008.4]
  input  [2:0] io_wPort_3_banks_0, // @[:@20008.4]
  input  [8:0] io_wPort_3_ofs_0, // @[:@20008.4]
  input  [7:0] io_wPort_3_data_0, // @[:@20008.4]
  input        io_wPort_3_en_0, // @[:@20008.4]
  input  [2:0] io_wPort_2_banks_1, // @[:@20008.4]
  input  [2:0] io_wPort_2_banks_0, // @[:@20008.4]
  input  [8:0] io_wPort_2_ofs_0, // @[:@20008.4]
  input  [7:0] io_wPort_2_data_0, // @[:@20008.4]
  input        io_wPort_2_en_0, // @[:@20008.4]
  input  [2:0] io_wPort_1_banks_1, // @[:@20008.4]
  input  [2:0] io_wPort_1_banks_0, // @[:@20008.4]
  input  [8:0] io_wPort_1_ofs_0, // @[:@20008.4]
  input  [7:0] io_wPort_1_data_0, // @[:@20008.4]
  input        io_wPort_1_en_0, // @[:@20008.4]
  input  [2:0] io_wPort_0_banks_1, // @[:@20008.4]
  input  [2:0] io_wPort_0_banks_0, // @[:@20008.4]
  input  [8:0] io_wPort_0_ofs_0, // @[:@20008.4]
  input  [7:0] io_wPort_0_data_0, // @[:@20008.4]
  input        io_wPort_0_en_0 // @[:@20008.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@20151.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@20151.4]
  wire [8:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20151.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20151.4]
  wire [8:0] Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20151.4]
  wire [7:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@20151.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@20151.4]
  wire [7:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@20151.4]
  wire  Mem1D_1_clock; // @[MemPrimitives.scala 64:21:@20167.4]
  wire  Mem1D_1_reset; // @[MemPrimitives.scala 64:21:@20167.4]
  wire [8:0] Mem1D_1_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20167.4]
  wire  Mem1D_1_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20167.4]
  wire [8:0] Mem1D_1_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20167.4]
  wire [7:0] Mem1D_1_io_w_data_0; // @[MemPrimitives.scala 64:21:@20167.4]
  wire  Mem1D_1_io_w_en_0; // @[MemPrimitives.scala 64:21:@20167.4]
  wire [7:0] Mem1D_1_io_output; // @[MemPrimitives.scala 64:21:@20167.4]
  wire  Mem1D_2_clock; // @[MemPrimitives.scala 64:21:@20183.4]
  wire  Mem1D_2_reset; // @[MemPrimitives.scala 64:21:@20183.4]
  wire [8:0] Mem1D_2_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20183.4]
  wire  Mem1D_2_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20183.4]
  wire [8:0] Mem1D_2_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20183.4]
  wire [7:0] Mem1D_2_io_w_data_0; // @[MemPrimitives.scala 64:21:@20183.4]
  wire  Mem1D_2_io_w_en_0; // @[MemPrimitives.scala 64:21:@20183.4]
  wire [7:0] Mem1D_2_io_output; // @[MemPrimitives.scala 64:21:@20183.4]
  wire  Mem1D_3_clock; // @[MemPrimitives.scala 64:21:@20199.4]
  wire  Mem1D_3_reset; // @[MemPrimitives.scala 64:21:@20199.4]
  wire [8:0] Mem1D_3_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20199.4]
  wire  Mem1D_3_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20199.4]
  wire [8:0] Mem1D_3_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20199.4]
  wire [7:0] Mem1D_3_io_w_data_0; // @[MemPrimitives.scala 64:21:@20199.4]
  wire  Mem1D_3_io_w_en_0; // @[MemPrimitives.scala 64:21:@20199.4]
  wire [7:0] Mem1D_3_io_output; // @[MemPrimitives.scala 64:21:@20199.4]
  wire  Mem1D_4_clock; // @[MemPrimitives.scala 64:21:@20215.4]
  wire  Mem1D_4_reset; // @[MemPrimitives.scala 64:21:@20215.4]
  wire [8:0] Mem1D_4_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20215.4]
  wire  Mem1D_4_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20215.4]
  wire [8:0] Mem1D_4_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20215.4]
  wire [7:0] Mem1D_4_io_w_data_0; // @[MemPrimitives.scala 64:21:@20215.4]
  wire  Mem1D_4_io_w_en_0; // @[MemPrimitives.scala 64:21:@20215.4]
  wire [7:0] Mem1D_4_io_output; // @[MemPrimitives.scala 64:21:@20215.4]
  wire  Mem1D_5_clock; // @[MemPrimitives.scala 64:21:@20231.4]
  wire  Mem1D_5_reset; // @[MemPrimitives.scala 64:21:@20231.4]
  wire [8:0] Mem1D_5_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20231.4]
  wire  Mem1D_5_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20231.4]
  wire [8:0] Mem1D_5_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20231.4]
  wire [7:0] Mem1D_5_io_w_data_0; // @[MemPrimitives.scala 64:21:@20231.4]
  wire  Mem1D_5_io_w_en_0; // @[MemPrimitives.scala 64:21:@20231.4]
  wire [7:0] Mem1D_5_io_output; // @[MemPrimitives.scala 64:21:@20231.4]
  wire  Mem1D_6_clock; // @[MemPrimitives.scala 64:21:@20247.4]
  wire  Mem1D_6_reset; // @[MemPrimitives.scala 64:21:@20247.4]
  wire [8:0] Mem1D_6_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20247.4]
  wire  Mem1D_6_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20247.4]
  wire [8:0] Mem1D_6_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20247.4]
  wire [7:0] Mem1D_6_io_w_data_0; // @[MemPrimitives.scala 64:21:@20247.4]
  wire  Mem1D_6_io_w_en_0; // @[MemPrimitives.scala 64:21:@20247.4]
  wire [7:0] Mem1D_6_io_output; // @[MemPrimitives.scala 64:21:@20247.4]
  wire  Mem1D_7_clock; // @[MemPrimitives.scala 64:21:@20263.4]
  wire  Mem1D_7_reset; // @[MemPrimitives.scala 64:21:@20263.4]
  wire [8:0] Mem1D_7_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20263.4]
  wire  Mem1D_7_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20263.4]
  wire [8:0] Mem1D_7_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20263.4]
  wire [7:0] Mem1D_7_io_w_data_0; // @[MemPrimitives.scala 64:21:@20263.4]
  wire  Mem1D_7_io_w_en_0; // @[MemPrimitives.scala 64:21:@20263.4]
  wire [7:0] Mem1D_7_io_output; // @[MemPrimitives.scala 64:21:@20263.4]
  wire  Mem1D_8_clock; // @[MemPrimitives.scala 64:21:@20279.4]
  wire  Mem1D_8_reset; // @[MemPrimitives.scala 64:21:@20279.4]
  wire [8:0] Mem1D_8_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20279.4]
  wire  Mem1D_8_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20279.4]
  wire [8:0] Mem1D_8_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20279.4]
  wire [7:0] Mem1D_8_io_w_data_0; // @[MemPrimitives.scala 64:21:@20279.4]
  wire  Mem1D_8_io_w_en_0; // @[MemPrimitives.scala 64:21:@20279.4]
  wire [7:0] Mem1D_8_io_output; // @[MemPrimitives.scala 64:21:@20279.4]
  wire  Mem1D_9_clock; // @[MemPrimitives.scala 64:21:@20295.4]
  wire  Mem1D_9_reset; // @[MemPrimitives.scala 64:21:@20295.4]
  wire [8:0] Mem1D_9_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20295.4]
  wire  Mem1D_9_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20295.4]
  wire [8:0] Mem1D_9_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20295.4]
  wire [7:0] Mem1D_9_io_w_data_0; // @[MemPrimitives.scala 64:21:@20295.4]
  wire  Mem1D_9_io_w_en_0; // @[MemPrimitives.scala 64:21:@20295.4]
  wire [7:0] Mem1D_9_io_output; // @[MemPrimitives.scala 64:21:@20295.4]
  wire  Mem1D_10_clock; // @[MemPrimitives.scala 64:21:@20311.4]
  wire  Mem1D_10_reset; // @[MemPrimitives.scala 64:21:@20311.4]
  wire [8:0] Mem1D_10_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20311.4]
  wire  Mem1D_10_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20311.4]
  wire [8:0] Mem1D_10_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20311.4]
  wire [7:0] Mem1D_10_io_w_data_0; // @[MemPrimitives.scala 64:21:@20311.4]
  wire  Mem1D_10_io_w_en_0; // @[MemPrimitives.scala 64:21:@20311.4]
  wire [7:0] Mem1D_10_io_output; // @[MemPrimitives.scala 64:21:@20311.4]
  wire  Mem1D_11_clock; // @[MemPrimitives.scala 64:21:@20327.4]
  wire  Mem1D_11_reset; // @[MemPrimitives.scala 64:21:@20327.4]
  wire [8:0] Mem1D_11_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20327.4]
  wire  Mem1D_11_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20327.4]
  wire [8:0] Mem1D_11_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20327.4]
  wire [7:0] Mem1D_11_io_w_data_0; // @[MemPrimitives.scala 64:21:@20327.4]
  wire  Mem1D_11_io_w_en_0; // @[MemPrimitives.scala 64:21:@20327.4]
  wire [7:0] Mem1D_11_io_output; // @[MemPrimitives.scala 64:21:@20327.4]
  wire  Mem1D_12_clock; // @[MemPrimitives.scala 64:21:@20343.4]
  wire  Mem1D_12_reset; // @[MemPrimitives.scala 64:21:@20343.4]
  wire [8:0] Mem1D_12_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20343.4]
  wire  Mem1D_12_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20343.4]
  wire [8:0] Mem1D_12_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20343.4]
  wire [7:0] Mem1D_12_io_w_data_0; // @[MemPrimitives.scala 64:21:@20343.4]
  wire  Mem1D_12_io_w_en_0; // @[MemPrimitives.scala 64:21:@20343.4]
  wire [7:0] Mem1D_12_io_output; // @[MemPrimitives.scala 64:21:@20343.4]
  wire  Mem1D_13_clock; // @[MemPrimitives.scala 64:21:@20359.4]
  wire  Mem1D_13_reset; // @[MemPrimitives.scala 64:21:@20359.4]
  wire [8:0] Mem1D_13_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20359.4]
  wire  Mem1D_13_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20359.4]
  wire [8:0] Mem1D_13_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20359.4]
  wire [7:0] Mem1D_13_io_w_data_0; // @[MemPrimitives.scala 64:21:@20359.4]
  wire  Mem1D_13_io_w_en_0; // @[MemPrimitives.scala 64:21:@20359.4]
  wire [7:0] Mem1D_13_io_output; // @[MemPrimitives.scala 64:21:@20359.4]
  wire  Mem1D_14_clock; // @[MemPrimitives.scala 64:21:@20375.4]
  wire  Mem1D_14_reset; // @[MemPrimitives.scala 64:21:@20375.4]
  wire [8:0] Mem1D_14_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20375.4]
  wire  Mem1D_14_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20375.4]
  wire [8:0] Mem1D_14_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20375.4]
  wire [7:0] Mem1D_14_io_w_data_0; // @[MemPrimitives.scala 64:21:@20375.4]
  wire  Mem1D_14_io_w_en_0; // @[MemPrimitives.scala 64:21:@20375.4]
  wire [7:0] Mem1D_14_io_output; // @[MemPrimitives.scala 64:21:@20375.4]
  wire  Mem1D_15_clock; // @[MemPrimitives.scala 64:21:@20391.4]
  wire  Mem1D_15_reset; // @[MemPrimitives.scala 64:21:@20391.4]
  wire [8:0] Mem1D_15_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20391.4]
  wire  Mem1D_15_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20391.4]
  wire [8:0] Mem1D_15_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20391.4]
  wire [7:0] Mem1D_15_io_w_data_0; // @[MemPrimitives.scala 64:21:@20391.4]
  wire  Mem1D_15_io_w_en_0; // @[MemPrimitives.scala 64:21:@20391.4]
  wire [7:0] Mem1D_15_io_output; // @[MemPrimitives.scala 64:21:@20391.4]
  wire  Mem1D_16_clock; // @[MemPrimitives.scala 64:21:@20407.4]
  wire  Mem1D_16_reset; // @[MemPrimitives.scala 64:21:@20407.4]
  wire [8:0] Mem1D_16_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20407.4]
  wire  Mem1D_16_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20407.4]
  wire [8:0] Mem1D_16_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20407.4]
  wire [7:0] Mem1D_16_io_w_data_0; // @[MemPrimitives.scala 64:21:@20407.4]
  wire  Mem1D_16_io_w_en_0; // @[MemPrimitives.scala 64:21:@20407.4]
  wire [7:0] Mem1D_16_io_output; // @[MemPrimitives.scala 64:21:@20407.4]
  wire  Mem1D_17_clock; // @[MemPrimitives.scala 64:21:@20423.4]
  wire  Mem1D_17_reset; // @[MemPrimitives.scala 64:21:@20423.4]
  wire [8:0] Mem1D_17_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20423.4]
  wire  Mem1D_17_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20423.4]
  wire [8:0] Mem1D_17_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20423.4]
  wire [7:0] Mem1D_17_io_w_data_0; // @[MemPrimitives.scala 64:21:@20423.4]
  wire  Mem1D_17_io_w_en_0; // @[MemPrimitives.scala 64:21:@20423.4]
  wire [7:0] Mem1D_17_io_output; // @[MemPrimitives.scala 64:21:@20423.4]
  wire  Mem1D_18_clock; // @[MemPrimitives.scala 64:21:@20439.4]
  wire  Mem1D_18_reset; // @[MemPrimitives.scala 64:21:@20439.4]
  wire [8:0] Mem1D_18_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20439.4]
  wire  Mem1D_18_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20439.4]
  wire [8:0] Mem1D_18_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20439.4]
  wire [7:0] Mem1D_18_io_w_data_0; // @[MemPrimitives.scala 64:21:@20439.4]
  wire  Mem1D_18_io_w_en_0; // @[MemPrimitives.scala 64:21:@20439.4]
  wire [7:0] Mem1D_18_io_output; // @[MemPrimitives.scala 64:21:@20439.4]
  wire  Mem1D_19_clock; // @[MemPrimitives.scala 64:21:@20455.4]
  wire  Mem1D_19_reset; // @[MemPrimitives.scala 64:21:@20455.4]
  wire [8:0] Mem1D_19_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20455.4]
  wire  Mem1D_19_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20455.4]
  wire [8:0] Mem1D_19_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20455.4]
  wire [7:0] Mem1D_19_io_w_data_0; // @[MemPrimitives.scala 64:21:@20455.4]
  wire  Mem1D_19_io_w_en_0; // @[MemPrimitives.scala 64:21:@20455.4]
  wire [7:0] Mem1D_19_io_output; // @[MemPrimitives.scala 64:21:@20455.4]
  wire  Mem1D_20_clock; // @[MemPrimitives.scala 64:21:@20471.4]
  wire  Mem1D_20_reset; // @[MemPrimitives.scala 64:21:@20471.4]
  wire [8:0] Mem1D_20_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20471.4]
  wire  Mem1D_20_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20471.4]
  wire [8:0] Mem1D_20_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20471.4]
  wire [7:0] Mem1D_20_io_w_data_0; // @[MemPrimitives.scala 64:21:@20471.4]
  wire  Mem1D_20_io_w_en_0; // @[MemPrimitives.scala 64:21:@20471.4]
  wire [7:0] Mem1D_20_io_output; // @[MemPrimitives.scala 64:21:@20471.4]
  wire  Mem1D_21_clock; // @[MemPrimitives.scala 64:21:@20487.4]
  wire  Mem1D_21_reset; // @[MemPrimitives.scala 64:21:@20487.4]
  wire [8:0] Mem1D_21_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20487.4]
  wire  Mem1D_21_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20487.4]
  wire [8:0] Mem1D_21_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20487.4]
  wire [7:0] Mem1D_21_io_w_data_0; // @[MemPrimitives.scala 64:21:@20487.4]
  wire  Mem1D_21_io_w_en_0; // @[MemPrimitives.scala 64:21:@20487.4]
  wire [7:0] Mem1D_21_io_output; // @[MemPrimitives.scala 64:21:@20487.4]
  wire  Mem1D_22_clock; // @[MemPrimitives.scala 64:21:@20503.4]
  wire  Mem1D_22_reset; // @[MemPrimitives.scala 64:21:@20503.4]
  wire [8:0] Mem1D_22_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20503.4]
  wire  Mem1D_22_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20503.4]
  wire [8:0] Mem1D_22_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20503.4]
  wire [7:0] Mem1D_22_io_w_data_0; // @[MemPrimitives.scala 64:21:@20503.4]
  wire  Mem1D_22_io_w_en_0; // @[MemPrimitives.scala 64:21:@20503.4]
  wire [7:0] Mem1D_22_io_output; // @[MemPrimitives.scala 64:21:@20503.4]
  wire  Mem1D_23_clock; // @[MemPrimitives.scala 64:21:@20519.4]
  wire  Mem1D_23_reset; // @[MemPrimitives.scala 64:21:@20519.4]
  wire [8:0] Mem1D_23_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20519.4]
  wire  Mem1D_23_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20519.4]
  wire [8:0] Mem1D_23_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20519.4]
  wire [7:0] Mem1D_23_io_w_data_0; // @[MemPrimitives.scala 64:21:@20519.4]
  wire  Mem1D_23_io_w_en_0; // @[MemPrimitives.scala 64:21:@20519.4]
  wire [7:0] Mem1D_23_io_output; // @[MemPrimitives.scala 64:21:@20519.4]
  wire  StickySelects_clock; // @[MemPrimitives.scala 121:29:@21027.4]
  wire  StickySelects_reset; // @[MemPrimitives.scala 121:29:@21027.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 121:29:@21027.4]
  wire  StickySelects_io_ins_1; // @[MemPrimitives.scala 121:29:@21027.4]
  wire  StickySelects_io_ins_2; // @[MemPrimitives.scala 121:29:@21027.4]
  wire  StickySelects_io_ins_3; // @[MemPrimitives.scala 121:29:@21027.4]
  wire  StickySelects_io_ins_4; // @[MemPrimitives.scala 121:29:@21027.4]
  wire  StickySelects_io_ins_5; // @[MemPrimitives.scala 121:29:@21027.4]
  wire  StickySelects_io_ins_6; // @[MemPrimitives.scala 121:29:@21027.4]
  wire  StickySelects_io_ins_7; // @[MemPrimitives.scala 121:29:@21027.4]
  wire  StickySelects_io_ins_8; // @[MemPrimitives.scala 121:29:@21027.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 121:29:@21027.4]
  wire  StickySelects_io_outs_1; // @[MemPrimitives.scala 121:29:@21027.4]
  wire  StickySelects_io_outs_2; // @[MemPrimitives.scala 121:29:@21027.4]
  wire  StickySelects_io_outs_3; // @[MemPrimitives.scala 121:29:@21027.4]
  wire  StickySelects_io_outs_4; // @[MemPrimitives.scala 121:29:@21027.4]
  wire  StickySelects_io_outs_5; // @[MemPrimitives.scala 121:29:@21027.4]
  wire  StickySelects_io_outs_6; // @[MemPrimitives.scala 121:29:@21027.4]
  wire  StickySelects_io_outs_7; // @[MemPrimitives.scala 121:29:@21027.4]
  wire  StickySelects_io_outs_8; // @[MemPrimitives.scala 121:29:@21027.4]
  wire  StickySelects_1_clock; // @[MemPrimitives.scala 121:29:@21116.4]
  wire  StickySelects_1_reset; // @[MemPrimitives.scala 121:29:@21116.4]
  wire  StickySelects_1_io_ins_0; // @[MemPrimitives.scala 121:29:@21116.4]
  wire  StickySelects_1_io_ins_1; // @[MemPrimitives.scala 121:29:@21116.4]
  wire  StickySelects_1_io_ins_2; // @[MemPrimitives.scala 121:29:@21116.4]
  wire  StickySelects_1_io_ins_3; // @[MemPrimitives.scala 121:29:@21116.4]
  wire  StickySelects_1_io_ins_4; // @[MemPrimitives.scala 121:29:@21116.4]
  wire  StickySelects_1_io_ins_5; // @[MemPrimitives.scala 121:29:@21116.4]
  wire  StickySelects_1_io_ins_6; // @[MemPrimitives.scala 121:29:@21116.4]
  wire  StickySelects_1_io_ins_7; // @[MemPrimitives.scala 121:29:@21116.4]
  wire  StickySelects_1_io_ins_8; // @[MemPrimitives.scala 121:29:@21116.4]
  wire  StickySelects_1_io_outs_0; // @[MemPrimitives.scala 121:29:@21116.4]
  wire  StickySelects_1_io_outs_1; // @[MemPrimitives.scala 121:29:@21116.4]
  wire  StickySelects_1_io_outs_2; // @[MemPrimitives.scala 121:29:@21116.4]
  wire  StickySelects_1_io_outs_3; // @[MemPrimitives.scala 121:29:@21116.4]
  wire  StickySelects_1_io_outs_4; // @[MemPrimitives.scala 121:29:@21116.4]
  wire  StickySelects_1_io_outs_5; // @[MemPrimitives.scala 121:29:@21116.4]
  wire  StickySelects_1_io_outs_6; // @[MemPrimitives.scala 121:29:@21116.4]
  wire  StickySelects_1_io_outs_7; // @[MemPrimitives.scala 121:29:@21116.4]
  wire  StickySelects_1_io_outs_8; // @[MemPrimitives.scala 121:29:@21116.4]
  wire  StickySelects_2_clock; // @[MemPrimitives.scala 121:29:@21205.4]
  wire  StickySelects_2_reset; // @[MemPrimitives.scala 121:29:@21205.4]
  wire  StickySelects_2_io_ins_0; // @[MemPrimitives.scala 121:29:@21205.4]
  wire  StickySelects_2_io_ins_1; // @[MemPrimitives.scala 121:29:@21205.4]
  wire  StickySelects_2_io_ins_2; // @[MemPrimitives.scala 121:29:@21205.4]
  wire  StickySelects_2_io_ins_3; // @[MemPrimitives.scala 121:29:@21205.4]
  wire  StickySelects_2_io_ins_4; // @[MemPrimitives.scala 121:29:@21205.4]
  wire  StickySelects_2_io_ins_5; // @[MemPrimitives.scala 121:29:@21205.4]
  wire  StickySelects_2_io_ins_6; // @[MemPrimitives.scala 121:29:@21205.4]
  wire  StickySelects_2_io_ins_7; // @[MemPrimitives.scala 121:29:@21205.4]
  wire  StickySelects_2_io_ins_8; // @[MemPrimitives.scala 121:29:@21205.4]
  wire  StickySelects_2_io_outs_0; // @[MemPrimitives.scala 121:29:@21205.4]
  wire  StickySelects_2_io_outs_1; // @[MemPrimitives.scala 121:29:@21205.4]
  wire  StickySelects_2_io_outs_2; // @[MemPrimitives.scala 121:29:@21205.4]
  wire  StickySelects_2_io_outs_3; // @[MemPrimitives.scala 121:29:@21205.4]
  wire  StickySelects_2_io_outs_4; // @[MemPrimitives.scala 121:29:@21205.4]
  wire  StickySelects_2_io_outs_5; // @[MemPrimitives.scala 121:29:@21205.4]
  wire  StickySelects_2_io_outs_6; // @[MemPrimitives.scala 121:29:@21205.4]
  wire  StickySelects_2_io_outs_7; // @[MemPrimitives.scala 121:29:@21205.4]
  wire  StickySelects_2_io_outs_8; // @[MemPrimitives.scala 121:29:@21205.4]
  wire  StickySelects_3_clock; // @[MemPrimitives.scala 121:29:@21294.4]
  wire  StickySelects_3_reset; // @[MemPrimitives.scala 121:29:@21294.4]
  wire  StickySelects_3_io_ins_0; // @[MemPrimitives.scala 121:29:@21294.4]
  wire  StickySelects_3_io_ins_1; // @[MemPrimitives.scala 121:29:@21294.4]
  wire  StickySelects_3_io_ins_2; // @[MemPrimitives.scala 121:29:@21294.4]
  wire  StickySelects_3_io_ins_3; // @[MemPrimitives.scala 121:29:@21294.4]
  wire  StickySelects_3_io_ins_4; // @[MemPrimitives.scala 121:29:@21294.4]
  wire  StickySelects_3_io_ins_5; // @[MemPrimitives.scala 121:29:@21294.4]
  wire  StickySelects_3_io_ins_6; // @[MemPrimitives.scala 121:29:@21294.4]
  wire  StickySelects_3_io_ins_7; // @[MemPrimitives.scala 121:29:@21294.4]
  wire  StickySelects_3_io_ins_8; // @[MemPrimitives.scala 121:29:@21294.4]
  wire  StickySelects_3_io_outs_0; // @[MemPrimitives.scala 121:29:@21294.4]
  wire  StickySelects_3_io_outs_1; // @[MemPrimitives.scala 121:29:@21294.4]
  wire  StickySelects_3_io_outs_2; // @[MemPrimitives.scala 121:29:@21294.4]
  wire  StickySelects_3_io_outs_3; // @[MemPrimitives.scala 121:29:@21294.4]
  wire  StickySelects_3_io_outs_4; // @[MemPrimitives.scala 121:29:@21294.4]
  wire  StickySelects_3_io_outs_5; // @[MemPrimitives.scala 121:29:@21294.4]
  wire  StickySelects_3_io_outs_6; // @[MemPrimitives.scala 121:29:@21294.4]
  wire  StickySelects_3_io_outs_7; // @[MemPrimitives.scala 121:29:@21294.4]
  wire  StickySelects_3_io_outs_8; // @[MemPrimitives.scala 121:29:@21294.4]
  wire  StickySelects_4_clock; // @[MemPrimitives.scala 121:29:@21383.4]
  wire  StickySelects_4_reset; // @[MemPrimitives.scala 121:29:@21383.4]
  wire  StickySelects_4_io_ins_0; // @[MemPrimitives.scala 121:29:@21383.4]
  wire  StickySelects_4_io_ins_1; // @[MemPrimitives.scala 121:29:@21383.4]
  wire  StickySelects_4_io_ins_2; // @[MemPrimitives.scala 121:29:@21383.4]
  wire  StickySelects_4_io_ins_3; // @[MemPrimitives.scala 121:29:@21383.4]
  wire  StickySelects_4_io_ins_4; // @[MemPrimitives.scala 121:29:@21383.4]
  wire  StickySelects_4_io_ins_5; // @[MemPrimitives.scala 121:29:@21383.4]
  wire  StickySelects_4_io_ins_6; // @[MemPrimitives.scala 121:29:@21383.4]
  wire  StickySelects_4_io_ins_7; // @[MemPrimitives.scala 121:29:@21383.4]
  wire  StickySelects_4_io_ins_8; // @[MemPrimitives.scala 121:29:@21383.4]
  wire  StickySelects_4_io_outs_0; // @[MemPrimitives.scala 121:29:@21383.4]
  wire  StickySelects_4_io_outs_1; // @[MemPrimitives.scala 121:29:@21383.4]
  wire  StickySelects_4_io_outs_2; // @[MemPrimitives.scala 121:29:@21383.4]
  wire  StickySelects_4_io_outs_3; // @[MemPrimitives.scala 121:29:@21383.4]
  wire  StickySelects_4_io_outs_4; // @[MemPrimitives.scala 121:29:@21383.4]
  wire  StickySelects_4_io_outs_5; // @[MemPrimitives.scala 121:29:@21383.4]
  wire  StickySelects_4_io_outs_6; // @[MemPrimitives.scala 121:29:@21383.4]
  wire  StickySelects_4_io_outs_7; // @[MemPrimitives.scala 121:29:@21383.4]
  wire  StickySelects_4_io_outs_8; // @[MemPrimitives.scala 121:29:@21383.4]
  wire  StickySelects_5_clock; // @[MemPrimitives.scala 121:29:@21472.4]
  wire  StickySelects_5_reset; // @[MemPrimitives.scala 121:29:@21472.4]
  wire  StickySelects_5_io_ins_0; // @[MemPrimitives.scala 121:29:@21472.4]
  wire  StickySelects_5_io_ins_1; // @[MemPrimitives.scala 121:29:@21472.4]
  wire  StickySelects_5_io_ins_2; // @[MemPrimitives.scala 121:29:@21472.4]
  wire  StickySelects_5_io_ins_3; // @[MemPrimitives.scala 121:29:@21472.4]
  wire  StickySelects_5_io_ins_4; // @[MemPrimitives.scala 121:29:@21472.4]
  wire  StickySelects_5_io_ins_5; // @[MemPrimitives.scala 121:29:@21472.4]
  wire  StickySelects_5_io_ins_6; // @[MemPrimitives.scala 121:29:@21472.4]
  wire  StickySelects_5_io_ins_7; // @[MemPrimitives.scala 121:29:@21472.4]
  wire  StickySelects_5_io_ins_8; // @[MemPrimitives.scala 121:29:@21472.4]
  wire  StickySelects_5_io_outs_0; // @[MemPrimitives.scala 121:29:@21472.4]
  wire  StickySelects_5_io_outs_1; // @[MemPrimitives.scala 121:29:@21472.4]
  wire  StickySelects_5_io_outs_2; // @[MemPrimitives.scala 121:29:@21472.4]
  wire  StickySelects_5_io_outs_3; // @[MemPrimitives.scala 121:29:@21472.4]
  wire  StickySelects_5_io_outs_4; // @[MemPrimitives.scala 121:29:@21472.4]
  wire  StickySelects_5_io_outs_5; // @[MemPrimitives.scala 121:29:@21472.4]
  wire  StickySelects_5_io_outs_6; // @[MemPrimitives.scala 121:29:@21472.4]
  wire  StickySelects_5_io_outs_7; // @[MemPrimitives.scala 121:29:@21472.4]
  wire  StickySelects_5_io_outs_8; // @[MemPrimitives.scala 121:29:@21472.4]
  wire  StickySelects_6_clock; // @[MemPrimitives.scala 121:29:@21561.4]
  wire  StickySelects_6_reset; // @[MemPrimitives.scala 121:29:@21561.4]
  wire  StickySelects_6_io_ins_0; // @[MemPrimitives.scala 121:29:@21561.4]
  wire  StickySelects_6_io_ins_1; // @[MemPrimitives.scala 121:29:@21561.4]
  wire  StickySelects_6_io_ins_2; // @[MemPrimitives.scala 121:29:@21561.4]
  wire  StickySelects_6_io_ins_3; // @[MemPrimitives.scala 121:29:@21561.4]
  wire  StickySelects_6_io_ins_4; // @[MemPrimitives.scala 121:29:@21561.4]
  wire  StickySelects_6_io_ins_5; // @[MemPrimitives.scala 121:29:@21561.4]
  wire  StickySelects_6_io_ins_6; // @[MemPrimitives.scala 121:29:@21561.4]
  wire  StickySelects_6_io_ins_7; // @[MemPrimitives.scala 121:29:@21561.4]
  wire  StickySelects_6_io_ins_8; // @[MemPrimitives.scala 121:29:@21561.4]
  wire  StickySelects_6_io_outs_0; // @[MemPrimitives.scala 121:29:@21561.4]
  wire  StickySelects_6_io_outs_1; // @[MemPrimitives.scala 121:29:@21561.4]
  wire  StickySelects_6_io_outs_2; // @[MemPrimitives.scala 121:29:@21561.4]
  wire  StickySelects_6_io_outs_3; // @[MemPrimitives.scala 121:29:@21561.4]
  wire  StickySelects_6_io_outs_4; // @[MemPrimitives.scala 121:29:@21561.4]
  wire  StickySelects_6_io_outs_5; // @[MemPrimitives.scala 121:29:@21561.4]
  wire  StickySelects_6_io_outs_6; // @[MemPrimitives.scala 121:29:@21561.4]
  wire  StickySelects_6_io_outs_7; // @[MemPrimitives.scala 121:29:@21561.4]
  wire  StickySelects_6_io_outs_8; // @[MemPrimitives.scala 121:29:@21561.4]
  wire  StickySelects_7_clock; // @[MemPrimitives.scala 121:29:@21650.4]
  wire  StickySelects_7_reset; // @[MemPrimitives.scala 121:29:@21650.4]
  wire  StickySelects_7_io_ins_0; // @[MemPrimitives.scala 121:29:@21650.4]
  wire  StickySelects_7_io_ins_1; // @[MemPrimitives.scala 121:29:@21650.4]
  wire  StickySelects_7_io_ins_2; // @[MemPrimitives.scala 121:29:@21650.4]
  wire  StickySelects_7_io_ins_3; // @[MemPrimitives.scala 121:29:@21650.4]
  wire  StickySelects_7_io_ins_4; // @[MemPrimitives.scala 121:29:@21650.4]
  wire  StickySelects_7_io_ins_5; // @[MemPrimitives.scala 121:29:@21650.4]
  wire  StickySelects_7_io_ins_6; // @[MemPrimitives.scala 121:29:@21650.4]
  wire  StickySelects_7_io_ins_7; // @[MemPrimitives.scala 121:29:@21650.4]
  wire  StickySelects_7_io_ins_8; // @[MemPrimitives.scala 121:29:@21650.4]
  wire  StickySelects_7_io_outs_0; // @[MemPrimitives.scala 121:29:@21650.4]
  wire  StickySelects_7_io_outs_1; // @[MemPrimitives.scala 121:29:@21650.4]
  wire  StickySelects_7_io_outs_2; // @[MemPrimitives.scala 121:29:@21650.4]
  wire  StickySelects_7_io_outs_3; // @[MemPrimitives.scala 121:29:@21650.4]
  wire  StickySelects_7_io_outs_4; // @[MemPrimitives.scala 121:29:@21650.4]
  wire  StickySelects_7_io_outs_5; // @[MemPrimitives.scala 121:29:@21650.4]
  wire  StickySelects_7_io_outs_6; // @[MemPrimitives.scala 121:29:@21650.4]
  wire  StickySelects_7_io_outs_7; // @[MemPrimitives.scala 121:29:@21650.4]
  wire  StickySelects_7_io_outs_8; // @[MemPrimitives.scala 121:29:@21650.4]
  wire  StickySelects_8_clock; // @[MemPrimitives.scala 121:29:@21739.4]
  wire  StickySelects_8_reset; // @[MemPrimitives.scala 121:29:@21739.4]
  wire  StickySelects_8_io_ins_0; // @[MemPrimitives.scala 121:29:@21739.4]
  wire  StickySelects_8_io_ins_1; // @[MemPrimitives.scala 121:29:@21739.4]
  wire  StickySelects_8_io_ins_2; // @[MemPrimitives.scala 121:29:@21739.4]
  wire  StickySelects_8_io_ins_3; // @[MemPrimitives.scala 121:29:@21739.4]
  wire  StickySelects_8_io_ins_4; // @[MemPrimitives.scala 121:29:@21739.4]
  wire  StickySelects_8_io_ins_5; // @[MemPrimitives.scala 121:29:@21739.4]
  wire  StickySelects_8_io_ins_6; // @[MemPrimitives.scala 121:29:@21739.4]
  wire  StickySelects_8_io_ins_7; // @[MemPrimitives.scala 121:29:@21739.4]
  wire  StickySelects_8_io_ins_8; // @[MemPrimitives.scala 121:29:@21739.4]
  wire  StickySelects_8_io_outs_0; // @[MemPrimitives.scala 121:29:@21739.4]
  wire  StickySelects_8_io_outs_1; // @[MemPrimitives.scala 121:29:@21739.4]
  wire  StickySelects_8_io_outs_2; // @[MemPrimitives.scala 121:29:@21739.4]
  wire  StickySelects_8_io_outs_3; // @[MemPrimitives.scala 121:29:@21739.4]
  wire  StickySelects_8_io_outs_4; // @[MemPrimitives.scala 121:29:@21739.4]
  wire  StickySelects_8_io_outs_5; // @[MemPrimitives.scala 121:29:@21739.4]
  wire  StickySelects_8_io_outs_6; // @[MemPrimitives.scala 121:29:@21739.4]
  wire  StickySelects_8_io_outs_7; // @[MemPrimitives.scala 121:29:@21739.4]
  wire  StickySelects_8_io_outs_8; // @[MemPrimitives.scala 121:29:@21739.4]
  wire  StickySelects_9_clock; // @[MemPrimitives.scala 121:29:@21828.4]
  wire  StickySelects_9_reset; // @[MemPrimitives.scala 121:29:@21828.4]
  wire  StickySelects_9_io_ins_0; // @[MemPrimitives.scala 121:29:@21828.4]
  wire  StickySelects_9_io_ins_1; // @[MemPrimitives.scala 121:29:@21828.4]
  wire  StickySelects_9_io_ins_2; // @[MemPrimitives.scala 121:29:@21828.4]
  wire  StickySelects_9_io_ins_3; // @[MemPrimitives.scala 121:29:@21828.4]
  wire  StickySelects_9_io_ins_4; // @[MemPrimitives.scala 121:29:@21828.4]
  wire  StickySelects_9_io_ins_5; // @[MemPrimitives.scala 121:29:@21828.4]
  wire  StickySelects_9_io_ins_6; // @[MemPrimitives.scala 121:29:@21828.4]
  wire  StickySelects_9_io_ins_7; // @[MemPrimitives.scala 121:29:@21828.4]
  wire  StickySelects_9_io_ins_8; // @[MemPrimitives.scala 121:29:@21828.4]
  wire  StickySelects_9_io_outs_0; // @[MemPrimitives.scala 121:29:@21828.4]
  wire  StickySelects_9_io_outs_1; // @[MemPrimitives.scala 121:29:@21828.4]
  wire  StickySelects_9_io_outs_2; // @[MemPrimitives.scala 121:29:@21828.4]
  wire  StickySelects_9_io_outs_3; // @[MemPrimitives.scala 121:29:@21828.4]
  wire  StickySelects_9_io_outs_4; // @[MemPrimitives.scala 121:29:@21828.4]
  wire  StickySelects_9_io_outs_5; // @[MemPrimitives.scala 121:29:@21828.4]
  wire  StickySelects_9_io_outs_6; // @[MemPrimitives.scala 121:29:@21828.4]
  wire  StickySelects_9_io_outs_7; // @[MemPrimitives.scala 121:29:@21828.4]
  wire  StickySelects_9_io_outs_8; // @[MemPrimitives.scala 121:29:@21828.4]
  wire  StickySelects_10_clock; // @[MemPrimitives.scala 121:29:@21917.4]
  wire  StickySelects_10_reset; // @[MemPrimitives.scala 121:29:@21917.4]
  wire  StickySelects_10_io_ins_0; // @[MemPrimitives.scala 121:29:@21917.4]
  wire  StickySelects_10_io_ins_1; // @[MemPrimitives.scala 121:29:@21917.4]
  wire  StickySelects_10_io_ins_2; // @[MemPrimitives.scala 121:29:@21917.4]
  wire  StickySelects_10_io_ins_3; // @[MemPrimitives.scala 121:29:@21917.4]
  wire  StickySelects_10_io_ins_4; // @[MemPrimitives.scala 121:29:@21917.4]
  wire  StickySelects_10_io_ins_5; // @[MemPrimitives.scala 121:29:@21917.4]
  wire  StickySelects_10_io_ins_6; // @[MemPrimitives.scala 121:29:@21917.4]
  wire  StickySelects_10_io_ins_7; // @[MemPrimitives.scala 121:29:@21917.4]
  wire  StickySelects_10_io_ins_8; // @[MemPrimitives.scala 121:29:@21917.4]
  wire  StickySelects_10_io_outs_0; // @[MemPrimitives.scala 121:29:@21917.4]
  wire  StickySelects_10_io_outs_1; // @[MemPrimitives.scala 121:29:@21917.4]
  wire  StickySelects_10_io_outs_2; // @[MemPrimitives.scala 121:29:@21917.4]
  wire  StickySelects_10_io_outs_3; // @[MemPrimitives.scala 121:29:@21917.4]
  wire  StickySelects_10_io_outs_4; // @[MemPrimitives.scala 121:29:@21917.4]
  wire  StickySelects_10_io_outs_5; // @[MemPrimitives.scala 121:29:@21917.4]
  wire  StickySelects_10_io_outs_6; // @[MemPrimitives.scala 121:29:@21917.4]
  wire  StickySelects_10_io_outs_7; // @[MemPrimitives.scala 121:29:@21917.4]
  wire  StickySelects_10_io_outs_8; // @[MemPrimitives.scala 121:29:@21917.4]
  wire  StickySelects_11_clock; // @[MemPrimitives.scala 121:29:@22006.4]
  wire  StickySelects_11_reset; // @[MemPrimitives.scala 121:29:@22006.4]
  wire  StickySelects_11_io_ins_0; // @[MemPrimitives.scala 121:29:@22006.4]
  wire  StickySelects_11_io_ins_1; // @[MemPrimitives.scala 121:29:@22006.4]
  wire  StickySelects_11_io_ins_2; // @[MemPrimitives.scala 121:29:@22006.4]
  wire  StickySelects_11_io_ins_3; // @[MemPrimitives.scala 121:29:@22006.4]
  wire  StickySelects_11_io_ins_4; // @[MemPrimitives.scala 121:29:@22006.4]
  wire  StickySelects_11_io_ins_5; // @[MemPrimitives.scala 121:29:@22006.4]
  wire  StickySelects_11_io_ins_6; // @[MemPrimitives.scala 121:29:@22006.4]
  wire  StickySelects_11_io_ins_7; // @[MemPrimitives.scala 121:29:@22006.4]
  wire  StickySelects_11_io_ins_8; // @[MemPrimitives.scala 121:29:@22006.4]
  wire  StickySelects_11_io_outs_0; // @[MemPrimitives.scala 121:29:@22006.4]
  wire  StickySelects_11_io_outs_1; // @[MemPrimitives.scala 121:29:@22006.4]
  wire  StickySelects_11_io_outs_2; // @[MemPrimitives.scala 121:29:@22006.4]
  wire  StickySelects_11_io_outs_3; // @[MemPrimitives.scala 121:29:@22006.4]
  wire  StickySelects_11_io_outs_4; // @[MemPrimitives.scala 121:29:@22006.4]
  wire  StickySelects_11_io_outs_5; // @[MemPrimitives.scala 121:29:@22006.4]
  wire  StickySelects_11_io_outs_6; // @[MemPrimitives.scala 121:29:@22006.4]
  wire  StickySelects_11_io_outs_7; // @[MemPrimitives.scala 121:29:@22006.4]
  wire  StickySelects_11_io_outs_8; // @[MemPrimitives.scala 121:29:@22006.4]
  wire  StickySelects_12_clock; // @[MemPrimitives.scala 121:29:@22095.4]
  wire  StickySelects_12_reset; // @[MemPrimitives.scala 121:29:@22095.4]
  wire  StickySelects_12_io_ins_0; // @[MemPrimitives.scala 121:29:@22095.4]
  wire  StickySelects_12_io_ins_1; // @[MemPrimitives.scala 121:29:@22095.4]
  wire  StickySelects_12_io_ins_2; // @[MemPrimitives.scala 121:29:@22095.4]
  wire  StickySelects_12_io_ins_3; // @[MemPrimitives.scala 121:29:@22095.4]
  wire  StickySelects_12_io_ins_4; // @[MemPrimitives.scala 121:29:@22095.4]
  wire  StickySelects_12_io_ins_5; // @[MemPrimitives.scala 121:29:@22095.4]
  wire  StickySelects_12_io_ins_6; // @[MemPrimitives.scala 121:29:@22095.4]
  wire  StickySelects_12_io_ins_7; // @[MemPrimitives.scala 121:29:@22095.4]
  wire  StickySelects_12_io_ins_8; // @[MemPrimitives.scala 121:29:@22095.4]
  wire  StickySelects_12_io_outs_0; // @[MemPrimitives.scala 121:29:@22095.4]
  wire  StickySelects_12_io_outs_1; // @[MemPrimitives.scala 121:29:@22095.4]
  wire  StickySelects_12_io_outs_2; // @[MemPrimitives.scala 121:29:@22095.4]
  wire  StickySelects_12_io_outs_3; // @[MemPrimitives.scala 121:29:@22095.4]
  wire  StickySelects_12_io_outs_4; // @[MemPrimitives.scala 121:29:@22095.4]
  wire  StickySelects_12_io_outs_5; // @[MemPrimitives.scala 121:29:@22095.4]
  wire  StickySelects_12_io_outs_6; // @[MemPrimitives.scala 121:29:@22095.4]
  wire  StickySelects_12_io_outs_7; // @[MemPrimitives.scala 121:29:@22095.4]
  wire  StickySelects_12_io_outs_8; // @[MemPrimitives.scala 121:29:@22095.4]
  wire  StickySelects_13_clock; // @[MemPrimitives.scala 121:29:@22184.4]
  wire  StickySelects_13_reset; // @[MemPrimitives.scala 121:29:@22184.4]
  wire  StickySelects_13_io_ins_0; // @[MemPrimitives.scala 121:29:@22184.4]
  wire  StickySelects_13_io_ins_1; // @[MemPrimitives.scala 121:29:@22184.4]
  wire  StickySelects_13_io_ins_2; // @[MemPrimitives.scala 121:29:@22184.4]
  wire  StickySelects_13_io_ins_3; // @[MemPrimitives.scala 121:29:@22184.4]
  wire  StickySelects_13_io_ins_4; // @[MemPrimitives.scala 121:29:@22184.4]
  wire  StickySelects_13_io_ins_5; // @[MemPrimitives.scala 121:29:@22184.4]
  wire  StickySelects_13_io_ins_6; // @[MemPrimitives.scala 121:29:@22184.4]
  wire  StickySelects_13_io_ins_7; // @[MemPrimitives.scala 121:29:@22184.4]
  wire  StickySelects_13_io_ins_8; // @[MemPrimitives.scala 121:29:@22184.4]
  wire  StickySelects_13_io_outs_0; // @[MemPrimitives.scala 121:29:@22184.4]
  wire  StickySelects_13_io_outs_1; // @[MemPrimitives.scala 121:29:@22184.4]
  wire  StickySelects_13_io_outs_2; // @[MemPrimitives.scala 121:29:@22184.4]
  wire  StickySelects_13_io_outs_3; // @[MemPrimitives.scala 121:29:@22184.4]
  wire  StickySelects_13_io_outs_4; // @[MemPrimitives.scala 121:29:@22184.4]
  wire  StickySelects_13_io_outs_5; // @[MemPrimitives.scala 121:29:@22184.4]
  wire  StickySelects_13_io_outs_6; // @[MemPrimitives.scala 121:29:@22184.4]
  wire  StickySelects_13_io_outs_7; // @[MemPrimitives.scala 121:29:@22184.4]
  wire  StickySelects_13_io_outs_8; // @[MemPrimitives.scala 121:29:@22184.4]
  wire  StickySelects_14_clock; // @[MemPrimitives.scala 121:29:@22273.4]
  wire  StickySelects_14_reset; // @[MemPrimitives.scala 121:29:@22273.4]
  wire  StickySelects_14_io_ins_0; // @[MemPrimitives.scala 121:29:@22273.4]
  wire  StickySelects_14_io_ins_1; // @[MemPrimitives.scala 121:29:@22273.4]
  wire  StickySelects_14_io_ins_2; // @[MemPrimitives.scala 121:29:@22273.4]
  wire  StickySelects_14_io_ins_3; // @[MemPrimitives.scala 121:29:@22273.4]
  wire  StickySelects_14_io_ins_4; // @[MemPrimitives.scala 121:29:@22273.4]
  wire  StickySelects_14_io_ins_5; // @[MemPrimitives.scala 121:29:@22273.4]
  wire  StickySelects_14_io_ins_6; // @[MemPrimitives.scala 121:29:@22273.4]
  wire  StickySelects_14_io_ins_7; // @[MemPrimitives.scala 121:29:@22273.4]
  wire  StickySelects_14_io_ins_8; // @[MemPrimitives.scala 121:29:@22273.4]
  wire  StickySelects_14_io_outs_0; // @[MemPrimitives.scala 121:29:@22273.4]
  wire  StickySelects_14_io_outs_1; // @[MemPrimitives.scala 121:29:@22273.4]
  wire  StickySelects_14_io_outs_2; // @[MemPrimitives.scala 121:29:@22273.4]
  wire  StickySelects_14_io_outs_3; // @[MemPrimitives.scala 121:29:@22273.4]
  wire  StickySelects_14_io_outs_4; // @[MemPrimitives.scala 121:29:@22273.4]
  wire  StickySelects_14_io_outs_5; // @[MemPrimitives.scala 121:29:@22273.4]
  wire  StickySelects_14_io_outs_6; // @[MemPrimitives.scala 121:29:@22273.4]
  wire  StickySelects_14_io_outs_7; // @[MemPrimitives.scala 121:29:@22273.4]
  wire  StickySelects_14_io_outs_8; // @[MemPrimitives.scala 121:29:@22273.4]
  wire  StickySelects_15_clock; // @[MemPrimitives.scala 121:29:@22362.4]
  wire  StickySelects_15_reset; // @[MemPrimitives.scala 121:29:@22362.4]
  wire  StickySelects_15_io_ins_0; // @[MemPrimitives.scala 121:29:@22362.4]
  wire  StickySelects_15_io_ins_1; // @[MemPrimitives.scala 121:29:@22362.4]
  wire  StickySelects_15_io_ins_2; // @[MemPrimitives.scala 121:29:@22362.4]
  wire  StickySelects_15_io_ins_3; // @[MemPrimitives.scala 121:29:@22362.4]
  wire  StickySelects_15_io_ins_4; // @[MemPrimitives.scala 121:29:@22362.4]
  wire  StickySelects_15_io_ins_5; // @[MemPrimitives.scala 121:29:@22362.4]
  wire  StickySelects_15_io_ins_6; // @[MemPrimitives.scala 121:29:@22362.4]
  wire  StickySelects_15_io_ins_7; // @[MemPrimitives.scala 121:29:@22362.4]
  wire  StickySelects_15_io_ins_8; // @[MemPrimitives.scala 121:29:@22362.4]
  wire  StickySelects_15_io_outs_0; // @[MemPrimitives.scala 121:29:@22362.4]
  wire  StickySelects_15_io_outs_1; // @[MemPrimitives.scala 121:29:@22362.4]
  wire  StickySelects_15_io_outs_2; // @[MemPrimitives.scala 121:29:@22362.4]
  wire  StickySelects_15_io_outs_3; // @[MemPrimitives.scala 121:29:@22362.4]
  wire  StickySelects_15_io_outs_4; // @[MemPrimitives.scala 121:29:@22362.4]
  wire  StickySelects_15_io_outs_5; // @[MemPrimitives.scala 121:29:@22362.4]
  wire  StickySelects_15_io_outs_6; // @[MemPrimitives.scala 121:29:@22362.4]
  wire  StickySelects_15_io_outs_7; // @[MemPrimitives.scala 121:29:@22362.4]
  wire  StickySelects_15_io_outs_8; // @[MemPrimitives.scala 121:29:@22362.4]
  wire  StickySelects_16_clock; // @[MemPrimitives.scala 121:29:@22451.4]
  wire  StickySelects_16_reset; // @[MemPrimitives.scala 121:29:@22451.4]
  wire  StickySelects_16_io_ins_0; // @[MemPrimitives.scala 121:29:@22451.4]
  wire  StickySelects_16_io_ins_1; // @[MemPrimitives.scala 121:29:@22451.4]
  wire  StickySelects_16_io_ins_2; // @[MemPrimitives.scala 121:29:@22451.4]
  wire  StickySelects_16_io_ins_3; // @[MemPrimitives.scala 121:29:@22451.4]
  wire  StickySelects_16_io_ins_4; // @[MemPrimitives.scala 121:29:@22451.4]
  wire  StickySelects_16_io_ins_5; // @[MemPrimitives.scala 121:29:@22451.4]
  wire  StickySelects_16_io_ins_6; // @[MemPrimitives.scala 121:29:@22451.4]
  wire  StickySelects_16_io_ins_7; // @[MemPrimitives.scala 121:29:@22451.4]
  wire  StickySelects_16_io_ins_8; // @[MemPrimitives.scala 121:29:@22451.4]
  wire  StickySelects_16_io_outs_0; // @[MemPrimitives.scala 121:29:@22451.4]
  wire  StickySelects_16_io_outs_1; // @[MemPrimitives.scala 121:29:@22451.4]
  wire  StickySelects_16_io_outs_2; // @[MemPrimitives.scala 121:29:@22451.4]
  wire  StickySelects_16_io_outs_3; // @[MemPrimitives.scala 121:29:@22451.4]
  wire  StickySelects_16_io_outs_4; // @[MemPrimitives.scala 121:29:@22451.4]
  wire  StickySelects_16_io_outs_5; // @[MemPrimitives.scala 121:29:@22451.4]
  wire  StickySelects_16_io_outs_6; // @[MemPrimitives.scala 121:29:@22451.4]
  wire  StickySelects_16_io_outs_7; // @[MemPrimitives.scala 121:29:@22451.4]
  wire  StickySelects_16_io_outs_8; // @[MemPrimitives.scala 121:29:@22451.4]
  wire  StickySelects_17_clock; // @[MemPrimitives.scala 121:29:@22540.4]
  wire  StickySelects_17_reset; // @[MemPrimitives.scala 121:29:@22540.4]
  wire  StickySelects_17_io_ins_0; // @[MemPrimitives.scala 121:29:@22540.4]
  wire  StickySelects_17_io_ins_1; // @[MemPrimitives.scala 121:29:@22540.4]
  wire  StickySelects_17_io_ins_2; // @[MemPrimitives.scala 121:29:@22540.4]
  wire  StickySelects_17_io_ins_3; // @[MemPrimitives.scala 121:29:@22540.4]
  wire  StickySelects_17_io_ins_4; // @[MemPrimitives.scala 121:29:@22540.4]
  wire  StickySelects_17_io_ins_5; // @[MemPrimitives.scala 121:29:@22540.4]
  wire  StickySelects_17_io_ins_6; // @[MemPrimitives.scala 121:29:@22540.4]
  wire  StickySelects_17_io_ins_7; // @[MemPrimitives.scala 121:29:@22540.4]
  wire  StickySelects_17_io_ins_8; // @[MemPrimitives.scala 121:29:@22540.4]
  wire  StickySelects_17_io_outs_0; // @[MemPrimitives.scala 121:29:@22540.4]
  wire  StickySelects_17_io_outs_1; // @[MemPrimitives.scala 121:29:@22540.4]
  wire  StickySelects_17_io_outs_2; // @[MemPrimitives.scala 121:29:@22540.4]
  wire  StickySelects_17_io_outs_3; // @[MemPrimitives.scala 121:29:@22540.4]
  wire  StickySelects_17_io_outs_4; // @[MemPrimitives.scala 121:29:@22540.4]
  wire  StickySelects_17_io_outs_5; // @[MemPrimitives.scala 121:29:@22540.4]
  wire  StickySelects_17_io_outs_6; // @[MemPrimitives.scala 121:29:@22540.4]
  wire  StickySelects_17_io_outs_7; // @[MemPrimitives.scala 121:29:@22540.4]
  wire  StickySelects_17_io_outs_8; // @[MemPrimitives.scala 121:29:@22540.4]
  wire  StickySelects_18_clock; // @[MemPrimitives.scala 121:29:@22629.4]
  wire  StickySelects_18_reset; // @[MemPrimitives.scala 121:29:@22629.4]
  wire  StickySelects_18_io_ins_0; // @[MemPrimitives.scala 121:29:@22629.4]
  wire  StickySelects_18_io_ins_1; // @[MemPrimitives.scala 121:29:@22629.4]
  wire  StickySelects_18_io_ins_2; // @[MemPrimitives.scala 121:29:@22629.4]
  wire  StickySelects_18_io_ins_3; // @[MemPrimitives.scala 121:29:@22629.4]
  wire  StickySelects_18_io_ins_4; // @[MemPrimitives.scala 121:29:@22629.4]
  wire  StickySelects_18_io_ins_5; // @[MemPrimitives.scala 121:29:@22629.4]
  wire  StickySelects_18_io_ins_6; // @[MemPrimitives.scala 121:29:@22629.4]
  wire  StickySelects_18_io_ins_7; // @[MemPrimitives.scala 121:29:@22629.4]
  wire  StickySelects_18_io_ins_8; // @[MemPrimitives.scala 121:29:@22629.4]
  wire  StickySelects_18_io_outs_0; // @[MemPrimitives.scala 121:29:@22629.4]
  wire  StickySelects_18_io_outs_1; // @[MemPrimitives.scala 121:29:@22629.4]
  wire  StickySelects_18_io_outs_2; // @[MemPrimitives.scala 121:29:@22629.4]
  wire  StickySelects_18_io_outs_3; // @[MemPrimitives.scala 121:29:@22629.4]
  wire  StickySelects_18_io_outs_4; // @[MemPrimitives.scala 121:29:@22629.4]
  wire  StickySelects_18_io_outs_5; // @[MemPrimitives.scala 121:29:@22629.4]
  wire  StickySelects_18_io_outs_6; // @[MemPrimitives.scala 121:29:@22629.4]
  wire  StickySelects_18_io_outs_7; // @[MemPrimitives.scala 121:29:@22629.4]
  wire  StickySelects_18_io_outs_8; // @[MemPrimitives.scala 121:29:@22629.4]
  wire  StickySelects_19_clock; // @[MemPrimitives.scala 121:29:@22718.4]
  wire  StickySelects_19_reset; // @[MemPrimitives.scala 121:29:@22718.4]
  wire  StickySelects_19_io_ins_0; // @[MemPrimitives.scala 121:29:@22718.4]
  wire  StickySelects_19_io_ins_1; // @[MemPrimitives.scala 121:29:@22718.4]
  wire  StickySelects_19_io_ins_2; // @[MemPrimitives.scala 121:29:@22718.4]
  wire  StickySelects_19_io_ins_3; // @[MemPrimitives.scala 121:29:@22718.4]
  wire  StickySelects_19_io_ins_4; // @[MemPrimitives.scala 121:29:@22718.4]
  wire  StickySelects_19_io_ins_5; // @[MemPrimitives.scala 121:29:@22718.4]
  wire  StickySelects_19_io_ins_6; // @[MemPrimitives.scala 121:29:@22718.4]
  wire  StickySelects_19_io_ins_7; // @[MemPrimitives.scala 121:29:@22718.4]
  wire  StickySelects_19_io_ins_8; // @[MemPrimitives.scala 121:29:@22718.4]
  wire  StickySelects_19_io_outs_0; // @[MemPrimitives.scala 121:29:@22718.4]
  wire  StickySelects_19_io_outs_1; // @[MemPrimitives.scala 121:29:@22718.4]
  wire  StickySelects_19_io_outs_2; // @[MemPrimitives.scala 121:29:@22718.4]
  wire  StickySelects_19_io_outs_3; // @[MemPrimitives.scala 121:29:@22718.4]
  wire  StickySelects_19_io_outs_4; // @[MemPrimitives.scala 121:29:@22718.4]
  wire  StickySelects_19_io_outs_5; // @[MemPrimitives.scala 121:29:@22718.4]
  wire  StickySelects_19_io_outs_6; // @[MemPrimitives.scala 121:29:@22718.4]
  wire  StickySelects_19_io_outs_7; // @[MemPrimitives.scala 121:29:@22718.4]
  wire  StickySelects_19_io_outs_8; // @[MemPrimitives.scala 121:29:@22718.4]
  wire  StickySelects_20_clock; // @[MemPrimitives.scala 121:29:@22807.4]
  wire  StickySelects_20_reset; // @[MemPrimitives.scala 121:29:@22807.4]
  wire  StickySelects_20_io_ins_0; // @[MemPrimitives.scala 121:29:@22807.4]
  wire  StickySelects_20_io_ins_1; // @[MemPrimitives.scala 121:29:@22807.4]
  wire  StickySelects_20_io_ins_2; // @[MemPrimitives.scala 121:29:@22807.4]
  wire  StickySelects_20_io_ins_3; // @[MemPrimitives.scala 121:29:@22807.4]
  wire  StickySelects_20_io_ins_4; // @[MemPrimitives.scala 121:29:@22807.4]
  wire  StickySelects_20_io_ins_5; // @[MemPrimitives.scala 121:29:@22807.4]
  wire  StickySelects_20_io_ins_6; // @[MemPrimitives.scala 121:29:@22807.4]
  wire  StickySelects_20_io_ins_7; // @[MemPrimitives.scala 121:29:@22807.4]
  wire  StickySelects_20_io_ins_8; // @[MemPrimitives.scala 121:29:@22807.4]
  wire  StickySelects_20_io_outs_0; // @[MemPrimitives.scala 121:29:@22807.4]
  wire  StickySelects_20_io_outs_1; // @[MemPrimitives.scala 121:29:@22807.4]
  wire  StickySelects_20_io_outs_2; // @[MemPrimitives.scala 121:29:@22807.4]
  wire  StickySelects_20_io_outs_3; // @[MemPrimitives.scala 121:29:@22807.4]
  wire  StickySelects_20_io_outs_4; // @[MemPrimitives.scala 121:29:@22807.4]
  wire  StickySelects_20_io_outs_5; // @[MemPrimitives.scala 121:29:@22807.4]
  wire  StickySelects_20_io_outs_6; // @[MemPrimitives.scala 121:29:@22807.4]
  wire  StickySelects_20_io_outs_7; // @[MemPrimitives.scala 121:29:@22807.4]
  wire  StickySelects_20_io_outs_8; // @[MemPrimitives.scala 121:29:@22807.4]
  wire  StickySelects_21_clock; // @[MemPrimitives.scala 121:29:@22896.4]
  wire  StickySelects_21_reset; // @[MemPrimitives.scala 121:29:@22896.4]
  wire  StickySelects_21_io_ins_0; // @[MemPrimitives.scala 121:29:@22896.4]
  wire  StickySelects_21_io_ins_1; // @[MemPrimitives.scala 121:29:@22896.4]
  wire  StickySelects_21_io_ins_2; // @[MemPrimitives.scala 121:29:@22896.4]
  wire  StickySelects_21_io_ins_3; // @[MemPrimitives.scala 121:29:@22896.4]
  wire  StickySelects_21_io_ins_4; // @[MemPrimitives.scala 121:29:@22896.4]
  wire  StickySelects_21_io_ins_5; // @[MemPrimitives.scala 121:29:@22896.4]
  wire  StickySelects_21_io_ins_6; // @[MemPrimitives.scala 121:29:@22896.4]
  wire  StickySelects_21_io_ins_7; // @[MemPrimitives.scala 121:29:@22896.4]
  wire  StickySelects_21_io_ins_8; // @[MemPrimitives.scala 121:29:@22896.4]
  wire  StickySelects_21_io_outs_0; // @[MemPrimitives.scala 121:29:@22896.4]
  wire  StickySelects_21_io_outs_1; // @[MemPrimitives.scala 121:29:@22896.4]
  wire  StickySelects_21_io_outs_2; // @[MemPrimitives.scala 121:29:@22896.4]
  wire  StickySelects_21_io_outs_3; // @[MemPrimitives.scala 121:29:@22896.4]
  wire  StickySelects_21_io_outs_4; // @[MemPrimitives.scala 121:29:@22896.4]
  wire  StickySelects_21_io_outs_5; // @[MemPrimitives.scala 121:29:@22896.4]
  wire  StickySelects_21_io_outs_6; // @[MemPrimitives.scala 121:29:@22896.4]
  wire  StickySelects_21_io_outs_7; // @[MemPrimitives.scala 121:29:@22896.4]
  wire  StickySelects_21_io_outs_8; // @[MemPrimitives.scala 121:29:@22896.4]
  wire  StickySelects_22_clock; // @[MemPrimitives.scala 121:29:@22985.4]
  wire  StickySelects_22_reset; // @[MemPrimitives.scala 121:29:@22985.4]
  wire  StickySelects_22_io_ins_0; // @[MemPrimitives.scala 121:29:@22985.4]
  wire  StickySelects_22_io_ins_1; // @[MemPrimitives.scala 121:29:@22985.4]
  wire  StickySelects_22_io_ins_2; // @[MemPrimitives.scala 121:29:@22985.4]
  wire  StickySelects_22_io_ins_3; // @[MemPrimitives.scala 121:29:@22985.4]
  wire  StickySelects_22_io_ins_4; // @[MemPrimitives.scala 121:29:@22985.4]
  wire  StickySelects_22_io_ins_5; // @[MemPrimitives.scala 121:29:@22985.4]
  wire  StickySelects_22_io_ins_6; // @[MemPrimitives.scala 121:29:@22985.4]
  wire  StickySelects_22_io_ins_7; // @[MemPrimitives.scala 121:29:@22985.4]
  wire  StickySelects_22_io_ins_8; // @[MemPrimitives.scala 121:29:@22985.4]
  wire  StickySelects_22_io_outs_0; // @[MemPrimitives.scala 121:29:@22985.4]
  wire  StickySelects_22_io_outs_1; // @[MemPrimitives.scala 121:29:@22985.4]
  wire  StickySelects_22_io_outs_2; // @[MemPrimitives.scala 121:29:@22985.4]
  wire  StickySelects_22_io_outs_3; // @[MemPrimitives.scala 121:29:@22985.4]
  wire  StickySelects_22_io_outs_4; // @[MemPrimitives.scala 121:29:@22985.4]
  wire  StickySelects_22_io_outs_5; // @[MemPrimitives.scala 121:29:@22985.4]
  wire  StickySelects_22_io_outs_6; // @[MemPrimitives.scala 121:29:@22985.4]
  wire  StickySelects_22_io_outs_7; // @[MemPrimitives.scala 121:29:@22985.4]
  wire  StickySelects_22_io_outs_8; // @[MemPrimitives.scala 121:29:@22985.4]
  wire  StickySelects_23_clock; // @[MemPrimitives.scala 121:29:@23074.4]
  wire  StickySelects_23_reset; // @[MemPrimitives.scala 121:29:@23074.4]
  wire  StickySelects_23_io_ins_0; // @[MemPrimitives.scala 121:29:@23074.4]
  wire  StickySelects_23_io_ins_1; // @[MemPrimitives.scala 121:29:@23074.4]
  wire  StickySelects_23_io_ins_2; // @[MemPrimitives.scala 121:29:@23074.4]
  wire  StickySelects_23_io_ins_3; // @[MemPrimitives.scala 121:29:@23074.4]
  wire  StickySelects_23_io_ins_4; // @[MemPrimitives.scala 121:29:@23074.4]
  wire  StickySelects_23_io_ins_5; // @[MemPrimitives.scala 121:29:@23074.4]
  wire  StickySelects_23_io_ins_6; // @[MemPrimitives.scala 121:29:@23074.4]
  wire  StickySelects_23_io_ins_7; // @[MemPrimitives.scala 121:29:@23074.4]
  wire  StickySelects_23_io_ins_8; // @[MemPrimitives.scala 121:29:@23074.4]
  wire  StickySelects_23_io_outs_0; // @[MemPrimitives.scala 121:29:@23074.4]
  wire  StickySelects_23_io_outs_1; // @[MemPrimitives.scala 121:29:@23074.4]
  wire  StickySelects_23_io_outs_2; // @[MemPrimitives.scala 121:29:@23074.4]
  wire  StickySelects_23_io_outs_3; // @[MemPrimitives.scala 121:29:@23074.4]
  wire  StickySelects_23_io_outs_4; // @[MemPrimitives.scala 121:29:@23074.4]
  wire  StickySelects_23_io_outs_5; // @[MemPrimitives.scala 121:29:@23074.4]
  wire  StickySelects_23_io_outs_6; // @[MemPrimitives.scala 121:29:@23074.4]
  wire  StickySelects_23_io_outs_7; // @[MemPrimitives.scala 121:29:@23074.4]
  wire  StickySelects_23_io_outs_8; // @[MemPrimitives.scala 121:29:@23074.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@23164.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@23164.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@23164.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@23164.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@23164.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@23172.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@23172.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@23172.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@23172.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@23172.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@23180.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@23180.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@23180.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@23180.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@23180.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@23188.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@23188.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@23188.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@23188.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@23188.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@23196.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@23196.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@23196.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@23196.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@23196.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@23204.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@23204.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@23204.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@23204.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@23204.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@23212.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@23212.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@23212.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@23212.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@23212.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@23220.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@23220.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@23220.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@23220.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@23220.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@23228.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@23228.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@23228.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@23228.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@23228.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@23236.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@23236.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@23236.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@23236.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@23236.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@23244.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@23244.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@23244.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@23244.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@23244.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@23252.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@23252.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@23252.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@23252.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@23252.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@23308.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@23308.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@23308.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@23308.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@23308.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@23316.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@23316.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@23316.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@23316.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@23316.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@23324.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@23324.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@23324.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@23324.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@23324.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@23332.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@23332.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@23332.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@23332.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@23332.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@23340.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@23340.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@23340.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@23340.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@23340.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@23348.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@23348.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@23348.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@23348.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@23348.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@23356.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@23356.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@23356.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@23356.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@23356.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@23364.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@23364.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@23364.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@23364.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@23364.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@23372.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@23372.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@23372.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@23372.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@23372.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@23380.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@23380.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@23380.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@23380.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@23380.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@23388.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@23388.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@23388.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@23388.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@23388.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@23396.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@23396.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@23396.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@23396.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@23396.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@23452.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@23452.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@23452.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@23452.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@23452.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@23460.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@23460.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@23460.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@23460.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@23460.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@23468.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@23468.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@23468.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@23468.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@23468.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@23476.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@23476.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@23476.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@23476.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@23476.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@23484.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@23484.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@23484.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@23484.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@23484.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@23492.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@23492.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@23492.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@23492.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@23492.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@23500.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@23500.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@23500.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@23500.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@23500.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@23508.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@23508.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@23508.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@23508.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@23508.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@23516.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@23516.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@23516.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@23516.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@23516.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@23524.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@23524.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@23524.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@23524.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@23524.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@23532.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@23532.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@23532.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@23532.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@23532.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@23540.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@23540.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@23540.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@23540.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@23540.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@23596.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@23596.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@23596.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@23596.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@23596.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@23604.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@23604.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@23604.4]
  wire  RetimeWrapper_37_io_in; // @[package.scala 93:22:@23604.4]
  wire  RetimeWrapper_37_io_out; // @[package.scala 93:22:@23604.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@23612.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@23612.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@23612.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@23612.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@23612.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@23620.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@23620.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@23620.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@23620.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@23620.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@23628.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@23628.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@23628.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@23628.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@23628.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@23636.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@23636.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@23636.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@23636.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@23636.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@23644.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@23644.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@23644.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@23644.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@23644.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@23652.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@23652.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@23652.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@23652.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@23652.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@23660.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@23660.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@23660.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@23660.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@23660.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@23668.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@23668.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@23668.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@23668.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@23668.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@23676.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@23676.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@23676.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@23676.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@23676.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@23684.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@23684.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@23684.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@23684.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@23684.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@23740.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@23740.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@23740.4]
  wire  RetimeWrapper_48_io_in; // @[package.scala 93:22:@23740.4]
  wire  RetimeWrapper_48_io_out; // @[package.scala 93:22:@23740.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@23748.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@23748.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@23748.4]
  wire  RetimeWrapper_49_io_in; // @[package.scala 93:22:@23748.4]
  wire  RetimeWrapper_49_io_out; // @[package.scala 93:22:@23748.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@23756.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@23756.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@23756.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@23756.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@23756.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@23764.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@23764.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@23764.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@23764.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@23764.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@23772.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@23772.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@23772.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@23772.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@23772.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@23780.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@23780.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@23780.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@23780.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@23780.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@23788.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@23788.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@23788.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@23788.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@23788.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@23796.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@23796.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@23796.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@23796.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@23796.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@23804.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@23804.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@23804.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@23804.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@23804.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@23812.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@23812.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@23812.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@23812.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@23812.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@23820.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@23820.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@23820.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@23820.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@23820.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@23828.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@23828.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@23828.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@23828.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@23828.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@23884.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@23884.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@23884.4]
  wire  RetimeWrapper_60_io_in; // @[package.scala 93:22:@23884.4]
  wire  RetimeWrapper_60_io_out; // @[package.scala 93:22:@23884.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@23892.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@23892.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@23892.4]
  wire  RetimeWrapper_61_io_in; // @[package.scala 93:22:@23892.4]
  wire  RetimeWrapper_61_io_out; // @[package.scala 93:22:@23892.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@23900.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@23900.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@23900.4]
  wire  RetimeWrapper_62_io_in; // @[package.scala 93:22:@23900.4]
  wire  RetimeWrapper_62_io_out; // @[package.scala 93:22:@23900.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@23908.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@23908.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@23908.4]
  wire  RetimeWrapper_63_io_in; // @[package.scala 93:22:@23908.4]
  wire  RetimeWrapper_63_io_out; // @[package.scala 93:22:@23908.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@23916.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@23916.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@23916.4]
  wire  RetimeWrapper_64_io_in; // @[package.scala 93:22:@23916.4]
  wire  RetimeWrapper_64_io_out; // @[package.scala 93:22:@23916.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@23924.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@23924.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@23924.4]
  wire  RetimeWrapper_65_io_in; // @[package.scala 93:22:@23924.4]
  wire  RetimeWrapper_65_io_out; // @[package.scala 93:22:@23924.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@23932.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@23932.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@23932.4]
  wire  RetimeWrapper_66_io_in; // @[package.scala 93:22:@23932.4]
  wire  RetimeWrapper_66_io_out; // @[package.scala 93:22:@23932.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@23940.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@23940.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@23940.4]
  wire  RetimeWrapper_67_io_in; // @[package.scala 93:22:@23940.4]
  wire  RetimeWrapper_67_io_out; // @[package.scala 93:22:@23940.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@23948.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@23948.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@23948.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@23948.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@23948.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@23956.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@23956.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@23956.4]
  wire  RetimeWrapper_69_io_in; // @[package.scala 93:22:@23956.4]
  wire  RetimeWrapper_69_io_out; // @[package.scala 93:22:@23956.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@23964.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@23964.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@23964.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@23964.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@23964.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@23972.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@23972.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@23972.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@23972.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@23972.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@24028.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@24028.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@24028.4]
  wire  RetimeWrapper_72_io_in; // @[package.scala 93:22:@24028.4]
  wire  RetimeWrapper_72_io_out; // @[package.scala 93:22:@24028.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@24036.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@24036.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@24036.4]
  wire  RetimeWrapper_73_io_in; // @[package.scala 93:22:@24036.4]
  wire  RetimeWrapper_73_io_out; // @[package.scala 93:22:@24036.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@24044.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@24044.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@24044.4]
  wire  RetimeWrapper_74_io_in; // @[package.scala 93:22:@24044.4]
  wire  RetimeWrapper_74_io_out; // @[package.scala 93:22:@24044.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@24052.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@24052.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@24052.4]
  wire  RetimeWrapper_75_io_in; // @[package.scala 93:22:@24052.4]
  wire  RetimeWrapper_75_io_out; // @[package.scala 93:22:@24052.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@24060.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@24060.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@24060.4]
  wire  RetimeWrapper_76_io_in; // @[package.scala 93:22:@24060.4]
  wire  RetimeWrapper_76_io_out; // @[package.scala 93:22:@24060.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@24068.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@24068.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@24068.4]
  wire  RetimeWrapper_77_io_in; // @[package.scala 93:22:@24068.4]
  wire  RetimeWrapper_77_io_out; // @[package.scala 93:22:@24068.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@24076.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@24076.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@24076.4]
  wire  RetimeWrapper_78_io_in; // @[package.scala 93:22:@24076.4]
  wire  RetimeWrapper_78_io_out; // @[package.scala 93:22:@24076.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@24084.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@24084.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@24084.4]
  wire  RetimeWrapper_79_io_in; // @[package.scala 93:22:@24084.4]
  wire  RetimeWrapper_79_io_out; // @[package.scala 93:22:@24084.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@24092.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@24092.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@24092.4]
  wire  RetimeWrapper_80_io_in; // @[package.scala 93:22:@24092.4]
  wire  RetimeWrapper_80_io_out; // @[package.scala 93:22:@24092.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@24100.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@24100.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@24100.4]
  wire  RetimeWrapper_81_io_in; // @[package.scala 93:22:@24100.4]
  wire  RetimeWrapper_81_io_out; // @[package.scala 93:22:@24100.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@24108.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@24108.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@24108.4]
  wire  RetimeWrapper_82_io_in; // @[package.scala 93:22:@24108.4]
  wire  RetimeWrapper_82_io_out; // @[package.scala 93:22:@24108.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@24116.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@24116.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@24116.4]
  wire  RetimeWrapper_83_io_in; // @[package.scala 93:22:@24116.4]
  wire  RetimeWrapper_83_io_out; // @[package.scala 93:22:@24116.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@24172.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@24172.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@24172.4]
  wire  RetimeWrapper_84_io_in; // @[package.scala 93:22:@24172.4]
  wire  RetimeWrapper_84_io_out; // @[package.scala 93:22:@24172.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@24180.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@24180.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@24180.4]
  wire  RetimeWrapper_85_io_in; // @[package.scala 93:22:@24180.4]
  wire  RetimeWrapper_85_io_out; // @[package.scala 93:22:@24180.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@24188.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@24188.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@24188.4]
  wire  RetimeWrapper_86_io_in; // @[package.scala 93:22:@24188.4]
  wire  RetimeWrapper_86_io_out; // @[package.scala 93:22:@24188.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@24196.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@24196.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@24196.4]
  wire  RetimeWrapper_87_io_in; // @[package.scala 93:22:@24196.4]
  wire  RetimeWrapper_87_io_out; // @[package.scala 93:22:@24196.4]
  wire  RetimeWrapper_88_clock; // @[package.scala 93:22:@24204.4]
  wire  RetimeWrapper_88_reset; // @[package.scala 93:22:@24204.4]
  wire  RetimeWrapper_88_io_flow; // @[package.scala 93:22:@24204.4]
  wire  RetimeWrapper_88_io_in; // @[package.scala 93:22:@24204.4]
  wire  RetimeWrapper_88_io_out; // @[package.scala 93:22:@24204.4]
  wire  RetimeWrapper_89_clock; // @[package.scala 93:22:@24212.4]
  wire  RetimeWrapper_89_reset; // @[package.scala 93:22:@24212.4]
  wire  RetimeWrapper_89_io_flow; // @[package.scala 93:22:@24212.4]
  wire  RetimeWrapper_89_io_in; // @[package.scala 93:22:@24212.4]
  wire  RetimeWrapper_89_io_out; // @[package.scala 93:22:@24212.4]
  wire  RetimeWrapper_90_clock; // @[package.scala 93:22:@24220.4]
  wire  RetimeWrapper_90_reset; // @[package.scala 93:22:@24220.4]
  wire  RetimeWrapper_90_io_flow; // @[package.scala 93:22:@24220.4]
  wire  RetimeWrapper_90_io_in; // @[package.scala 93:22:@24220.4]
  wire  RetimeWrapper_90_io_out; // @[package.scala 93:22:@24220.4]
  wire  RetimeWrapper_91_clock; // @[package.scala 93:22:@24228.4]
  wire  RetimeWrapper_91_reset; // @[package.scala 93:22:@24228.4]
  wire  RetimeWrapper_91_io_flow; // @[package.scala 93:22:@24228.4]
  wire  RetimeWrapper_91_io_in; // @[package.scala 93:22:@24228.4]
  wire  RetimeWrapper_91_io_out; // @[package.scala 93:22:@24228.4]
  wire  RetimeWrapper_92_clock; // @[package.scala 93:22:@24236.4]
  wire  RetimeWrapper_92_reset; // @[package.scala 93:22:@24236.4]
  wire  RetimeWrapper_92_io_flow; // @[package.scala 93:22:@24236.4]
  wire  RetimeWrapper_92_io_in; // @[package.scala 93:22:@24236.4]
  wire  RetimeWrapper_92_io_out; // @[package.scala 93:22:@24236.4]
  wire  RetimeWrapper_93_clock; // @[package.scala 93:22:@24244.4]
  wire  RetimeWrapper_93_reset; // @[package.scala 93:22:@24244.4]
  wire  RetimeWrapper_93_io_flow; // @[package.scala 93:22:@24244.4]
  wire  RetimeWrapper_93_io_in; // @[package.scala 93:22:@24244.4]
  wire  RetimeWrapper_93_io_out; // @[package.scala 93:22:@24244.4]
  wire  RetimeWrapper_94_clock; // @[package.scala 93:22:@24252.4]
  wire  RetimeWrapper_94_reset; // @[package.scala 93:22:@24252.4]
  wire  RetimeWrapper_94_io_flow; // @[package.scala 93:22:@24252.4]
  wire  RetimeWrapper_94_io_in; // @[package.scala 93:22:@24252.4]
  wire  RetimeWrapper_94_io_out; // @[package.scala 93:22:@24252.4]
  wire  RetimeWrapper_95_clock; // @[package.scala 93:22:@24260.4]
  wire  RetimeWrapper_95_reset; // @[package.scala 93:22:@24260.4]
  wire  RetimeWrapper_95_io_flow; // @[package.scala 93:22:@24260.4]
  wire  RetimeWrapper_95_io_in; // @[package.scala 93:22:@24260.4]
  wire  RetimeWrapper_95_io_out; // @[package.scala 93:22:@24260.4]
  wire  RetimeWrapper_96_clock; // @[package.scala 93:22:@24316.4]
  wire  RetimeWrapper_96_reset; // @[package.scala 93:22:@24316.4]
  wire  RetimeWrapper_96_io_flow; // @[package.scala 93:22:@24316.4]
  wire  RetimeWrapper_96_io_in; // @[package.scala 93:22:@24316.4]
  wire  RetimeWrapper_96_io_out; // @[package.scala 93:22:@24316.4]
  wire  RetimeWrapper_97_clock; // @[package.scala 93:22:@24324.4]
  wire  RetimeWrapper_97_reset; // @[package.scala 93:22:@24324.4]
  wire  RetimeWrapper_97_io_flow; // @[package.scala 93:22:@24324.4]
  wire  RetimeWrapper_97_io_in; // @[package.scala 93:22:@24324.4]
  wire  RetimeWrapper_97_io_out; // @[package.scala 93:22:@24324.4]
  wire  RetimeWrapper_98_clock; // @[package.scala 93:22:@24332.4]
  wire  RetimeWrapper_98_reset; // @[package.scala 93:22:@24332.4]
  wire  RetimeWrapper_98_io_flow; // @[package.scala 93:22:@24332.4]
  wire  RetimeWrapper_98_io_in; // @[package.scala 93:22:@24332.4]
  wire  RetimeWrapper_98_io_out; // @[package.scala 93:22:@24332.4]
  wire  RetimeWrapper_99_clock; // @[package.scala 93:22:@24340.4]
  wire  RetimeWrapper_99_reset; // @[package.scala 93:22:@24340.4]
  wire  RetimeWrapper_99_io_flow; // @[package.scala 93:22:@24340.4]
  wire  RetimeWrapper_99_io_in; // @[package.scala 93:22:@24340.4]
  wire  RetimeWrapper_99_io_out; // @[package.scala 93:22:@24340.4]
  wire  RetimeWrapper_100_clock; // @[package.scala 93:22:@24348.4]
  wire  RetimeWrapper_100_reset; // @[package.scala 93:22:@24348.4]
  wire  RetimeWrapper_100_io_flow; // @[package.scala 93:22:@24348.4]
  wire  RetimeWrapper_100_io_in; // @[package.scala 93:22:@24348.4]
  wire  RetimeWrapper_100_io_out; // @[package.scala 93:22:@24348.4]
  wire  RetimeWrapper_101_clock; // @[package.scala 93:22:@24356.4]
  wire  RetimeWrapper_101_reset; // @[package.scala 93:22:@24356.4]
  wire  RetimeWrapper_101_io_flow; // @[package.scala 93:22:@24356.4]
  wire  RetimeWrapper_101_io_in; // @[package.scala 93:22:@24356.4]
  wire  RetimeWrapper_101_io_out; // @[package.scala 93:22:@24356.4]
  wire  RetimeWrapper_102_clock; // @[package.scala 93:22:@24364.4]
  wire  RetimeWrapper_102_reset; // @[package.scala 93:22:@24364.4]
  wire  RetimeWrapper_102_io_flow; // @[package.scala 93:22:@24364.4]
  wire  RetimeWrapper_102_io_in; // @[package.scala 93:22:@24364.4]
  wire  RetimeWrapper_102_io_out; // @[package.scala 93:22:@24364.4]
  wire  RetimeWrapper_103_clock; // @[package.scala 93:22:@24372.4]
  wire  RetimeWrapper_103_reset; // @[package.scala 93:22:@24372.4]
  wire  RetimeWrapper_103_io_flow; // @[package.scala 93:22:@24372.4]
  wire  RetimeWrapper_103_io_in; // @[package.scala 93:22:@24372.4]
  wire  RetimeWrapper_103_io_out; // @[package.scala 93:22:@24372.4]
  wire  RetimeWrapper_104_clock; // @[package.scala 93:22:@24380.4]
  wire  RetimeWrapper_104_reset; // @[package.scala 93:22:@24380.4]
  wire  RetimeWrapper_104_io_flow; // @[package.scala 93:22:@24380.4]
  wire  RetimeWrapper_104_io_in; // @[package.scala 93:22:@24380.4]
  wire  RetimeWrapper_104_io_out; // @[package.scala 93:22:@24380.4]
  wire  RetimeWrapper_105_clock; // @[package.scala 93:22:@24388.4]
  wire  RetimeWrapper_105_reset; // @[package.scala 93:22:@24388.4]
  wire  RetimeWrapper_105_io_flow; // @[package.scala 93:22:@24388.4]
  wire  RetimeWrapper_105_io_in; // @[package.scala 93:22:@24388.4]
  wire  RetimeWrapper_105_io_out; // @[package.scala 93:22:@24388.4]
  wire  RetimeWrapper_106_clock; // @[package.scala 93:22:@24396.4]
  wire  RetimeWrapper_106_reset; // @[package.scala 93:22:@24396.4]
  wire  RetimeWrapper_106_io_flow; // @[package.scala 93:22:@24396.4]
  wire  RetimeWrapper_106_io_in; // @[package.scala 93:22:@24396.4]
  wire  RetimeWrapper_106_io_out; // @[package.scala 93:22:@24396.4]
  wire  RetimeWrapper_107_clock; // @[package.scala 93:22:@24404.4]
  wire  RetimeWrapper_107_reset; // @[package.scala 93:22:@24404.4]
  wire  RetimeWrapper_107_io_flow; // @[package.scala 93:22:@24404.4]
  wire  RetimeWrapper_107_io_in; // @[package.scala 93:22:@24404.4]
  wire  RetimeWrapper_107_io_out; // @[package.scala 93:22:@24404.4]
  wire  RetimeWrapper_108_clock; // @[package.scala 93:22:@24460.4]
  wire  RetimeWrapper_108_reset; // @[package.scala 93:22:@24460.4]
  wire  RetimeWrapper_108_io_flow; // @[package.scala 93:22:@24460.4]
  wire  RetimeWrapper_108_io_in; // @[package.scala 93:22:@24460.4]
  wire  RetimeWrapper_108_io_out; // @[package.scala 93:22:@24460.4]
  wire  RetimeWrapper_109_clock; // @[package.scala 93:22:@24468.4]
  wire  RetimeWrapper_109_reset; // @[package.scala 93:22:@24468.4]
  wire  RetimeWrapper_109_io_flow; // @[package.scala 93:22:@24468.4]
  wire  RetimeWrapper_109_io_in; // @[package.scala 93:22:@24468.4]
  wire  RetimeWrapper_109_io_out; // @[package.scala 93:22:@24468.4]
  wire  RetimeWrapper_110_clock; // @[package.scala 93:22:@24476.4]
  wire  RetimeWrapper_110_reset; // @[package.scala 93:22:@24476.4]
  wire  RetimeWrapper_110_io_flow; // @[package.scala 93:22:@24476.4]
  wire  RetimeWrapper_110_io_in; // @[package.scala 93:22:@24476.4]
  wire  RetimeWrapper_110_io_out; // @[package.scala 93:22:@24476.4]
  wire  RetimeWrapper_111_clock; // @[package.scala 93:22:@24484.4]
  wire  RetimeWrapper_111_reset; // @[package.scala 93:22:@24484.4]
  wire  RetimeWrapper_111_io_flow; // @[package.scala 93:22:@24484.4]
  wire  RetimeWrapper_111_io_in; // @[package.scala 93:22:@24484.4]
  wire  RetimeWrapper_111_io_out; // @[package.scala 93:22:@24484.4]
  wire  RetimeWrapper_112_clock; // @[package.scala 93:22:@24492.4]
  wire  RetimeWrapper_112_reset; // @[package.scala 93:22:@24492.4]
  wire  RetimeWrapper_112_io_flow; // @[package.scala 93:22:@24492.4]
  wire  RetimeWrapper_112_io_in; // @[package.scala 93:22:@24492.4]
  wire  RetimeWrapper_112_io_out; // @[package.scala 93:22:@24492.4]
  wire  RetimeWrapper_113_clock; // @[package.scala 93:22:@24500.4]
  wire  RetimeWrapper_113_reset; // @[package.scala 93:22:@24500.4]
  wire  RetimeWrapper_113_io_flow; // @[package.scala 93:22:@24500.4]
  wire  RetimeWrapper_113_io_in; // @[package.scala 93:22:@24500.4]
  wire  RetimeWrapper_113_io_out; // @[package.scala 93:22:@24500.4]
  wire  RetimeWrapper_114_clock; // @[package.scala 93:22:@24508.4]
  wire  RetimeWrapper_114_reset; // @[package.scala 93:22:@24508.4]
  wire  RetimeWrapper_114_io_flow; // @[package.scala 93:22:@24508.4]
  wire  RetimeWrapper_114_io_in; // @[package.scala 93:22:@24508.4]
  wire  RetimeWrapper_114_io_out; // @[package.scala 93:22:@24508.4]
  wire  RetimeWrapper_115_clock; // @[package.scala 93:22:@24516.4]
  wire  RetimeWrapper_115_reset; // @[package.scala 93:22:@24516.4]
  wire  RetimeWrapper_115_io_flow; // @[package.scala 93:22:@24516.4]
  wire  RetimeWrapper_115_io_in; // @[package.scala 93:22:@24516.4]
  wire  RetimeWrapper_115_io_out; // @[package.scala 93:22:@24516.4]
  wire  RetimeWrapper_116_clock; // @[package.scala 93:22:@24524.4]
  wire  RetimeWrapper_116_reset; // @[package.scala 93:22:@24524.4]
  wire  RetimeWrapper_116_io_flow; // @[package.scala 93:22:@24524.4]
  wire  RetimeWrapper_116_io_in; // @[package.scala 93:22:@24524.4]
  wire  RetimeWrapper_116_io_out; // @[package.scala 93:22:@24524.4]
  wire  RetimeWrapper_117_clock; // @[package.scala 93:22:@24532.4]
  wire  RetimeWrapper_117_reset; // @[package.scala 93:22:@24532.4]
  wire  RetimeWrapper_117_io_flow; // @[package.scala 93:22:@24532.4]
  wire  RetimeWrapper_117_io_in; // @[package.scala 93:22:@24532.4]
  wire  RetimeWrapper_117_io_out; // @[package.scala 93:22:@24532.4]
  wire  RetimeWrapper_118_clock; // @[package.scala 93:22:@24540.4]
  wire  RetimeWrapper_118_reset; // @[package.scala 93:22:@24540.4]
  wire  RetimeWrapper_118_io_flow; // @[package.scala 93:22:@24540.4]
  wire  RetimeWrapper_118_io_in; // @[package.scala 93:22:@24540.4]
  wire  RetimeWrapper_118_io_out; // @[package.scala 93:22:@24540.4]
  wire  RetimeWrapper_119_clock; // @[package.scala 93:22:@24548.4]
  wire  RetimeWrapper_119_reset; // @[package.scala 93:22:@24548.4]
  wire  RetimeWrapper_119_io_flow; // @[package.scala 93:22:@24548.4]
  wire  RetimeWrapper_119_io_in; // @[package.scala 93:22:@24548.4]
  wire  RetimeWrapper_119_io_out; // @[package.scala 93:22:@24548.4]
  wire  RetimeWrapper_120_clock; // @[package.scala 93:22:@24604.4]
  wire  RetimeWrapper_120_reset; // @[package.scala 93:22:@24604.4]
  wire  RetimeWrapper_120_io_flow; // @[package.scala 93:22:@24604.4]
  wire  RetimeWrapper_120_io_in; // @[package.scala 93:22:@24604.4]
  wire  RetimeWrapper_120_io_out; // @[package.scala 93:22:@24604.4]
  wire  RetimeWrapper_121_clock; // @[package.scala 93:22:@24612.4]
  wire  RetimeWrapper_121_reset; // @[package.scala 93:22:@24612.4]
  wire  RetimeWrapper_121_io_flow; // @[package.scala 93:22:@24612.4]
  wire  RetimeWrapper_121_io_in; // @[package.scala 93:22:@24612.4]
  wire  RetimeWrapper_121_io_out; // @[package.scala 93:22:@24612.4]
  wire  RetimeWrapper_122_clock; // @[package.scala 93:22:@24620.4]
  wire  RetimeWrapper_122_reset; // @[package.scala 93:22:@24620.4]
  wire  RetimeWrapper_122_io_flow; // @[package.scala 93:22:@24620.4]
  wire  RetimeWrapper_122_io_in; // @[package.scala 93:22:@24620.4]
  wire  RetimeWrapper_122_io_out; // @[package.scala 93:22:@24620.4]
  wire  RetimeWrapper_123_clock; // @[package.scala 93:22:@24628.4]
  wire  RetimeWrapper_123_reset; // @[package.scala 93:22:@24628.4]
  wire  RetimeWrapper_123_io_flow; // @[package.scala 93:22:@24628.4]
  wire  RetimeWrapper_123_io_in; // @[package.scala 93:22:@24628.4]
  wire  RetimeWrapper_123_io_out; // @[package.scala 93:22:@24628.4]
  wire  RetimeWrapper_124_clock; // @[package.scala 93:22:@24636.4]
  wire  RetimeWrapper_124_reset; // @[package.scala 93:22:@24636.4]
  wire  RetimeWrapper_124_io_flow; // @[package.scala 93:22:@24636.4]
  wire  RetimeWrapper_124_io_in; // @[package.scala 93:22:@24636.4]
  wire  RetimeWrapper_124_io_out; // @[package.scala 93:22:@24636.4]
  wire  RetimeWrapper_125_clock; // @[package.scala 93:22:@24644.4]
  wire  RetimeWrapper_125_reset; // @[package.scala 93:22:@24644.4]
  wire  RetimeWrapper_125_io_flow; // @[package.scala 93:22:@24644.4]
  wire  RetimeWrapper_125_io_in; // @[package.scala 93:22:@24644.4]
  wire  RetimeWrapper_125_io_out; // @[package.scala 93:22:@24644.4]
  wire  RetimeWrapper_126_clock; // @[package.scala 93:22:@24652.4]
  wire  RetimeWrapper_126_reset; // @[package.scala 93:22:@24652.4]
  wire  RetimeWrapper_126_io_flow; // @[package.scala 93:22:@24652.4]
  wire  RetimeWrapper_126_io_in; // @[package.scala 93:22:@24652.4]
  wire  RetimeWrapper_126_io_out; // @[package.scala 93:22:@24652.4]
  wire  RetimeWrapper_127_clock; // @[package.scala 93:22:@24660.4]
  wire  RetimeWrapper_127_reset; // @[package.scala 93:22:@24660.4]
  wire  RetimeWrapper_127_io_flow; // @[package.scala 93:22:@24660.4]
  wire  RetimeWrapper_127_io_in; // @[package.scala 93:22:@24660.4]
  wire  RetimeWrapper_127_io_out; // @[package.scala 93:22:@24660.4]
  wire  RetimeWrapper_128_clock; // @[package.scala 93:22:@24668.4]
  wire  RetimeWrapper_128_reset; // @[package.scala 93:22:@24668.4]
  wire  RetimeWrapper_128_io_flow; // @[package.scala 93:22:@24668.4]
  wire  RetimeWrapper_128_io_in; // @[package.scala 93:22:@24668.4]
  wire  RetimeWrapper_128_io_out; // @[package.scala 93:22:@24668.4]
  wire  RetimeWrapper_129_clock; // @[package.scala 93:22:@24676.4]
  wire  RetimeWrapper_129_reset; // @[package.scala 93:22:@24676.4]
  wire  RetimeWrapper_129_io_flow; // @[package.scala 93:22:@24676.4]
  wire  RetimeWrapper_129_io_in; // @[package.scala 93:22:@24676.4]
  wire  RetimeWrapper_129_io_out; // @[package.scala 93:22:@24676.4]
  wire  RetimeWrapper_130_clock; // @[package.scala 93:22:@24684.4]
  wire  RetimeWrapper_130_reset; // @[package.scala 93:22:@24684.4]
  wire  RetimeWrapper_130_io_flow; // @[package.scala 93:22:@24684.4]
  wire  RetimeWrapper_130_io_in; // @[package.scala 93:22:@24684.4]
  wire  RetimeWrapper_130_io_out; // @[package.scala 93:22:@24684.4]
  wire  RetimeWrapper_131_clock; // @[package.scala 93:22:@24692.4]
  wire  RetimeWrapper_131_reset; // @[package.scala 93:22:@24692.4]
  wire  RetimeWrapper_131_io_flow; // @[package.scala 93:22:@24692.4]
  wire  RetimeWrapper_131_io_in; // @[package.scala 93:22:@24692.4]
  wire  RetimeWrapper_131_io_out; // @[package.scala 93:22:@24692.4]
  wire  RetimeWrapper_132_clock; // @[package.scala 93:22:@24748.4]
  wire  RetimeWrapper_132_reset; // @[package.scala 93:22:@24748.4]
  wire  RetimeWrapper_132_io_flow; // @[package.scala 93:22:@24748.4]
  wire  RetimeWrapper_132_io_in; // @[package.scala 93:22:@24748.4]
  wire  RetimeWrapper_132_io_out; // @[package.scala 93:22:@24748.4]
  wire  RetimeWrapper_133_clock; // @[package.scala 93:22:@24756.4]
  wire  RetimeWrapper_133_reset; // @[package.scala 93:22:@24756.4]
  wire  RetimeWrapper_133_io_flow; // @[package.scala 93:22:@24756.4]
  wire  RetimeWrapper_133_io_in; // @[package.scala 93:22:@24756.4]
  wire  RetimeWrapper_133_io_out; // @[package.scala 93:22:@24756.4]
  wire  RetimeWrapper_134_clock; // @[package.scala 93:22:@24764.4]
  wire  RetimeWrapper_134_reset; // @[package.scala 93:22:@24764.4]
  wire  RetimeWrapper_134_io_flow; // @[package.scala 93:22:@24764.4]
  wire  RetimeWrapper_134_io_in; // @[package.scala 93:22:@24764.4]
  wire  RetimeWrapper_134_io_out; // @[package.scala 93:22:@24764.4]
  wire  RetimeWrapper_135_clock; // @[package.scala 93:22:@24772.4]
  wire  RetimeWrapper_135_reset; // @[package.scala 93:22:@24772.4]
  wire  RetimeWrapper_135_io_flow; // @[package.scala 93:22:@24772.4]
  wire  RetimeWrapper_135_io_in; // @[package.scala 93:22:@24772.4]
  wire  RetimeWrapper_135_io_out; // @[package.scala 93:22:@24772.4]
  wire  RetimeWrapper_136_clock; // @[package.scala 93:22:@24780.4]
  wire  RetimeWrapper_136_reset; // @[package.scala 93:22:@24780.4]
  wire  RetimeWrapper_136_io_flow; // @[package.scala 93:22:@24780.4]
  wire  RetimeWrapper_136_io_in; // @[package.scala 93:22:@24780.4]
  wire  RetimeWrapper_136_io_out; // @[package.scala 93:22:@24780.4]
  wire  RetimeWrapper_137_clock; // @[package.scala 93:22:@24788.4]
  wire  RetimeWrapper_137_reset; // @[package.scala 93:22:@24788.4]
  wire  RetimeWrapper_137_io_flow; // @[package.scala 93:22:@24788.4]
  wire  RetimeWrapper_137_io_in; // @[package.scala 93:22:@24788.4]
  wire  RetimeWrapper_137_io_out; // @[package.scala 93:22:@24788.4]
  wire  RetimeWrapper_138_clock; // @[package.scala 93:22:@24796.4]
  wire  RetimeWrapper_138_reset; // @[package.scala 93:22:@24796.4]
  wire  RetimeWrapper_138_io_flow; // @[package.scala 93:22:@24796.4]
  wire  RetimeWrapper_138_io_in; // @[package.scala 93:22:@24796.4]
  wire  RetimeWrapper_138_io_out; // @[package.scala 93:22:@24796.4]
  wire  RetimeWrapper_139_clock; // @[package.scala 93:22:@24804.4]
  wire  RetimeWrapper_139_reset; // @[package.scala 93:22:@24804.4]
  wire  RetimeWrapper_139_io_flow; // @[package.scala 93:22:@24804.4]
  wire  RetimeWrapper_139_io_in; // @[package.scala 93:22:@24804.4]
  wire  RetimeWrapper_139_io_out; // @[package.scala 93:22:@24804.4]
  wire  RetimeWrapper_140_clock; // @[package.scala 93:22:@24812.4]
  wire  RetimeWrapper_140_reset; // @[package.scala 93:22:@24812.4]
  wire  RetimeWrapper_140_io_flow; // @[package.scala 93:22:@24812.4]
  wire  RetimeWrapper_140_io_in; // @[package.scala 93:22:@24812.4]
  wire  RetimeWrapper_140_io_out; // @[package.scala 93:22:@24812.4]
  wire  RetimeWrapper_141_clock; // @[package.scala 93:22:@24820.4]
  wire  RetimeWrapper_141_reset; // @[package.scala 93:22:@24820.4]
  wire  RetimeWrapper_141_io_flow; // @[package.scala 93:22:@24820.4]
  wire  RetimeWrapper_141_io_in; // @[package.scala 93:22:@24820.4]
  wire  RetimeWrapper_141_io_out; // @[package.scala 93:22:@24820.4]
  wire  RetimeWrapper_142_clock; // @[package.scala 93:22:@24828.4]
  wire  RetimeWrapper_142_reset; // @[package.scala 93:22:@24828.4]
  wire  RetimeWrapper_142_io_flow; // @[package.scala 93:22:@24828.4]
  wire  RetimeWrapper_142_io_in; // @[package.scala 93:22:@24828.4]
  wire  RetimeWrapper_142_io_out; // @[package.scala 93:22:@24828.4]
  wire  RetimeWrapper_143_clock; // @[package.scala 93:22:@24836.4]
  wire  RetimeWrapper_143_reset; // @[package.scala 93:22:@24836.4]
  wire  RetimeWrapper_143_io_flow; // @[package.scala 93:22:@24836.4]
  wire  RetimeWrapper_143_io_in; // @[package.scala 93:22:@24836.4]
  wire  RetimeWrapper_143_io_out; // @[package.scala 93:22:@24836.4]
  wire  RetimeWrapper_144_clock; // @[package.scala 93:22:@24892.4]
  wire  RetimeWrapper_144_reset; // @[package.scala 93:22:@24892.4]
  wire  RetimeWrapper_144_io_flow; // @[package.scala 93:22:@24892.4]
  wire  RetimeWrapper_144_io_in; // @[package.scala 93:22:@24892.4]
  wire  RetimeWrapper_144_io_out; // @[package.scala 93:22:@24892.4]
  wire  RetimeWrapper_145_clock; // @[package.scala 93:22:@24900.4]
  wire  RetimeWrapper_145_reset; // @[package.scala 93:22:@24900.4]
  wire  RetimeWrapper_145_io_flow; // @[package.scala 93:22:@24900.4]
  wire  RetimeWrapper_145_io_in; // @[package.scala 93:22:@24900.4]
  wire  RetimeWrapper_145_io_out; // @[package.scala 93:22:@24900.4]
  wire  RetimeWrapper_146_clock; // @[package.scala 93:22:@24908.4]
  wire  RetimeWrapper_146_reset; // @[package.scala 93:22:@24908.4]
  wire  RetimeWrapper_146_io_flow; // @[package.scala 93:22:@24908.4]
  wire  RetimeWrapper_146_io_in; // @[package.scala 93:22:@24908.4]
  wire  RetimeWrapper_146_io_out; // @[package.scala 93:22:@24908.4]
  wire  RetimeWrapper_147_clock; // @[package.scala 93:22:@24916.4]
  wire  RetimeWrapper_147_reset; // @[package.scala 93:22:@24916.4]
  wire  RetimeWrapper_147_io_flow; // @[package.scala 93:22:@24916.4]
  wire  RetimeWrapper_147_io_in; // @[package.scala 93:22:@24916.4]
  wire  RetimeWrapper_147_io_out; // @[package.scala 93:22:@24916.4]
  wire  RetimeWrapper_148_clock; // @[package.scala 93:22:@24924.4]
  wire  RetimeWrapper_148_reset; // @[package.scala 93:22:@24924.4]
  wire  RetimeWrapper_148_io_flow; // @[package.scala 93:22:@24924.4]
  wire  RetimeWrapper_148_io_in; // @[package.scala 93:22:@24924.4]
  wire  RetimeWrapper_148_io_out; // @[package.scala 93:22:@24924.4]
  wire  RetimeWrapper_149_clock; // @[package.scala 93:22:@24932.4]
  wire  RetimeWrapper_149_reset; // @[package.scala 93:22:@24932.4]
  wire  RetimeWrapper_149_io_flow; // @[package.scala 93:22:@24932.4]
  wire  RetimeWrapper_149_io_in; // @[package.scala 93:22:@24932.4]
  wire  RetimeWrapper_149_io_out; // @[package.scala 93:22:@24932.4]
  wire  RetimeWrapper_150_clock; // @[package.scala 93:22:@24940.4]
  wire  RetimeWrapper_150_reset; // @[package.scala 93:22:@24940.4]
  wire  RetimeWrapper_150_io_flow; // @[package.scala 93:22:@24940.4]
  wire  RetimeWrapper_150_io_in; // @[package.scala 93:22:@24940.4]
  wire  RetimeWrapper_150_io_out; // @[package.scala 93:22:@24940.4]
  wire  RetimeWrapper_151_clock; // @[package.scala 93:22:@24948.4]
  wire  RetimeWrapper_151_reset; // @[package.scala 93:22:@24948.4]
  wire  RetimeWrapper_151_io_flow; // @[package.scala 93:22:@24948.4]
  wire  RetimeWrapper_151_io_in; // @[package.scala 93:22:@24948.4]
  wire  RetimeWrapper_151_io_out; // @[package.scala 93:22:@24948.4]
  wire  RetimeWrapper_152_clock; // @[package.scala 93:22:@24956.4]
  wire  RetimeWrapper_152_reset; // @[package.scala 93:22:@24956.4]
  wire  RetimeWrapper_152_io_flow; // @[package.scala 93:22:@24956.4]
  wire  RetimeWrapper_152_io_in; // @[package.scala 93:22:@24956.4]
  wire  RetimeWrapper_152_io_out; // @[package.scala 93:22:@24956.4]
  wire  RetimeWrapper_153_clock; // @[package.scala 93:22:@24964.4]
  wire  RetimeWrapper_153_reset; // @[package.scala 93:22:@24964.4]
  wire  RetimeWrapper_153_io_flow; // @[package.scala 93:22:@24964.4]
  wire  RetimeWrapper_153_io_in; // @[package.scala 93:22:@24964.4]
  wire  RetimeWrapper_153_io_out; // @[package.scala 93:22:@24964.4]
  wire  RetimeWrapper_154_clock; // @[package.scala 93:22:@24972.4]
  wire  RetimeWrapper_154_reset; // @[package.scala 93:22:@24972.4]
  wire  RetimeWrapper_154_io_flow; // @[package.scala 93:22:@24972.4]
  wire  RetimeWrapper_154_io_in; // @[package.scala 93:22:@24972.4]
  wire  RetimeWrapper_154_io_out; // @[package.scala 93:22:@24972.4]
  wire  RetimeWrapper_155_clock; // @[package.scala 93:22:@24980.4]
  wire  RetimeWrapper_155_reset; // @[package.scala 93:22:@24980.4]
  wire  RetimeWrapper_155_io_flow; // @[package.scala 93:22:@24980.4]
  wire  RetimeWrapper_155_io_in; // @[package.scala 93:22:@24980.4]
  wire  RetimeWrapper_155_io_out; // @[package.scala 93:22:@24980.4]
  wire  RetimeWrapper_156_clock; // @[package.scala 93:22:@25036.4]
  wire  RetimeWrapper_156_reset; // @[package.scala 93:22:@25036.4]
  wire  RetimeWrapper_156_io_flow; // @[package.scala 93:22:@25036.4]
  wire  RetimeWrapper_156_io_in; // @[package.scala 93:22:@25036.4]
  wire  RetimeWrapper_156_io_out; // @[package.scala 93:22:@25036.4]
  wire  RetimeWrapper_157_clock; // @[package.scala 93:22:@25044.4]
  wire  RetimeWrapper_157_reset; // @[package.scala 93:22:@25044.4]
  wire  RetimeWrapper_157_io_flow; // @[package.scala 93:22:@25044.4]
  wire  RetimeWrapper_157_io_in; // @[package.scala 93:22:@25044.4]
  wire  RetimeWrapper_157_io_out; // @[package.scala 93:22:@25044.4]
  wire  RetimeWrapper_158_clock; // @[package.scala 93:22:@25052.4]
  wire  RetimeWrapper_158_reset; // @[package.scala 93:22:@25052.4]
  wire  RetimeWrapper_158_io_flow; // @[package.scala 93:22:@25052.4]
  wire  RetimeWrapper_158_io_in; // @[package.scala 93:22:@25052.4]
  wire  RetimeWrapper_158_io_out; // @[package.scala 93:22:@25052.4]
  wire  RetimeWrapper_159_clock; // @[package.scala 93:22:@25060.4]
  wire  RetimeWrapper_159_reset; // @[package.scala 93:22:@25060.4]
  wire  RetimeWrapper_159_io_flow; // @[package.scala 93:22:@25060.4]
  wire  RetimeWrapper_159_io_in; // @[package.scala 93:22:@25060.4]
  wire  RetimeWrapper_159_io_out; // @[package.scala 93:22:@25060.4]
  wire  RetimeWrapper_160_clock; // @[package.scala 93:22:@25068.4]
  wire  RetimeWrapper_160_reset; // @[package.scala 93:22:@25068.4]
  wire  RetimeWrapper_160_io_flow; // @[package.scala 93:22:@25068.4]
  wire  RetimeWrapper_160_io_in; // @[package.scala 93:22:@25068.4]
  wire  RetimeWrapper_160_io_out; // @[package.scala 93:22:@25068.4]
  wire  RetimeWrapper_161_clock; // @[package.scala 93:22:@25076.4]
  wire  RetimeWrapper_161_reset; // @[package.scala 93:22:@25076.4]
  wire  RetimeWrapper_161_io_flow; // @[package.scala 93:22:@25076.4]
  wire  RetimeWrapper_161_io_in; // @[package.scala 93:22:@25076.4]
  wire  RetimeWrapper_161_io_out; // @[package.scala 93:22:@25076.4]
  wire  RetimeWrapper_162_clock; // @[package.scala 93:22:@25084.4]
  wire  RetimeWrapper_162_reset; // @[package.scala 93:22:@25084.4]
  wire  RetimeWrapper_162_io_flow; // @[package.scala 93:22:@25084.4]
  wire  RetimeWrapper_162_io_in; // @[package.scala 93:22:@25084.4]
  wire  RetimeWrapper_162_io_out; // @[package.scala 93:22:@25084.4]
  wire  RetimeWrapper_163_clock; // @[package.scala 93:22:@25092.4]
  wire  RetimeWrapper_163_reset; // @[package.scala 93:22:@25092.4]
  wire  RetimeWrapper_163_io_flow; // @[package.scala 93:22:@25092.4]
  wire  RetimeWrapper_163_io_in; // @[package.scala 93:22:@25092.4]
  wire  RetimeWrapper_163_io_out; // @[package.scala 93:22:@25092.4]
  wire  RetimeWrapper_164_clock; // @[package.scala 93:22:@25100.4]
  wire  RetimeWrapper_164_reset; // @[package.scala 93:22:@25100.4]
  wire  RetimeWrapper_164_io_flow; // @[package.scala 93:22:@25100.4]
  wire  RetimeWrapper_164_io_in; // @[package.scala 93:22:@25100.4]
  wire  RetimeWrapper_164_io_out; // @[package.scala 93:22:@25100.4]
  wire  RetimeWrapper_165_clock; // @[package.scala 93:22:@25108.4]
  wire  RetimeWrapper_165_reset; // @[package.scala 93:22:@25108.4]
  wire  RetimeWrapper_165_io_flow; // @[package.scala 93:22:@25108.4]
  wire  RetimeWrapper_165_io_in; // @[package.scala 93:22:@25108.4]
  wire  RetimeWrapper_165_io_out; // @[package.scala 93:22:@25108.4]
  wire  RetimeWrapper_166_clock; // @[package.scala 93:22:@25116.4]
  wire  RetimeWrapper_166_reset; // @[package.scala 93:22:@25116.4]
  wire  RetimeWrapper_166_io_flow; // @[package.scala 93:22:@25116.4]
  wire  RetimeWrapper_166_io_in; // @[package.scala 93:22:@25116.4]
  wire  RetimeWrapper_166_io_out; // @[package.scala 93:22:@25116.4]
  wire  RetimeWrapper_167_clock; // @[package.scala 93:22:@25124.4]
  wire  RetimeWrapper_167_reset; // @[package.scala 93:22:@25124.4]
  wire  RetimeWrapper_167_io_flow; // @[package.scala 93:22:@25124.4]
  wire  RetimeWrapper_167_io_in; // @[package.scala 93:22:@25124.4]
  wire  RetimeWrapper_167_io_out; // @[package.scala 93:22:@25124.4]
  wire  RetimeWrapper_168_clock; // @[package.scala 93:22:@25180.4]
  wire  RetimeWrapper_168_reset; // @[package.scala 93:22:@25180.4]
  wire  RetimeWrapper_168_io_flow; // @[package.scala 93:22:@25180.4]
  wire  RetimeWrapper_168_io_in; // @[package.scala 93:22:@25180.4]
  wire  RetimeWrapper_168_io_out; // @[package.scala 93:22:@25180.4]
  wire  RetimeWrapper_169_clock; // @[package.scala 93:22:@25188.4]
  wire  RetimeWrapper_169_reset; // @[package.scala 93:22:@25188.4]
  wire  RetimeWrapper_169_io_flow; // @[package.scala 93:22:@25188.4]
  wire  RetimeWrapper_169_io_in; // @[package.scala 93:22:@25188.4]
  wire  RetimeWrapper_169_io_out; // @[package.scala 93:22:@25188.4]
  wire  RetimeWrapper_170_clock; // @[package.scala 93:22:@25196.4]
  wire  RetimeWrapper_170_reset; // @[package.scala 93:22:@25196.4]
  wire  RetimeWrapper_170_io_flow; // @[package.scala 93:22:@25196.4]
  wire  RetimeWrapper_170_io_in; // @[package.scala 93:22:@25196.4]
  wire  RetimeWrapper_170_io_out; // @[package.scala 93:22:@25196.4]
  wire  RetimeWrapper_171_clock; // @[package.scala 93:22:@25204.4]
  wire  RetimeWrapper_171_reset; // @[package.scala 93:22:@25204.4]
  wire  RetimeWrapper_171_io_flow; // @[package.scala 93:22:@25204.4]
  wire  RetimeWrapper_171_io_in; // @[package.scala 93:22:@25204.4]
  wire  RetimeWrapper_171_io_out; // @[package.scala 93:22:@25204.4]
  wire  RetimeWrapper_172_clock; // @[package.scala 93:22:@25212.4]
  wire  RetimeWrapper_172_reset; // @[package.scala 93:22:@25212.4]
  wire  RetimeWrapper_172_io_flow; // @[package.scala 93:22:@25212.4]
  wire  RetimeWrapper_172_io_in; // @[package.scala 93:22:@25212.4]
  wire  RetimeWrapper_172_io_out; // @[package.scala 93:22:@25212.4]
  wire  RetimeWrapper_173_clock; // @[package.scala 93:22:@25220.4]
  wire  RetimeWrapper_173_reset; // @[package.scala 93:22:@25220.4]
  wire  RetimeWrapper_173_io_flow; // @[package.scala 93:22:@25220.4]
  wire  RetimeWrapper_173_io_in; // @[package.scala 93:22:@25220.4]
  wire  RetimeWrapper_173_io_out; // @[package.scala 93:22:@25220.4]
  wire  RetimeWrapper_174_clock; // @[package.scala 93:22:@25228.4]
  wire  RetimeWrapper_174_reset; // @[package.scala 93:22:@25228.4]
  wire  RetimeWrapper_174_io_flow; // @[package.scala 93:22:@25228.4]
  wire  RetimeWrapper_174_io_in; // @[package.scala 93:22:@25228.4]
  wire  RetimeWrapper_174_io_out; // @[package.scala 93:22:@25228.4]
  wire  RetimeWrapper_175_clock; // @[package.scala 93:22:@25236.4]
  wire  RetimeWrapper_175_reset; // @[package.scala 93:22:@25236.4]
  wire  RetimeWrapper_175_io_flow; // @[package.scala 93:22:@25236.4]
  wire  RetimeWrapper_175_io_in; // @[package.scala 93:22:@25236.4]
  wire  RetimeWrapper_175_io_out; // @[package.scala 93:22:@25236.4]
  wire  RetimeWrapper_176_clock; // @[package.scala 93:22:@25244.4]
  wire  RetimeWrapper_176_reset; // @[package.scala 93:22:@25244.4]
  wire  RetimeWrapper_176_io_flow; // @[package.scala 93:22:@25244.4]
  wire  RetimeWrapper_176_io_in; // @[package.scala 93:22:@25244.4]
  wire  RetimeWrapper_176_io_out; // @[package.scala 93:22:@25244.4]
  wire  RetimeWrapper_177_clock; // @[package.scala 93:22:@25252.4]
  wire  RetimeWrapper_177_reset; // @[package.scala 93:22:@25252.4]
  wire  RetimeWrapper_177_io_flow; // @[package.scala 93:22:@25252.4]
  wire  RetimeWrapper_177_io_in; // @[package.scala 93:22:@25252.4]
  wire  RetimeWrapper_177_io_out; // @[package.scala 93:22:@25252.4]
  wire  RetimeWrapper_178_clock; // @[package.scala 93:22:@25260.4]
  wire  RetimeWrapper_178_reset; // @[package.scala 93:22:@25260.4]
  wire  RetimeWrapper_178_io_flow; // @[package.scala 93:22:@25260.4]
  wire  RetimeWrapper_178_io_in; // @[package.scala 93:22:@25260.4]
  wire  RetimeWrapper_178_io_out; // @[package.scala 93:22:@25260.4]
  wire  RetimeWrapper_179_clock; // @[package.scala 93:22:@25268.4]
  wire  RetimeWrapper_179_reset; // @[package.scala 93:22:@25268.4]
  wire  RetimeWrapper_179_io_flow; // @[package.scala 93:22:@25268.4]
  wire  RetimeWrapper_179_io_in; // @[package.scala 93:22:@25268.4]
  wire  RetimeWrapper_179_io_out; // @[package.scala 93:22:@25268.4]
  wire  RetimeWrapper_180_clock; // @[package.scala 93:22:@25324.4]
  wire  RetimeWrapper_180_reset; // @[package.scala 93:22:@25324.4]
  wire  RetimeWrapper_180_io_flow; // @[package.scala 93:22:@25324.4]
  wire  RetimeWrapper_180_io_in; // @[package.scala 93:22:@25324.4]
  wire  RetimeWrapper_180_io_out; // @[package.scala 93:22:@25324.4]
  wire  RetimeWrapper_181_clock; // @[package.scala 93:22:@25332.4]
  wire  RetimeWrapper_181_reset; // @[package.scala 93:22:@25332.4]
  wire  RetimeWrapper_181_io_flow; // @[package.scala 93:22:@25332.4]
  wire  RetimeWrapper_181_io_in; // @[package.scala 93:22:@25332.4]
  wire  RetimeWrapper_181_io_out; // @[package.scala 93:22:@25332.4]
  wire  RetimeWrapper_182_clock; // @[package.scala 93:22:@25340.4]
  wire  RetimeWrapper_182_reset; // @[package.scala 93:22:@25340.4]
  wire  RetimeWrapper_182_io_flow; // @[package.scala 93:22:@25340.4]
  wire  RetimeWrapper_182_io_in; // @[package.scala 93:22:@25340.4]
  wire  RetimeWrapper_182_io_out; // @[package.scala 93:22:@25340.4]
  wire  RetimeWrapper_183_clock; // @[package.scala 93:22:@25348.4]
  wire  RetimeWrapper_183_reset; // @[package.scala 93:22:@25348.4]
  wire  RetimeWrapper_183_io_flow; // @[package.scala 93:22:@25348.4]
  wire  RetimeWrapper_183_io_in; // @[package.scala 93:22:@25348.4]
  wire  RetimeWrapper_183_io_out; // @[package.scala 93:22:@25348.4]
  wire  RetimeWrapper_184_clock; // @[package.scala 93:22:@25356.4]
  wire  RetimeWrapper_184_reset; // @[package.scala 93:22:@25356.4]
  wire  RetimeWrapper_184_io_flow; // @[package.scala 93:22:@25356.4]
  wire  RetimeWrapper_184_io_in; // @[package.scala 93:22:@25356.4]
  wire  RetimeWrapper_184_io_out; // @[package.scala 93:22:@25356.4]
  wire  RetimeWrapper_185_clock; // @[package.scala 93:22:@25364.4]
  wire  RetimeWrapper_185_reset; // @[package.scala 93:22:@25364.4]
  wire  RetimeWrapper_185_io_flow; // @[package.scala 93:22:@25364.4]
  wire  RetimeWrapper_185_io_in; // @[package.scala 93:22:@25364.4]
  wire  RetimeWrapper_185_io_out; // @[package.scala 93:22:@25364.4]
  wire  RetimeWrapper_186_clock; // @[package.scala 93:22:@25372.4]
  wire  RetimeWrapper_186_reset; // @[package.scala 93:22:@25372.4]
  wire  RetimeWrapper_186_io_flow; // @[package.scala 93:22:@25372.4]
  wire  RetimeWrapper_186_io_in; // @[package.scala 93:22:@25372.4]
  wire  RetimeWrapper_186_io_out; // @[package.scala 93:22:@25372.4]
  wire  RetimeWrapper_187_clock; // @[package.scala 93:22:@25380.4]
  wire  RetimeWrapper_187_reset; // @[package.scala 93:22:@25380.4]
  wire  RetimeWrapper_187_io_flow; // @[package.scala 93:22:@25380.4]
  wire  RetimeWrapper_187_io_in; // @[package.scala 93:22:@25380.4]
  wire  RetimeWrapper_187_io_out; // @[package.scala 93:22:@25380.4]
  wire  RetimeWrapper_188_clock; // @[package.scala 93:22:@25388.4]
  wire  RetimeWrapper_188_reset; // @[package.scala 93:22:@25388.4]
  wire  RetimeWrapper_188_io_flow; // @[package.scala 93:22:@25388.4]
  wire  RetimeWrapper_188_io_in; // @[package.scala 93:22:@25388.4]
  wire  RetimeWrapper_188_io_out; // @[package.scala 93:22:@25388.4]
  wire  RetimeWrapper_189_clock; // @[package.scala 93:22:@25396.4]
  wire  RetimeWrapper_189_reset; // @[package.scala 93:22:@25396.4]
  wire  RetimeWrapper_189_io_flow; // @[package.scala 93:22:@25396.4]
  wire  RetimeWrapper_189_io_in; // @[package.scala 93:22:@25396.4]
  wire  RetimeWrapper_189_io_out; // @[package.scala 93:22:@25396.4]
  wire  RetimeWrapper_190_clock; // @[package.scala 93:22:@25404.4]
  wire  RetimeWrapper_190_reset; // @[package.scala 93:22:@25404.4]
  wire  RetimeWrapper_190_io_flow; // @[package.scala 93:22:@25404.4]
  wire  RetimeWrapper_190_io_in; // @[package.scala 93:22:@25404.4]
  wire  RetimeWrapper_190_io_out; // @[package.scala 93:22:@25404.4]
  wire  RetimeWrapper_191_clock; // @[package.scala 93:22:@25412.4]
  wire  RetimeWrapper_191_reset; // @[package.scala 93:22:@25412.4]
  wire  RetimeWrapper_191_io_flow; // @[package.scala 93:22:@25412.4]
  wire  RetimeWrapper_191_io_in; // @[package.scala 93:22:@25412.4]
  wire  RetimeWrapper_191_io_out; // @[package.scala 93:22:@25412.4]
  wire  RetimeWrapper_192_clock; // @[package.scala 93:22:@25468.4]
  wire  RetimeWrapper_192_reset; // @[package.scala 93:22:@25468.4]
  wire  RetimeWrapper_192_io_flow; // @[package.scala 93:22:@25468.4]
  wire  RetimeWrapper_192_io_in; // @[package.scala 93:22:@25468.4]
  wire  RetimeWrapper_192_io_out; // @[package.scala 93:22:@25468.4]
  wire  RetimeWrapper_193_clock; // @[package.scala 93:22:@25476.4]
  wire  RetimeWrapper_193_reset; // @[package.scala 93:22:@25476.4]
  wire  RetimeWrapper_193_io_flow; // @[package.scala 93:22:@25476.4]
  wire  RetimeWrapper_193_io_in; // @[package.scala 93:22:@25476.4]
  wire  RetimeWrapper_193_io_out; // @[package.scala 93:22:@25476.4]
  wire  RetimeWrapper_194_clock; // @[package.scala 93:22:@25484.4]
  wire  RetimeWrapper_194_reset; // @[package.scala 93:22:@25484.4]
  wire  RetimeWrapper_194_io_flow; // @[package.scala 93:22:@25484.4]
  wire  RetimeWrapper_194_io_in; // @[package.scala 93:22:@25484.4]
  wire  RetimeWrapper_194_io_out; // @[package.scala 93:22:@25484.4]
  wire  RetimeWrapper_195_clock; // @[package.scala 93:22:@25492.4]
  wire  RetimeWrapper_195_reset; // @[package.scala 93:22:@25492.4]
  wire  RetimeWrapper_195_io_flow; // @[package.scala 93:22:@25492.4]
  wire  RetimeWrapper_195_io_in; // @[package.scala 93:22:@25492.4]
  wire  RetimeWrapper_195_io_out; // @[package.scala 93:22:@25492.4]
  wire  RetimeWrapper_196_clock; // @[package.scala 93:22:@25500.4]
  wire  RetimeWrapper_196_reset; // @[package.scala 93:22:@25500.4]
  wire  RetimeWrapper_196_io_flow; // @[package.scala 93:22:@25500.4]
  wire  RetimeWrapper_196_io_in; // @[package.scala 93:22:@25500.4]
  wire  RetimeWrapper_196_io_out; // @[package.scala 93:22:@25500.4]
  wire  RetimeWrapper_197_clock; // @[package.scala 93:22:@25508.4]
  wire  RetimeWrapper_197_reset; // @[package.scala 93:22:@25508.4]
  wire  RetimeWrapper_197_io_flow; // @[package.scala 93:22:@25508.4]
  wire  RetimeWrapper_197_io_in; // @[package.scala 93:22:@25508.4]
  wire  RetimeWrapper_197_io_out; // @[package.scala 93:22:@25508.4]
  wire  RetimeWrapper_198_clock; // @[package.scala 93:22:@25516.4]
  wire  RetimeWrapper_198_reset; // @[package.scala 93:22:@25516.4]
  wire  RetimeWrapper_198_io_flow; // @[package.scala 93:22:@25516.4]
  wire  RetimeWrapper_198_io_in; // @[package.scala 93:22:@25516.4]
  wire  RetimeWrapper_198_io_out; // @[package.scala 93:22:@25516.4]
  wire  RetimeWrapper_199_clock; // @[package.scala 93:22:@25524.4]
  wire  RetimeWrapper_199_reset; // @[package.scala 93:22:@25524.4]
  wire  RetimeWrapper_199_io_flow; // @[package.scala 93:22:@25524.4]
  wire  RetimeWrapper_199_io_in; // @[package.scala 93:22:@25524.4]
  wire  RetimeWrapper_199_io_out; // @[package.scala 93:22:@25524.4]
  wire  RetimeWrapper_200_clock; // @[package.scala 93:22:@25532.4]
  wire  RetimeWrapper_200_reset; // @[package.scala 93:22:@25532.4]
  wire  RetimeWrapper_200_io_flow; // @[package.scala 93:22:@25532.4]
  wire  RetimeWrapper_200_io_in; // @[package.scala 93:22:@25532.4]
  wire  RetimeWrapper_200_io_out; // @[package.scala 93:22:@25532.4]
  wire  RetimeWrapper_201_clock; // @[package.scala 93:22:@25540.4]
  wire  RetimeWrapper_201_reset; // @[package.scala 93:22:@25540.4]
  wire  RetimeWrapper_201_io_flow; // @[package.scala 93:22:@25540.4]
  wire  RetimeWrapper_201_io_in; // @[package.scala 93:22:@25540.4]
  wire  RetimeWrapper_201_io_out; // @[package.scala 93:22:@25540.4]
  wire  RetimeWrapper_202_clock; // @[package.scala 93:22:@25548.4]
  wire  RetimeWrapper_202_reset; // @[package.scala 93:22:@25548.4]
  wire  RetimeWrapper_202_io_flow; // @[package.scala 93:22:@25548.4]
  wire  RetimeWrapper_202_io_in; // @[package.scala 93:22:@25548.4]
  wire  RetimeWrapper_202_io_out; // @[package.scala 93:22:@25548.4]
  wire  RetimeWrapper_203_clock; // @[package.scala 93:22:@25556.4]
  wire  RetimeWrapper_203_reset; // @[package.scala 93:22:@25556.4]
  wire  RetimeWrapper_203_io_flow; // @[package.scala 93:22:@25556.4]
  wire  RetimeWrapper_203_io_in; // @[package.scala 93:22:@25556.4]
  wire  RetimeWrapper_203_io_out; // @[package.scala 93:22:@25556.4]
  wire  RetimeWrapper_204_clock; // @[package.scala 93:22:@25612.4]
  wire  RetimeWrapper_204_reset; // @[package.scala 93:22:@25612.4]
  wire  RetimeWrapper_204_io_flow; // @[package.scala 93:22:@25612.4]
  wire  RetimeWrapper_204_io_in; // @[package.scala 93:22:@25612.4]
  wire  RetimeWrapper_204_io_out; // @[package.scala 93:22:@25612.4]
  wire  RetimeWrapper_205_clock; // @[package.scala 93:22:@25620.4]
  wire  RetimeWrapper_205_reset; // @[package.scala 93:22:@25620.4]
  wire  RetimeWrapper_205_io_flow; // @[package.scala 93:22:@25620.4]
  wire  RetimeWrapper_205_io_in; // @[package.scala 93:22:@25620.4]
  wire  RetimeWrapper_205_io_out; // @[package.scala 93:22:@25620.4]
  wire  RetimeWrapper_206_clock; // @[package.scala 93:22:@25628.4]
  wire  RetimeWrapper_206_reset; // @[package.scala 93:22:@25628.4]
  wire  RetimeWrapper_206_io_flow; // @[package.scala 93:22:@25628.4]
  wire  RetimeWrapper_206_io_in; // @[package.scala 93:22:@25628.4]
  wire  RetimeWrapper_206_io_out; // @[package.scala 93:22:@25628.4]
  wire  RetimeWrapper_207_clock; // @[package.scala 93:22:@25636.4]
  wire  RetimeWrapper_207_reset; // @[package.scala 93:22:@25636.4]
  wire  RetimeWrapper_207_io_flow; // @[package.scala 93:22:@25636.4]
  wire  RetimeWrapper_207_io_in; // @[package.scala 93:22:@25636.4]
  wire  RetimeWrapper_207_io_out; // @[package.scala 93:22:@25636.4]
  wire  RetimeWrapper_208_clock; // @[package.scala 93:22:@25644.4]
  wire  RetimeWrapper_208_reset; // @[package.scala 93:22:@25644.4]
  wire  RetimeWrapper_208_io_flow; // @[package.scala 93:22:@25644.4]
  wire  RetimeWrapper_208_io_in; // @[package.scala 93:22:@25644.4]
  wire  RetimeWrapper_208_io_out; // @[package.scala 93:22:@25644.4]
  wire  RetimeWrapper_209_clock; // @[package.scala 93:22:@25652.4]
  wire  RetimeWrapper_209_reset; // @[package.scala 93:22:@25652.4]
  wire  RetimeWrapper_209_io_flow; // @[package.scala 93:22:@25652.4]
  wire  RetimeWrapper_209_io_in; // @[package.scala 93:22:@25652.4]
  wire  RetimeWrapper_209_io_out; // @[package.scala 93:22:@25652.4]
  wire  RetimeWrapper_210_clock; // @[package.scala 93:22:@25660.4]
  wire  RetimeWrapper_210_reset; // @[package.scala 93:22:@25660.4]
  wire  RetimeWrapper_210_io_flow; // @[package.scala 93:22:@25660.4]
  wire  RetimeWrapper_210_io_in; // @[package.scala 93:22:@25660.4]
  wire  RetimeWrapper_210_io_out; // @[package.scala 93:22:@25660.4]
  wire  RetimeWrapper_211_clock; // @[package.scala 93:22:@25668.4]
  wire  RetimeWrapper_211_reset; // @[package.scala 93:22:@25668.4]
  wire  RetimeWrapper_211_io_flow; // @[package.scala 93:22:@25668.4]
  wire  RetimeWrapper_211_io_in; // @[package.scala 93:22:@25668.4]
  wire  RetimeWrapper_211_io_out; // @[package.scala 93:22:@25668.4]
  wire  RetimeWrapper_212_clock; // @[package.scala 93:22:@25676.4]
  wire  RetimeWrapper_212_reset; // @[package.scala 93:22:@25676.4]
  wire  RetimeWrapper_212_io_flow; // @[package.scala 93:22:@25676.4]
  wire  RetimeWrapper_212_io_in; // @[package.scala 93:22:@25676.4]
  wire  RetimeWrapper_212_io_out; // @[package.scala 93:22:@25676.4]
  wire  RetimeWrapper_213_clock; // @[package.scala 93:22:@25684.4]
  wire  RetimeWrapper_213_reset; // @[package.scala 93:22:@25684.4]
  wire  RetimeWrapper_213_io_flow; // @[package.scala 93:22:@25684.4]
  wire  RetimeWrapper_213_io_in; // @[package.scala 93:22:@25684.4]
  wire  RetimeWrapper_213_io_out; // @[package.scala 93:22:@25684.4]
  wire  RetimeWrapper_214_clock; // @[package.scala 93:22:@25692.4]
  wire  RetimeWrapper_214_reset; // @[package.scala 93:22:@25692.4]
  wire  RetimeWrapper_214_io_flow; // @[package.scala 93:22:@25692.4]
  wire  RetimeWrapper_214_io_in; // @[package.scala 93:22:@25692.4]
  wire  RetimeWrapper_214_io_out; // @[package.scala 93:22:@25692.4]
  wire  RetimeWrapper_215_clock; // @[package.scala 93:22:@25700.4]
  wire  RetimeWrapper_215_reset; // @[package.scala 93:22:@25700.4]
  wire  RetimeWrapper_215_io_flow; // @[package.scala 93:22:@25700.4]
  wire  RetimeWrapper_215_io_in; // @[package.scala 93:22:@25700.4]
  wire  RetimeWrapper_215_io_out; // @[package.scala 93:22:@25700.4]
  wire  _T_700; // @[MemPrimitives.scala 82:210:@20535.4]
  wire  _T_702; // @[MemPrimitives.scala 82:210:@20536.4]
  wire  _T_703; // @[MemPrimitives.scala 82:228:@20537.4]
  wire  _T_704; // @[MemPrimitives.scala 83:102:@20538.4]
  wire  _T_706; // @[MemPrimitives.scala 82:210:@20539.4]
  wire  _T_708; // @[MemPrimitives.scala 82:210:@20540.4]
  wire  _T_709; // @[MemPrimitives.scala 82:228:@20541.4]
  wire  _T_710; // @[MemPrimitives.scala 83:102:@20542.4]
  wire [17:0] _T_712; // @[Cat.scala 30:58:@20544.4]
  wire [17:0] _T_714; // @[Cat.scala 30:58:@20546.4]
  wire [17:0] _T_715; // @[Mux.scala 31:69:@20547.4]
  wire  _T_720; // @[MemPrimitives.scala 82:210:@20554.4]
  wire  _T_722; // @[MemPrimitives.scala 82:210:@20555.4]
  wire  _T_723; // @[MemPrimitives.scala 82:228:@20556.4]
  wire  _T_724; // @[MemPrimitives.scala 83:102:@20557.4]
  wire  _T_726; // @[MemPrimitives.scala 82:210:@20558.4]
  wire  _T_728; // @[MemPrimitives.scala 82:210:@20559.4]
  wire  _T_729; // @[MemPrimitives.scala 82:228:@20560.4]
  wire  _T_730; // @[MemPrimitives.scala 83:102:@20561.4]
  wire [17:0] _T_732; // @[Cat.scala 30:58:@20563.4]
  wire [17:0] _T_734; // @[Cat.scala 30:58:@20565.4]
  wire [17:0] _T_735; // @[Mux.scala 31:69:@20566.4]
  wire  _T_742; // @[MemPrimitives.scala 82:210:@20574.4]
  wire  _T_743; // @[MemPrimitives.scala 82:228:@20575.4]
  wire  _T_744; // @[MemPrimitives.scala 83:102:@20576.4]
  wire  _T_748; // @[MemPrimitives.scala 82:210:@20578.4]
  wire  _T_749; // @[MemPrimitives.scala 82:228:@20579.4]
  wire  _T_750; // @[MemPrimitives.scala 83:102:@20580.4]
  wire [17:0] _T_752; // @[Cat.scala 30:58:@20582.4]
  wire [17:0] _T_754; // @[Cat.scala 30:58:@20584.4]
  wire [17:0] _T_755; // @[Mux.scala 31:69:@20585.4]
  wire  _T_762; // @[MemPrimitives.scala 82:210:@20593.4]
  wire  _T_763; // @[MemPrimitives.scala 82:228:@20594.4]
  wire  _T_764; // @[MemPrimitives.scala 83:102:@20595.4]
  wire  _T_768; // @[MemPrimitives.scala 82:210:@20597.4]
  wire  _T_769; // @[MemPrimitives.scala 82:228:@20598.4]
  wire  _T_770; // @[MemPrimitives.scala 83:102:@20599.4]
  wire [17:0] _T_772; // @[Cat.scala 30:58:@20601.4]
  wire [17:0] _T_774; // @[Cat.scala 30:58:@20603.4]
  wire [17:0] _T_775; // @[Mux.scala 31:69:@20604.4]
  wire  _T_782; // @[MemPrimitives.scala 82:210:@20612.4]
  wire  _T_783; // @[MemPrimitives.scala 82:228:@20613.4]
  wire  _T_784; // @[MemPrimitives.scala 83:102:@20614.4]
  wire  _T_788; // @[MemPrimitives.scala 82:210:@20616.4]
  wire  _T_789; // @[MemPrimitives.scala 82:228:@20617.4]
  wire  _T_790; // @[MemPrimitives.scala 83:102:@20618.4]
  wire [17:0] _T_792; // @[Cat.scala 30:58:@20620.4]
  wire [17:0] _T_794; // @[Cat.scala 30:58:@20622.4]
  wire [17:0] _T_795; // @[Mux.scala 31:69:@20623.4]
  wire  _T_802; // @[MemPrimitives.scala 82:210:@20631.4]
  wire  _T_803; // @[MemPrimitives.scala 82:228:@20632.4]
  wire  _T_804; // @[MemPrimitives.scala 83:102:@20633.4]
  wire  _T_808; // @[MemPrimitives.scala 82:210:@20635.4]
  wire  _T_809; // @[MemPrimitives.scala 82:228:@20636.4]
  wire  _T_810; // @[MemPrimitives.scala 83:102:@20637.4]
  wire [17:0] _T_812; // @[Cat.scala 30:58:@20639.4]
  wire [17:0] _T_814; // @[Cat.scala 30:58:@20641.4]
  wire [17:0] _T_815; // @[Mux.scala 31:69:@20642.4]
  wire  _T_820; // @[MemPrimitives.scala 82:210:@20649.4]
  wire  _T_823; // @[MemPrimitives.scala 82:228:@20651.4]
  wire  _T_824; // @[MemPrimitives.scala 83:102:@20652.4]
  wire  _T_826; // @[MemPrimitives.scala 82:210:@20653.4]
  wire  _T_829; // @[MemPrimitives.scala 82:228:@20655.4]
  wire  _T_830; // @[MemPrimitives.scala 83:102:@20656.4]
  wire [17:0] _T_832; // @[Cat.scala 30:58:@20658.4]
  wire [17:0] _T_834; // @[Cat.scala 30:58:@20660.4]
  wire [17:0] _T_835; // @[Mux.scala 31:69:@20661.4]
  wire  _T_840; // @[MemPrimitives.scala 82:210:@20668.4]
  wire  _T_843; // @[MemPrimitives.scala 82:228:@20670.4]
  wire  _T_844; // @[MemPrimitives.scala 83:102:@20671.4]
  wire  _T_846; // @[MemPrimitives.scala 82:210:@20672.4]
  wire  _T_849; // @[MemPrimitives.scala 82:228:@20674.4]
  wire  _T_850; // @[MemPrimitives.scala 83:102:@20675.4]
  wire [17:0] _T_852; // @[Cat.scala 30:58:@20677.4]
  wire [17:0] _T_854; // @[Cat.scala 30:58:@20679.4]
  wire [17:0] _T_855; // @[Mux.scala 31:69:@20680.4]
  wire  _T_863; // @[MemPrimitives.scala 82:228:@20689.4]
  wire  _T_864; // @[MemPrimitives.scala 83:102:@20690.4]
  wire  _T_869; // @[MemPrimitives.scala 82:228:@20693.4]
  wire  _T_870; // @[MemPrimitives.scala 83:102:@20694.4]
  wire [17:0] _T_872; // @[Cat.scala 30:58:@20696.4]
  wire [17:0] _T_874; // @[Cat.scala 30:58:@20698.4]
  wire [17:0] _T_875; // @[Mux.scala 31:69:@20699.4]
  wire  _T_883; // @[MemPrimitives.scala 82:228:@20708.4]
  wire  _T_884; // @[MemPrimitives.scala 83:102:@20709.4]
  wire  _T_889; // @[MemPrimitives.scala 82:228:@20712.4]
  wire  _T_890; // @[MemPrimitives.scala 83:102:@20713.4]
  wire [17:0] _T_892; // @[Cat.scala 30:58:@20715.4]
  wire [17:0] _T_894; // @[Cat.scala 30:58:@20717.4]
  wire [17:0] _T_895; // @[Mux.scala 31:69:@20718.4]
  wire  _T_903; // @[MemPrimitives.scala 82:228:@20727.4]
  wire  _T_904; // @[MemPrimitives.scala 83:102:@20728.4]
  wire  _T_909; // @[MemPrimitives.scala 82:228:@20731.4]
  wire  _T_910; // @[MemPrimitives.scala 83:102:@20732.4]
  wire [17:0] _T_912; // @[Cat.scala 30:58:@20734.4]
  wire [17:0] _T_914; // @[Cat.scala 30:58:@20736.4]
  wire [17:0] _T_915; // @[Mux.scala 31:69:@20737.4]
  wire  _T_923; // @[MemPrimitives.scala 82:228:@20746.4]
  wire  _T_924; // @[MemPrimitives.scala 83:102:@20747.4]
  wire  _T_929; // @[MemPrimitives.scala 82:228:@20750.4]
  wire  _T_930; // @[MemPrimitives.scala 83:102:@20751.4]
  wire [17:0] _T_932; // @[Cat.scala 30:58:@20753.4]
  wire [17:0] _T_934; // @[Cat.scala 30:58:@20755.4]
  wire [17:0] _T_935; // @[Mux.scala 31:69:@20756.4]
  wire  _T_940; // @[MemPrimitives.scala 82:210:@20763.4]
  wire  _T_943; // @[MemPrimitives.scala 82:228:@20765.4]
  wire  _T_944; // @[MemPrimitives.scala 83:102:@20766.4]
  wire  _T_946; // @[MemPrimitives.scala 82:210:@20767.4]
  wire  _T_949; // @[MemPrimitives.scala 82:228:@20769.4]
  wire  _T_950; // @[MemPrimitives.scala 83:102:@20770.4]
  wire [17:0] _T_952; // @[Cat.scala 30:58:@20772.4]
  wire [17:0] _T_954; // @[Cat.scala 30:58:@20774.4]
  wire [17:0] _T_955; // @[Mux.scala 31:69:@20775.4]
  wire  _T_960; // @[MemPrimitives.scala 82:210:@20782.4]
  wire  _T_963; // @[MemPrimitives.scala 82:228:@20784.4]
  wire  _T_964; // @[MemPrimitives.scala 83:102:@20785.4]
  wire  _T_966; // @[MemPrimitives.scala 82:210:@20786.4]
  wire  _T_969; // @[MemPrimitives.scala 82:228:@20788.4]
  wire  _T_970; // @[MemPrimitives.scala 83:102:@20789.4]
  wire [17:0] _T_972; // @[Cat.scala 30:58:@20791.4]
  wire [17:0] _T_974; // @[Cat.scala 30:58:@20793.4]
  wire [17:0] _T_975; // @[Mux.scala 31:69:@20794.4]
  wire  _T_983; // @[MemPrimitives.scala 82:228:@20803.4]
  wire  _T_984; // @[MemPrimitives.scala 83:102:@20804.4]
  wire  _T_989; // @[MemPrimitives.scala 82:228:@20807.4]
  wire  _T_990; // @[MemPrimitives.scala 83:102:@20808.4]
  wire [17:0] _T_992; // @[Cat.scala 30:58:@20810.4]
  wire [17:0] _T_994; // @[Cat.scala 30:58:@20812.4]
  wire [17:0] _T_995; // @[Mux.scala 31:69:@20813.4]
  wire  _T_1003; // @[MemPrimitives.scala 82:228:@20822.4]
  wire  _T_1004; // @[MemPrimitives.scala 83:102:@20823.4]
  wire  _T_1009; // @[MemPrimitives.scala 82:228:@20826.4]
  wire  _T_1010; // @[MemPrimitives.scala 83:102:@20827.4]
  wire [17:0] _T_1012; // @[Cat.scala 30:58:@20829.4]
  wire [17:0] _T_1014; // @[Cat.scala 30:58:@20831.4]
  wire [17:0] _T_1015; // @[Mux.scala 31:69:@20832.4]
  wire  _T_1023; // @[MemPrimitives.scala 82:228:@20841.4]
  wire  _T_1024; // @[MemPrimitives.scala 83:102:@20842.4]
  wire  _T_1029; // @[MemPrimitives.scala 82:228:@20845.4]
  wire  _T_1030; // @[MemPrimitives.scala 83:102:@20846.4]
  wire [17:0] _T_1032; // @[Cat.scala 30:58:@20848.4]
  wire [17:0] _T_1034; // @[Cat.scala 30:58:@20850.4]
  wire [17:0] _T_1035; // @[Mux.scala 31:69:@20851.4]
  wire  _T_1043; // @[MemPrimitives.scala 82:228:@20860.4]
  wire  _T_1044; // @[MemPrimitives.scala 83:102:@20861.4]
  wire  _T_1049; // @[MemPrimitives.scala 82:228:@20864.4]
  wire  _T_1050; // @[MemPrimitives.scala 83:102:@20865.4]
  wire [17:0] _T_1052; // @[Cat.scala 30:58:@20867.4]
  wire [17:0] _T_1054; // @[Cat.scala 30:58:@20869.4]
  wire [17:0] _T_1055; // @[Mux.scala 31:69:@20870.4]
  wire  _T_1060; // @[MemPrimitives.scala 82:210:@20877.4]
  wire  _T_1063; // @[MemPrimitives.scala 82:228:@20879.4]
  wire  _T_1064; // @[MemPrimitives.scala 83:102:@20880.4]
  wire  _T_1066; // @[MemPrimitives.scala 82:210:@20881.4]
  wire  _T_1069; // @[MemPrimitives.scala 82:228:@20883.4]
  wire  _T_1070; // @[MemPrimitives.scala 83:102:@20884.4]
  wire [17:0] _T_1072; // @[Cat.scala 30:58:@20886.4]
  wire [17:0] _T_1074; // @[Cat.scala 30:58:@20888.4]
  wire [17:0] _T_1075; // @[Mux.scala 31:69:@20889.4]
  wire  _T_1080; // @[MemPrimitives.scala 82:210:@20896.4]
  wire  _T_1083; // @[MemPrimitives.scala 82:228:@20898.4]
  wire  _T_1084; // @[MemPrimitives.scala 83:102:@20899.4]
  wire  _T_1086; // @[MemPrimitives.scala 82:210:@20900.4]
  wire  _T_1089; // @[MemPrimitives.scala 82:228:@20902.4]
  wire  _T_1090; // @[MemPrimitives.scala 83:102:@20903.4]
  wire [17:0] _T_1092; // @[Cat.scala 30:58:@20905.4]
  wire [17:0] _T_1094; // @[Cat.scala 30:58:@20907.4]
  wire [17:0] _T_1095; // @[Mux.scala 31:69:@20908.4]
  wire  _T_1103; // @[MemPrimitives.scala 82:228:@20917.4]
  wire  _T_1104; // @[MemPrimitives.scala 83:102:@20918.4]
  wire  _T_1109; // @[MemPrimitives.scala 82:228:@20921.4]
  wire  _T_1110; // @[MemPrimitives.scala 83:102:@20922.4]
  wire [17:0] _T_1112; // @[Cat.scala 30:58:@20924.4]
  wire [17:0] _T_1114; // @[Cat.scala 30:58:@20926.4]
  wire [17:0] _T_1115; // @[Mux.scala 31:69:@20927.4]
  wire  _T_1123; // @[MemPrimitives.scala 82:228:@20936.4]
  wire  _T_1124; // @[MemPrimitives.scala 83:102:@20937.4]
  wire  _T_1129; // @[MemPrimitives.scala 82:228:@20940.4]
  wire  _T_1130; // @[MemPrimitives.scala 83:102:@20941.4]
  wire [17:0] _T_1132; // @[Cat.scala 30:58:@20943.4]
  wire [17:0] _T_1134; // @[Cat.scala 30:58:@20945.4]
  wire [17:0] _T_1135; // @[Mux.scala 31:69:@20946.4]
  wire  _T_1143; // @[MemPrimitives.scala 82:228:@20955.4]
  wire  _T_1144; // @[MemPrimitives.scala 83:102:@20956.4]
  wire  _T_1149; // @[MemPrimitives.scala 82:228:@20959.4]
  wire  _T_1150; // @[MemPrimitives.scala 83:102:@20960.4]
  wire [17:0] _T_1152; // @[Cat.scala 30:58:@20962.4]
  wire [17:0] _T_1154; // @[Cat.scala 30:58:@20964.4]
  wire [17:0] _T_1155; // @[Mux.scala 31:69:@20965.4]
  wire  _T_1163; // @[MemPrimitives.scala 82:228:@20974.4]
  wire  _T_1164; // @[MemPrimitives.scala 83:102:@20975.4]
  wire  _T_1169; // @[MemPrimitives.scala 82:228:@20978.4]
  wire  _T_1170; // @[MemPrimitives.scala 83:102:@20979.4]
  wire [17:0] _T_1172; // @[Cat.scala 30:58:@20981.4]
  wire [17:0] _T_1174; // @[Cat.scala 30:58:@20983.4]
  wire [17:0] _T_1175; // @[Mux.scala 31:69:@20984.4]
  wire  _T_1180; // @[MemPrimitives.scala 110:210:@20991.4]
  wire  _T_1182; // @[MemPrimitives.scala 110:210:@20992.4]
  wire  _T_1183; // @[MemPrimitives.scala 110:228:@20993.4]
  wire  _T_1186; // @[MemPrimitives.scala 110:210:@20995.4]
  wire  _T_1188; // @[MemPrimitives.scala 110:210:@20996.4]
  wire  _T_1189; // @[MemPrimitives.scala 110:228:@20997.4]
  wire  _T_1192; // @[MemPrimitives.scala 110:210:@20999.4]
  wire  _T_1194; // @[MemPrimitives.scala 110:210:@21000.4]
  wire  _T_1195; // @[MemPrimitives.scala 110:228:@21001.4]
  wire  _T_1198; // @[MemPrimitives.scala 110:210:@21003.4]
  wire  _T_1200; // @[MemPrimitives.scala 110:210:@21004.4]
  wire  _T_1201; // @[MemPrimitives.scala 110:228:@21005.4]
  wire  _T_1204; // @[MemPrimitives.scala 110:210:@21007.4]
  wire  _T_1206; // @[MemPrimitives.scala 110:210:@21008.4]
  wire  _T_1207; // @[MemPrimitives.scala 110:228:@21009.4]
  wire  _T_1210; // @[MemPrimitives.scala 110:210:@21011.4]
  wire  _T_1212; // @[MemPrimitives.scala 110:210:@21012.4]
  wire  _T_1213; // @[MemPrimitives.scala 110:228:@21013.4]
  wire  _T_1216; // @[MemPrimitives.scala 110:210:@21015.4]
  wire  _T_1218; // @[MemPrimitives.scala 110:210:@21016.4]
  wire  _T_1219; // @[MemPrimitives.scala 110:228:@21017.4]
  wire  _T_1222; // @[MemPrimitives.scala 110:210:@21019.4]
  wire  _T_1224; // @[MemPrimitives.scala 110:210:@21020.4]
  wire  _T_1225; // @[MemPrimitives.scala 110:228:@21021.4]
  wire  _T_1228; // @[MemPrimitives.scala 110:210:@21023.4]
  wire  _T_1230; // @[MemPrimitives.scala 110:210:@21024.4]
  wire  _T_1231; // @[MemPrimitives.scala 110:228:@21025.4]
  wire  _T_1233; // @[MemPrimitives.scala 123:41:@21039.4]
  wire  _T_1234; // @[MemPrimitives.scala 123:41:@21040.4]
  wire  _T_1235; // @[MemPrimitives.scala 123:41:@21041.4]
  wire  _T_1236; // @[MemPrimitives.scala 123:41:@21042.4]
  wire  _T_1237; // @[MemPrimitives.scala 123:41:@21043.4]
  wire  _T_1238; // @[MemPrimitives.scala 123:41:@21044.4]
  wire  _T_1239; // @[MemPrimitives.scala 123:41:@21045.4]
  wire  _T_1240; // @[MemPrimitives.scala 123:41:@21046.4]
  wire  _T_1241; // @[MemPrimitives.scala 123:41:@21047.4]
  wire [10:0] _T_1243; // @[Cat.scala 30:58:@21049.4]
  wire [10:0] _T_1245; // @[Cat.scala 30:58:@21051.4]
  wire [10:0] _T_1247; // @[Cat.scala 30:58:@21053.4]
  wire [10:0] _T_1249; // @[Cat.scala 30:58:@21055.4]
  wire [10:0] _T_1251; // @[Cat.scala 30:58:@21057.4]
  wire [10:0] _T_1253; // @[Cat.scala 30:58:@21059.4]
  wire [10:0] _T_1255; // @[Cat.scala 30:58:@21061.4]
  wire [10:0] _T_1257; // @[Cat.scala 30:58:@21063.4]
  wire [10:0] _T_1259; // @[Cat.scala 30:58:@21065.4]
  wire [10:0] _T_1260; // @[Mux.scala 31:69:@21066.4]
  wire [10:0] _T_1261; // @[Mux.scala 31:69:@21067.4]
  wire [10:0] _T_1262; // @[Mux.scala 31:69:@21068.4]
  wire [10:0] _T_1263; // @[Mux.scala 31:69:@21069.4]
  wire [10:0] _T_1264; // @[Mux.scala 31:69:@21070.4]
  wire [10:0] _T_1265; // @[Mux.scala 31:69:@21071.4]
  wire [10:0] _T_1266; // @[Mux.scala 31:69:@21072.4]
  wire [10:0] _T_1267; // @[Mux.scala 31:69:@21073.4]
  wire  _T_1272; // @[MemPrimitives.scala 110:210:@21080.4]
  wire  _T_1274; // @[MemPrimitives.scala 110:210:@21081.4]
  wire  _T_1275; // @[MemPrimitives.scala 110:228:@21082.4]
  wire  _T_1278; // @[MemPrimitives.scala 110:210:@21084.4]
  wire  _T_1280; // @[MemPrimitives.scala 110:210:@21085.4]
  wire  _T_1281; // @[MemPrimitives.scala 110:228:@21086.4]
  wire  _T_1284; // @[MemPrimitives.scala 110:210:@21088.4]
  wire  _T_1286; // @[MemPrimitives.scala 110:210:@21089.4]
  wire  _T_1287; // @[MemPrimitives.scala 110:228:@21090.4]
  wire  _T_1290; // @[MemPrimitives.scala 110:210:@21092.4]
  wire  _T_1292; // @[MemPrimitives.scala 110:210:@21093.4]
  wire  _T_1293; // @[MemPrimitives.scala 110:228:@21094.4]
  wire  _T_1296; // @[MemPrimitives.scala 110:210:@21096.4]
  wire  _T_1298; // @[MemPrimitives.scala 110:210:@21097.4]
  wire  _T_1299; // @[MemPrimitives.scala 110:228:@21098.4]
  wire  _T_1302; // @[MemPrimitives.scala 110:210:@21100.4]
  wire  _T_1304; // @[MemPrimitives.scala 110:210:@21101.4]
  wire  _T_1305; // @[MemPrimitives.scala 110:228:@21102.4]
  wire  _T_1308; // @[MemPrimitives.scala 110:210:@21104.4]
  wire  _T_1310; // @[MemPrimitives.scala 110:210:@21105.4]
  wire  _T_1311; // @[MemPrimitives.scala 110:228:@21106.4]
  wire  _T_1314; // @[MemPrimitives.scala 110:210:@21108.4]
  wire  _T_1316; // @[MemPrimitives.scala 110:210:@21109.4]
  wire  _T_1317; // @[MemPrimitives.scala 110:228:@21110.4]
  wire  _T_1320; // @[MemPrimitives.scala 110:210:@21112.4]
  wire  _T_1322; // @[MemPrimitives.scala 110:210:@21113.4]
  wire  _T_1323; // @[MemPrimitives.scala 110:228:@21114.4]
  wire  _T_1325; // @[MemPrimitives.scala 123:41:@21128.4]
  wire  _T_1326; // @[MemPrimitives.scala 123:41:@21129.4]
  wire  _T_1327; // @[MemPrimitives.scala 123:41:@21130.4]
  wire  _T_1328; // @[MemPrimitives.scala 123:41:@21131.4]
  wire  _T_1329; // @[MemPrimitives.scala 123:41:@21132.4]
  wire  _T_1330; // @[MemPrimitives.scala 123:41:@21133.4]
  wire  _T_1331; // @[MemPrimitives.scala 123:41:@21134.4]
  wire  _T_1332; // @[MemPrimitives.scala 123:41:@21135.4]
  wire  _T_1333; // @[MemPrimitives.scala 123:41:@21136.4]
  wire [10:0] _T_1335; // @[Cat.scala 30:58:@21138.4]
  wire [10:0] _T_1337; // @[Cat.scala 30:58:@21140.4]
  wire [10:0] _T_1339; // @[Cat.scala 30:58:@21142.4]
  wire [10:0] _T_1341; // @[Cat.scala 30:58:@21144.4]
  wire [10:0] _T_1343; // @[Cat.scala 30:58:@21146.4]
  wire [10:0] _T_1345; // @[Cat.scala 30:58:@21148.4]
  wire [10:0] _T_1347; // @[Cat.scala 30:58:@21150.4]
  wire [10:0] _T_1349; // @[Cat.scala 30:58:@21152.4]
  wire [10:0] _T_1351; // @[Cat.scala 30:58:@21154.4]
  wire [10:0] _T_1352; // @[Mux.scala 31:69:@21155.4]
  wire [10:0] _T_1353; // @[Mux.scala 31:69:@21156.4]
  wire [10:0] _T_1354; // @[Mux.scala 31:69:@21157.4]
  wire [10:0] _T_1355; // @[Mux.scala 31:69:@21158.4]
  wire [10:0] _T_1356; // @[Mux.scala 31:69:@21159.4]
  wire [10:0] _T_1357; // @[Mux.scala 31:69:@21160.4]
  wire [10:0] _T_1358; // @[Mux.scala 31:69:@21161.4]
  wire [10:0] _T_1359; // @[Mux.scala 31:69:@21162.4]
  wire  _T_1366; // @[MemPrimitives.scala 110:210:@21170.4]
  wire  _T_1367; // @[MemPrimitives.scala 110:228:@21171.4]
  wire  _T_1372; // @[MemPrimitives.scala 110:210:@21174.4]
  wire  _T_1373; // @[MemPrimitives.scala 110:228:@21175.4]
  wire  _T_1378; // @[MemPrimitives.scala 110:210:@21178.4]
  wire  _T_1379; // @[MemPrimitives.scala 110:228:@21179.4]
  wire  _T_1384; // @[MemPrimitives.scala 110:210:@21182.4]
  wire  _T_1385; // @[MemPrimitives.scala 110:228:@21183.4]
  wire  _T_1390; // @[MemPrimitives.scala 110:210:@21186.4]
  wire  _T_1391; // @[MemPrimitives.scala 110:228:@21187.4]
  wire  _T_1396; // @[MemPrimitives.scala 110:210:@21190.4]
  wire  _T_1397; // @[MemPrimitives.scala 110:228:@21191.4]
  wire  _T_1402; // @[MemPrimitives.scala 110:210:@21194.4]
  wire  _T_1403; // @[MemPrimitives.scala 110:228:@21195.4]
  wire  _T_1408; // @[MemPrimitives.scala 110:210:@21198.4]
  wire  _T_1409; // @[MemPrimitives.scala 110:228:@21199.4]
  wire  _T_1414; // @[MemPrimitives.scala 110:210:@21202.4]
  wire  _T_1415; // @[MemPrimitives.scala 110:228:@21203.4]
  wire  _T_1417; // @[MemPrimitives.scala 123:41:@21217.4]
  wire  _T_1418; // @[MemPrimitives.scala 123:41:@21218.4]
  wire  _T_1419; // @[MemPrimitives.scala 123:41:@21219.4]
  wire  _T_1420; // @[MemPrimitives.scala 123:41:@21220.4]
  wire  _T_1421; // @[MemPrimitives.scala 123:41:@21221.4]
  wire  _T_1422; // @[MemPrimitives.scala 123:41:@21222.4]
  wire  _T_1423; // @[MemPrimitives.scala 123:41:@21223.4]
  wire  _T_1424; // @[MemPrimitives.scala 123:41:@21224.4]
  wire  _T_1425; // @[MemPrimitives.scala 123:41:@21225.4]
  wire [10:0] _T_1427; // @[Cat.scala 30:58:@21227.4]
  wire [10:0] _T_1429; // @[Cat.scala 30:58:@21229.4]
  wire [10:0] _T_1431; // @[Cat.scala 30:58:@21231.4]
  wire [10:0] _T_1433; // @[Cat.scala 30:58:@21233.4]
  wire [10:0] _T_1435; // @[Cat.scala 30:58:@21235.4]
  wire [10:0] _T_1437; // @[Cat.scala 30:58:@21237.4]
  wire [10:0] _T_1439; // @[Cat.scala 30:58:@21239.4]
  wire [10:0] _T_1441; // @[Cat.scala 30:58:@21241.4]
  wire [10:0] _T_1443; // @[Cat.scala 30:58:@21243.4]
  wire [10:0] _T_1444; // @[Mux.scala 31:69:@21244.4]
  wire [10:0] _T_1445; // @[Mux.scala 31:69:@21245.4]
  wire [10:0] _T_1446; // @[Mux.scala 31:69:@21246.4]
  wire [10:0] _T_1447; // @[Mux.scala 31:69:@21247.4]
  wire [10:0] _T_1448; // @[Mux.scala 31:69:@21248.4]
  wire [10:0] _T_1449; // @[Mux.scala 31:69:@21249.4]
  wire [10:0] _T_1450; // @[Mux.scala 31:69:@21250.4]
  wire [10:0] _T_1451; // @[Mux.scala 31:69:@21251.4]
  wire  _T_1458; // @[MemPrimitives.scala 110:210:@21259.4]
  wire  _T_1459; // @[MemPrimitives.scala 110:228:@21260.4]
  wire  _T_1464; // @[MemPrimitives.scala 110:210:@21263.4]
  wire  _T_1465; // @[MemPrimitives.scala 110:228:@21264.4]
  wire  _T_1470; // @[MemPrimitives.scala 110:210:@21267.4]
  wire  _T_1471; // @[MemPrimitives.scala 110:228:@21268.4]
  wire  _T_1476; // @[MemPrimitives.scala 110:210:@21271.4]
  wire  _T_1477; // @[MemPrimitives.scala 110:228:@21272.4]
  wire  _T_1482; // @[MemPrimitives.scala 110:210:@21275.4]
  wire  _T_1483; // @[MemPrimitives.scala 110:228:@21276.4]
  wire  _T_1488; // @[MemPrimitives.scala 110:210:@21279.4]
  wire  _T_1489; // @[MemPrimitives.scala 110:228:@21280.4]
  wire  _T_1494; // @[MemPrimitives.scala 110:210:@21283.4]
  wire  _T_1495; // @[MemPrimitives.scala 110:228:@21284.4]
  wire  _T_1500; // @[MemPrimitives.scala 110:210:@21287.4]
  wire  _T_1501; // @[MemPrimitives.scala 110:228:@21288.4]
  wire  _T_1506; // @[MemPrimitives.scala 110:210:@21291.4]
  wire  _T_1507; // @[MemPrimitives.scala 110:228:@21292.4]
  wire  _T_1509; // @[MemPrimitives.scala 123:41:@21306.4]
  wire  _T_1510; // @[MemPrimitives.scala 123:41:@21307.4]
  wire  _T_1511; // @[MemPrimitives.scala 123:41:@21308.4]
  wire  _T_1512; // @[MemPrimitives.scala 123:41:@21309.4]
  wire  _T_1513; // @[MemPrimitives.scala 123:41:@21310.4]
  wire  _T_1514; // @[MemPrimitives.scala 123:41:@21311.4]
  wire  _T_1515; // @[MemPrimitives.scala 123:41:@21312.4]
  wire  _T_1516; // @[MemPrimitives.scala 123:41:@21313.4]
  wire  _T_1517; // @[MemPrimitives.scala 123:41:@21314.4]
  wire [10:0] _T_1519; // @[Cat.scala 30:58:@21316.4]
  wire [10:0] _T_1521; // @[Cat.scala 30:58:@21318.4]
  wire [10:0] _T_1523; // @[Cat.scala 30:58:@21320.4]
  wire [10:0] _T_1525; // @[Cat.scala 30:58:@21322.4]
  wire [10:0] _T_1527; // @[Cat.scala 30:58:@21324.4]
  wire [10:0] _T_1529; // @[Cat.scala 30:58:@21326.4]
  wire [10:0] _T_1531; // @[Cat.scala 30:58:@21328.4]
  wire [10:0] _T_1533; // @[Cat.scala 30:58:@21330.4]
  wire [10:0] _T_1535; // @[Cat.scala 30:58:@21332.4]
  wire [10:0] _T_1536; // @[Mux.scala 31:69:@21333.4]
  wire [10:0] _T_1537; // @[Mux.scala 31:69:@21334.4]
  wire [10:0] _T_1538; // @[Mux.scala 31:69:@21335.4]
  wire [10:0] _T_1539; // @[Mux.scala 31:69:@21336.4]
  wire [10:0] _T_1540; // @[Mux.scala 31:69:@21337.4]
  wire [10:0] _T_1541; // @[Mux.scala 31:69:@21338.4]
  wire [10:0] _T_1542; // @[Mux.scala 31:69:@21339.4]
  wire [10:0] _T_1543; // @[Mux.scala 31:69:@21340.4]
  wire  _T_1550; // @[MemPrimitives.scala 110:210:@21348.4]
  wire  _T_1551; // @[MemPrimitives.scala 110:228:@21349.4]
  wire  _T_1556; // @[MemPrimitives.scala 110:210:@21352.4]
  wire  _T_1557; // @[MemPrimitives.scala 110:228:@21353.4]
  wire  _T_1562; // @[MemPrimitives.scala 110:210:@21356.4]
  wire  _T_1563; // @[MemPrimitives.scala 110:228:@21357.4]
  wire  _T_1568; // @[MemPrimitives.scala 110:210:@21360.4]
  wire  _T_1569; // @[MemPrimitives.scala 110:228:@21361.4]
  wire  _T_1574; // @[MemPrimitives.scala 110:210:@21364.4]
  wire  _T_1575; // @[MemPrimitives.scala 110:228:@21365.4]
  wire  _T_1580; // @[MemPrimitives.scala 110:210:@21368.4]
  wire  _T_1581; // @[MemPrimitives.scala 110:228:@21369.4]
  wire  _T_1586; // @[MemPrimitives.scala 110:210:@21372.4]
  wire  _T_1587; // @[MemPrimitives.scala 110:228:@21373.4]
  wire  _T_1592; // @[MemPrimitives.scala 110:210:@21376.4]
  wire  _T_1593; // @[MemPrimitives.scala 110:228:@21377.4]
  wire  _T_1598; // @[MemPrimitives.scala 110:210:@21380.4]
  wire  _T_1599; // @[MemPrimitives.scala 110:228:@21381.4]
  wire  _T_1601; // @[MemPrimitives.scala 123:41:@21395.4]
  wire  _T_1602; // @[MemPrimitives.scala 123:41:@21396.4]
  wire  _T_1603; // @[MemPrimitives.scala 123:41:@21397.4]
  wire  _T_1604; // @[MemPrimitives.scala 123:41:@21398.4]
  wire  _T_1605; // @[MemPrimitives.scala 123:41:@21399.4]
  wire  _T_1606; // @[MemPrimitives.scala 123:41:@21400.4]
  wire  _T_1607; // @[MemPrimitives.scala 123:41:@21401.4]
  wire  _T_1608; // @[MemPrimitives.scala 123:41:@21402.4]
  wire  _T_1609; // @[MemPrimitives.scala 123:41:@21403.4]
  wire [10:0] _T_1611; // @[Cat.scala 30:58:@21405.4]
  wire [10:0] _T_1613; // @[Cat.scala 30:58:@21407.4]
  wire [10:0] _T_1615; // @[Cat.scala 30:58:@21409.4]
  wire [10:0] _T_1617; // @[Cat.scala 30:58:@21411.4]
  wire [10:0] _T_1619; // @[Cat.scala 30:58:@21413.4]
  wire [10:0] _T_1621; // @[Cat.scala 30:58:@21415.4]
  wire [10:0] _T_1623; // @[Cat.scala 30:58:@21417.4]
  wire [10:0] _T_1625; // @[Cat.scala 30:58:@21419.4]
  wire [10:0] _T_1627; // @[Cat.scala 30:58:@21421.4]
  wire [10:0] _T_1628; // @[Mux.scala 31:69:@21422.4]
  wire [10:0] _T_1629; // @[Mux.scala 31:69:@21423.4]
  wire [10:0] _T_1630; // @[Mux.scala 31:69:@21424.4]
  wire [10:0] _T_1631; // @[Mux.scala 31:69:@21425.4]
  wire [10:0] _T_1632; // @[Mux.scala 31:69:@21426.4]
  wire [10:0] _T_1633; // @[Mux.scala 31:69:@21427.4]
  wire [10:0] _T_1634; // @[Mux.scala 31:69:@21428.4]
  wire [10:0] _T_1635; // @[Mux.scala 31:69:@21429.4]
  wire  _T_1642; // @[MemPrimitives.scala 110:210:@21437.4]
  wire  _T_1643; // @[MemPrimitives.scala 110:228:@21438.4]
  wire  _T_1648; // @[MemPrimitives.scala 110:210:@21441.4]
  wire  _T_1649; // @[MemPrimitives.scala 110:228:@21442.4]
  wire  _T_1654; // @[MemPrimitives.scala 110:210:@21445.4]
  wire  _T_1655; // @[MemPrimitives.scala 110:228:@21446.4]
  wire  _T_1660; // @[MemPrimitives.scala 110:210:@21449.4]
  wire  _T_1661; // @[MemPrimitives.scala 110:228:@21450.4]
  wire  _T_1666; // @[MemPrimitives.scala 110:210:@21453.4]
  wire  _T_1667; // @[MemPrimitives.scala 110:228:@21454.4]
  wire  _T_1672; // @[MemPrimitives.scala 110:210:@21457.4]
  wire  _T_1673; // @[MemPrimitives.scala 110:228:@21458.4]
  wire  _T_1678; // @[MemPrimitives.scala 110:210:@21461.4]
  wire  _T_1679; // @[MemPrimitives.scala 110:228:@21462.4]
  wire  _T_1684; // @[MemPrimitives.scala 110:210:@21465.4]
  wire  _T_1685; // @[MemPrimitives.scala 110:228:@21466.4]
  wire  _T_1690; // @[MemPrimitives.scala 110:210:@21469.4]
  wire  _T_1691; // @[MemPrimitives.scala 110:228:@21470.4]
  wire  _T_1693; // @[MemPrimitives.scala 123:41:@21484.4]
  wire  _T_1694; // @[MemPrimitives.scala 123:41:@21485.4]
  wire  _T_1695; // @[MemPrimitives.scala 123:41:@21486.4]
  wire  _T_1696; // @[MemPrimitives.scala 123:41:@21487.4]
  wire  _T_1697; // @[MemPrimitives.scala 123:41:@21488.4]
  wire  _T_1698; // @[MemPrimitives.scala 123:41:@21489.4]
  wire  _T_1699; // @[MemPrimitives.scala 123:41:@21490.4]
  wire  _T_1700; // @[MemPrimitives.scala 123:41:@21491.4]
  wire  _T_1701; // @[MemPrimitives.scala 123:41:@21492.4]
  wire [10:0] _T_1703; // @[Cat.scala 30:58:@21494.4]
  wire [10:0] _T_1705; // @[Cat.scala 30:58:@21496.4]
  wire [10:0] _T_1707; // @[Cat.scala 30:58:@21498.4]
  wire [10:0] _T_1709; // @[Cat.scala 30:58:@21500.4]
  wire [10:0] _T_1711; // @[Cat.scala 30:58:@21502.4]
  wire [10:0] _T_1713; // @[Cat.scala 30:58:@21504.4]
  wire [10:0] _T_1715; // @[Cat.scala 30:58:@21506.4]
  wire [10:0] _T_1717; // @[Cat.scala 30:58:@21508.4]
  wire [10:0] _T_1719; // @[Cat.scala 30:58:@21510.4]
  wire [10:0] _T_1720; // @[Mux.scala 31:69:@21511.4]
  wire [10:0] _T_1721; // @[Mux.scala 31:69:@21512.4]
  wire [10:0] _T_1722; // @[Mux.scala 31:69:@21513.4]
  wire [10:0] _T_1723; // @[Mux.scala 31:69:@21514.4]
  wire [10:0] _T_1724; // @[Mux.scala 31:69:@21515.4]
  wire [10:0] _T_1725; // @[Mux.scala 31:69:@21516.4]
  wire [10:0] _T_1726; // @[Mux.scala 31:69:@21517.4]
  wire [10:0] _T_1727; // @[Mux.scala 31:69:@21518.4]
  wire  _T_1732; // @[MemPrimitives.scala 110:210:@21525.4]
  wire  _T_1735; // @[MemPrimitives.scala 110:228:@21527.4]
  wire  _T_1738; // @[MemPrimitives.scala 110:210:@21529.4]
  wire  _T_1741; // @[MemPrimitives.scala 110:228:@21531.4]
  wire  _T_1744; // @[MemPrimitives.scala 110:210:@21533.4]
  wire  _T_1747; // @[MemPrimitives.scala 110:228:@21535.4]
  wire  _T_1750; // @[MemPrimitives.scala 110:210:@21537.4]
  wire  _T_1753; // @[MemPrimitives.scala 110:228:@21539.4]
  wire  _T_1756; // @[MemPrimitives.scala 110:210:@21541.4]
  wire  _T_1759; // @[MemPrimitives.scala 110:228:@21543.4]
  wire  _T_1762; // @[MemPrimitives.scala 110:210:@21545.4]
  wire  _T_1765; // @[MemPrimitives.scala 110:228:@21547.4]
  wire  _T_1768; // @[MemPrimitives.scala 110:210:@21549.4]
  wire  _T_1771; // @[MemPrimitives.scala 110:228:@21551.4]
  wire  _T_1774; // @[MemPrimitives.scala 110:210:@21553.4]
  wire  _T_1777; // @[MemPrimitives.scala 110:228:@21555.4]
  wire  _T_1780; // @[MemPrimitives.scala 110:210:@21557.4]
  wire  _T_1783; // @[MemPrimitives.scala 110:228:@21559.4]
  wire  _T_1785; // @[MemPrimitives.scala 123:41:@21573.4]
  wire  _T_1786; // @[MemPrimitives.scala 123:41:@21574.4]
  wire  _T_1787; // @[MemPrimitives.scala 123:41:@21575.4]
  wire  _T_1788; // @[MemPrimitives.scala 123:41:@21576.4]
  wire  _T_1789; // @[MemPrimitives.scala 123:41:@21577.4]
  wire  _T_1790; // @[MemPrimitives.scala 123:41:@21578.4]
  wire  _T_1791; // @[MemPrimitives.scala 123:41:@21579.4]
  wire  _T_1792; // @[MemPrimitives.scala 123:41:@21580.4]
  wire  _T_1793; // @[MemPrimitives.scala 123:41:@21581.4]
  wire [10:0] _T_1795; // @[Cat.scala 30:58:@21583.4]
  wire [10:0] _T_1797; // @[Cat.scala 30:58:@21585.4]
  wire [10:0] _T_1799; // @[Cat.scala 30:58:@21587.4]
  wire [10:0] _T_1801; // @[Cat.scala 30:58:@21589.4]
  wire [10:0] _T_1803; // @[Cat.scala 30:58:@21591.4]
  wire [10:0] _T_1805; // @[Cat.scala 30:58:@21593.4]
  wire [10:0] _T_1807; // @[Cat.scala 30:58:@21595.4]
  wire [10:0] _T_1809; // @[Cat.scala 30:58:@21597.4]
  wire [10:0] _T_1811; // @[Cat.scala 30:58:@21599.4]
  wire [10:0] _T_1812; // @[Mux.scala 31:69:@21600.4]
  wire [10:0] _T_1813; // @[Mux.scala 31:69:@21601.4]
  wire [10:0] _T_1814; // @[Mux.scala 31:69:@21602.4]
  wire [10:0] _T_1815; // @[Mux.scala 31:69:@21603.4]
  wire [10:0] _T_1816; // @[Mux.scala 31:69:@21604.4]
  wire [10:0] _T_1817; // @[Mux.scala 31:69:@21605.4]
  wire [10:0] _T_1818; // @[Mux.scala 31:69:@21606.4]
  wire [10:0] _T_1819; // @[Mux.scala 31:69:@21607.4]
  wire  _T_1824; // @[MemPrimitives.scala 110:210:@21614.4]
  wire  _T_1827; // @[MemPrimitives.scala 110:228:@21616.4]
  wire  _T_1830; // @[MemPrimitives.scala 110:210:@21618.4]
  wire  _T_1833; // @[MemPrimitives.scala 110:228:@21620.4]
  wire  _T_1836; // @[MemPrimitives.scala 110:210:@21622.4]
  wire  _T_1839; // @[MemPrimitives.scala 110:228:@21624.4]
  wire  _T_1842; // @[MemPrimitives.scala 110:210:@21626.4]
  wire  _T_1845; // @[MemPrimitives.scala 110:228:@21628.4]
  wire  _T_1848; // @[MemPrimitives.scala 110:210:@21630.4]
  wire  _T_1851; // @[MemPrimitives.scala 110:228:@21632.4]
  wire  _T_1854; // @[MemPrimitives.scala 110:210:@21634.4]
  wire  _T_1857; // @[MemPrimitives.scala 110:228:@21636.4]
  wire  _T_1860; // @[MemPrimitives.scala 110:210:@21638.4]
  wire  _T_1863; // @[MemPrimitives.scala 110:228:@21640.4]
  wire  _T_1866; // @[MemPrimitives.scala 110:210:@21642.4]
  wire  _T_1869; // @[MemPrimitives.scala 110:228:@21644.4]
  wire  _T_1872; // @[MemPrimitives.scala 110:210:@21646.4]
  wire  _T_1875; // @[MemPrimitives.scala 110:228:@21648.4]
  wire  _T_1877; // @[MemPrimitives.scala 123:41:@21662.4]
  wire  _T_1878; // @[MemPrimitives.scala 123:41:@21663.4]
  wire  _T_1879; // @[MemPrimitives.scala 123:41:@21664.4]
  wire  _T_1880; // @[MemPrimitives.scala 123:41:@21665.4]
  wire  _T_1881; // @[MemPrimitives.scala 123:41:@21666.4]
  wire  _T_1882; // @[MemPrimitives.scala 123:41:@21667.4]
  wire  _T_1883; // @[MemPrimitives.scala 123:41:@21668.4]
  wire  _T_1884; // @[MemPrimitives.scala 123:41:@21669.4]
  wire  _T_1885; // @[MemPrimitives.scala 123:41:@21670.4]
  wire [10:0] _T_1887; // @[Cat.scala 30:58:@21672.4]
  wire [10:0] _T_1889; // @[Cat.scala 30:58:@21674.4]
  wire [10:0] _T_1891; // @[Cat.scala 30:58:@21676.4]
  wire [10:0] _T_1893; // @[Cat.scala 30:58:@21678.4]
  wire [10:0] _T_1895; // @[Cat.scala 30:58:@21680.4]
  wire [10:0] _T_1897; // @[Cat.scala 30:58:@21682.4]
  wire [10:0] _T_1899; // @[Cat.scala 30:58:@21684.4]
  wire [10:0] _T_1901; // @[Cat.scala 30:58:@21686.4]
  wire [10:0] _T_1903; // @[Cat.scala 30:58:@21688.4]
  wire [10:0] _T_1904; // @[Mux.scala 31:69:@21689.4]
  wire [10:0] _T_1905; // @[Mux.scala 31:69:@21690.4]
  wire [10:0] _T_1906; // @[Mux.scala 31:69:@21691.4]
  wire [10:0] _T_1907; // @[Mux.scala 31:69:@21692.4]
  wire [10:0] _T_1908; // @[Mux.scala 31:69:@21693.4]
  wire [10:0] _T_1909; // @[Mux.scala 31:69:@21694.4]
  wire [10:0] _T_1910; // @[Mux.scala 31:69:@21695.4]
  wire [10:0] _T_1911; // @[Mux.scala 31:69:@21696.4]
  wire  _T_1919; // @[MemPrimitives.scala 110:228:@21705.4]
  wire  _T_1925; // @[MemPrimitives.scala 110:228:@21709.4]
  wire  _T_1931; // @[MemPrimitives.scala 110:228:@21713.4]
  wire  _T_1937; // @[MemPrimitives.scala 110:228:@21717.4]
  wire  _T_1943; // @[MemPrimitives.scala 110:228:@21721.4]
  wire  _T_1949; // @[MemPrimitives.scala 110:228:@21725.4]
  wire  _T_1955; // @[MemPrimitives.scala 110:228:@21729.4]
  wire  _T_1961; // @[MemPrimitives.scala 110:228:@21733.4]
  wire  _T_1967; // @[MemPrimitives.scala 110:228:@21737.4]
  wire  _T_1969; // @[MemPrimitives.scala 123:41:@21751.4]
  wire  _T_1970; // @[MemPrimitives.scala 123:41:@21752.4]
  wire  _T_1971; // @[MemPrimitives.scala 123:41:@21753.4]
  wire  _T_1972; // @[MemPrimitives.scala 123:41:@21754.4]
  wire  _T_1973; // @[MemPrimitives.scala 123:41:@21755.4]
  wire  _T_1974; // @[MemPrimitives.scala 123:41:@21756.4]
  wire  _T_1975; // @[MemPrimitives.scala 123:41:@21757.4]
  wire  _T_1976; // @[MemPrimitives.scala 123:41:@21758.4]
  wire  _T_1977; // @[MemPrimitives.scala 123:41:@21759.4]
  wire [10:0] _T_1979; // @[Cat.scala 30:58:@21761.4]
  wire [10:0] _T_1981; // @[Cat.scala 30:58:@21763.4]
  wire [10:0] _T_1983; // @[Cat.scala 30:58:@21765.4]
  wire [10:0] _T_1985; // @[Cat.scala 30:58:@21767.4]
  wire [10:0] _T_1987; // @[Cat.scala 30:58:@21769.4]
  wire [10:0] _T_1989; // @[Cat.scala 30:58:@21771.4]
  wire [10:0] _T_1991; // @[Cat.scala 30:58:@21773.4]
  wire [10:0] _T_1993; // @[Cat.scala 30:58:@21775.4]
  wire [10:0] _T_1995; // @[Cat.scala 30:58:@21777.4]
  wire [10:0] _T_1996; // @[Mux.scala 31:69:@21778.4]
  wire [10:0] _T_1997; // @[Mux.scala 31:69:@21779.4]
  wire [10:0] _T_1998; // @[Mux.scala 31:69:@21780.4]
  wire [10:0] _T_1999; // @[Mux.scala 31:69:@21781.4]
  wire [10:0] _T_2000; // @[Mux.scala 31:69:@21782.4]
  wire [10:0] _T_2001; // @[Mux.scala 31:69:@21783.4]
  wire [10:0] _T_2002; // @[Mux.scala 31:69:@21784.4]
  wire [10:0] _T_2003; // @[Mux.scala 31:69:@21785.4]
  wire  _T_2011; // @[MemPrimitives.scala 110:228:@21794.4]
  wire  _T_2017; // @[MemPrimitives.scala 110:228:@21798.4]
  wire  _T_2023; // @[MemPrimitives.scala 110:228:@21802.4]
  wire  _T_2029; // @[MemPrimitives.scala 110:228:@21806.4]
  wire  _T_2035; // @[MemPrimitives.scala 110:228:@21810.4]
  wire  _T_2041; // @[MemPrimitives.scala 110:228:@21814.4]
  wire  _T_2047; // @[MemPrimitives.scala 110:228:@21818.4]
  wire  _T_2053; // @[MemPrimitives.scala 110:228:@21822.4]
  wire  _T_2059; // @[MemPrimitives.scala 110:228:@21826.4]
  wire  _T_2061; // @[MemPrimitives.scala 123:41:@21840.4]
  wire  _T_2062; // @[MemPrimitives.scala 123:41:@21841.4]
  wire  _T_2063; // @[MemPrimitives.scala 123:41:@21842.4]
  wire  _T_2064; // @[MemPrimitives.scala 123:41:@21843.4]
  wire  _T_2065; // @[MemPrimitives.scala 123:41:@21844.4]
  wire  _T_2066; // @[MemPrimitives.scala 123:41:@21845.4]
  wire  _T_2067; // @[MemPrimitives.scala 123:41:@21846.4]
  wire  _T_2068; // @[MemPrimitives.scala 123:41:@21847.4]
  wire  _T_2069; // @[MemPrimitives.scala 123:41:@21848.4]
  wire [10:0] _T_2071; // @[Cat.scala 30:58:@21850.4]
  wire [10:0] _T_2073; // @[Cat.scala 30:58:@21852.4]
  wire [10:0] _T_2075; // @[Cat.scala 30:58:@21854.4]
  wire [10:0] _T_2077; // @[Cat.scala 30:58:@21856.4]
  wire [10:0] _T_2079; // @[Cat.scala 30:58:@21858.4]
  wire [10:0] _T_2081; // @[Cat.scala 30:58:@21860.4]
  wire [10:0] _T_2083; // @[Cat.scala 30:58:@21862.4]
  wire [10:0] _T_2085; // @[Cat.scala 30:58:@21864.4]
  wire [10:0] _T_2087; // @[Cat.scala 30:58:@21866.4]
  wire [10:0] _T_2088; // @[Mux.scala 31:69:@21867.4]
  wire [10:0] _T_2089; // @[Mux.scala 31:69:@21868.4]
  wire [10:0] _T_2090; // @[Mux.scala 31:69:@21869.4]
  wire [10:0] _T_2091; // @[Mux.scala 31:69:@21870.4]
  wire [10:0] _T_2092; // @[Mux.scala 31:69:@21871.4]
  wire [10:0] _T_2093; // @[Mux.scala 31:69:@21872.4]
  wire [10:0] _T_2094; // @[Mux.scala 31:69:@21873.4]
  wire [10:0] _T_2095; // @[Mux.scala 31:69:@21874.4]
  wire  _T_2103; // @[MemPrimitives.scala 110:228:@21883.4]
  wire  _T_2109; // @[MemPrimitives.scala 110:228:@21887.4]
  wire  _T_2115; // @[MemPrimitives.scala 110:228:@21891.4]
  wire  _T_2121; // @[MemPrimitives.scala 110:228:@21895.4]
  wire  _T_2127; // @[MemPrimitives.scala 110:228:@21899.4]
  wire  _T_2133; // @[MemPrimitives.scala 110:228:@21903.4]
  wire  _T_2139; // @[MemPrimitives.scala 110:228:@21907.4]
  wire  _T_2145; // @[MemPrimitives.scala 110:228:@21911.4]
  wire  _T_2151; // @[MemPrimitives.scala 110:228:@21915.4]
  wire  _T_2153; // @[MemPrimitives.scala 123:41:@21929.4]
  wire  _T_2154; // @[MemPrimitives.scala 123:41:@21930.4]
  wire  _T_2155; // @[MemPrimitives.scala 123:41:@21931.4]
  wire  _T_2156; // @[MemPrimitives.scala 123:41:@21932.4]
  wire  _T_2157; // @[MemPrimitives.scala 123:41:@21933.4]
  wire  _T_2158; // @[MemPrimitives.scala 123:41:@21934.4]
  wire  _T_2159; // @[MemPrimitives.scala 123:41:@21935.4]
  wire  _T_2160; // @[MemPrimitives.scala 123:41:@21936.4]
  wire  _T_2161; // @[MemPrimitives.scala 123:41:@21937.4]
  wire [10:0] _T_2163; // @[Cat.scala 30:58:@21939.4]
  wire [10:0] _T_2165; // @[Cat.scala 30:58:@21941.4]
  wire [10:0] _T_2167; // @[Cat.scala 30:58:@21943.4]
  wire [10:0] _T_2169; // @[Cat.scala 30:58:@21945.4]
  wire [10:0] _T_2171; // @[Cat.scala 30:58:@21947.4]
  wire [10:0] _T_2173; // @[Cat.scala 30:58:@21949.4]
  wire [10:0] _T_2175; // @[Cat.scala 30:58:@21951.4]
  wire [10:0] _T_2177; // @[Cat.scala 30:58:@21953.4]
  wire [10:0] _T_2179; // @[Cat.scala 30:58:@21955.4]
  wire [10:0] _T_2180; // @[Mux.scala 31:69:@21956.4]
  wire [10:0] _T_2181; // @[Mux.scala 31:69:@21957.4]
  wire [10:0] _T_2182; // @[Mux.scala 31:69:@21958.4]
  wire [10:0] _T_2183; // @[Mux.scala 31:69:@21959.4]
  wire [10:0] _T_2184; // @[Mux.scala 31:69:@21960.4]
  wire [10:0] _T_2185; // @[Mux.scala 31:69:@21961.4]
  wire [10:0] _T_2186; // @[Mux.scala 31:69:@21962.4]
  wire [10:0] _T_2187; // @[Mux.scala 31:69:@21963.4]
  wire  _T_2195; // @[MemPrimitives.scala 110:228:@21972.4]
  wire  _T_2201; // @[MemPrimitives.scala 110:228:@21976.4]
  wire  _T_2207; // @[MemPrimitives.scala 110:228:@21980.4]
  wire  _T_2213; // @[MemPrimitives.scala 110:228:@21984.4]
  wire  _T_2219; // @[MemPrimitives.scala 110:228:@21988.4]
  wire  _T_2225; // @[MemPrimitives.scala 110:228:@21992.4]
  wire  _T_2231; // @[MemPrimitives.scala 110:228:@21996.4]
  wire  _T_2237; // @[MemPrimitives.scala 110:228:@22000.4]
  wire  _T_2243; // @[MemPrimitives.scala 110:228:@22004.4]
  wire  _T_2245; // @[MemPrimitives.scala 123:41:@22018.4]
  wire  _T_2246; // @[MemPrimitives.scala 123:41:@22019.4]
  wire  _T_2247; // @[MemPrimitives.scala 123:41:@22020.4]
  wire  _T_2248; // @[MemPrimitives.scala 123:41:@22021.4]
  wire  _T_2249; // @[MemPrimitives.scala 123:41:@22022.4]
  wire  _T_2250; // @[MemPrimitives.scala 123:41:@22023.4]
  wire  _T_2251; // @[MemPrimitives.scala 123:41:@22024.4]
  wire  _T_2252; // @[MemPrimitives.scala 123:41:@22025.4]
  wire  _T_2253; // @[MemPrimitives.scala 123:41:@22026.4]
  wire [10:0] _T_2255; // @[Cat.scala 30:58:@22028.4]
  wire [10:0] _T_2257; // @[Cat.scala 30:58:@22030.4]
  wire [10:0] _T_2259; // @[Cat.scala 30:58:@22032.4]
  wire [10:0] _T_2261; // @[Cat.scala 30:58:@22034.4]
  wire [10:0] _T_2263; // @[Cat.scala 30:58:@22036.4]
  wire [10:0] _T_2265; // @[Cat.scala 30:58:@22038.4]
  wire [10:0] _T_2267; // @[Cat.scala 30:58:@22040.4]
  wire [10:0] _T_2269; // @[Cat.scala 30:58:@22042.4]
  wire [10:0] _T_2271; // @[Cat.scala 30:58:@22044.4]
  wire [10:0] _T_2272; // @[Mux.scala 31:69:@22045.4]
  wire [10:0] _T_2273; // @[Mux.scala 31:69:@22046.4]
  wire [10:0] _T_2274; // @[Mux.scala 31:69:@22047.4]
  wire [10:0] _T_2275; // @[Mux.scala 31:69:@22048.4]
  wire [10:0] _T_2276; // @[Mux.scala 31:69:@22049.4]
  wire [10:0] _T_2277; // @[Mux.scala 31:69:@22050.4]
  wire [10:0] _T_2278; // @[Mux.scala 31:69:@22051.4]
  wire [10:0] _T_2279; // @[Mux.scala 31:69:@22052.4]
  wire  _T_2284; // @[MemPrimitives.scala 110:210:@22059.4]
  wire  _T_2287; // @[MemPrimitives.scala 110:228:@22061.4]
  wire  _T_2290; // @[MemPrimitives.scala 110:210:@22063.4]
  wire  _T_2293; // @[MemPrimitives.scala 110:228:@22065.4]
  wire  _T_2296; // @[MemPrimitives.scala 110:210:@22067.4]
  wire  _T_2299; // @[MemPrimitives.scala 110:228:@22069.4]
  wire  _T_2302; // @[MemPrimitives.scala 110:210:@22071.4]
  wire  _T_2305; // @[MemPrimitives.scala 110:228:@22073.4]
  wire  _T_2308; // @[MemPrimitives.scala 110:210:@22075.4]
  wire  _T_2311; // @[MemPrimitives.scala 110:228:@22077.4]
  wire  _T_2314; // @[MemPrimitives.scala 110:210:@22079.4]
  wire  _T_2317; // @[MemPrimitives.scala 110:228:@22081.4]
  wire  _T_2320; // @[MemPrimitives.scala 110:210:@22083.4]
  wire  _T_2323; // @[MemPrimitives.scala 110:228:@22085.4]
  wire  _T_2326; // @[MemPrimitives.scala 110:210:@22087.4]
  wire  _T_2329; // @[MemPrimitives.scala 110:228:@22089.4]
  wire  _T_2332; // @[MemPrimitives.scala 110:210:@22091.4]
  wire  _T_2335; // @[MemPrimitives.scala 110:228:@22093.4]
  wire  _T_2337; // @[MemPrimitives.scala 123:41:@22107.4]
  wire  _T_2338; // @[MemPrimitives.scala 123:41:@22108.4]
  wire  _T_2339; // @[MemPrimitives.scala 123:41:@22109.4]
  wire  _T_2340; // @[MemPrimitives.scala 123:41:@22110.4]
  wire  _T_2341; // @[MemPrimitives.scala 123:41:@22111.4]
  wire  _T_2342; // @[MemPrimitives.scala 123:41:@22112.4]
  wire  _T_2343; // @[MemPrimitives.scala 123:41:@22113.4]
  wire  _T_2344; // @[MemPrimitives.scala 123:41:@22114.4]
  wire  _T_2345; // @[MemPrimitives.scala 123:41:@22115.4]
  wire [10:0] _T_2347; // @[Cat.scala 30:58:@22117.4]
  wire [10:0] _T_2349; // @[Cat.scala 30:58:@22119.4]
  wire [10:0] _T_2351; // @[Cat.scala 30:58:@22121.4]
  wire [10:0] _T_2353; // @[Cat.scala 30:58:@22123.4]
  wire [10:0] _T_2355; // @[Cat.scala 30:58:@22125.4]
  wire [10:0] _T_2357; // @[Cat.scala 30:58:@22127.4]
  wire [10:0] _T_2359; // @[Cat.scala 30:58:@22129.4]
  wire [10:0] _T_2361; // @[Cat.scala 30:58:@22131.4]
  wire [10:0] _T_2363; // @[Cat.scala 30:58:@22133.4]
  wire [10:0] _T_2364; // @[Mux.scala 31:69:@22134.4]
  wire [10:0] _T_2365; // @[Mux.scala 31:69:@22135.4]
  wire [10:0] _T_2366; // @[Mux.scala 31:69:@22136.4]
  wire [10:0] _T_2367; // @[Mux.scala 31:69:@22137.4]
  wire [10:0] _T_2368; // @[Mux.scala 31:69:@22138.4]
  wire [10:0] _T_2369; // @[Mux.scala 31:69:@22139.4]
  wire [10:0] _T_2370; // @[Mux.scala 31:69:@22140.4]
  wire [10:0] _T_2371; // @[Mux.scala 31:69:@22141.4]
  wire  _T_2376; // @[MemPrimitives.scala 110:210:@22148.4]
  wire  _T_2379; // @[MemPrimitives.scala 110:228:@22150.4]
  wire  _T_2382; // @[MemPrimitives.scala 110:210:@22152.4]
  wire  _T_2385; // @[MemPrimitives.scala 110:228:@22154.4]
  wire  _T_2388; // @[MemPrimitives.scala 110:210:@22156.4]
  wire  _T_2391; // @[MemPrimitives.scala 110:228:@22158.4]
  wire  _T_2394; // @[MemPrimitives.scala 110:210:@22160.4]
  wire  _T_2397; // @[MemPrimitives.scala 110:228:@22162.4]
  wire  _T_2400; // @[MemPrimitives.scala 110:210:@22164.4]
  wire  _T_2403; // @[MemPrimitives.scala 110:228:@22166.4]
  wire  _T_2406; // @[MemPrimitives.scala 110:210:@22168.4]
  wire  _T_2409; // @[MemPrimitives.scala 110:228:@22170.4]
  wire  _T_2412; // @[MemPrimitives.scala 110:210:@22172.4]
  wire  _T_2415; // @[MemPrimitives.scala 110:228:@22174.4]
  wire  _T_2418; // @[MemPrimitives.scala 110:210:@22176.4]
  wire  _T_2421; // @[MemPrimitives.scala 110:228:@22178.4]
  wire  _T_2424; // @[MemPrimitives.scala 110:210:@22180.4]
  wire  _T_2427; // @[MemPrimitives.scala 110:228:@22182.4]
  wire  _T_2429; // @[MemPrimitives.scala 123:41:@22196.4]
  wire  _T_2430; // @[MemPrimitives.scala 123:41:@22197.4]
  wire  _T_2431; // @[MemPrimitives.scala 123:41:@22198.4]
  wire  _T_2432; // @[MemPrimitives.scala 123:41:@22199.4]
  wire  _T_2433; // @[MemPrimitives.scala 123:41:@22200.4]
  wire  _T_2434; // @[MemPrimitives.scala 123:41:@22201.4]
  wire  _T_2435; // @[MemPrimitives.scala 123:41:@22202.4]
  wire  _T_2436; // @[MemPrimitives.scala 123:41:@22203.4]
  wire  _T_2437; // @[MemPrimitives.scala 123:41:@22204.4]
  wire [10:0] _T_2439; // @[Cat.scala 30:58:@22206.4]
  wire [10:0] _T_2441; // @[Cat.scala 30:58:@22208.4]
  wire [10:0] _T_2443; // @[Cat.scala 30:58:@22210.4]
  wire [10:0] _T_2445; // @[Cat.scala 30:58:@22212.4]
  wire [10:0] _T_2447; // @[Cat.scala 30:58:@22214.4]
  wire [10:0] _T_2449; // @[Cat.scala 30:58:@22216.4]
  wire [10:0] _T_2451; // @[Cat.scala 30:58:@22218.4]
  wire [10:0] _T_2453; // @[Cat.scala 30:58:@22220.4]
  wire [10:0] _T_2455; // @[Cat.scala 30:58:@22222.4]
  wire [10:0] _T_2456; // @[Mux.scala 31:69:@22223.4]
  wire [10:0] _T_2457; // @[Mux.scala 31:69:@22224.4]
  wire [10:0] _T_2458; // @[Mux.scala 31:69:@22225.4]
  wire [10:0] _T_2459; // @[Mux.scala 31:69:@22226.4]
  wire [10:0] _T_2460; // @[Mux.scala 31:69:@22227.4]
  wire [10:0] _T_2461; // @[Mux.scala 31:69:@22228.4]
  wire [10:0] _T_2462; // @[Mux.scala 31:69:@22229.4]
  wire [10:0] _T_2463; // @[Mux.scala 31:69:@22230.4]
  wire  _T_2471; // @[MemPrimitives.scala 110:228:@22239.4]
  wire  _T_2477; // @[MemPrimitives.scala 110:228:@22243.4]
  wire  _T_2483; // @[MemPrimitives.scala 110:228:@22247.4]
  wire  _T_2489; // @[MemPrimitives.scala 110:228:@22251.4]
  wire  _T_2495; // @[MemPrimitives.scala 110:228:@22255.4]
  wire  _T_2501; // @[MemPrimitives.scala 110:228:@22259.4]
  wire  _T_2507; // @[MemPrimitives.scala 110:228:@22263.4]
  wire  _T_2513; // @[MemPrimitives.scala 110:228:@22267.4]
  wire  _T_2519; // @[MemPrimitives.scala 110:228:@22271.4]
  wire  _T_2521; // @[MemPrimitives.scala 123:41:@22285.4]
  wire  _T_2522; // @[MemPrimitives.scala 123:41:@22286.4]
  wire  _T_2523; // @[MemPrimitives.scala 123:41:@22287.4]
  wire  _T_2524; // @[MemPrimitives.scala 123:41:@22288.4]
  wire  _T_2525; // @[MemPrimitives.scala 123:41:@22289.4]
  wire  _T_2526; // @[MemPrimitives.scala 123:41:@22290.4]
  wire  _T_2527; // @[MemPrimitives.scala 123:41:@22291.4]
  wire  _T_2528; // @[MemPrimitives.scala 123:41:@22292.4]
  wire  _T_2529; // @[MemPrimitives.scala 123:41:@22293.4]
  wire [10:0] _T_2531; // @[Cat.scala 30:58:@22295.4]
  wire [10:0] _T_2533; // @[Cat.scala 30:58:@22297.4]
  wire [10:0] _T_2535; // @[Cat.scala 30:58:@22299.4]
  wire [10:0] _T_2537; // @[Cat.scala 30:58:@22301.4]
  wire [10:0] _T_2539; // @[Cat.scala 30:58:@22303.4]
  wire [10:0] _T_2541; // @[Cat.scala 30:58:@22305.4]
  wire [10:0] _T_2543; // @[Cat.scala 30:58:@22307.4]
  wire [10:0] _T_2545; // @[Cat.scala 30:58:@22309.4]
  wire [10:0] _T_2547; // @[Cat.scala 30:58:@22311.4]
  wire [10:0] _T_2548; // @[Mux.scala 31:69:@22312.4]
  wire [10:0] _T_2549; // @[Mux.scala 31:69:@22313.4]
  wire [10:0] _T_2550; // @[Mux.scala 31:69:@22314.4]
  wire [10:0] _T_2551; // @[Mux.scala 31:69:@22315.4]
  wire [10:0] _T_2552; // @[Mux.scala 31:69:@22316.4]
  wire [10:0] _T_2553; // @[Mux.scala 31:69:@22317.4]
  wire [10:0] _T_2554; // @[Mux.scala 31:69:@22318.4]
  wire [10:0] _T_2555; // @[Mux.scala 31:69:@22319.4]
  wire  _T_2563; // @[MemPrimitives.scala 110:228:@22328.4]
  wire  _T_2569; // @[MemPrimitives.scala 110:228:@22332.4]
  wire  _T_2575; // @[MemPrimitives.scala 110:228:@22336.4]
  wire  _T_2581; // @[MemPrimitives.scala 110:228:@22340.4]
  wire  _T_2587; // @[MemPrimitives.scala 110:228:@22344.4]
  wire  _T_2593; // @[MemPrimitives.scala 110:228:@22348.4]
  wire  _T_2599; // @[MemPrimitives.scala 110:228:@22352.4]
  wire  _T_2605; // @[MemPrimitives.scala 110:228:@22356.4]
  wire  _T_2611; // @[MemPrimitives.scala 110:228:@22360.4]
  wire  _T_2613; // @[MemPrimitives.scala 123:41:@22374.4]
  wire  _T_2614; // @[MemPrimitives.scala 123:41:@22375.4]
  wire  _T_2615; // @[MemPrimitives.scala 123:41:@22376.4]
  wire  _T_2616; // @[MemPrimitives.scala 123:41:@22377.4]
  wire  _T_2617; // @[MemPrimitives.scala 123:41:@22378.4]
  wire  _T_2618; // @[MemPrimitives.scala 123:41:@22379.4]
  wire  _T_2619; // @[MemPrimitives.scala 123:41:@22380.4]
  wire  _T_2620; // @[MemPrimitives.scala 123:41:@22381.4]
  wire  _T_2621; // @[MemPrimitives.scala 123:41:@22382.4]
  wire [10:0] _T_2623; // @[Cat.scala 30:58:@22384.4]
  wire [10:0] _T_2625; // @[Cat.scala 30:58:@22386.4]
  wire [10:0] _T_2627; // @[Cat.scala 30:58:@22388.4]
  wire [10:0] _T_2629; // @[Cat.scala 30:58:@22390.4]
  wire [10:0] _T_2631; // @[Cat.scala 30:58:@22392.4]
  wire [10:0] _T_2633; // @[Cat.scala 30:58:@22394.4]
  wire [10:0] _T_2635; // @[Cat.scala 30:58:@22396.4]
  wire [10:0] _T_2637; // @[Cat.scala 30:58:@22398.4]
  wire [10:0] _T_2639; // @[Cat.scala 30:58:@22400.4]
  wire [10:0] _T_2640; // @[Mux.scala 31:69:@22401.4]
  wire [10:0] _T_2641; // @[Mux.scala 31:69:@22402.4]
  wire [10:0] _T_2642; // @[Mux.scala 31:69:@22403.4]
  wire [10:0] _T_2643; // @[Mux.scala 31:69:@22404.4]
  wire [10:0] _T_2644; // @[Mux.scala 31:69:@22405.4]
  wire [10:0] _T_2645; // @[Mux.scala 31:69:@22406.4]
  wire [10:0] _T_2646; // @[Mux.scala 31:69:@22407.4]
  wire [10:0] _T_2647; // @[Mux.scala 31:69:@22408.4]
  wire  _T_2655; // @[MemPrimitives.scala 110:228:@22417.4]
  wire  _T_2661; // @[MemPrimitives.scala 110:228:@22421.4]
  wire  _T_2667; // @[MemPrimitives.scala 110:228:@22425.4]
  wire  _T_2673; // @[MemPrimitives.scala 110:228:@22429.4]
  wire  _T_2679; // @[MemPrimitives.scala 110:228:@22433.4]
  wire  _T_2685; // @[MemPrimitives.scala 110:228:@22437.4]
  wire  _T_2691; // @[MemPrimitives.scala 110:228:@22441.4]
  wire  _T_2697; // @[MemPrimitives.scala 110:228:@22445.4]
  wire  _T_2703; // @[MemPrimitives.scala 110:228:@22449.4]
  wire  _T_2705; // @[MemPrimitives.scala 123:41:@22463.4]
  wire  _T_2706; // @[MemPrimitives.scala 123:41:@22464.4]
  wire  _T_2707; // @[MemPrimitives.scala 123:41:@22465.4]
  wire  _T_2708; // @[MemPrimitives.scala 123:41:@22466.4]
  wire  _T_2709; // @[MemPrimitives.scala 123:41:@22467.4]
  wire  _T_2710; // @[MemPrimitives.scala 123:41:@22468.4]
  wire  _T_2711; // @[MemPrimitives.scala 123:41:@22469.4]
  wire  _T_2712; // @[MemPrimitives.scala 123:41:@22470.4]
  wire  _T_2713; // @[MemPrimitives.scala 123:41:@22471.4]
  wire [10:0] _T_2715; // @[Cat.scala 30:58:@22473.4]
  wire [10:0] _T_2717; // @[Cat.scala 30:58:@22475.4]
  wire [10:0] _T_2719; // @[Cat.scala 30:58:@22477.4]
  wire [10:0] _T_2721; // @[Cat.scala 30:58:@22479.4]
  wire [10:0] _T_2723; // @[Cat.scala 30:58:@22481.4]
  wire [10:0] _T_2725; // @[Cat.scala 30:58:@22483.4]
  wire [10:0] _T_2727; // @[Cat.scala 30:58:@22485.4]
  wire [10:0] _T_2729; // @[Cat.scala 30:58:@22487.4]
  wire [10:0] _T_2731; // @[Cat.scala 30:58:@22489.4]
  wire [10:0] _T_2732; // @[Mux.scala 31:69:@22490.4]
  wire [10:0] _T_2733; // @[Mux.scala 31:69:@22491.4]
  wire [10:0] _T_2734; // @[Mux.scala 31:69:@22492.4]
  wire [10:0] _T_2735; // @[Mux.scala 31:69:@22493.4]
  wire [10:0] _T_2736; // @[Mux.scala 31:69:@22494.4]
  wire [10:0] _T_2737; // @[Mux.scala 31:69:@22495.4]
  wire [10:0] _T_2738; // @[Mux.scala 31:69:@22496.4]
  wire [10:0] _T_2739; // @[Mux.scala 31:69:@22497.4]
  wire  _T_2747; // @[MemPrimitives.scala 110:228:@22506.4]
  wire  _T_2753; // @[MemPrimitives.scala 110:228:@22510.4]
  wire  _T_2759; // @[MemPrimitives.scala 110:228:@22514.4]
  wire  _T_2765; // @[MemPrimitives.scala 110:228:@22518.4]
  wire  _T_2771; // @[MemPrimitives.scala 110:228:@22522.4]
  wire  _T_2777; // @[MemPrimitives.scala 110:228:@22526.4]
  wire  _T_2783; // @[MemPrimitives.scala 110:228:@22530.4]
  wire  _T_2789; // @[MemPrimitives.scala 110:228:@22534.4]
  wire  _T_2795; // @[MemPrimitives.scala 110:228:@22538.4]
  wire  _T_2797; // @[MemPrimitives.scala 123:41:@22552.4]
  wire  _T_2798; // @[MemPrimitives.scala 123:41:@22553.4]
  wire  _T_2799; // @[MemPrimitives.scala 123:41:@22554.4]
  wire  _T_2800; // @[MemPrimitives.scala 123:41:@22555.4]
  wire  _T_2801; // @[MemPrimitives.scala 123:41:@22556.4]
  wire  _T_2802; // @[MemPrimitives.scala 123:41:@22557.4]
  wire  _T_2803; // @[MemPrimitives.scala 123:41:@22558.4]
  wire  _T_2804; // @[MemPrimitives.scala 123:41:@22559.4]
  wire  _T_2805; // @[MemPrimitives.scala 123:41:@22560.4]
  wire [10:0] _T_2807; // @[Cat.scala 30:58:@22562.4]
  wire [10:0] _T_2809; // @[Cat.scala 30:58:@22564.4]
  wire [10:0] _T_2811; // @[Cat.scala 30:58:@22566.4]
  wire [10:0] _T_2813; // @[Cat.scala 30:58:@22568.4]
  wire [10:0] _T_2815; // @[Cat.scala 30:58:@22570.4]
  wire [10:0] _T_2817; // @[Cat.scala 30:58:@22572.4]
  wire [10:0] _T_2819; // @[Cat.scala 30:58:@22574.4]
  wire [10:0] _T_2821; // @[Cat.scala 30:58:@22576.4]
  wire [10:0] _T_2823; // @[Cat.scala 30:58:@22578.4]
  wire [10:0] _T_2824; // @[Mux.scala 31:69:@22579.4]
  wire [10:0] _T_2825; // @[Mux.scala 31:69:@22580.4]
  wire [10:0] _T_2826; // @[Mux.scala 31:69:@22581.4]
  wire [10:0] _T_2827; // @[Mux.scala 31:69:@22582.4]
  wire [10:0] _T_2828; // @[Mux.scala 31:69:@22583.4]
  wire [10:0] _T_2829; // @[Mux.scala 31:69:@22584.4]
  wire [10:0] _T_2830; // @[Mux.scala 31:69:@22585.4]
  wire [10:0] _T_2831; // @[Mux.scala 31:69:@22586.4]
  wire  _T_2836; // @[MemPrimitives.scala 110:210:@22593.4]
  wire  _T_2839; // @[MemPrimitives.scala 110:228:@22595.4]
  wire  _T_2842; // @[MemPrimitives.scala 110:210:@22597.4]
  wire  _T_2845; // @[MemPrimitives.scala 110:228:@22599.4]
  wire  _T_2848; // @[MemPrimitives.scala 110:210:@22601.4]
  wire  _T_2851; // @[MemPrimitives.scala 110:228:@22603.4]
  wire  _T_2854; // @[MemPrimitives.scala 110:210:@22605.4]
  wire  _T_2857; // @[MemPrimitives.scala 110:228:@22607.4]
  wire  _T_2860; // @[MemPrimitives.scala 110:210:@22609.4]
  wire  _T_2863; // @[MemPrimitives.scala 110:228:@22611.4]
  wire  _T_2866; // @[MemPrimitives.scala 110:210:@22613.4]
  wire  _T_2869; // @[MemPrimitives.scala 110:228:@22615.4]
  wire  _T_2872; // @[MemPrimitives.scala 110:210:@22617.4]
  wire  _T_2875; // @[MemPrimitives.scala 110:228:@22619.4]
  wire  _T_2878; // @[MemPrimitives.scala 110:210:@22621.4]
  wire  _T_2881; // @[MemPrimitives.scala 110:228:@22623.4]
  wire  _T_2884; // @[MemPrimitives.scala 110:210:@22625.4]
  wire  _T_2887; // @[MemPrimitives.scala 110:228:@22627.4]
  wire  _T_2889; // @[MemPrimitives.scala 123:41:@22641.4]
  wire  _T_2890; // @[MemPrimitives.scala 123:41:@22642.4]
  wire  _T_2891; // @[MemPrimitives.scala 123:41:@22643.4]
  wire  _T_2892; // @[MemPrimitives.scala 123:41:@22644.4]
  wire  _T_2893; // @[MemPrimitives.scala 123:41:@22645.4]
  wire  _T_2894; // @[MemPrimitives.scala 123:41:@22646.4]
  wire  _T_2895; // @[MemPrimitives.scala 123:41:@22647.4]
  wire  _T_2896; // @[MemPrimitives.scala 123:41:@22648.4]
  wire  _T_2897; // @[MemPrimitives.scala 123:41:@22649.4]
  wire [10:0] _T_2899; // @[Cat.scala 30:58:@22651.4]
  wire [10:0] _T_2901; // @[Cat.scala 30:58:@22653.4]
  wire [10:0] _T_2903; // @[Cat.scala 30:58:@22655.4]
  wire [10:0] _T_2905; // @[Cat.scala 30:58:@22657.4]
  wire [10:0] _T_2907; // @[Cat.scala 30:58:@22659.4]
  wire [10:0] _T_2909; // @[Cat.scala 30:58:@22661.4]
  wire [10:0] _T_2911; // @[Cat.scala 30:58:@22663.4]
  wire [10:0] _T_2913; // @[Cat.scala 30:58:@22665.4]
  wire [10:0] _T_2915; // @[Cat.scala 30:58:@22667.4]
  wire [10:0] _T_2916; // @[Mux.scala 31:69:@22668.4]
  wire [10:0] _T_2917; // @[Mux.scala 31:69:@22669.4]
  wire [10:0] _T_2918; // @[Mux.scala 31:69:@22670.4]
  wire [10:0] _T_2919; // @[Mux.scala 31:69:@22671.4]
  wire [10:0] _T_2920; // @[Mux.scala 31:69:@22672.4]
  wire [10:0] _T_2921; // @[Mux.scala 31:69:@22673.4]
  wire [10:0] _T_2922; // @[Mux.scala 31:69:@22674.4]
  wire [10:0] _T_2923; // @[Mux.scala 31:69:@22675.4]
  wire  _T_2928; // @[MemPrimitives.scala 110:210:@22682.4]
  wire  _T_2931; // @[MemPrimitives.scala 110:228:@22684.4]
  wire  _T_2934; // @[MemPrimitives.scala 110:210:@22686.4]
  wire  _T_2937; // @[MemPrimitives.scala 110:228:@22688.4]
  wire  _T_2940; // @[MemPrimitives.scala 110:210:@22690.4]
  wire  _T_2943; // @[MemPrimitives.scala 110:228:@22692.4]
  wire  _T_2946; // @[MemPrimitives.scala 110:210:@22694.4]
  wire  _T_2949; // @[MemPrimitives.scala 110:228:@22696.4]
  wire  _T_2952; // @[MemPrimitives.scala 110:210:@22698.4]
  wire  _T_2955; // @[MemPrimitives.scala 110:228:@22700.4]
  wire  _T_2958; // @[MemPrimitives.scala 110:210:@22702.4]
  wire  _T_2961; // @[MemPrimitives.scala 110:228:@22704.4]
  wire  _T_2964; // @[MemPrimitives.scala 110:210:@22706.4]
  wire  _T_2967; // @[MemPrimitives.scala 110:228:@22708.4]
  wire  _T_2970; // @[MemPrimitives.scala 110:210:@22710.4]
  wire  _T_2973; // @[MemPrimitives.scala 110:228:@22712.4]
  wire  _T_2976; // @[MemPrimitives.scala 110:210:@22714.4]
  wire  _T_2979; // @[MemPrimitives.scala 110:228:@22716.4]
  wire  _T_2981; // @[MemPrimitives.scala 123:41:@22730.4]
  wire  _T_2982; // @[MemPrimitives.scala 123:41:@22731.4]
  wire  _T_2983; // @[MemPrimitives.scala 123:41:@22732.4]
  wire  _T_2984; // @[MemPrimitives.scala 123:41:@22733.4]
  wire  _T_2985; // @[MemPrimitives.scala 123:41:@22734.4]
  wire  _T_2986; // @[MemPrimitives.scala 123:41:@22735.4]
  wire  _T_2987; // @[MemPrimitives.scala 123:41:@22736.4]
  wire  _T_2988; // @[MemPrimitives.scala 123:41:@22737.4]
  wire  _T_2989; // @[MemPrimitives.scala 123:41:@22738.4]
  wire [10:0] _T_2991; // @[Cat.scala 30:58:@22740.4]
  wire [10:0] _T_2993; // @[Cat.scala 30:58:@22742.4]
  wire [10:0] _T_2995; // @[Cat.scala 30:58:@22744.4]
  wire [10:0] _T_2997; // @[Cat.scala 30:58:@22746.4]
  wire [10:0] _T_2999; // @[Cat.scala 30:58:@22748.4]
  wire [10:0] _T_3001; // @[Cat.scala 30:58:@22750.4]
  wire [10:0] _T_3003; // @[Cat.scala 30:58:@22752.4]
  wire [10:0] _T_3005; // @[Cat.scala 30:58:@22754.4]
  wire [10:0] _T_3007; // @[Cat.scala 30:58:@22756.4]
  wire [10:0] _T_3008; // @[Mux.scala 31:69:@22757.4]
  wire [10:0] _T_3009; // @[Mux.scala 31:69:@22758.4]
  wire [10:0] _T_3010; // @[Mux.scala 31:69:@22759.4]
  wire [10:0] _T_3011; // @[Mux.scala 31:69:@22760.4]
  wire [10:0] _T_3012; // @[Mux.scala 31:69:@22761.4]
  wire [10:0] _T_3013; // @[Mux.scala 31:69:@22762.4]
  wire [10:0] _T_3014; // @[Mux.scala 31:69:@22763.4]
  wire [10:0] _T_3015; // @[Mux.scala 31:69:@22764.4]
  wire  _T_3023; // @[MemPrimitives.scala 110:228:@22773.4]
  wire  _T_3029; // @[MemPrimitives.scala 110:228:@22777.4]
  wire  _T_3035; // @[MemPrimitives.scala 110:228:@22781.4]
  wire  _T_3041; // @[MemPrimitives.scala 110:228:@22785.4]
  wire  _T_3047; // @[MemPrimitives.scala 110:228:@22789.4]
  wire  _T_3053; // @[MemPrimitives.scala 110:228:@22793.4]
  wire  _T_3059; // @[MemPrimitives.scala 110:228:@22797.4]
  wire  _T_3065; // @[MemPrimitives.scala 110:228:@22801.4]
  wire  _T_3071; // @[MemPrimitives.scala 110:228:@22805.4]
  wire  _T_3073; // @[MemPrimitives.scala 123:41:@22819.4]
  wire  _T_3074; // @[MemPrimitives.scala 123:41:@22820.4]
  wire  _T_3075; // @[MemPrimitives.scala 123:41:@22821.4]
  wire  _T_3076; // @[MemPrimitives.scala 123:41:@22822.4]
  wire  _T_3077; // @[MemPrimitives.scala 123:41:@22823.4]
  wire  _T_3078; // @[MemPrimitives.scala 123:41:@22824.4]
  wire  _T_3079; // @[MemPrimitives.scala 123:41:@22825.4]
  wire  _T_3080; // @[MemPrimitives.scala 123:41:@22826.4]
  wire  _T_3081; // @[MemPrimitives.scala 123:41:@22827.4]
  wire [10:0] _T_3083; // @[Cat.scala 30:58:@22829.4]
  wire [10:0] _T_3085; // @[Cat.scala 30:58:@22831.4]
  wire [10:0] _T_3087; // @[Cat.scala 30:58:@22833.4]
  wire [10:0] _T_3089; // @[Cat.scala 30:58:@22835.4]
  wire [10:0] _T_3091; // @[Cat.scala 30:58:@22837.4]
  wire [10:0] _T_3093; // @[Cat.scala 30:58:@22839.4]
  wire [10:0] _T_3095; // @[Cat.scala 30:58:@22841.4]
  wire [10:0] _T_3097; // @[Cat.scala 30:58:@22843.4]
  wire [10:0] _T_3099; // @[Cat.scala 30:58:@22845.4]
  wire [10:0] _T_3100; // @[Mux.scala 31:69:@22846.4]
  wire [10:0] _T_3101; // @[Mux.scala 31:69:@22847.4]
  wire [10:0] _T_3102; // @[Mux.scala 31:69:@22848.4]
  wire [10:0] _T_3103; // @[Mux.scala 31:69:@22849.4]
  wire [10:0] _T_3104; // @[Mux.scala 31:69:@22850.4]
  wire [10:0] _T_3105; // @[Mux.scala 31:69:@22851.4]
  wire [10:0] _T_3106; // @[Mux.scala 31:69:@22852.4]
  wire [10:0] _T_3107; // @[Mux.scala 31:69:@22853.4]
  wire  _T_3115; // @[MemPrimitives.scala 110:228:@22862.4]
  wire  _T_3121; // @[MemPrimitives.scala 110:228:@22866.4]
  wire  _T_3127; // @[MemPrimitives.scala 110:228:@22870.4]
  wire  _T_3133; // @[MemPrimitives.scala 110:228:@22874.4]
  wire  _T_3139; // @[MemPrimitives.scala 110:228:@22878.4]
  wire  _T_3145; // @[MemPrimitives.scala 110:228:@22882.4]
  wire  _T_3151; // @[MemPrimitives.scala 110:228:@22886.4]
  wire  _T_3157; // @[MemPrimitives.scala 110:228:@22890.4]
  wire  _T_3163; // @[MemPrimitives.scala 110:228:@22894.4]
  wire  _T_3165; // @[MemPrimitives.scala 123:41:@22908.4]
  wire  _T_3166; // @[MemPrimitives.scala 123:41:@22909.4]
  wire  _T_3167; // @[MemPrimitives.scala 123:41:@22910.4]
  wire  _T_3168; // @[MemPrimitives.scala 123:41:@22911.4]
  wire  _T_3169; // @[MemPrimitives.scala 123:41:@22912.4]
  wire  _T_3170; // @[MemPrimitives.scala 123:41:@22913.4]
  wire  _T_3171; // @[MemPrimitives.scala 123:41:@22914.4]
  wire  _T_3172; // @[MemPrimitives.scala 123:41:@22915.4]
  wire  _T_3173; // @[MemPrimitives.scala 123:41:@22916.4]
  wire [10:0] _T_3175; // @[Cat.scala 30:58:@22918.4]
  wire [10:0] _T_3177; // @[Cat.scala 30:58:@22920.4]
  wire [10:0] _T_3179; // @[Cat.scala 30:58:@22922.4]
  wire [10:0] _T_3181; // @[Cat.scala 30:58:@22924.4]
  wire [10:0] _T_3183; // @[Cat.scala 30:58:@22926.4]
  wire [10:0] _T_3185; // @[Cat.scala 30:58:@22928.4]
  wire [10:0] _T_3187; // @[Cat.scala 30:58:@22930.4]
  wire [10:0] _T_3189; // @[Cat.scala 30:58:@22932.4]
  wire [10:0] _T_3191; // @[Cat.scala 30:58:@22934.4]
  wire [10:0] _T_3192; // @[Mux.scala 31:69:@22935.4]
  wire [10:0] _T_3193; // @[Mux.scala 31:69:@22936.4]
  wire [10:0] _T_3194; // @[Mux.scala 31:69:@22937.4]
  wire [10:0] _T_3195; // @[Mux.scala 31:69:@22938.4]
  wire [10:0] _T_3196; // @[Mux.scala 31:69:@22939.4]
  wire [10:0] _T_3197; // @[Mux.scala 31:69:@22940.4]
  wire [10:0] _T_3198; // @[Mux.scala 31:69:@22941.4]
  wire [10:0] _T_3199; // @[Mux.scala 31:69:@22942.4]
  wire  _T_3207; // @[MemPrimitives.scala 110:228:@22951.4]
  wire  _T_3213; // @[MemPrimitives.scala 110:228:@22955.4]
  wire  _T_3219; // @[MemPrimitives.scala 110:228:@22959.4]
  wire  _T_3225; // @[MemPrimitives.scala 110:228:@22963.4]
  wire  _T_3231; // @[MemPrimitives.scala 110:228:@22967.4]
  wire  _T_3237; // @[MemPrimitives.scala 110:228:@22971.4]
  wire  _T_3243; // @[MemPrimitives.scala 110:228:@22975.4]
  wire  _T_3249; // @[MemPrimitives.scala 110:228:@22979.4]
  wire  _T_3255; // @[MemPrimitives.scala 110:228:@22983.4]
  wire  _T_3257; // @[MemPrimitives.scala 123:41:@22997.4]
  wire  _T_3258; // @[MemPrimitives.scala 123:41:@22998.4]
  wire  _T_3259; // @[MemPrimitives.scala 123:41:@22999.4]
  wire  _T_3260; // @[MemPrimitives.scala 123:41:@23000.4]
  wire  _T_3261; // @[MemPrimitives.scala 123:41:@23001.4]
  wire  _T_3262; // @[MemPrimitives.scala 123:41:@23002.4]
  wire  _T_3263; // @[MemPrimitives.scala 123:41:@23003.4]
  wire  _T_3264; // @[MemPrimitives.scala 123:41:@23004.4]
  wire  _T_3265; // @[MemPrimitives.scala 123:41:@23005.4]
  wire [10:0] _T_3267; // @[Cat.scala 30:58:@23007.4]
  wire [10:0] _T_3269; // @[Cat.scala 30:58:@23009.4]
  wire [10:0] _T_3271; // @[Cat.scala 30:58:@23011.4]
  wire [10:0] _T_3273; // @[Cat.scala 30:58:@23013.4]
  wire [10:0] _T_3275; // @[Cat.scala 30:58:@23015.4]
  wire [10:0] _T_3277; // @[Cat.scala 30:58:@23017.4]
  wire [10:0] _T_3279; // @[Cat.scala 30:58:@23019.4]
  wire [10:0] _T_3281; // @[Cat.scala 30:58:@23021.4]
  wire [10:0] _T_3283; // @[Cat.scala 30:58:@23023.4]
  wire [10:0] _T_3284; // @[Mux.scala 31:69:@23024.4]
  wire [10:0] _T_3285; // @[Mux.scala 31:69:@23025.4]
  wire [10:0] _T_3286; // @[Mux.scala 31:69:@23026.4]
  wire [10:0] _T_3287; // @[Mux.scala 31:69:@23027.4]
  wire [10:0] _T_3288; // @[Mux.scala 31:69:@23028.4]
  wire [10:0] _T_3289; // @[Mux.scala 31:69:@23029.4]
  wire [10:0] _T_3290; // @[Mux.scala 31:69:@23030.4]
  wire [10:0] _T_3291; // @[Mux.scala 31:69:@23031.4]
  wire  _T_3299; // @[MemPrimitives.scala 110:228:@23040.4]
  wire  _T_3305; // @[MemPrimitives.scala 110:228:@23044.4]
  wire  _T_3311; // @[MemPrimitives.scala 110:228:@23048.4]
  wire  _T_3317; // @[MemPrimitives.scala 110:228:@23052.4]
  wire  _T_3323; // @[MemPrimitives.scala 110:228:@23056.4]
  wire  _T_3329; // @[MemPrimitives.scala 110:228:@23060.4]
  wire  _T_3335; // @[MemPrimitives.scala 110:228:@23064.4]
  wire  _T_3341; // @[MemPrimitives.scala 110:228:@23068.4]
  wire  _T_3347; // @[MemPrimitives.scala 110:228:@23072.4]
  wire  _T_3349; // @[MemPrimitives.scala 123:41:@23086.4]
  wire  _T_3350; // @[MemPrimitives.scala 123:41:@23087.4]
  wire  _T_3351; // @[MemPrimitives.scala 123:41:@23088.4]
  wire  _T_3352; // @[MemPrimitives.scala 123:41:@23089.4]
  wire  _T_3353; // @[MemPrimitives.scala 123:41:@23090.4]
  wire  _T_3354; // @[MemPrimitives.scala 123:41:@23091.4]
  wire  _T_3355; // @[MemPrimitives.scala 123:41:@23092.4]
  wire  _T_3356; // @[MemPrimitives.scala 123:41:@23093.4]
  wire  _T_3357; // @[MemPrimitives.scala 123:41:@23094.4]
  wire [10:0] _T_3359; // @[Cat.scala 30:58:@23096.4]
  wire [10:0] _T_3361; // @[Cat.scala 30:58:@23098.4]
  wire [10:0] _T_3363; // @[Cat.scala 30:58:@23100.4]
  wire [10:0] _T_3365; // @[Cat.scala 30:58:@23102.4]
  wire [10:0] _T_3367; // @[Cat.scala 30:58:@23104.4]
  wire [10:0] _T_3369; // @[Cat.scala 30:58:@23106.4]
  wire [10:0] _T_3371; // @[Cat.scala 30:58:@23108.4]
  wire [10:0] _T_3373; // @[Cat.scala 30:58:@23110.4]
  wire [10:0] _T_3375; // @[Cat.scala 30:58:@23112.4]
  wire [10:0] _T_3376; // @[Mux.scala 31:69:@23113.4]
  wire [10:0] _T_3377; // @[Mux.scala 31:69:@23114.4]
  wire [10:0] _T_3378; // @[Mux.scala 31:69:@23115.4]
  wire [10:0] _T_3379; // @[Mux.scala 31:69:@23116.4]
  wire [10:0] _T_3380; // @[Mux.scala 31:69:@23117.4]
  wire [10:0] _T_3381; // @[Mux.scala 31:69:@23118.4]
  wire [10:0] _T_3382; // @[Mux.scala 31:69:@23119.4]
  wire [10:0] _T_3383; // @[Mux.scala 31:69:@23120.4]
  wire  _T_3479; // @[package.scala 96:25:@23249.4 package.scala 96:25:@23250.4]
  wire [7:0] _T_3483; // @[Mux.scala 31:69:@23259.4]
  wire  _T_3476; // @[package.scala 96:25:@23241.4 package.scala 96:25:@23242.4]
  wire [7:0] _T_3484; // @[Mux.scala 31:69:@23260.4]
  wire  _T_3473; // @[package.scala 96:25:@23233.4 package.scala 96:25:@23234.4]
  wire [7:0] _T_3485; // @[Mux.scala 31:69:@23261.4]
  wire  _T_3470; // @[package.scala 96:25:@23225.4 package.scala 96:25:@23226.4]
  wire [7:0] _T_3486; // @[Mux.scala 31:69:@23262.4]
  wire  _T_3467; // @[package.scala 96:25:@23217.4 package.scala 96:25:@23218.4]
  wire [7:0] _T_3487; // @[Mux.scala 31:69:@23263.4]
  wire  _T_3464; // @[package.scala 96:25:@23209.4 package.scala 96:25:@23210.4]
  wire [7:0] _T_3488; // @[Mux.scala 31:69:@23264.4]
  wire  _T_3461; // @[package.scala 96:25:@23201.4 package.scala 96:25:@23202.4]
  wire [7:0] _T_3489; // @[Mux.scala 31:69:@23265.4]
  wire  _T_3458; // @[package.scala 96:25:@23193.4 package.scala 96:25:@23194.4]
  wire [7:0] _T_3490; // @[Mux.scala 31:69:@23266.4]
  wire  _T_3455; // @[package.scala 96:25:@23185.4 package.scala 96:25:@23186.4]
  wire [7:0] _T_3491; // @[Mux.scala 31:69:@23267.4]
  wire  _T_3452; // @[package.scala 96:25:@23177.4 package.scala 96:25:@23178.4]
  wire [7:0] _T_3492; // @[Mux.scala 31:69:@23268.4]
  wire  _T_3449; // @[package.scala 96:25:@23169.4 package.scala 96:25:@23170.4]
  wire  _T_3586; // @[package.scala 96:25:@23393.4 package.scala 96:25:@23394.4]
  wire [7:0] _T_3590; // @[Mux.scala 31:69:@23403.4]
  wire  _T_3583; // @[package.scala 96:25:@23385.4 package.scala 96:25:@23386.4]
  wire [7:0] _T_3591; // @[Mux.scala 31:69:@23404.4]
  wire  _T_3580; // @[package.scala 96:25:@23377.4 package.scala 96:25:@23378.4]
  wire [7:0] _T_3592; // @[Mux.scala 31:69:@23405.4]
  wire  _T_3577; // @[package.scala 96:25:@23369.4 package.scala 96:25:@23370.4]
  wire [7:0] _T_3593; // @[Mux.scala 31:69:@23406.4]
  wire  _T_3574; // @[package.scala 96:25:@23361.4 package.scala 96:25:@23362.4]
  wire [7:0] _T_3594; // @[Mux.scala 31:69:@23407.4]
  wire  _T_3571; // @[package.scala 96:25:@23353.4 package.scala 96:25:@23354.4]
  wire [7:0] _T_3595; // @[Mux.scala 31:69:@23408.4]
  wire  _T_3568; // @[package.scala 96:25:@23345.4 package.scala 96:25:@23346.4]
  wire [7:0] _T_3596; // @[Mux.scala 31:69:@23409.4]
  wire  _T_3565; // @[package.scala 96:25:@23337.4 package.scala 96:25:@23338.4]
  wire [7:0] _T_3597; // @[Mux.scala 31:69:@23410.4]
  wire  _T_3562; // @[package.scala 96:25:@23329.4 package.scala 96:25:@23330.4]
  wire [7:0] _T_3598; // @[Mux.scala 31:69:@23411.4]
  wire  _T_3559; // @[package.scala 96:25:@23321.4 package.scala 96:25:@23322.4]
  wire [7:0] _T_3599; // @[Mux.scala 31:69:@23412.4]
  wire  _T_3556; // @[package.scala 96:25:@23313.4 package.scala 96:25:@23314.4]
  wire  _T_3693; // @[package.scala 96:25:@23537.4 package.scala 96:25:@23538.4]
  wire [7:0] _T_3697; // @[Mux.scala 31:69:@23547.4]
  wire  _T_3690; // @[package.scala 96:25:@23529.4 package.scala 96:25:@23530.4]
  wire [7:0] _T_3698; // @[Mux.scala 31:69:@23548.4]
  wire  _T_3687; // @[package.scala 96:25:@23521.4 package.scala 96:25:@23522.4]
  wire [7:0] _T_3699; // @[Mux.scala 31:69:@23549.4]
  wire  _T_3684; // @[package.scala 96:25:@23513.4 package.scala 96:25:@23514.4]
  wire [7:0] _T_3700; // @[Mux.scala 31:69:@23550.4]
  wire  _T_3681; // @[package.scala 96:25:@23505.4 package.scala 96:25:@23506.4]
  wire [7:0] _T_3701; // @[Mux.scala 31:69:@23551.4]
  wire  _T_3678; // @[package.scala 96:25:@23497.4 package.scala 96:25:@23498.4]
  wire [7:0] _T_3702; // @[Mux.scala 31:69:@23552.4]
  wire  _T_3675; // @[package.scala 96:25:@23489.4 package.scala 96:25:@23490.4]
  wire [7:0] _T_3703; // @[Mux.scala 31:69:@23553.4]
  wire  _T_3672; // @[package.scala 96:25:@23481.4 package.scala 96:25:@23482.4]
  wire [7:0] _T_3704; // @[Mux.scala 31:69:@23554.4]
  wire  _T_3669; // @[package.scala 96:25:@23473.4 package.scala 96:25:@23474.4]
  wire [7:0] _T_3705; // @[Mux.scala 31:69:@23555.4]
  wire  _T_3666; // @[package.scala 96:25:@23465.4 package.scala 96:25:@23466.4]
  wire [7:0] _T_3706; // @[Mux.scala 31:69:@23556.4]
  wire  _T_3663; // @[package.scala 96:25:@23457.4 package.scala 96:25:@23458.4]
  wire  _T_3800; // @[package.scala 96:25:@23681.4 package.scala 96:25:@23682.4]
  wire [7:0] _T_3804; // @[Mux.scala 31:69:@23691.4]
  wire  _T_3797; // @[package.scala 96:25:@23673.4 package.scala 96:25:@23674.4]
  wire [7:0] _T_3805; // @[Mux.scala 31:69:@23692.4]
  wire  _T_3794; // @[package.scala 96:25:@23665.4 package.scala 96:25:@23666.4]
  wire [7:0] _T_3806; // @[Mux.scala 31:69:@23693.4]
  wire  _T_3791; // @[package.scala 96:25:@23657.4 package.scala 96:25:@23658.4]
  wire [7:0] _T_3807; // @[Mux.scala 31:69:@23694.4]
  wire  _T_3788; // @[package.scala 96:25:@23649.4 package.scala 96:25:@23650.4]
  wire [7:0] _T_3808; // @[Mux.scala 31:69:@23695.4]
  wire  _T_3785; // @[package.scala 96:25:@23641.4 package.scala 96:25:@23642.4]
  wire [7:0] _T_3809; // @[Mux.scala 31:69:@23696.4]
  wire  _T_3782; // @[package.scala 96:25:@23633.4 package.scala 96:25:@23634.4]
  wire [7:0] _T_3810; // @[Mux.scala 31:69:@23697.4]
  wire  _T_3779; // @[package.scala 96:25:@23625.4 package.scala 96:25:@23626.4]
  wire [7:0] _T_3811; // @[Mux.scala 31:69:@23698.4]
  wire  _T_3776; // @[package.scala 96:25:@23617.4 package.scala 96:25:@23618.4]
  wire [7:0] _T_3812; // @[Mux.scala 31:69:@23699.4]
  wire  _T_3773; // @[package.scala 96:25:@23609.4 package.scala 96:25:@23610.4]
  wire [7:0] _T_3813; // @[Mux.scala 31:69:@23700.4]
  wire  _T_3770; // @[package.scala 96:25:@23601.4 package.scala 96:25:@23602.4]
  wire  _T_3907; // @[package.scala 96:25:@23825.4 package.scala 96:25:@23826.4]
  wire [7:0] _T_3911; // @[Mux.scala 31:69:@23835.4]
  wire  _T_3904; // @[package.scala 96:25:@23817.4 package.scala 96:25:@23818.4]
  wire [7:0] _T_3912; // @[Mux.scala 31:69:@23836.4]
  wire  _T_3901; // @[package.scala 96:25:@23809.4 package.scala 96:25:@23810.4]
  wire [7:0] _T_3913; // @[Mux.scala 31:69:@23837.4]
  wire  _T_3898; // @[package.scala 96:25:@23801.4 package.scala 96:25:@23802.4]
  wire [7:0] _T_3914; // @[Mux.scala 31:69:@23838.4]
  wire  _T_3895; // @[package.scala 96:25:@23793.4 package.scala 96:25:@23794.4]
  wire [7:0] _T_3915; // @[Mux.scala 31:69:@23839.4]
  wire  _T_3892; // @[package.scala 96:25:@23785.4 package.scala 96:25:@23786.4]
  wire [7:0] _T_3916; // @[Mux.scala 31:69:@23840.4]
  wire  _T_3889; // @[package.scala 96:25:@23777.4 package.scala 96:25:@23778.4]
  wire [7:0] _T_3917; // @[Mux.scala 31:69:@23841.4]
  wire  _T_3886; // @[package.scala 96:25:@23769.4 package.scala 96:25:@23770.4]
  wire [7:0] _T_3918; // @[Mux.scala 31:69:@23842.4]
  wire  _T_3883; // @[package.scala 96:25:@23761.4 package.scala 96:25:@23762.4]
  wire [7:0] _T_3919; // @[Mux.scala 31:69:@23843.4]
  wire  _T_3880; // @[package.scala 96:25:@23753.4 package.scala 96:25:@23754.4]
  wire [7:0] _T_3920; // @[Mux.scala 31:69:@23844.4]
  wire  _T_3877; // @[package.scala 96:25:@23745.4 package.scala 96:25:@23746.4]
  wire  _T_4014; // @[package.scala 96:25:@23969.4 package.scala 96:25:@23970.4]
  wire [7:0] _T_4018; // @[Mux.scala 31:69:@23979.4]
  wire  _T_4011; // @[package.scala 96:25:@23961.4 package.scala 96:25:@23962.4]
  wire [7:0] _T_4019; // @[Mux.scala 31:69:@23980.4]
  wire  _T_4008; // @[package.scala 96:25:@23953.4 package.scala 96:25:@23954.4]
  wire [7:0] _T_4020; // @[Mux.scala 31:69:@23981.4]
  wire  _T_4005; // @[package.scala 96:25:@23945.4 package.scala 96:25:@23946.4]
  wire [7:0] _T_4021; // @[Mux.scala 31:69:@23982.4]
  wire  _T_4002; // @[package.scala 96:25:@23937.4 package.scala 96:25:@23938.4]
  wire [7:0] _T_4022; // @[Mux.scala 31:69:@23983.4]
  wire  _T_3999; // @[package.scala 96:25:@23929.4 package.scala 96:25:@23930.4]
  wire [7:0] _T_4023; // @[Mux.scala 31:69:@23984.4]
  wire  _T_3996; // @[package.scala 96:25:@23921.4 package.scala 96:25:@23922.4]
  wire [7:0] _T_4024; // @[Mux.scala 31:69:@23985.4]
  wire  _T_3993; // @[package.scala 96:25:@23913.4 package.scala 96:25:@23914.4]
  wire [7:0] _T_4025; // @[Mux.scala 31:69:@23986.4]
  wire  _T_3990; // @[package.scala 96:25:@23905.4 package.scala 96:25:@23906.4]
  wire [7:0] _T_4026; // @[Mux.scala 31:69:@23987.4]
  wire  _T_3987; // @[package.scala 96:25:@23897.4 package.scala 96:25:@23898.4]
  wire [7:0] _T_4027; // @[Mux.scala 31:69:@23988.4]
  wire  _T_3984; // @[package.scala 96:25:@23889.4 package.scala 96:25:@23890.4]
  wire  _T_4121; // @[package.scala 96:25:@24113.4 package.scala 96:25:@24114.4]
  wire [7:0] _T_4125; // @[Mux.scala 31:69:@24123.4]
  wire  _T_4118; // @[package.scala 96:25:@24105.4 package.scala 96:25:@24106.4]
  wire [7:0] _T_4126; // @[Mux.scala 31:69:@24124.4]
  wire  _T_4115; // @[package.scala 96:25:@24097.4 package.scala 96:25:@24098.4]
  wire [7:0] _T_4127; // @[Mux.scala 31:69:@24125.4]
  wire  _T_4112; // @[package.scala 96:25:@24089.4 package.scala 96:25:@24090.4]
  wire [7:0] _T_4128; // @[Mux.scala 31:69:@24126.4]
  wire  _T_4109; // @[package.scala 96:25:@24081.4 package.scala 96:25:@24082.4]
  wire [7:0] _T_4129; // @[Mux.scala 31:69:@24127.4]
  wire  _T_4106; // @[package.scala 96:25:@24073.4 package.scala 96:25:@24074.4]
  wire [7:0] _T_4130; // @[Mux.scala 31:69:@24128.4]
  wire  _T_4103; // @[package.scala 96:25:@24065.4 package.scala 96:25:@24066.4]
  wire [7:0] _T_4131; // @[Mux.scala 31:69:@24129.4]
  wire  _T_4100; // @[package.scala 96:25:@24057.4 package.scala 96:25:@24058.4]
  wire [7:0] _T_4132; // @[Mux.scala 31:69:@24130.4]
  wire  _T_4097; // @[package.scala 96:25:@24049.4 package.scala 96:25:@24050.4]
  wire [7:0] _T_4133; // @[Mux.scala 31:69:@24131.4]
  wire  _T_4094; // @[package.scala 96:25:@24041.4 package.scala 96:25:@24042.4]
  wire [7:0] _T_4134; // @[Mux.scala 31:69:@24132.4]
  wire  _T_4091; // @[package.scala 96:25:@24033.4 package.scala 96:25:@24034.4]
  wire  _T_4228; // @[package.scala 96:25:@24257.4 package.scala 96:25:@24258.4]
  wire [7:0] _T_4232; // @[Mux.scala 31:69:@24267.4]
  wire  _T_4225; // @[package.scala 96:25:@24249.4 package.scala 96:25:@24250.4]
  wire [7:0] _T_4233; // @[Mux.scala 31:69:@24268.4]
  wire  _T_4222; // @[package.scala 96:25:@24241.4 package.scala 96:25:@24242.4]
  wire [7:0] _T_4234; // @[Mux.scala 31:69:@24269.4]
  wire  _T_4219; // @[package.scala 96:25:@24233.4 package.scala 96:25:@24234.4]
  wire [7:0] _T_4235; // @[Mux.scala 31:69:@24270.4]
  wire  _T_4216; // @[package.scala 96:25:@24225.4 package.scala 96:25:@24226.4]
  wire [7:0] _T_4236; // @[Mux.scala 31:69:@24271.4]
  wire  _T_4213; // @[package.scala 96:25:@24217.4 package.scala 96:25:@24218.4]
  wire [7:0] _T_4237; // @[Mux.scala 31:69:@24272.4]
  wire  _T_4210; // @[package.scala 96:25:@24209.4 package.scala 96:25:@24210.4]
  wire [7:0] _T_4238; // @[Mux.scala 31:69:@24273.4]
  wire  _T_4207; // @[package.scala 96:25:@24201.4 package.scala 96:25:@24202.4]
  wire [7:0] _T_4239; // @[Mux.scala 31:69:@24274.4]
  wire  _T_4204; // @[package.scala 96:25:@24193.4 package.scala 96:25:@24194.4]
  wire [7:0] _T_4240; // @[Mux.scala 31:69:@24275.4]
  wire  _T_4201; // @[package.scala 96:25:@24185.4 package.scala 96:25:@24186.4]
  wire [7:0] _T_4241; // @[Mux.scala 31:69:@24276.4]
  wire  _T_4198; // @[package.scala 96:25:@24177.4 package.scala 96:25:@24178.4]
  wire  _T_4335; // @[package.scala 96:25:@24401.4 package.scala 96:25:@24402.4]
  wire [7:0] _T_4339; // @[Mux.scala 31:69:@24411.4]
  wire  _T_4332; // @[package.scala 96:25:@24393.4 package.scala 96:25:@24394.4]
  wire [7:0] _T_4340; // @[Mux.scala 31:69:@24412.4]
  wire  _T_4329; // @[package.scala 96:25:@24385.4 package.scala 96:25:@24386.4]
  wire [7:0] _T_4341; // @[Mux.scala 31:69:@24413.4]
  wire  _T_4326; // @[package.scala 96:25:@24377.4 package.scala 96:25:@24378.4]
  wire [7:0] _T_4342; // @[Mux.scala 31:69:@24414.4]
  wire  _T_4323; // @[package.scala 96:25:@24369.4 package.scala 96:25:@24370.4]
  wire [7:0] _T_4343; // @[Mux.scala 31:69:@24415.4]
  wire  _T_4320; // @[package.scala 96:25:@24361.4 package.scala 96:25:@24362.4]
  wire [7:0] _T_4344; // @[Mux.scala 31:69:@24416.4]
  wire  _T_4317; // @[package.scala 96:25:@24353.4 package.scala 96:25:@24354.4]
  wire [7:0] _T_4345; // @[Mux.scala 31:69:@24417.4]
  wire  _T_4314; // @[package.scala 96:25:@24345.4 package.scala 96:25:@24346.4]
  wire [7:0] _T_4346; // @[Mux.scala 31:69:@24418.4]
  wire  _T_4311; // @[package.scala 96:25:@24337.4 package.scala 96:25:@24338.4]
  wire [7:0] _T_4347; // @[Mux.scala 31:69:@24419.4]
  wire  _T_4308; // @[package.scala 96:25:@24329.4 package.scala 96:25:@24330.4]
  wire [7:0] _T_4348; // @[Mux.scala 31:69:@24420.4]
  wire  _T_4305; // @[package.scala 96:25:@24321.4 package.scala 96:25:@24322.4]
  wire  _T_4442; // @[package.scala 96:25:@24545.4 package.scala 96:25:@24546.4]
  wire [7:0] _T_4446; // @[Mux.scala 31:69:@24555.4]
  wire  _T_4439; // @[package.scala 96:25:@24537.4 package.scala 96:25:@24538.4]
  wire [7:0] _T_4447; // @[Mux.scala 31:69:@24556.4]
  wire  _T_4436; // @[package.scala 96:25:@24529.4 package.scala 96:25:@24530.4]
  wire [7:0] _T_4448; // @[Mux.scala 31:69:@24557.4]
  wire  _T_4433; // @[package.scala 96:25:@24521.4 package.scala 96:25:@24522.4]
  wire [7:0] _T_4449; // @[Mux.scala 31:69:@24558.4]
  wire  _T_4430; // @[package.scala 96:25:@24513.4 package.scala 96:25:@24514.4]
  wire [7:0] _T_4450; // @[Mux.scala 31:69:@24559.4]
  wire  _T_4427; // @[package.scala 96:25:@24505.4 package.scala 96:25:@24506.4]
  wire [7:0] _T_4451; // @[Mux.scala 31:69:@24560.4]
  wire  _T_4424; // @[package.scala 96:25:@24497.4 package.scala 96:25:@24498.4]
  wire [7:0] _T_4452; // @[Mux.scala 31:69:@24561.4]
  wire  _T_4421; // @[package.scala 96:25:@24489.4 package.scala 96:25:@24490.4]
  wire [7:0] _T_4453; // @[Mux.scala 31:69:@24562.4]
  wire  _T_4418; // @[package.scala 96:25:@24481.4 package.scala 96:25:@24482.4]
  wire [7:0] _T_4454; // @[Mux.scala 31:69:@24563.4]
  wire  _T_4415; // @[package.scala 96:25:@24473.4 package.scala 96:25:@24474.4]
  wire [7:0] _T_4455; // @[Mux.scala 31:69:@24564.4]
  wire  _T_4412; // @[package.scala 96:25:@24465.4 package.scala 96:25:@24466.4]
  wire  _T_4549; // @[package.scala 96:25:@24689.4 package.scala 96:25:@24690.4]
  wire [7:0] _T_4553; // @[Mux.scala 31:69:@24699.4]
  wire  _T_4546; // @[package.scala 96:25:@24681.4 package.scala 96:25:@24682.4]
  wire [7:0] _T_4554; // @[Mux.scala 31:69:@24700.4]
  wire  _T_4543; // @[package.scala 96:25:@24673.4 package.scala 96:25:@24674.4]
  wire [7:0] _T_4555; // @[Mux.scala 31:69:@24701.4]
  wire  _T_4540; // @[package.scala 96:25:@24665.4 package.scala 96:25:@24666.4]
  wire [7:0] _T_4556; // @[Mux.scala 31:69:@24702.4]
  wire  _T_4537; // @[package.scala 96:25:@24657.4 package.scala 96:25:@24658.4]
  wire [7:0] _T_4557; // @[Mux.scala 31:69:@24703.4]
  wire  _T_4534; // @[package.scala 96:25:@24649.4 package.scala 96:25:@24650.4]
  wire [7:0] _T_4558; // @[Mux.scala 31:69:@24704.4]
  wire  _T_4531; // @[package.scala 96:25:@24641.4 package.scala 96:25:@24642.4]
  wire [7:0] _T_4559; // @[Mux.scala 31:69:@24705.4]
  wire  _T_4528; // @[package.scala 96:25:@24633.4 package.scala 96:25:@24634.4]
  wire [7:0] _T_4560; // @[Mux.scala 31:69:@24706.4]
  wire  _T_4525; // @[package.scala 96:25:@24625.4 package.scala 96:25:@24626.4]
  wire [7:0] _T_4561; // @[Mux.scala 31:69:@24707.4]
  wire  _T_4522; // @[package.scala 96:25:@24617.4 package.scala 96:25:@24618.4]
  wire [7:0] _T_4562; // @[Mux.scala 31:69:@24708.4]
  wire  _T_4519; // @[package.scala 96:25:@24609.4 package.scala 96:25:@24610.4]
  wire  _T_4656; // @[package.scala 96:25:@24833.4 package.scala 96:25:@24834.4]
  wire [7:0] _T_4660; // @[Mux.scala 31:69:@24843.4]
  wire  _T_4653; // @[package.scala 96:25:@24825.4 package.scala 96:25:@24826.4]
  wire [7:0] _T_4661; // @[Mux.scala 31:69:@24844.4]
  wire  _T_4650; // @[package.scala 96:25:@24817.4 package.scala 96:25:@24818.4]
  wire [7:0] _T_4662; // @[Mux.scala 31:69:@24845.4]
  wire  _T_4647; // @[package.scala 96:25:@24809.4 package.scala 96:25:@24810.4]
  wire [7:0] _T_4663; // @[Mux.scala 31:69:@24846.4]
  wire  _T_4644; // @[package.scala 96:25:@24801.4 package.scala 96:25:@24802.4]
  wire [7:0] _T_4664; // @[Mux.scala 31:69:@24847.4]
  wire  _T_4641; // @[package.scala 96:25:@24793.4 package.scala 96:25:@24794.4]
  wire [7:0] _T_4665; // @[Mux.scala 31:69:@24848.4]
  wire  _T_4638; // @[package.scala 96:25:@24785.4 package.scala 96:25:@24786.4]
  wire [7:0] _T_4666; // @[Mux.scala 31:69:@24849.4]
  wire  _T_4635; // @[package.scala 96:25:@24777.4 package.scala 96:25:@24778.4]
  wire [7:0] _T_4667; // @[Mux.scala 31:69:@24850.4]
  wire  _T_4632; // @[package.scala 96:25:@24769.4 package.scala 96:25:@24770.4]
  wire [7:0] _T_4668; // @[Mux.scala 31:69:@24851.4]
  wire  _T_4629; // @[package.scala 96:25:@24761.4 package.scala 96:25:@24762.4]
  wire [7:0] _T_4669; // @[Mux.scala 31:69:@24852.4]
  wire  _T_4626; // @[package.scala 96:25:@24753.4 package.scala 96:25:@24754.4]
  wire  _T_4763; // @[package.scala 96:25:@24977.4 package.scala 96:25:@24978.4]
  wire [7:0] _T_4767; // @[Mux.scala 31:69:@24987.4]
  wire  _T_4760; // @[package.scala 96:25:@24969.4 package.scala 96:25:@24970.4]
  wire [7:0] _T_4768; // @[Mux.scala 31:69:@24988.4]
  wire  _T_4757; // @[package.scala 96:25:@24961.4 package.scala 96:25:@24962.4]
  wire [7:0] _T_4769; // @[Mux.scala 31:69:@24989.4]
  wire  _T_4754; // @[package.scala 96:25:@24953.4 package.scala 96:25:@24954.4]
  wire [7:0] _T_4770; // @[Mux.scala 31:69:@24990.4]
  wire  _T_4751; // @[package.scala 96:25:@24945.4 package.scala 96:25:@24946.4]
  wire [7:0] _T_4771; // @[Mux.scala 31:69:@24991.4]
  wire  _T_4748; // @[package.scala 96:25:@24937.4 package.scala 96:25:@24938.4]
  wire [7:0] _T_4772; // @[Mux.scala 31:69:@24992.4]
  wire  _T_4745; // @[package.scala 96:25:@24929.4 package.scala 96:25:@24930.4]
  wire [7:0] _T_4773; // @[Mux.scala 31:69:@24993.4]
  wire  _T_4742; // @[package.scala 96:25:@24921.4 package.scala 96:25:@24922.4]
  wire [7:0] _T_4774; // @[Mux.scala 31:69:@24994.4]
  wire  _T_4739; // @[package.scala 96:25:@24913.4 package.scala 96:25:@24914.4]
  wire [7:0] _T_4775; // @[Mux.scala 31:69:@24995.4]
  wire  _T_4736; // @[package.scala 96:25:@24905.4 package.scala 96:25:@24906.4]
  wire [7:0] _T_4776; // @[Mux.scala 31:69:@24996.4]
  wire  _T_4733; // @[package.scala 96:25:@24897.4 package.scala 96:25:@24898.4]
  wire  _T_4870; // @[package.scala 96:25:@25121.4 package.scala 96:25:@25122.4]
  wire [7:0] _T_4874; // @[Mux.scala 31:69:@25131.4]
  wire  _T_4867; // @[package.scala 96:25:@25113.4 package.scala 96:25:@25114.4]
  wire [7:0] _T_4875; // @[Mux.scala 31:69:@25132.4]
  wire  _T_4864; // @[package.scala 96:25:@25105.4 package.scala 96:25:@25106.4]
  wire [7:0] _T_4876; // @[Mux.scala 31:69:@25133.4]
  wire  _T_4861; // @[package.scala 96:25:@25097.4 package.scala 96:25:@25098.4]
  wire [7:0] _T_4877; // @[Mux.scala 31:69:@25134.4]
  wire  _T_4858; // @[package.scala 96:25:@25089.4 package.scala 96:25:@25090.4]
  wire [7:0] _T_4878; // @[Mux.scala 31:69:@25135.4]
  wire  _T_4855; // @[package.scala 96:25:@25081.4 package.scala 96:25:@25082.4]
  wire [7:0] _T_4879; // @[Mux.scala 31:69:@25136.4]
  wire  _T_4852; // @[package.scala 96:25:@25073.4 package.scala 96:25:@25074.4]
  wire [7:0] _T_4880; // @[Mux.scala 31:69:@25137.4]
  wire  _T_4849; // @[package.scala 96:25:@25065.4 package.scala 96:25:@25066.4]
  wire [7:0] _T_4881; // @[Mux.scala 31:69:@25138.4]
  wire  _T_4846; // @[package.scala 96:25:@25057.4 package.scala 96:25:@25058.4]
  wire [7:0] _T_4882; // @[Mux.scala 31:69:@25139.4]
  wire  _T_4843; // @[package.scala 96:25:@25049.4 package.scala 96:25:@25050.4]
  wire [7:0] _T_4883; // @[Mux.scala 31:69:@25140.4]
  wire  _T_4840; // @[package.scala 96:25:@25041.4 package.scala 96:25:@25042.4]
  wire  _T_4977; // @[package.scala 96:25:@25265.4 package.scala 96:25:@25266.4]
  wire [7:0] _T_4981; // @[Mux.scala 31:69:@25275.4]
  wire  _T_4974; // @[package.scala 96:25:@25257.4 package.scala 96:25:@25258.4]
  wire [7:0] _T_4982; // @[Mux.scala 31:69:@25276.4]
  wire  _T_4971; // @[package.scala 96:25:@25249.4 package.scala 96:25:@25250.4]
  wire [7:0] _T_4983; // @[Mux.scala 31:69:@25277.4]
  wire  _T_4968; // @[package.scala 96:25:@25241.4 package.scala 96:25:@25242.4]
  wire [7:0] _T_4984; // @[Mux.scala 31:69:@25278.4]
  wire  _T_4965; // @[package.scala 96:25:@25233.4 package.scala 96:25:@25234.4]
  wire [7:0] _T_4985; // @[Mux.scala 31:69:@25279.4]
  wire  _T_4962; // @[package.scala 96:25:@25225.4 package.scala 96:25:@25226.4]
  wire [7:0] _T_4986; // @[Mux.scala 31:69:@25280.4]
  wire  _T_4959; // @[package.scala 96:25:@25217.4 package.scala 96:25:@25218.4]
  wire [7:0] _T_4987; // @[Mux.scala 31:69:@25281.4]
  wire  _T_4956; // @[package.scala 96:25:@25209.4 package.scala 96:25:@25210.4]
  wire [7:0] _T_4988; // @[Mux.scala 31:69:@25282.4]
  wire  _T_4953; // @[package.scala 96:25:@25201.4 package.scala 96:25:@25202.4]
  wire [7:0] _T_4989; // @[Mux.scala 31:69:@25283.4]
  wire  _T_4950; // @[package.scala 96:25:@25193.4 package.scala 96:25:@25194.4]
  wire [7:0] _T_4990; // @[Mux.scala 31:69:@25284.4]
  wire  _T_4947; // @[package.scala 96:25:@25185.4 package.scala 96:25:@25186.4]
  wire  _T_5084; // @[package.scala 96:25:@25409.4 package.scala 96:25:@25410.4]
  wire [7:0] _T_5088; // @[Mux.scala 31:69:@25419.4]
  wire  _T_5081; // @[package.scala 96:25:@25401.4 package.scala 96:25:@25402.4]
  wire [7:0] _T_5089; // @[Mux.scala 31:69:@25420.4]
  wire  _T_5078; // @[package.scala 96:25:@25393.4 package.scala 96:25:@25394.4]
  wire [7:0] _T_5090; // @[Mux.scala 31:69:@25421.4]
  wire  _T_5075; // @[package.scala 96:25:@25385.4 package.scala 96:25:@25386.4]
  wire [7:0] _T_5091; // @[Mux.scala 31:69:@25422.4]
  wire  _T_5072; // @[package.scala 96:25:@25377.4 package.scala 96:25:@25378.4]
  wire [7:0] _T_5092; // @[Mux.scala 31:69:@25423.4]
  wire  _T_5069; // @[package.scala 96:25:@25369.4 package.scala 96:25:@25370.4]
  wire [7:0] _T_5093; // @[Mux.scala 31:69:@25424.4]
  wire  _T_5066; // @[package.scala 96:25:@25361.4 package.scala 96:25:@25362.4]
  wire [7:0] _T_5094; // @[Mux.scala 31:69:@25425.4]
  wire  _T_5063; // @[package.scala 96:25:@25353.4 package.scala 96:25:@25354.4]
  wire [7:0] _T_5095; // @[Mux.scala 31:69:@25426.4]
  wire  _T_5060; // @[package.scala 96:25:@25345.4 package.scala 96:25:@25346.4]
  wire [7:0] _T_5096; // @[Mux.scala 31:69:@25427.4]
  wire  _T_5057; // @[package.scala 96:25:@25337.4 package.scala 96:25:@25338.4]
  wire [7:0] _T_5097; // @[Mux.scala 31:69:@25428.4]
  wire  _T_5054; // @[package.scala 96:25:@25329.4 package.scala 96:25:@25330.4]
  wire  _T_5191; // @[package.scala 96:25:@25553.4 package.scala 96:25:@25554.4]
  wire [7:0] _T_5195; // @[Mux.scala 31:69:@25563.4]
  wire  _T_5188; // @[package.scala 96:25:@25545.4 package.scala 96:25:@25546.4]
  wire [7:0] _T_5196; // @[Mux.scala 31:69:@25564.4]
  wire  _T_5185; // @[package.scala 96:25:@25537.4 package.scala 96:25:@25538.4]
  wire [7:0] _T_5197; // @[Mux.scala 31:69:@25565.4]
  wire  _T_5182; // @[package.scala 96:25:@25529.4 package.scala 96:25:@25530.4]
  wire [7:0] _T_5198; // @[Mux.scala 31:69:@25566.4]
  wire  _T_5179; // @[package.scala 96:25:@25521.4 package.scala 96:25:@25522.4]
  wire [7:0] _T_5199; // @[Mux.scala 31:69:@25567.4]
  wire  _T_5176; // @[package.scala 96:25:@25513.4 package.scala 96:25:@25514.4]
  wire [7:0] _T_5200; // @[Mux.scala 31:69:@25568.4]
  wire  _T_5173; // @[package.scala 96:25:@25505.4 package.scala 96:25:@25506.4]
  wire [7:0] _T_5201; // @[Mux.scala 31:69:@25569.4]
  wire  _T_5170; // @[package.scala 96:25:@25497.4 package.scala 96:25:@25498.4]
  wire [7:0] _T_5202; // @[Mux.scala 31:69:@25570.4]
  wire  _T_5167; // @[package.scala 96:25:@25489.4 package.scala 96:25:@25490.4]
  wire [7:0] _T_5203; // @[Mux.scala 31:69:@25571.4]
  wire  _T_5164; // @[package.scala 96:25:@25481.4 package.scala 96:25:@25482.4]
  wire [7:0] _T_5204; // @[Mux.scala 31:69:@25572.4]
  wire  _T_5161; // @[package.scala 96:25:@25473.4 package.scala 96:25:@25474.4]
  wire  _T_5298; // @[package.scala 96:25:@25697.4 package.scala 96:25:@25698.4]
  wire [7:0] _T_5302; // @[Mux.scala 31:69:@25707.4]
  wire  _T_5295; // @[package.scala 96:25:@25689.4 package.scala 96:25:@25690.4]
  wire [7:0] _T_5303; // @[Mux.scala 31:69:@25708.4]
  wire  _T_5292; // @[package.scala 96:25:@25681.4 package.scala 96:25:@25682.4]
  wire [7:0] _T_5304; // @[Mux.scala 31:69:@25709.4]
  wire  _T_5289; // @[package.scala 96:25:@25673.4 package.scala 96:25:@25674.4]
  wire [7:0] _T_5305; // @[Mux.scala 31:69:@25710.4]
  wire  _T_5286; // @[package.scala 96:25:@25665.4 package.scala 96:25:@25666.4]
  wire [7:0] _T_5306; // @[Mux.scala 31:69:@25711.4]
  wire  _T_5283; // @[package.scala 96:25:@25657.4 package.scala 96:25:@25658.4]
  wire [7:0] _T_5307; // @[Mux.scala 31:69:@25712.4]
  wire  _T_5280; // @[package.scala 96:25:@25649.4 package.scala 96:25:@25650.4]
  wire [7:0] _T_5308; // @[Mux.scala 31:69:@25713.4]
  wire  _T_5277; // @[package.scala 96:25:@25641.4 package.scala 96:25:@25642.4]
  wire [7:0] _T_5309; // @[Mux.scala 31:69:@25714.4]
  wire  _T_5274; // @[package.scala 96:25:@25633.4 package.scala 96:25:@25634.4]
  wire [7:0] _T_5310; // @[Mux.scala 31:69:@25715.4]
  wire  _T_5271; // @[package.scala 96:25:@25625.4 package.scala 96:25:@25626.4]
  wire [7:0] _T_5311; // @[Mux.scala 31:69:@25716.4]
  wire  _T_5268; // @[package.scala 96:25:@25617.4 package.scala 96:25:@25618.4]
  Mem1D_5 Mem1D ( // @[MemPrimitives.scala 64:21:@20151.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  Mem1D_5 Mem1D_1 ( // @[MemPrimitives.scala 64:21:@20167.4]
    .clock(Mem1D_1_clock),
    .reset(Mem1D_1_reset),
    .io_r_ofs_0(Mem1D_1_io_r_ofs_0),
    .io_r_backpressure(Mem1D_1_io_r_backpressure),
    .io_w_ofs_0(Mem1D_1_io_w_ofs_0),
    .io_w_data_0(Mem1D_1_io_w_data_0),
    .io_w_en_0(Mem1D_1_io_w_en_0),
    .io_output(Mem1D_1_io_output)
  );
  Mem1D_5 Mem1D_2 ( // @[MemPrimitives.scala 64:21:@20183.4]
    .clock(Mem1D_2_clock),
    .reset(Mem1D_2_reset),
    .io_r_ofs_0(Mem1D_2_io_r_ofs_0),
    .io_r_backpressure(Mem1D_2_io_r_backpressure),
    .io_w_ofs_0(Mem1D_2_io_w_ofs_0),
    .io_w_data_0(Mem1D_2_io_w_data_0),
    .io_w_en_0(Mem1D_2_io_w_en_0),
    .io_output(Mem1D_2_io_output)
  );
  Mem1D_5 Mem1D_3 ( // @[MemPrimitives.scala 64:21:@20199.4]
    .clock(Mem1D_3_clock),
    .reset(Mem1D_3_reset),
    .io_r_ofs_0(Mem1D_3_io_r_ofs_0),
    .io_r_backpressure(Mem1D_3_io_r_backpressure),
    .io_w_ofs_0(Mem1D_3_io_w_ofs_0),
    .io_w_data_0(Mem1D_3_io_w_data_0),
    .io_w_en_0(Mem1D_3_io_w_en_0),
    .io_output(Mem1D_3_io_output)
  );
  Mem1D_5 Mem1D_4 ( // @[MemPrimitives.scala 64:21:@20215.4]
    .clock(Mem1D_4_clock),
    .reset(Mem1D_4_reset),
    .io_r_ofs_0(Mem1D_4_io_r_ofs_0),
    .io_r_backpressure(Mem1D_4_io_r_backpressure),
    .io_w_ofs_0(Mem1D_4_io_w_ofs_0),
    .io_w_data_0(Mem1D_4_io_w_data_0),
    .io_w_en_0(Mem1D_4_io_w_en_0),
    .io_output(Mem1D_4_io_output)
  );
  Mem1D_5 Mem1D_5 ( // @[MemPrimitives.scala 64:21:@20231.4]
    .clock(Mem1D_5_clock),
    .reset(Mem1D_5_reset),
    .io_r_ofs_0(Mem1D_5_io_r_ofs_0),
    .io_r_backpressure(Mem1D_5_io_r_backpressure),
    .io_w_ofs_0(Mem1D_5_io_w_ofs_0),
    .io_w_data_0(Mem1D_5_io_w_data_0),
    .io_w_en_0(Mem1D_5_io_w_en_0),
    .io_output(Mem1D_5_io_output)
  );
  Mem1D_5 Mem1D_6 ( // @[MemPrimitives.scala 64:21:@20247.4]
    .clock(Mem1D_6_clock),
    .reset(Mem1D_6_reset),
    .io_r_ofs_0(Mem1D_6_io_r_ofs_0),
    .io_r_backpressure(Mem1D_6_io_r_backpressure),
    .io_w_ofs_0(Mem1D_6_io_w_ofs_0),
    .io_w_data_0(Mem1D_6_io_w_data_0),
    .io_w_en_0(Mem1D_6_io_w_en_0),
    .io_output(Mem1D_6_io_output)
  );
  Mem1D_5 Mem1D_7 ( // @[MemPrimitives.scala 64:21:@20263.4]
    .clock(Mem1D_7_clock),
    .reset(Mem1D_7_reset),
    .io_r_ofs_0(Mem1D_7_io_r_ofs_0),
    .io_r_backpressure(Mem1D_7_io_r_backpressure),
    .io_w_ofs_0(Mem1D_7_io_w_ofs_0),
    .io_w_data_0(Mem1D_7_io_w_data_0),
    .io_w_en_0(Mem1D_7_io_w_en_0),
    .io_output(Mem1D_7_io_output)
  );
  Mem1D_5 Mem1D_8 ( // @[MemPrimitives.scala 64:21:@20279.4]
    .clock(Mem1D_8_clock),
    .reset(Mem1D_8_reset),
    .io_r_ofs_0(Mem1D_8_io_r_ofs_0),
    .io_r_backpressure(Mem1D_8_io_r_backpressure),
    .io_w_ofs_0(Mem1D_8_io_w_ofs_0),
    .io_w_data_0(Mem1D_8_io_w_data_0),
    .io_w_en_0(Mem1D_8_io_w_en_0),
    .io_output(Mem1D_8_io_output)
  );
  Mem1D_5 Mem1D_9 ( // @[MemPrimitives.scala 64:21:@20295.4]
    .clock(Mem1D_9_clock),
    .reset(Mem1D_9_reset),
    .io_r_ofs_0(Mem1D_9_io_r_ofs_0),
    .io_r_backpressure(Mem1D_9_io_r_backpressure),
    .io_w_ofs_0(Mem1D_9_io_w_ofs_0),
    .io_w_data_0(Mem1D_9_io_w_data_0),
    .io_w_en_0(Mem1D_9_io_w_en_0),
    .io_output(Mem1D_9_io_output)
  );
  Mem1D_5 Mem1D_10 ( // @[MemPrimitives.scala 64:21:@20311.4]
    .clock(Mem1D_10_clock),
    .reset(Mem1D_10_reset),
    .io_r_ofs_0(Mem1D_10_io_r_ofs_0),
    .io_r_backpressure(Mem1D_10_io_r_backpressure),
    .io_w_ofs_0(Mem1D_10_io_w_ofs_0),
    .io_w_data_0(Mem1D_10_io_w_data_0),
    .io_w_en_0(Mem1D_10_io_w_en_0),
    .io_output(Mem1D_10_io_output)
  );
  Mem1D_5 Mem1D_11 ( // @[MemPrimitives.scala 64:21:@20327.4]
    .clock(Mem1D_11_clock),
    .reset(Mem1D_11_reset),
    .io_r_ofs_0(Mem1D_11_io_r_ofs_0),
    .io_r_backpressure(Mem1D_11_io_r_backpressure),
    .io_w_ofs_0(Mem1D_11_io_w_ofs_0),
    .io_w_data_0(Mem1D_11_io_w_data_0),
    .io_w_en_0(Mem1D_11_io_w_en_0),
    .io_output(Mem1D_11_io_output)
  );
  Mem1D_5 Mem1D_12 ( // @[MemPrimitives.scala 64:21:@20343.4]
    .clock(Mem1D_12_clock),
    .reset(Mem1D_12_reset),
    .io_r_ofs_0(Mem1D_12_io_r_ofs_0),
    .io_r_backpressure(Mem1D_12_io_r_backpressure),
    .io_w_ofs_0(Mem1D_12_io_w_ofs_0),
    .io_w_data_0(Mem1D_12_io_w_data_0),
    .io_w_en_0(Mem1D_12_io_w_en_0),
    .io_output(Mem1D_12_io_output)
  );
  Mem1D_5 Mem1D_13 ( // @[MemPrimitives.scala 64:21:@20359.4]
    .clock(Mem1D_13_clock),
    .reset(Mem1D_13_reset),
    .io_r_ofs_0(Mem1D_13_io_r_ofs_0),
    .io_r_backpressure(Mem1D_13_io_r_backpressure),
    .io_w_ofs_0(Mem1D_13_io_w_ofs_0),
    .io_w_data_0(Mem1D_13_io_w_data_0),
    .io_w_en_0(Mem1D_13_io_w_en_0),
    .io_output(Mem1D_13_io_output)
  );
  Mem1D_5 Mem1D_14 ( // @[MemPrimitives.scala 64:21:@20375.4]
    .clock(Mem1D_14_clock),
    .reset(Mem1D_14_reset),
    .io_r_ofs_0(Mem1D_14_io_r_ofs_0),
    .io_r_backpressure(Mem1D_14_io_r_backpressure),
    .io_w_ofs_0(Mem1D_14_io_w_ofs_0),
    .io_w_data_0(Mem1D_14_io_w_data_0),
    .io_w_en_0(Mem1D_14_io_w_en_0),
    .io_output(Mem1D_14_io_output)
  );
  Mem1D_5 Mem1D_15 ( // @[MemPrimitives.scala 64:21:@20391.4]
    .clock(Mem1D_15_clock),
    .reset(Mem1D_15_reset),
    .io_r_ofs_0(Mem1D_15_io_r_ofs_0),
    .io_r_backpressure(Mem1D_15_io_r_backpressure),
    .io_w_ofs_0(Mem1D_15_io_w_ofs_0),
    .io_w_data_0(Mem1D_15_io_w_data_0),
    .io_w_en_0(Mem1D_15_io_w_en_0),
    .io_output(Mem1D_15_io_output)
  );
  Mem1D_5 Mem1D_16 ( // @[MemPrimitives.scala 64:21:@20407.4]
    .clock(Mem1D_16_clock),
    .reset(Mem1D_16_reset),
    .io_r_ofs_0(Mem1D_16_io_r_ofs_0),
    .io_r_backpressure(Mem1D_16_io_r_backpressure),
    .io_w_ofs_0(Mem1D_16_io_w_ofs_0),
    .io_w_data_0(Mem1D_16_io_w_data_0),
    .io_w_en_0(Mem1D_16_io_w_en_0),
    .io_output(Mem1D_16_io_output)
  );
  Mem1D_5 Mem1D_17 ( // @[MemPrimitives.scala 64:21:@20423.4]
    .clock(Mem1D_17_clock),
    .reset(Mem1D_17_reset),
    .io_r_ofs_0(Mem1D_17_io_r_ofs_0),
    .io_r_backpressure(Mem1D_17_io_r_backpressure),
    .io_w_ofs_0(Mem1D_17_io_w_ofs_0),
    .io_w_data_0(Mem1D_17_io_w_data_0),
    .io_w_en_0(Mem1D_17_io_w_en_0),
    .io_output(Mem1D_17_io_output)
  );
  Mem1D_5 Mem1D_18 ( // @[MemPrimitives.scala 64:21:@20439.4]
    .clock(Mem1D_18_clock),
    .reset(Mem1D_18_reset),
    .io_r_ofs_0(Mem1D_18_io_r_ofs_0),
    .io_r_backpressure(Mem1D_18_io_r_backpressure),
    .io_w_ofs_0(Mem1D_18_io_w_ofs_0),
    .io_w_data_0(Mem1D_18_io_w_data_0),
    .io_w_en_0(Mem1D_18_io_w_en_0),
    .io_output(Mem1D_18_io_output)
  );
  Mem1D_5 Mem1D_19 ( // @[MemPrimitives.scala 64:21:@20455.4]
    .clock(Mem1D_19_clock),
    .reset(Mem1D_19_reset),
    .io_r_ofs_0(Mem1D_19_io_r_ofs_0),
    .io_r_backpressure(Mem1D_19_io_r_backpressure),
    .io_w_ofs_0(Mem1D_19_io_w_ofs_0),
    .io_w_data_0(Mem1D_19_io_w_data_0),
    .io_w_en_0(Mem1D_19_io_w_en_0),
    .io_output(Mem1D_19_io_output)
  );
  Mem1D_5 Mem1D_20 ( // @[MemPrimitives.scala 64:21:@20471.4]
    .clock(Mem1D_20_clock),
    .reset(Mem1D_20_reset),
    .io_r_ofs_0(Mem1D_20_io_r_ofs_0),
    .io_r_backpressure(Mem1D_20_io_r_backpressure),
    .io_w_ofs_0(Mem1D_20_io_w_ofs_0),
    .io_w_data_0(Mem1D_20_io_w_data_0),
    .io_w_en_0(Mem1D_20_io_w_en_0),
    .io_output(Mem1D_20_io_output)
  );
  Mem1D_5 Mem1D_21 ( // @[MemPrimitives.scala 64:21:@20487.4]
    .clock(Mem1D_21_clock),
    .reset(Mem1D_21_reset),
    .io_r_ofs_0(Mem1D_21_io_r_ofs_0),
    .io_r_backpressure(Mem1D_21_io_r_backpressure),
    .io_w_ofs_0(Mem1D_21_io_w_ofs_0),
    .io_w_data_0(Mem1D_21_io_w_data_0),
    .io_w_en_0(Mem1D_21_io_w_en_0),
    .io_output(Mem1D_21_io_output)
  );
  Mem1D_5 Mem1D_22 ( // @[MemPrimitives.scala 64:21:@20503.4]
    .clock(Mem1D_22_clock),
    .reset(Mem1D_22_reset),
    .io_r_ofs_0(Mem1D_22_io_r_ofs_0),
    .io_r_backpressure(Mem1D_22_io_r_backpressure),
    .io_w_ofs_0(Mem1D_22_io_w_ofs_0),
    .io_w_data_0(Mem1D_22_io_w_data_0),
    .io_w_en_0(Mem1D_22_io_w_en_0),
    .io_output(Mem1D_22_io_output)
  );
  Mem1D_5 Mem1D_23 ( // @[MemPrimitives.scala 64:21:@20519.4]
    .clock(Mem1D_23_clock),
    .reset(Mem1D_23_reset),
    .io_r_ofs_0(Mem1D_23_io_r_ofs_0),
    .io_r_backpressure(Mem1D_23_io_r_backpressure),
    .io_w_ofs_0(Mem1D_23_io_w_ofs_0),
    .io_w_data_0(Mem1D_23_io_w_data_0),
    .io_w_en_0(Mem1D_23_io_w_en_0),
    .io_output(Mem1D_23_io_output)
  );
  StickySelects_1 StickySelects ( // @[MemPrimitives.scala 121:29:@21027.4]
    .clock(StickySelects_clock),
    .reset(StickySelects_reset),
    .io_ins_0(StickySelects_io_ins_0),
    .io_ins_1(StickySelects_io_ins_1),
    .io_ins_2(StickySelects_io_ins_2),
    .io_ins_3(StickySelects_io_ins_3),
    .io_ins_4(StickySelects_io_ins_4),
    .io_ins_5(StickySelects_io_ins_5),
    .io_ins_6(StickySelects_io_ins_6),
    .io_ins_7(StickySelects_io_ins_7),
    .io_ins_8(StickySelects_io_ins_8),
    .io_outs_0(StickySelects_io_outs_0),
    .io_outs_1(StickySelects_io_outs_1),
    .io_outs_2(StickySelects_io_outs_2),
    .io_outs_3(StickySelects_io_outs_3),
    .io_outs_4(StickySelects_io_outs_4),
    .io_outs_5(StickySelects_io_outs_5),
    .io_outs_6(StickySelects_io_outs_6),
    .io_outs_7(StickySelects_io_outs_7),
    .io_outs_8(StickySelects_io_outs_8)
  );
  StickySelects_1 StickySelects_1 ( // @[MemPrimitives.scala 121:29:@21116.4]
    .clock(StickySelects_1_clock),
    .reset(StickySelects_1_reset),
    .io_ins_0(StickySelects_1_io_ins_0),
    .io_ins_1(StickySelects_1_io_ins_1),
    .io_ins_2(StickySelects_1_io_ins_2),
    .io_ins_3(StickySelects_1_io_ins_3),
    .io_ins_4(StickySelects_1_io_ins_4),
    .io_ins_5(StickySelects_1_io_ins_5),
    .io_ins_6(StickySelects_1_io_ins_6),
    .io_ins_7(StickySelects_1_io_ins_7),
    .io_ins_8(StickySelects_1_io_ins_8),
    .io_outs_0(StickySelects_1_io_outs_0),
    .io_outs_1(StickySelects_1_io_outs_1),
    .io_outs_2(StickySelects_1_io_outs_2),
    .io_outs_3(StickySelects_1_io_outs_3),
    .io_outs_4(StickySelects_1_io_outs_4),
    .io_outs_5(StickySelects_1_io_outs_5),
    .io_outs_6(StickySelects_1_io_outs_6),
    .io_outs_7(StickySelects_1_io_outs_7),
    .io_outs_8(StickySelects_1_io_outs_8)
  );
  StickySelects_1 StickySelects_2 ( // @[MemPrimitives.scala 121:29:@21205.4]
    .clock(StickySelects_2_clock),
    .reset(StickySelects_2_reset),
    .io_ins_0(StickySelects_2_io_ins_0),
    .io_ins_1(StickySelects_2_io_ins_1),
    .io_ins_2(StickySelects_2_io_ins_2),
    .io_ins_3(StickySelects_2_io_ins_3),
    .io_ins_4(StickySelects_2_io_ins_4),
    .io_ins_5(StickySelects_2_io_ins_5),
    .io_ins_6(StickySelects_2_io_ins_6),
    .io_ins_7(StickySelects_2_io_ins_7),
    .io_ins_8(StickySelects_2_io_ins_8),
    .io_outs_0(StickySelects_2_io_outs_0),
    .io_outs_1(StickySelects_2_io_outs_1),
    .io_outs_2(StickySelects_2_io_outs_2),
    .io_outs_3(StickySelects_2_io_outs_3),
    .io_outs_4(StickySelects_2_io_outs_4),
    .io_outs_5(StickySelects_2_io_outs_5),
    .io_outs_6(StickySelects_2_io_outs_6),
    .io_outs_7(StickySelects_2_io_outs_7),
    .io_outs_8(StickySelects_2_io_outs_8)
  );
  StickySelects_1 StickySelects_3 ( // @[MemPrimitives.scala 121:29:@21294.4]
    .clock(StickySelects_3_clock),
    .reset(StickySelects_3_reset),
    .io_ins_0(StickySelects_3_io_ins_0),
    .io_ins_1(StickySelects_3_io_ins_1),
    .io_ins_2(StickySelects_3_io_ins_2),
    .io_ins_3(StickySelects_3_io_ins_3),
    .io_ins_4(StickySelects_3_io_ins_4),
    .io_ins_5(StickySelects_3_io_ins_5),
    .io_ins_6(StickySelects_3_io_ins_6),
    .io_ins_7(StickySelects_3_io_ins_7),
    .io_ins_8(StickySelects_3_io_ins_8),
    .io_outs_0(StickySelects_3_io_outs_0),
    .io_outs_1(StickySelects_3_io_outs_1),
    .io_outs_2(StickySelects_3_io_outs_2),
    .io_outs_3(StickySelects_3_io_outs_3),
    .io_outs_4(StickySelects_3_io_outs_4),
    .io_outs_5(StickySelects_3_io_outs_5),
    .io_outs_6(StickySelects_3_io_outs_6),
    .io_outs_7(StickySelects_3_io_outs_7),
    .io_outs_8(StickySelects_3_io_outs_8)
  );
  StickySelects_1 StickySelects_4 ( // @[MemPrimitives.scala 121:29:@21383.4]
    .clock(StickySelects_4_clock),
    .reset(StickySelects_4_reset),
    .io_ins_0(StickySelects_4_io_ins_0),
    .io_ins_1(StickySelects_4_io_ins_1),
    .io_ins_2(StickySelects_4_io_ins_2),
    .io_ins_3(StickySelects_4_io_ins_3),
    .io_ins_4(StickySelects_4_io_ins_4),
    .io_ins_5(StickySelects_4_io_ins_5),
    .io_ins_6(StickySelects_4_io_ins_6),
    .io_ins_7(StickySelects_4_io_ins_7),
    .io_ins_8(StickySelects_4_io_ins_8),
    .io_outs_0(StickySelects_4_io_outs_0),
    .io_outs_1(StickySelects_4_io_outs_1),
    .io_outs_2(StickySelects_4_io_outs_2),
    .io_outs_3(StickySelects_4_io_outs_3),
    .io_outs_4(StickySelects_4_io_outs_4),
    .io_outs_5(StickySelects_4_io_outs_5),
    .io_outs_6(StickySelects_4_io_outs_6),
    .io_outs_7(StickySelects_4_io_outs_7),
    .io_outs_8(StickySelects_4_io_outs_8)
  );
  StickySelects_1 StickySelects_5 ( // @[MemPrimitives.scala 121:29:@21472.4]
    .clock(StickySelects_5_clock),
    .reset(StickySelects_5_reset),
    .io_ins_0(StickySelects_5_io_ins_0),
    .io_ins_1(StickySelects_5_io_ins_1),
    .io_ins_2(StickySelects_5_io_ins_2),
    .io_ins_3(StickySelects_5_io_ins_3),
    .io_ins_4(StickySelects_5_io_ins_4),
    .io_ins_5(StickySelects_5_io_ins_5),
    .io_ins_6(StickySelects_5_io_ins_6),
    .io_ins_7(StickySelects_5_io_ins_7),
    .io_ins_8(StickySelects_5_io_ins_8),
    .io_outs_0(StickySelects_5_io_outs_0),
    .io_outs_1(StickySelects_5_io_outs_1),
    .io_outs_2(StickySelects_5_io_outs_2),
    .io_outs_3(StickySelects_5_io_outs_3),
    .io_outs_4(StickySelects_5_io_outs_4),
    .io_outs_5(StickySelects_5_io_outs_5),
    .io_outs_6(StickySelects_5_io_outs_6),
    .io_outs_7(StickySelects_5_io_outs_7),
    .io_outs_8(StickySelects_5_io_outs_8)
  );
  StickySelects_1 StickySelects_6 ( // @[MemPrimitives.scala 121:29:@21561.4]
    .clock(StickySelects_6_clock),
    .reset(StickySelects_6_reset),
    .io_ins_0(StickySelects_6_io_ins_0),
    .io_ins_1(StickySelects_6_io_ins_1),
    .io_ins_2(StickySelects_6_io_ins_2),
    .io_ins_3(StickySelects_6_io_ins_3),
    .io_ins_4(StickySelects_6_io_ins_4),
    .io_ins_5(StickySelects_6_io_ins_5),
    .io_ins_6(StickySelects_6_io_ins_6),
    .io_ins_7(StickySelects_6_io_ins_7),
    .io_ins_8(StickySelects_6_io_ins_8),
    .io_outs_0(StickySelects_6_io_outs_0),
    .io_outs_1(StickySelects_6_io_outs_1),
    .io_outs_2(StickySelects_6_io_outs_2),
    .io_outs_3(StickySelects_6_io_outs_3),
    .io_outs_4(StickySelects_6_io_outs_4),
    .io_outs_5(StickySelects_6_io_outs_5),
    .io_outs_6(StickySelects_6_io_outs_6),
    .io_outs_7(StickySelects_6_io_outs_7),
    .io_outs_8(StickySelects_6_io_outs_8)
  );
  StickySelects_1 StickySelects_7 ( // @[MemPrimitives.scala 121:29:@21650.4]
    .clock(StickySelects_7_clock),
    .reset(StickySelects_7_reset),
    .io_ins_0(StickySelects_7_io_ins_0),
    .io_ins_1(StickySelects_7_io_ins_1),
    .io_ins_2(StickySelects_7_io_ins_2),
    .io_ins_3(StickySelects_7_io_ins_3),
    .io_ins_4(StickySelects_7_io_ins_4),
    .io_ins_5(StickySelects_7_io_ins_5),
    .io_ins_6(StickySelects_7_io_ins_6),
    .io_ins_7(StickySelects_7_io_ins_7),
    .io_ins_8(StickySelects_7_io_ins_8),
    .io_outs_0(StickySelects_7_io_outs_0),
    .io_outs_1(StickySelects_7_io_outs_1),
    .io_outs_2(StickySelects_7_io_outs_2),
    .io_outs_3(StickySelects_7_io_outs_3),
    .io_outs_4(StickySelects_7_io_outs_4),
    .io_outs_5(StickySelects_7_io_outs_5),
    .io_outs_6(StickySelects_7_io_outs_6),
    .io_outs_7(StickySelects_7_io_outs_7),
    .io_outs_8(StickySelects_7_io_outs_8)
  );
  StickySelects_1 StickySelects_8 ( // @[MemPrimitives.scala 121:29:@21739.4]
    .clock(StickySelects_8_clock),
    .reset(StickySelects_8_reset),
    .io_ins_0(StickySelects_8_io_ins_0),
    .io_ins_1(StickySelects_8_io_ins_1),
    .io_ins_2(StickySelects_8_io_ins_2),
    .io_ins_3(StickySelects_8_io_ins_3),
    .io_ins_4(StickySelects_8_io_ins_4),
    .io_ins_5(StickySelects_8_io_ins_5),
    .io_ins_6(StickySelects_8_io_ins_6),
    .io_ins_7(StickySelects_8_io_ins_7),
    .io_ins_8(StickySelects_8_io_ins_8),
    .io_outs_0(StickySelects_8_io_outs_0),
    .io_outs_1(StickySelects_8_io_outs_1),
    .io_outs_2(StickySelects_8_io_outs_2),
    .io_outs_3(StickySelects_8_io_outs_3),
    .io_outs_4(StickySelects_8_io_outs_4),
    .io_outs_5(StickySelects_8_io_outs_5),
    .io_outs_6(StickySelects_8_io_outs_6),
    .io_outs_7(StickySelects_8_io_outs_7),
    .io_outs_8(StickySelects_8_io_outs_8)
  );
  StickySelects_1 StickySelects_9 ( // @[MemPrimitives.scala 121:29:@21828.4]
    .clock(StickySelects_9_clock),
    .reset(StickySelects_9_reset),
    .io_ins_0(StickySelects_9_io_ins_0),
    .io_ins_1(StickySelects_9_io_ins_1),
    .io_ins_2(StickySelects_9_io_ins_2),
    .io_ins_3(StickySelects_9_io_ins_3),
    .io_ins_4(StickySelects_9_io_ins_4),
    .io_ins_5(StickySelects_9_io_ins_5),
    .io_ins_6(StickySelects_9_io_ins_6),
    .io_ins_7(StickySelects_9_io_ins_7),
    .io_ins_8(StickySelects_9_io_ins_8),
    .io_outs_0(StickySelects_9_io_outs_0),
    .io_outs_1(StickySelects_9_io_outs_1),
    .io_outs_2(StickySelects_9_io_outs_2),
    .io_outs_3(StickySelects_9_io_outs_3),
    .io_outs_4(StickySelects_9_io_outs_4),
    .io_outs_5(StickySelects_9_io_outs_5),
    .io_outs_6(StickySelects_9_io_outs_6),
    .io_outs_7(StickySelects_9_io_outs_7),
    .io_outs_8(StickySelects_9_io_outs_8)
  );
  StickySelects_1 StickySelects_10 ( // @[MemPrimitives.scala 121:29:@21917.4]
    .clock(StickySelects_10_clock),
    .reset(StickySelects_10_reset),
    .io_ins_0(StickySelects_10_io_ins_0),
    .io_ins_1(StickySelects_10_io_ins_1),
    .io_ins_2(StickySelects_10_io_ins_2),
    .io_ins_3(StickySelects_10_io_ins_3),
    .io_ins_4(StickySelects_10_io_ins_4),
    .io_ins_5(StickySelects_10_io_ins_5),
    .io_ins_6(StickySelects_10_io_ins_6),
    .io_ins_7(StickySelects_10_io_ins_7),
    .io_ins_8(StickySelects_10_io_ins_8),
    .io_outs_0(StickySelects_10_io_outs_0),
    .io_outs_1(StickySelects_10_io_outs_1),
    .io_outs_2(StickySelects_10_io_outs_2),
    .io_outs_3(StickySelects_10_io_outs_3),
    .io_outs_4(StickySelects_10_io_outs_4),
    .io_outs_5(StickySelects_10_io_outs_5),
    .io_outs_6(StickySelects_10_io_outs_6),
    .io_outs_7(StickySelects_10_io_outs_7),
    .io_outs_8(StickySelects_10_io_outs_8)
  );
  StickySelects_1 StickySelects_11 ( // @[MemPrimitives.scala 121:29:@22006.4]
    .clock(StickySelects_11_clock),
    .reset(StickySelects_11_reset),
    .io_ins_0(StickySelects_11_io_ins_0),
    .io_ins_1(StickySelects_11_io_ins_1),
    .io_ins_2(StickySelects_11_io_ins_2),
    .io_ins_3(StickySelects_11_io_ins_3),
    .io_ins_4(StickySelects_11_io_ins_4),
    .io_ins_5(StickySelects_11_io_ins_5),
    .io_ins_6(StickySelects_11_io_ins_6),
    .io_ins_7(StickySelects_11_io_ins_7),
    .io_ins_8(StickySelects_11_io_ins_8),
    .io_outs_0(StickySelects_11_io_outs_0),
    .io_outs_1(StickySelects_11_io_outs_1),
    .io_outs_2(StickySelects_11_io_outs_2),
    .io_outs_3(StickySelects_11_io_outs_3),
    .io_outs_4(StickySelects_11_io_outs_4),
    .io_outs_5(StickySelects_11_io_outs_5),
    .io_outs_6(StickySelects_11_io_outs_6),
    .io_outs_7(StickySelects_11_io_outs_7),
    .io_outs_8(StickySelects_11_io_outs_8)
  );
  StickySelects_1 StickySelects_12 ( // @[MemPrimitives.scala 121:29:@22095.4]
    .clock(StickySelects_12_clock),
    .reset(StickySelects_12_reset),
    .io_ins_0(StickySelects_12_io_ins_0),
    .io_ins_1(StickySelects_12_io_ins_1),
    .io_ins_2(StickySelects_12_io_ins_2),
    .io_ins_3(StickySelects_12_io_ins_3),
    .io_ins_4(StickySelects_12_io_ins_4),
    .io_ins_5(StickySelects_12_io_ins_5),
    .io_ins_6(StickySelects_12_io_ins_6),
    .io_ins_7(StickySelects_12_io_ins_7),
    .io_ins_8(StickySelects_12_io_ins_8),
    .io_outs_0(StickySelects_12_io_outs_0),
    .io_outs_1(StickySelects_12_io_outs_1),
    .io_outs_2(StickySelects_12_io_outs_2),
    .io_outs_3(StickySelects_12_io_outs_3),
    .io_outs_4(StickySelects_12_io_outs_4),
    .io_outs_5(StickySelects_12_io_outs_5),
    .io_outs_6(StickySelects_12_io_outs_6),
    .io_outs_7(StickySelects_12_io_outs_7),
    .io_outs_8(StickySelects_12_io_outs_8)
  );
  StickySelects_1 StickySelects_13 ( // @[MemPrimitives.scala 121:29:@22184.4]
    .clock(StickySelects_13_clock),
    .reset(StickySelects_13_reset),
    .io_ins_0(StickySelects_13_io_ins_0),
    .io_ins_1(StickySelects_13_io_ins_1),
    .io_ins_2(StickySelects_13_io_ins_2),
    .io_ins_3(StickySelects_13_io_ins_3),
    .io_ins_4(StickySelects_13_io_ins_4),
    .io_ins_5(StickySelects_13_io_ins_5),
    .io_ins_6(StickySelects_13_io_ins_6),
    .io_ins_7(StickySelects_13_io_ins_7),
    .io_ins_8(StickySelects_13_io_ins_8),
    .io_outs_0(StickySelects_13_io_outs_0),
    .io_outs_1(StickySelects_13_io_outs_1),
    .io_outs_2(StickySelects_13_io_outs_2),
    .io_outs_3(StickySelects_13_io_outs_3),
    .io_outs_4(StickySelects_13_io_outs_4),
    .io_outs_5(StickySelects_13_io_outs_5),
    .io_outs_6(StickySelects_13_io_outs_6),
    .io_outs_7(StickySelects_13_io_outs_7),
    .io_outs_8(StickySelects_13_io_outs_8)
  );
  StickySelects_1 StickySelects_14 ( // @[MemPrimitives.scala 121:29:@22273.4]
    .clock(StickySelects_14_clock),
    .reset(StickySelects_14_reset),
    .io_ins_0(StickySelects_14_io_ins_0),
    .io_ins_1(StickySelects_14_io_ins_1),
    .io_ins_2(StickySelects_14_io_ins_2),
    .io_ins_3(StickySelects_14_io_ins_3),
    .io_ins_4(StickySelects_14_io_ins_4),
    .io_ins_5(StickySelects_14_io_ins_5),
    .io_ins_6(StickySelects_14_io_ins_6),
    .io_ins_7(StickySelects_14_io_ins_7),
    .io_ins_8(StickySelects_14_io_ins_8),
    .io_outs_0(StickySelects_14_io_outs_0),
    .io_outs_1(StickySelects_14_io_outs_1),
    .io_outs_2(StickySelects_14_io_outs_2),
    .io_outs_3(StickySelects_14_io_outs_3),
    .io_outs_4(StickySelects_14_io_outs_4),
    .io_outs_5(StickySelects_14_io_outs_5),
    .io_outs_6(StickySelects_14_io_outs_6),
    .io_outs_7(StickySelects_14_io_outs_7),
    .io_outs_8(StickySelects_14_io_outs_8)
  );
  StickySelects_1 StickySelects_15 ( // @[MemPrimitives.scala 121:29:@22362.4]
    .clock(StickySelects_15_clock),
    .reset(StickySelects_15_reset),
    .io_ins_0(StickySelects_15_io_ins_0),
    .io_ins_1(StickySelects_15_io_ins_1),
    .io_ins_2(StickySelects_15_io_ins_2),
    .io_ins_3(StickySelects_15_io_ins_3),
    .io_ins_4(StickySelects_15_io_ins_4),
    .io_ins_5(StickySelects_15_io_ins_5),
    .io_ins_6(StickySelects_15_io_ins_6),
    .io_ins_7(StickySelects_15_io_ins_7),
    .io_ins_8(StickySelects_15_io_ins_8),
    .io_outs_0(StickySelects_15_io_outs_0),
    .io_outs_1(StickySelects_15_io_outs_1),
    .io_outs_2(StickySelects_15_io_outs_2),
    .io_outs_3(StickySelects_15_io_outs_3),
    .io_outs_4(StickySelects_15_io_outs_4),
    .io_outs_5(StickySelects_15_io_outs_5),
    .io_outs_6(StickySelects_15_io_outs_6),
    .io_outs_7(StickySelects_15_io_outs_7),
    .io_outs_8(StickySelects_15_io_outs_8)
  );
  StickySelects_1 StickySelects_16 ( // @[MemPrimitives.scala 121:29:@22451.4]
    .clock(StickySelects_16_clock),
    .reset(StickySelects_16_reset),
    .io_ins_0(StickySelects_16_io_ins_0),
    .io_ins_1(StickySelects_16_io_ins_1),
    .io_ins_2(StickySelects_16_io_ins_2),
    .io_ins_3(StickySelects_16_io_ins_3),
    .io_ins_4(StickySelects_16_io_ins_4),
    .io_ins_5(StickySelects_16_io_ins_5),
    .io_ins_6(StickySelects_16_io_ins_6),
    .io_ins_7(StickySelects_16_io_ins_7),
    .io_ins_8(StickySelects_16_io_ins_8),
    .io_outs_0(StickySelects_16_io_outs_0),
    .io_outs_1(StickySelects_16_io_outs_1),
    .io_outs_2(StickySelects_16_io_outs_2),
    .io_outs_3(StickySelects_16_io_outs_3),
    .io_outs_4(StickySelects_16_io_outs_4),
    .io_outs_5(StickySelects_16_io_outs_5),
    .io_outs_6(StickySelects_16_io_outs_6),
    .io_outs_7(StickySelects_16_io_outs_7),
    .io_outs_8(StickySelects_16_io_outs_8)
  );
  StickySelects_1 StickySelects_17 ( // @[MemPrimitives.scala 121:29:@22540.4]
    .clock(StickySelects_17_clock),
    .reset(StickySelects_17_reset),
    .io_ins_0(StickySelects_17_io_ins_0),
    .io_ins_1(StickySelects_17_io_ins_1),
    .io_ins_2(StickySelects_17_io_ins_2),
    .io_ins_3(StickySelects_17_io_ins_3),
    .io_ins_4(StickySelects_17_io_ins_4),
    .io_ins_5(StickySelects_17_io_ins_5),
    .io_ins_6(StickySelects_17_io_ins_6),
    .io_ins_7(StickySelects_17_io_ins_7),
    .io_ins_8(StickySelects_17_io_ins_8),
    .io_outs_0(StickySelects_17_io_outs_0),
    .io_outs_1(StickySelects_17_io_outs_1),
    .io_outs_2(StickySelects_17_io_outs_2),
    .io_outs_3(StickySelects_17_io_outs_3),
    .io_outs_4(StickySelects_17_io_outs_4),
    .io_outs_5(StickySelects_17_io_outs_5),
    .io_outs_6(StickySelects_17_io_outs_6),
    .io_outs_7(StickySelects_17_io_outs_7),
    .io_outs_8(StickySelects_17_io_outs_8)
  );
  StickySelects_1 StickySelects_18 ( // @[MemPrimitives.scala 121:29:@22629.4]
    .clock(StickySelects_18_clock),
    .reset(StickySelects_18_reset),
    .io_ins_0(StickySelects_18_io_ins_0),
    .io_ins_1(StickySelects_18_io_ins_1),
    .io_ins_2(StickySelects_18_io_ins_2),
    .io_ins_3(StickySelects_18_io_ins_3),
    .io_ins_4(StickySelects_18_io_ins_4),
    .io_ins_5(StickySelects_18_io_ins_5),
    .io_ins_6(StickySelects_18_io_ins_6),
    .io_ins_7(StickySelects_18_io_ins_7),
    .io_ins_8(StickySelects_18_io_ins_8),
    .io_outs_0(StickySelects_18_io_outs_0),
    .io_outs_1(StickySelects_18_io_outs_1),
    .io_outs_2(StickySelects_18_io_outs_2),
    .io_outs_3(StickySelects_18_io_outs_3),
    .io_outs_4(StickySelects_18_io_outs_4),
    .io_outs_5(StickySelects_18_io_outs_5),
    .io_outs_6(StickySelects_18_io_outs_6),
    .io_outs_7(StickySelects_18_io_outs_7),
    .io_outs_8(StickySelects_18_io_outs_8)
  );
  StickySelects_1 StickySelects_19 ( // @[MemPrimitives.scala 121:29:@22718.4]
    .clock(StickySelects_19_clock),
    .reset(StickySelects_19_reset),
    .io_ins_0(StickySelects_19_io_ins_0),
    .io_ins_1(StickySelects_19_io_ins_1),
    .io_ins_2(StickySelects_19_io_ins_2),
    .io_ins_3(StickySelects_19_io_ins_3),
    .io_ins_4(StickySelects_19_io_ins_4),
    .io_ins_5(StickySelects_19_io_ins_5),
    .io_ins_6(StickySelects_19_io_ins_6),
    .io_ins_7(StickySelects_19_io_ins_7),
    .io_ins_8(StickySelects_19_io_ins_8),
    .io_outs_0(StickySelects_19_io_outs_0),
    .io_outs_1(StickySelects_19_io_outs_1),
    .io_outs_2(StickySelects_19_io_outs_2),
    .io_outs_3(StickySelects_19_io_outs_3),
    .io_outs_4(StickySelects_19_io_outs_4),
    .io_outs_5(StickySelects_19_io_outs_5),
    .io_outs_6(StickySelects_19_io_outs_6),
    .io_outs_7(StickySelects_19_io_outs_7),
    .io_outs_8(StickySelects_19_io_outs_8)
  );
  StickySelects_1 StickySelects_20 ( // @[MemPrimitives.scala 121:29:@22807.4]
    .clock(StickySelects_20_clock),
    .reset(StickySelects_20_reset),
    .io_ins_0(StickySelects_20_io_ins_0),
    .io_ins_1(StickySelects_20_io_ins_1),
    .io_ins_2(StickySelects_20_io_ins_2),
    .io_ins_3(StickySelects_20_io_ins_3),
    .io_ins_4(StickySelects_20_io_ins_4),
    .io_ins_5(StickySelects_20_io_ins_5),
    .io_ins_6(StickySelects_20_io_ins_6),
    .io_ins_7(StickySelects_20_io_ins_7),
    .io_ins_8(StickySelects_20_io_ins_8),
    .io_outs_0(StickySelects_20_io_outs_0),
    .io_outs_1(StickySelects_20_io_outs_1),
    .io_outs_2(StickySelects_20_io_outs_2),
    .io_outs_3(StickySelects_20_io_outs_3),
    .io_outs_4(StickySelects_20_io_outs_4),
    .io_outs_5(StickySelects_20_io_outs_5),
    .io_outs_6(StickySelects_20_io_outs_6),
    .io_outs_7(StickySelects_20_io_outs_7),
    .io_outs_8(StickySelects_20_io_outs_8)
  );
  StickySelects_1 StickySelects_21 ( // @[MemPrimitives.scala 121:29:@22896.4]
    .clock(StickySelects_21_clock),
    .reset(StickySelects_21_reset),
    .io_ins_0(StickySelects_21_io_ins_0),
    .io_ins_1(StickySelects_21_io_ins_1),
    .io_ins_2(StickySelects_21_io_ins_2),
    .io_ins_3(StickySelects_21_io_ins_3),
    .io_ins_4(StickySelects_21_io_ins_4),
    .io_ins_5(StickySelects_21_io_ins_5),
    .io_ins_6(StickySelects_21_io_ins_6),
    .io_ins_7(StickySelects_21_io_ins_7),
    .io_ins_8(StickySelects_21_io_ins_8),
    .io_outs_0(StickySelects_21_io_outs_0),
    .io_outs_1(StickySelects_21_io_outs_1),
    .io_outs_2(StickySelects_21_io_outs_2),
    .io_outs_3(StickySelects_21_io_outs_3),
    .io_outs_4(StickySelects_21_io_outs_4),
    .io_outs_5(StickySelects_21_io_outs_5),
    .io_outs_6(StickySelects_21_io_outs_6),
    .io_outs_7(StickySelects_21_io_outs_7),
    .io_outs_8(StickySelects_21_io_outs_8)
  );
  StickySelects_1 StickySelects_22 ( // @[MemPrimitives.scala 121:29:@22985.4]
    .clock(StickySelects_22_clock),
    .reset(StickySelects_22_reset),
    .io_ins_0(StickySelects_22_io_ins_0),
    .io_ins_1(StickySelects_22_io_ins_1),
    .io_ins_2(StickySelects_22_io_ins_2),
    .io_ins_3(StickySelects_22_io_ins_3),
    .io_ins_4(StickySelects_22_io_ins_4),
    .io_ins_5(StickySelects_22_io_ins_5),
    .io_ins_6(StickySelects_22_io_ins_6),
    .io_ins_7(StickySelects_22_io_ins_7),
    .io_ins_8(StickySelects_22_io_ins_8),
    .io_outs_0(StickySelects_22_io_outs_0),
    .io_outs_1(StickySelects_22_io_outs_1),
    .io_outs_2(StickySelects_22_io_outs_2),
    .io_outs_3(StickySelects_22_io_outs_3),
    .io_outs_4(StickySelects_22_io_outs_4),
    .io_outs_5(StickySelects_22_io_outs_5),
    .io_outs_6(StickySelects_22_io_outs_6),
    .io_outs_7(StickySelects_22_io_outs_7),
    .io_outs_8(StickySelects_22_io_outs_8)
  );
  StickySelects_1 StickySelects_23 ( // @[MemPrimitives.scala 121:29:@23074.4]
    .clock(StickySelects_23_clock),
    .reset(StickySelects_23_reset),
    .io_ins_0(StickySelects_23_io_ins_0),
    .io_ins_1(StickySelects_23_io_ins_1),
    .io_ins_2(StickySelects_23_io_ins_2),
    .io_ins_3(StickySelects_23_io_ins_3),
    .io_ins_4(StickySelects_23_io_ins_4),
    .io_ins_5(StickySelects_23_io_ins_5),
    .io_ins_6(StickySelects_23_io_ins_6),
    .io_ins_7(StickySelects_23_io_ins_7),
    .io_ins_8(StickySelects_23_io_ins_8),
    .io_outs_0(StickySelects_23_io_outs_0),
    .io_outs_1(StickySelects_23_io_outs_1),
    .io_outs_2(StickySelects_23_io_outs_2),
    .io_outs_3(StickySelects_23_io_outs_3),
    .io_outs_4(StickySelects_23_io_outs_4),
    .io_outs_5(StickySelects_23_io_outs_5),
    .io_outs_6(StickySelects_23_io_outs_6),
    .io_outs_7(StickySelects_23_io_outs_7),
    .io_outs_8(StickySelects_23_io_outs_8)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@23164.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@23172.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_2 ( // @[package.scala 93:22:@23180.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_3 ( // @[package.scala 93:22:@23188.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_4 ( // @[package.scala 93:22:@23196.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_5 ( // @[package.scala 93:22:@23204.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_6 ( // @[package.scala 93:22:@23212.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_7 ( // @[package.scala 93:22:@23220.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_8 ( // @[package.scala 93:22:@23228.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_9 ( // @[package.scala 93:22:@23236.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_10 ( // @[package.scala 93:22:@23244.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_11 ( // @[package.scala 93:22:@23252.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_12 ( // @[package.scala 93:22:@23308.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_13 ( // @[package.scala 93:22:@23316.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_14 ( // @[package.scala 93:22:@23324.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_15 ( // @[package.scala 93:22:@23332.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_16 ( // @[package.scala 93:22:@23340.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_17 ( // @[package.scala 93:22:@23348.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_18 ( // @[package.scala 93:22:@23356.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_19 ( // @[package.scala 93:22:@23364.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_20 ( // @[package.scala 93:22:@23372.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_21 ( // @[package.scala 93:22:@23380.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_22 ( // @[package.scala 93:22:@23388.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_23 ( // @[package.scala 93:22:@23396.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_24 ( // @[package.scala 93:22:@23452.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_25 ( // @[package.scala 93:22:@23460.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_26 ( // @[package.scala 93:22:@23468.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_27 ( // @[package.scala 93:22:@23476.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_28 ( // @[package.scala 93:22:@23484.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_29 ( // @[package.scala 93:22:@23492.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_30 ( // @[package.scala 93:22:@23500.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_31 ( // @[package.scala 93:22:@23508.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_32 ( // @[package.scala 93:22:@23516.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_33 ( // @[package.scala 93:22:@23524.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_34 ( // @[package.scala 93:22:@23532.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_35 ( // @[package.scala 93:22:@23540.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_36 ( // @[package.scala 93:22:@23596.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_37 ( // @[package.scala 93:22:@23604.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_38 ( // @[package.scala 93:22:@23612.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_39 ( // @[package.scala 93:22:@23620.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_40 ( // @[package.scala 93:22:@23628.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_41 ( // @[package.scala 93:22:@23636.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_42 ( // @[package.scala 93:22:@23644.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_43 ( // @[package.scala 93:22:@23652.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_44 ( // @[package.scala 93:22:@23660.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_45 ( // @[package.scala 93:22:@23668.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_46 ( // @[package.scala 93:22:@23676.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_47 ( // @[package.scala 93:22:@23684.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_48 ( // @[package.scala 93:22:@23740.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_49 ( // @[package.scala 93:22:@23748.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_50 ( // @[package.scala 93:22:@23756.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_51 ( // @[package.scala 93:22:@23764.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_52 ( // @[package.scala 93:22:@23772.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_53 ( // @[package.scala 93:22:@23780.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_54 ( // @[package.scala 93:22:@23788.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_55 ( // @[package.scala 93:22:@23796.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_56 ( // @[package.scala 93:22:@23804.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_57 ( // @[package.scala 93:22:@23812.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_58 ( // @[package.scala 93:22:@23820.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_59 ( // @[package.scala 93:22:@23828.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_60 ( // @[package.scala 93:22:@23884.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_61 ( // @[package.scala 93:22:@23892.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_62 ( // @[package.scala 93:22:@23900.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_63 ( // @[package.scala 93:22:@23908.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_64 ( // @[package.scala 93:22:@23916.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_65 ( // @[package.scala 93:22:@23924.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_66 ( // @[package.scala 93:22:@23932.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_67 ( // @[package.scala 93:22:@23940.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_68 ( // @[package.scala 93:22:@23948.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_69 ( // @[package.scala 93:22:@23956.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_70 ( // @[package.scala 93:22:@23964.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_71 ( // @[package.scala 93:22:@23972.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_72 ( // @[package.scala 93:22:@24028.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_73 ( // @[package.scala 93:22:@24036.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_74 ( // @[package.scala 93:22:@24044.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_75 ( // @[package.scala 93:22:@24052.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_76 ( // @[package.scala 93:22:@24060.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_77 ( // @[package.scala 93:22:@24068.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_78 ( // @[package.scala 93:22:@24076.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_79 ( // @[package.scala 93:22:@24084.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_80 ( // @[package.scala 93:22:@24092.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_81 ( // @[package.scala 93:22:@24100.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_82 ( // @[package.scala 93:22:@24108.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_83 ( // @[package.scala 93:22:@24116.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_84 ( // @[package.scala 93:22:@24172.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_85 ( // @[package.scala 93:22:@24180.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_86 ( // @[package.scala 93:22:@24188.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_87 ( // @[package.scala 93:22:@24196.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_88 ( // @[package.scala 93:22:@24204.4]
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_89 ( // @[package.scala 93:22:@24212.4]
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_90 ( // @[package.scala 93:22:@24220.4]
    .clock(RetimeWrapper_90_clock),
    .reset(RetimeWrapper_90_reset),
    .io_flow(RetimeWrapper_90_io_flow),
    .io_in(RetimeWrapper_90_io_in),
    .io_out(RetimeWrapper_90_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_91 ( // @[package.scala 93:22:@24228.4]
    .clock(RetimeWrapper_91_clock),
    .reset(RetimeWrapper_91_reset),
    .io_flow(RetimeWrapper_91_io_flow),
    .io_in(RetimeWrapper_91_io_in),
    .io_out(RetimeWrapper_91_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_92 ( // @[package.scala 93:22:@24236.4]
    .clock(RetimeWrapper_92_clock),
    .reset(RetimeWrapper_92_reset),
    .io_flow(RetimeWrapper_92_io_flow),
    .io_in(RetimeWrapper_92_io_in),
    .io_out(RetimeWrapper_92_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_93 ( // @[package.scala 93:22:@24244.4]
    .clock(RetimeWrapper_93_clock),
    .reset(RetimeWrapper_93_reset),
    .io_flow(RetimeWrapper_93_io_flow),
    .io_in(RetimeWrapper_93_io_in),
    .io_out(RetimeWrapper_93_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_94 ( // @[package.scala 93:22:@24252.4]
    .clock(RetimeWrapper_94_clock),
    .reset(RetimeWrapper_94_reset),
    .io_flow(RetimeWrapper_94_io_flow),
    .io_in(RetimeWrapper_94_io_in),
    .io_out(RetimeWrapper_94_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_95 ( // @[package.scala 93:22:@24260.4]
    .clock(RetimeWrapper_95_clock),
    .reset(RetimeWrapper_95_reset),
    .io_flow(RetimeWrapper_95_io_flow),
    .io_in(RetimeWrapper_95_io_in),
    .io_out(RetimeWrapper_95_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_96 ( // @[package.scala 93:22:@24316.4]
    .clock(RetimeWrapper_96_clock),
    .reset(RetimeWrapper_96_reset),
    .io_flow(RetimeWrapper_96_io_flow),
    .io_in(RetimeWrapper_96_io_in),
    .io_out(RetimeWrapper_96_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_97 ( // @[package.scala 93:22:@24324.4]
    .clock(RetimeWrapper_97_clock),
    .reset(RetimeWrapper_97_reset),
    .io_flow(RetimeWrapper_97_io_flow),
    .io_in(RetimeWrapper_97_io_in),
    .io_out(RetimeWrapper_97_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_98 ( // @[package.scala 93:22:@24332.4]
    .clock(RetimeWrapper_98_clock),
    .reset(RetimeWrapper_98_reset),
    .io_flow(RetimeWrapper_98_io_flow),
    .io_in(RetimeWrapper_98_io_in),
    .io_out(RetimeWrapper_98_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_99 ( // @[package.scala 93:22:@24340.4]
    .clock(RetimeWrapper_99_clock),
    .reset(RetimeWrapper_99_reset),
    .io_flow(RetimeWrapper_99_io_flow),
    .io_in(RetimeWrapper_99_io_in),
    .io_out(RetimeWrapper_99_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_100 ( // @[package.scala 93:22:@24348.4]
    .clock(RetimeWrapper_100_clock),
    .reset(RetimeWrapper_100_reset),
    .io_flow(RetimeWrapper_100_io_flow),
    .io_in(RetimeWrapper_100_io_in),
    .io_out(RetimeWrapper_100_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_101 ( // @[package.scala 93:22:@24356.4]
    .clock(RetimeWrapper_101_clock),
    .reset(RetimeWrapper_101_reset),
    .io_flow(RetimeWrapper_101_io_flow),
    .io_in(RetimeWrapper_101_io_in),
    .io_out(RetimeWrapper_101_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_102 ( // @[package.scala 93:22:@24364.4]
    .clock(RetimeWrapper_102_clock),
    .reset(RetimeWrapper_102_reset),
    .io_flow(RetimeWrapper_102_io_flow),
    .io_in(RetimeWrapper_102_io_in),
    .io_out(RetimeWrapper_102_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_103 ( // @[package.scala 93:22:@24372.4]
    .clock(RetimeWrapper_103_clock),
    .reset(RetimeWrapper_103_reset),
    .io_flow(RetimeWrapper_103_io_flow),
    .io_in(RetimeWrapper_103_io_in),
    .io_out(RetimeWrapper_103_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_104 ( // @[package.scala 93:22:@24380.4]
    .clock(RetimeWrapper_104_clock),
    .reset(RetimeWrapper_104_reset),
    .io_flow(RetimeWrapper_104_io_flow),
    .io_in(RetimeWrapper_104_io_in),
    .io_out(RetimeWrapper_104_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_105 ( // @[package.scala 93:22:@24388.4]
    .clock(RetimeWrapper_105_clock),
    .reset(RetimeWrapper_105_reset),
    .io_flow(RetimeWrapper_105_io_flow),
    .io_in(RetimeWrapper_105_io_in),
    .io_out(RetimeWrapper_105_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_106 ( // @[package.scala 93:22:@24396.4]
    .clock(RetimeWrapper_106_clock),
    .reset(RetimeWrapper_106_reset),
    .io_flow(RetimeWrapper_106_io_flow),
    .io_in(RetimeWrapper_106_io_in),
    .io_out(RetimeWrapper_106_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_107 ( // @[package.scala 93:22:@24404.4]
    .clock(RetimeWrapper_107_clock),
    .reset(RetimeWrapper_107_reset),
    .io_flow(RetimeWrapper_107_io_flow),
    .io_in(RetimeWrapper_107_io_in),
    .io_out(RetimeWrapper_107_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_108 ( // @[package.scala 93:22:@24460.4]
    .clock(RetimeWrapper_108_clock),
    .reset(RetimeWrapper_108_reset),
    .io_flow(RetimeWrapper_108_io_flow),
    .io_in(RetimeWrapper_108_io_in),
    .io_out(RetimeWrapper_108_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_109 ( // @[package.scala 93:22:@24468.4]
    .clock(RetimeWrapper_109_clock),
    .reset(RetimeWrapper_109_reset),
    .io_flow(RetimeWrapper_109_io_flow),
    .io_in(RetimeWrapper_109_io_in),
    .io_out(RetimeWrapper_109_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_110 ( // @[package.scala 93:22:@24476.4]
    .clock(RetimeWrapper_110_clock),
    .reset(RetimeWrapper_110_reset),
    .io_flow(RetimeWrapper_110_io_flow),
    .io_in(RetimeWrapper_110_io_in),
    .io_out(RetimeWrapper_110_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_111 ( // @[package.scala 93:22:@24484.4]
    .clock(RetimeWrapper_111_clock),
    .reset(RetimeWrapper_111_reset),
    .io_flow(RetimeWrapper_111_io_flow),
    .io_in(RetimeWrapper_111_io_in),
    .io_out(RetimeWrapper_111_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_112 ( // @[package.scala 93:22:@24492.4]
    .clock(RetimeWrapper_112_clock),
    .reset(RetimeWrapper_112_reset),
    .io_flow(RetimeWrapper_112_io_flow),
    .io_in(RetimeWrapper_112_io_in),
    .io_out(RetimeWrapper_112_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_113 ( // @[package.scala 93:22:@24500.4]
    .clock(RetimeWrapper_113_clock),
    .reset(RetimeWrapper_113_reset),
    .io_flow(RetimeWrapper_113_io_flow),
    .io_in(RetimeWrapper_113_io_in),
    .io_out(RetimeWrapper_113_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_114 ( // @[package.scala 93:22:@24508.4]
    .clock(RetimeWrapper_114_clock),
    .reset(RetimeWrapper_114_reset),
    .io_flow(RetimeWrapper_114_io_flow),
    .io_in(RetimeWrapper_114_io_in),
    .io_out(RetimeWrapper_114_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_115 ( // @[package.scala 93:22:@24516.4]
    .clock(RetimeWrapper_115_clock),
    .reset(RetimeWrapper_115_reset),
    .io_flow(RetimeWrapper_115_io_flow),
    .io_in(RetimeWrapper_115_io_in),
    .io_out(RetimeWrapper_115_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_116 ( // @[package.scala 93:22:@24524.4]
    .clock(RetimeWrapper_116_clock),
    .reset(RetimeWrapper_116_reset),
    .io_flow(RetimeWrapper_116_io_flow),
    .io_in(RetimeWrapper_116_io_in),
    .io_out(RetimeWrapper_116_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_117 ( // @[package.scala 93:22:@24532.4]
    .clock(RetimeWrapper_117_clock),
    .reset(RetimeWrapper_117_reset),
    .io_flow(RetimeWrapper_117_io_flow),
    .io_in(RetimeWrapper_117_io_in),
    .io_out(RetimeWrapper_117_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_118 ( // @[package.scala 93:22:@24540.4]
    .clock(RetimeWrapper_118_clock),
    .reset(RetimeWrapper_118_reset),
    .io_flow(RetimeWrapper_118_io_flow),
    .io_in(RetimeWrapper_118_io_in),
    .io_out(RetimeWrapper_118_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_119 ( // @[package.scala 93:22:@24548.4]
    .clock(RetimeWrapper_119_clock),
    .reset(RetimeWrapper_119_reset),
    .io_flow(RetimeWrapper_119_io_flow),
    .io_in(RetimeWrapper_119_io_in),
    .io_out(RetimeWrapper_119_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_120 ( // @[package.scala 93:22:@24604.4]
    .clock(RetimeWrapper_120_clock),
    .reset(RetimeWrapper_120_reset),
    .io_flow(RetimeWrapper_120_io_flow),
    .io_in(RetimeWrapper_120_io_in),
    .io_out(RetimeWrapper_120_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_121 ( // @[package.scala 93:22:@24612.4]
    .clock(RetimeWrapper_121_clock),
    .reset(RetimeWrapper_121_reset),
    .io_flow(RetimeWrapper_121_io_flow),
    .io_in(RetimeWrapper_121_io_in),
    .io_out(RetimeWrapper_121_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_122 ( // @[package.scala 93:22:@24620.4]
    .clock(RetimeWrapper_122_clock),
    .reset(RetimeWrapper_122_reset),
    .io_flow(RetimeWrapper_122_io_flow),
    .io_in(RetimeWrapper_122_io_in),
    .io_out(RetimeWrapper_122_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_123 ( // @[package.scala 93:22:@24628.4]
    .clock(RetimeWrapper_123_clock),
    .reset(RetimeWrapper_123_reset),
    .io_flow(RetimeWrapper_123_io_flow),
    .io_in(RetimeWrapper_123_io_in),
    .io_out(RetimeWrapper_123_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_124 ( // @[package.scala 93:22:@24636.4]
    .clock(RetimeWrapper_124_clock),
    .reset(RetimeWrapper_124_reset),
    .io_flow(RetimeWrapper_124_io_flow),
    .io_in(RetimeWrapper_124_io_in),
    .io_out(RetimeWrapper_124_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_125 ( // @[package.scala 93:22:@24644.4]
    .clock(RetimeWrapper_125_clock),
    .reset(RetimeWrapper_125_reset),
    .io_flow(RetimeWrapper_125_io_flow),
    .io_in(RetimeWrapper_125_io_in),
    .io_out(RetimeWrapper_125_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_126 ( // @[package.scala 93:22:@24652.4]
    .clock(RetimeWrapper_126_clock),
    .reset(RetimeWrapper_126_reset),
    .io_flow(RetimeWrapper_126_io_flow),
    .io_in(RetimeWrapper_126_io_in),
    .io_out(RetimeWrapper_126_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_127 ( // @[package.scala 93:22:@24660.4]
    .clock(RetimeWrapper_127_clock),
    .reset(RetimeWrapper_127_reset),
    .io_flow(RetimeWrapper_127_io_flow),
    .io_in(RetimeWrapper_127_io_in),
    .io_out(RetimeWrapper_127_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_128 ( // @[package.scala 93:22:@24668.4]
    .clock(RetimeWrapper_128_clock),
    .reset(RetimeWrapper_128_reset),
    .io_flow(RetimeWrapper_128_io_flow),
    .io_in(RetimeWrapper_128_io_in),
    .io_out(RetimeWrapper_128_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_129 ( // @[package.scala 93:22:@24676.4]
    .clock(RetimeWrapper_129_clock),
    .reset(RetimeWrapper_129_reset),
    .io_flow(RetimeWrapper_129_io_flow),
    .io_in(RetimeWrapper_129_io_in),
    .io_out(RetimeWrapper_129_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_130 ( // @[package.scala 93:22:@24684.4]
    .clock(RetimeWrapper_130_clock),
    .reset(RetimeWrapper_130_reset),
    .io_flow(RetimeWrapper_130_io_flow),
    .io_in(RetimeWrapper_130_io_in),
    .io_out(RetimeWrapper_130_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_131 ( // @[package.scala 93:22:@24692.4]
    .clock(RetimeWrapper_131_clock),
    .reset(RetimeWrapper_131_reset),
    .io_flow(RetimeWrapper_131_io_flow),
    .io_in(RetimeWrapper_131_io_in),
    .io_out(RetimeWrapper_131_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_132 ( // @[package.scala 93:22:@24748.4]
    .clock(RetimeWrapper_132_clock),
    .reset(RetimeWrapper_132_reset),
    .io_flow(RetimeWrapper_132_io_flow),
    .io_in(RetimeWrapper_132_io_in),
    .io_out(RetimeWrapper_132_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_133 ( // @[package.scala 93:22:@24756.4]
    .clock(RetimeWrapper_133_clock),
    .reset(RetimeWrapper_133_reset),
    .io_flow(RetimeWrapper_133_io_flow),
    .io_in(RetimeWrapper_133_io_in),
    .io_out(RetimeWrapper_133_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_134 ( // @[package.scala 93:22:@24764.4]
    .clock(RetimeWrapper_134_clock),
    .reset(RetimeWrapper_134_reset),
    .io_flow(RetimeWrapper_134_io_flow),
    .io_in(RetimeWrapper_134_io_in),
    .io_out(RetimeWrapper_134_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_135 ( // @[package.scala 93:22:@24772.4]
    .clock(RetimeWrapper_135_clock),
    .reset(RetimeWrapper_135_reset),
    .io_flow(RetimeWrapper_135_io_flow),
    .io_in(RetimeWrapper_135_io_in),
    .io_out(RetimeWrapper_135_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_136 ( // @[package.scala 93:22:@24780.4]
    .clock(RetimeWrapper_136_clock),
    .reset(RetimeWrapper_136_reset),
    .io_flow(RetimeWrapper_136_io_flow),
    .io_in(RetimeWrapper_136_io_in),
    .io_out(RetimeWrapper_136_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_137 ( // @[package.scala 93:22:@24788.4]
    .clock(RetimeWrapper_137_clock),
    .reset(RetimeWrapper_137_reset),
    .io_flow(RetimeWrapper_137_io_flow),
    .io_in(RetimeWrapper_137_io_in),
    .io_out(RetimeWrapper_137_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_138 ( // @[package.scala 93:22:@24796.4]
    .clock(RetimeWrapper_138_clock),
    .reset(RetimeWrapper_138_reset),
    .io_flow(RetimeWrapper_138_io_flow),
    .io_in(RetimeWrapper_138_io_in),
    .io_out(RetimeWrapper_138_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_139 ( // @[package.scala 93:22:@24804.4]
    .clock(RetimeWrapper_139_clock),
    .reset(RetimeWrapper_139_reset),
    .io_flow(RetimeWrapper_139_io_flow),
    .io_in(RetimeWrapper_139_io_in),
    .io_out(RetimeWrapper_139_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_140 ( // @[package.scala 93:22:@24812.4]
    .clock(RetimeWrapper_140_clock),
    .reset(RetimeWrapper_140_reset),
    .io_flow(RetimeWrapper_140_io_flow),
    .io_in(RetimeWrapper_140_io_in),
    .io_out(RetimeWrapper_140_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_141 ( // @[package.scala 93:22:@24820.4]
    .clock(RetimeWrapper_141_clock),
    .reset(RetimeWrapper_141_reset),
    .io_flow(RetimeWrapper_141_io_flow),
    .io_in(RetimeWrapper_141_io_in),
    .io_out(RetimeWrapper_141_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_142 ( // @[package.scala 93:22:@24828.4]
    .clock(RetimeWrapper_142_clock),
    .reset(RetimeWrapper_142_reset),
    .io_flow(RetimeWrapper_142_io_flow),
    .io_in(RetimeWrapper_142_io_in),
    .io_out(RetimeWrapper_142_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_143 ( // @[package.scala 93:22:@24836.4]
    .clock(RetimeWrapper_143_clock),
    .reset(RetimeWrapper_143_reset),
    .io_flow(RetimeWrapper_143_io_flow),
    .io_in(RetimeWrapper_143_io_in),
    .io_out(RetimeWrapper_143_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_144 ( // @[package.scala 93:22:@24892.4]
    .clock(RetimeWrapper_144_clock),
    .reset(RetimeWrapper_144_reset),
    .io_flow(RetimeWrapper_144_io_flow),
    .io_in(RetimeWrapper_144_io_in),
    .io_out(RetimeWrapper_144_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_145 ( // @[package.scala 93:22:@24900.4]
    .clock(RetimeWrapper_145_clock),
    .reset(RetimeWrapper_145_reset),
    .io_flow(RetimeWrapper_145_io_flow),
    .io_in(RetimeWrapper_145_io_in),
    .io_out(RetimeWrapper_145_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_146 ( // @[package.scala 93:22:@24908.4]
    .clock(RetimeWrapper_146_clock),
    .reset(RetimeWrapper_146_reset),
    .io_flow(RetimeWrapper_146_io_flow),
    .io_in(RetimeWrapper_146_io_in),
    .io_out(RetimeWrapper_146_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_147 ( // @[package.scala 93:22:@24916.4]
    .clock(RetimeWrapper_147_clock),
    .reset(RetimeWrapper_147_reset),
    .io_flow(RetimeWrapper_147_io_flow),
    .io_in(RetimeWrapper_147_io_in),
    .io_out(RetimeWrapper_147_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_148 ( // @[package.scala 93:22:@24924.4]
    .clock(RetimeWrapper_148_clock),
    .reset(RetimeWrapper_148_reset),
    .io_flow(RetimeWrapper_148_io_flow),
    .io_in(RetimeWrapper_148_io_in),
    .io_out(RetimeWrapper_148_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_149 ( // @[package.scala 93:22:@24932.4]
    .clock(RetimeWrapper_149_clock),
    .reset(RetimeWrapper_149_reset),
    .io_flow(RetimeWrapper_149_io_flow),
    .io_in(RetimeWrapper_149_io_in),
    .io_out(RetimeWrapper_149_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_150 ( // @[package.scala 93:22:@24940.4]
    .clock(RetimeWrapper_150_clock),
    .reset(RetimeWrapper_150_reset),
    .io_flow(RetimeWrapper_150_io_flow),
    .io_in(RetimeWrapper_150_io_in),
    .io_out(RetimeWrapper_150_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_151 ( // @[package.scala 93:22:@24948.4]
    .clock(RetimeWrapper_151_clock),
    .reset(RetimeWrapper_151_reset),
    .io_flow(RetimeWrapper_151_io_flow),
    .io_in(RetimeWrapper_151_io_in),
    .io_out(RetimeWrapper_151_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_152 ( // @[package.scala 93:22:@24956.4]
    .clock(RetimeWrapper_152_clock),
    .reset(RetimeWrapper_152_reset),
    .io_flow(RetimeWrapper_152_io_flow),
    .io_in(RetimeWrapper_152_io_in),
    .io_out(RetimeWrapper_152_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_153 ( // @[package.scala 93:22:@24964.4]
    .clock(RetimeWrapper_153_clock),
    .reset(RetimeWrapper_153_reset),
    .io_flow(RetimeWrapper_153_io_flow),
    .io_in(RetimeWrapper_153_io_in),
    .io_out(RetimeWrapper_153_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_154 ( // @[package.scala 93:22:@24972.4]
    .clock(RetimeWrapper_154_clock),
    .reset(RetimeWrapper_154_reset),
    .io_flow(RetimeWrapper_154_io_flow),
    .io_in(RetimeWrapper_154_io_in),
    .io_out(RetimeWrapper_154_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_155 ( // @[package.scala 93:22:@24980.4]
    .clock(RetimeWrapper_155_clock),
    .reset(RetimeWrapper_155_reset),
    .io_flow(RetimeWrapper_155_io_flow),
    .io_in(RetimeWrapper_155_io_in),
    .io_out(RetimeWrapper_155_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_156 ( // @[package.scala 93:22:@25036.4]
    .clock(RetimeWrapper_156_clock),
    .reset(RetimeWrapper_156_reset),
    .io_flow(RetimeWrapper_156_io_flow),
    .io_in(RetimeWrapper_156_io_in),
    .io_out(RetimeWrapper_156_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_157 ( // @[package.scala 93:22:@25044.4]
    .clock(RetimeWrapper_157_clock),
    .reset(RetimeWrapper_157_reset),
    .io_flow(RetimeWrapper_157_io_flow),
    .io_in(RetimeWrapper_157_io_in),
    .io_out(RetimeWrapper_157_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_158 ( // @[package.scala 93:22:@25052.4]
    .clock(RetimeWrapper_158_clock),
    .reset(RetimeWrapper_158_reset),
    .io_flow(RetimeWrapper_158_io_flow),
    .io_in(RetimeWrapper_158_io_in),
    .io_out(RetimeWrapper_158_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_159 ( // @[package.scala 93:22:@25060.4]
    .clock(RetimeWrapper_159_clock),
    .reset(RetimeWrapper_159_reset),
    .io_flow(RetimeWrapper_159_io_flow),
    .io_in(RetimeWrapper_159_io_in),
    .io_out(RetimeWrapper_159_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_160 ( // @[package.scala 93:22:@25068.4]
    .clock(RetimeWrapper_160_clock),
    .reset(RetimeWrapper_160_reset),
    .io_flow(RetimeWrapper_160_io_flow),
    .io_in(RetimeWrapper_160_io_in),
    .io_out(RetimeWrapper_160_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_161 ( // @[package.scala 93:22:@25076.4]
    .clock(RetimeWrapper_161_clock),
    .reset(RetimeWrapper_161_reset),
    .io_flow(RetimeWrapper_161_io_flow),
    .io_in(RetimeWrapper_161_io_in),
    .io_out(RetimeWrapper_161_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_162 ( // @[package.scala 93:22:@25084.4]
    .clock(RetimeWrapper_162_clock),
    .reset(RetimeWrapper_162_reset),
    .io_flow(RetimeWrapper_162_io_flow),
    .io_in(RetimeWrapper_162_io_in),
    .io_out(RetimeWrapper_162_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_163 ( // @[package.scala 93:22:@25092.4]
    .clock(RetimeWrapper_163_clock),
    .reset(RetimeWrapper_163_reset),
    .io_flow(RetimeWrapper_163_io_flow),
    .io_in(RetimeWrapper_163_io_in),
    .io_out(RetimeWrapper_163_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_164 ( // @[package.scala 93:22:@25100.4]
    .clock(RetimeWrapper_164_clock),
    .reset(RetimeWrapper_164_reset),
    .io_flow(RetimeWrapper_164_io_flow),
    .io_in(RetimeWrapper_164_io_in),
    .io_out(RetimeWrapper_164_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_165 ( // @[package.scala 93:22:@25108.4]
    .clock(RetimeWrapper_165_clock),
    .reset(RetimeWrapper_165_reset),
    .io_flow(RetimeWrapper_165_io_flow),
    .io_in(RetimeWrapper_165_io_in),
    .io_out(RetimeWrapper_165_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_166 ( // @[package.scala 93:22:@25116.4]
    .clock(RetimeWrapper_166_clock),
    .reset(RetimeWrapper_166_reset),
    .io_flow(RetimeWrapper_166_io_flow),
    .io_in(RetimeWrapper_166_io_in),
    .io_out(RetimeWrapper_166_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_167 ( // @[package.scala 93:22:@25124.4]
    .clock(RetimeWrapper_167_clock),
    .reset(RetimeWrapper_167_reset),
    .io_flow(RetimeWrapper_167_io_flow),
    .io_in(RetimeWrapper_167_io_in),
    .io_out(RetimeWrapper_167_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_168 ( // @[package.scala 93:22:@25180.4]
    .clock(RetimeWrapper_168_clock),
    .reset(RetimeWrapper_168_reset),
    .io_flow(RetimeWrapper_168_io_flow),
    .io_in(RetimeWrapper_168_io_in),
    .io_out(RetimeWrapper_168_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_169 ( // @[package.scala 93:22:@25188.4]
    .clock(RetimeWrapper_169_clock),
    .reset(RetimeWrapper_169_reset),
    .io_flow(RetimeWrapper_169_io_flow),
    .io_in(RetimeWrapper_169_io_in),
    .io_out(RetimeWrapper_169_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_170 ( // @[package.scala 93:22:@25196.4]
    .clock(RetimeWrapper_170_clock),
    .reset(RetimeWrapper_170_reset),
    .io_flow(RetimeWrapper_170_io_flow),
    .io_in(RetimeWrapper_170_io_in),
    .io_out(RetimeWrapper_170_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_171 ( // @[package.scala 93:22:@25204.4]
    .clock(RetimeWrapper_171_clock),
    .reset(RetimeWrapper_171_reset),
    .io_flow(RetimeWrapper_171_io_flow),
    .io_in(RetimeWrapper_171_io_in),
    .io_out(RetimeWrapper_171_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_172 ( // @[package.scala 93:22:@25212.4]
    .clock(RetimeWrapper_172_clock),
    .reset(RetimeWrapper_172_reset),
    .io_flow(RetimeWrapper_172_io_flow),
    .io_in(RetimeWrapper_172_io_in),
    .io_out(RetimeWrapper_172_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_173 ( // @[package.scala 93:22:@25220.4]
    .clock(RetimeWrapper_173_clock),
    .reset(RetimeWrapper_173_reset),
    .io_flow(RetimeWrapper_173_io_flow),
    .io_in(RetimeWrapper_173_io_in),
    .io_out(RetimeWrapper_173_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_174 ( // @[package.scala 93:22:@25228.4]
    .clock(RetimeWrapper_174_clock),
    .reset(RetimeWrapper_174_reset),
    .io_flow(RetimeWrapper_174_io_flow),
    .io_in(RetimeWrapper_174_io_in),
    .io_out(RetimeWrapper_174_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_175 ( // @[package.scala 93:22:@25236.4]
    .clock(RetimeWrapper_175_clock),
    .reset(RetimeWrapper_175_reset),
    .io_flow(RetimeWrapper_175_io_flow),
    .io_in(RetimeWrapper_175_io_in),
    .io_out(RetimeWrapper_175_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_176 ( // @[package.scala 93:22:@25244.4]
    .clock(RetimeWrapper_176_clock),
    .reset(RetimeWrapper_176_reset),
    .io_flow(RetimeWrapper_176_io_flow),
    .io_in(RetimeWrapper_176_io_in),
    .io_out(RetimeWrapper_176_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_177 ( // @[package.scala 93:22:@25252.4]
    .clock(RetimeWrapper_177_clock),
    .reset(RetimeWrapper_177_reset),
    .io_flow(RetimeWrapper_177_io_flow),
    .io_in(RetimeWrapper_177_io_in),
    .io_out(RetimeWrapper_177_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_178 ( // @[package.scala 93:22:@25260.4]
    .clock(RetimeWrapper_178_clock),
    .reset(RetimeWrapper_178_reset),
    .io_flow(RetimeWrapper_178_io_flow),
    .io_in(RetimeWrapper_178_io_in),
    .io_out(RetimeWrapper_178_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_179 ( // @[package.scala 93:22:@25268.4]
    .clock(RetimeWrapper_179_clock),
    .reset(RetimeWrapper_179_reset),
    .io_flow(RetimeWrapper_179_io_flow),
    .io_in(RetimeWrapper_179_io_in),
    .io_out(RetimeWrapper_179_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_180 ( // @[package.scala 93:22:@25324.4]
    .clock(RetimeWrapper_180_clock),
    .reset(RetimeWrapper_180_reset),
    .io_flow(RetimeWrapper_180_io_flow),
    .io_in(RetimeWrapper_180_io_in),
    .io_out(RetimeWrapper_180_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_181 ( // @[package.scala 93:22:@25332.4]
    .clock(RetimeWrapper_181_clock),
    .reset(RetimeWrapper_181_reset),
    .io_flow(RetimeWrapper_181_io_flow),
    .io_in(RetimeWrapper_181_io_in),
    .io_out(RetimeWrapper_181_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_182 ( // @[package.scala 93:22:@25340.4]
    .clock(RetimeWrapper_182_clock),
    .reset(RetimeWrapper_182_reset),
    .io_flow(RetimeWrapper_182_io_flow),
    .io_in(RetimeWrapper_182_io_in),
    .io_out(RetimeWrapper_182_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_183 ( // @[package.scala 93:22:@25348.4]
    .clock(RetimeWrapper_183_clock),
    .reset(RetimeWrapper_183_reset),
    .io_flow(RetimeWrapper_183_io_flow),
    .io_in(RetimeWrapper_183_io_in),
    .io_out(RetimeWrapper_183_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_184 ( // @[package.scala 93:22:@25356.4]
    .clock(RetimeWrapper_184_clock),
    .reset(RetimeWrapper_184_reset),
    .io_flow(RetimeWrapper_184_io_flow),
    .io_in(RetimeWrapper_184_io_in),
    .io_out(RetimeWrapper_184_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_185 ( // @[package.scala 93:22:@25364.4]
    .clock(RetimeWrapper_185_clock),
    .reset(RetimeWrapper_185_reset),
    .io_flow(RetimeWrapper_185_io_flow),
    .io_in(RetimeWrapper_185_io_in),
    .io_out(RetimeWrapper_185_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_186 ( // @[package.scala 93:22:@25372.4]
    .clock(RetimeWrapper_186_clock),
    .reset(RetimeWrapper_186_reset),
    .io_flow(RetimeWrapper_186_io_flow),
    .io_in(RetimeWrapper_186_io_in),
    .io_out(RetimeWrapper_186_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_187 ( // @[package.scala 93:22:@25380.4]
    .clock(RetimeWrapper_187_clock),
    .reset(RetimeWrapper_187_reset),
    .io_flow(RetimeWrapper_187_io_flow),
    .io_in(RetimeWrapper_187_io_in),
    .io_out(RetimeWrapper_187_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_188 ( // @[package.scala 93:22:@25388.4]
    .clock(RetimeWrapper_188_clock),
    .reset(RetimeWrapper_188_reset),
    .io_flow(RetimeWrapper_188_io_flow),
    .io_in(RetimeWrapper_188_io_in),
    .io_out(RetimeWrapper_188_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_189 ( // @[package.scala 93:22:@25396.4]
    .clock(RetimeWrapper_189_clock),
    .reset(RetimeWrapper_189_reset),
    .io_flow(RetimeWrapper_189_io_flow),
    .io_in(RetimeWrapper_189_io_in),
    .io_out(RetimeWrapper_189_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_190 ( // @[package.scala 93:22:@25404.4]
    .clock(RetimeWrapper_190_clock),
    .reset(RetimeWrapper_190_reset),
    .io_flow(RetimeWrapper_190_io_flow),
    .io_in(RetimeWrapper_190_io_in),
    .io_out(RetimeWrapper_190_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_191 ( // @[package.scala 93:22:@25412.4]
    .clock(RetimeWrapper_191_clock),
    .reset(RetimeWrapper_191_reset),
    .io_flow(RetimeWrapper_191_io_flow),
    .io_in(RetimeWrapper_191_io_in),
    .io_out(RetimeWrapper_191_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_192 ( // @[package.scala 93:22:@25468.4]
    .clock(RetimeWrapper_192_clock),
    .reset(RetimeWrapper_192_reset),
    .io_flow(RetimeWrapper_192_io_flow),
    .io_in(RetimeWrapper_192_io_in),
    .io_out(RetimeWrapper_192_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_193 ( // @[package.scala 93:22:@25476.4]
    .clock(RetimeWrapper_193_clock),
    .reset(RetimeWrapper_193_reset),
    .io_flow(RetimeWrapper_193_io_flow),
    .io_in(RetimeWrapper_193_io_in),
    .io_out(RetimeWrapper_193_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_194 ( // @[package.scala 93:22:@25484.4]
    .clock(RetimeWrapper_194_clock),
    .reset(RetimeWrapper_194_reset),
    .io_flow(RetimeWrapper_194_io_flow),
    .io_in(RetimeWrapper_194_io_in),
    .io_out(RetimeWrapper_194_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_195 ( // @[package.scala 93:22:@25492.4]
    .clock(RetimeWrapper_195_clock),
    .reset(RetimeWrapper_195_reset),
    .io_flow(RetimeWrapper_195_io_flow),
    .io_in(RetimeWrapper_195_io_in),
    .io_out(RetimeWrapper_195_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_196 ( // @[package.scala 93:22:@25500.4]
    .clock(RetimeWrapper_196_clock),
    .reset(RetimeWrapper_196_reset),
    .io_flow(RetimeWrapper_196_io_flow),
    .io_in(RetimeWrapper_196_io_in),
    .io_out(RetimeWrapper_196_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_197 ( // @[package.scala 93:22:@25508.4]
    .clock(RetimeWrapper_197_clock),
    .reset(RetimeWrapper_197_reset),
    .io_flow(RetimeWrapper_197_io_flow),
    .io_in(RetimeWrapper_197_io_in),
    .io_out(RetimeWrapper_197_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_198 ( // @[package.scala 93:22:@25516.4]
    .clock(RetimeWrapper_198_clock),
    .reset(RetimeWrapper_198_reset),
    .io_flow(RetimeWrapper_198_io_flow),
    .io_in(RetimeWrapper_198_io_in),
    .io_out(RetimeWrapper_198_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_199 ( // @[package.scala 93:22:@25524.4]
    .clock(RetimeWrapper_199_clock),
    .reset(RetimeWrapper_199_reset),
    .io_flow(RetimeWrapper_199_io_flow),
    .io_in(RetimeWrapper_199_io_in),
    .io_out(RetimeWrapper_199_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_200 ( // @[package.scala 93:22:@25532.4]
    .clock(RetimeWrapper_200_clock),
    .reset(RetimeWrapper_200_reset),
    .io_flow(RetimeWrapper_200_io_flow),
    .io_in(RetimeWrapper_200_io_in),
    .io_out(RetimeWrapper_200_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_201 ( // @[package.scala 93:22:@25540.4]
    .clock(RetimeWrapper_201_clock),
    .reset(RetimeWrapper_201_reset),
    .io_flow(RetimeWrapper_201_io_flow),
    .io_in(RetimeWrapper_201_io_in),
    .io_out(RetimeWrapper_201_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_202 ( // @[package.scala 93:22:@25548.4]
    .clock(RetimeWrapper_202_clock),
    .reset(RetimeWrapper_202_reset),
    .io_flow(RetimeWrapper_202_io_flow),
    .io_in(RetimeWrapper_202_io_in),
    .io_out(RetimeWrapper_202_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_203 ( // @[package.scala 93:22:@25556.4]
    .clock(RetimeWrapper_203_clock),
    .reset(RetimeWrapper_203_reset),
    .io_flow(RetimeWrapper_203_io_flow),
    .io_in(RetimeWrapper_203_io_in),
    .io_out(RetimeWrapper_203_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_204 ( // @[package.scala 93:22:@25612.4]
    .clock(RetimeWrapper_204_clock),
    .reset(RetimeWrapper_204_reset),
    .io_flow(RetimeWrapper_204_io_flow),
    .io_in(RetimeWrapper_204_io_in),
    .io_out(RetimeWrapper_204_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_205 ( // @[package.scala 93:22:@25620.4]
    .clock(RetimeWrapper_205_clock),
    .reset(RetimeWrapper_205_reset),
    .io_flow(RetimeWrapper_205_io_flow),
    .io_in(RetimeWrapper_205_io_in),
    .io_out(RetimeWrapper_205_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_206 ( // @[package.scala 93:22:@25628.4]
    .clock(RetimeWrapper_206_clock),
    .reset(RetimeWrapper_206_reset),
    .io_flow(RetimeWrapper_206_io_flow),
    .io_in(RetimeWrapper_206_io_in),
    .io_out(RetimeWrapper_206_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_207 ( // @[package.scala 93:22:@25636.4]
    .clock(RetimeWrapper_207_clock),
    .reset(RetimeWrapper_207_reset),
    .io_flow(RetimeWrapper_207_io_flow),
    .io_in(RetimeWrapper_207_io_in),
    .io_out(RetimeWrapper_207_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_208 ( // @[package.scala 93:22:@25644.4]
    .clock(RetimeWrapper_208_clock),
    .reset(RetimeWrapper_208_reset),
    .io_flow(RetimeWrapper_208_io_flow),
    .io_in(RetimeWrapper_208_io_in),
    .io_out(RetimeWrapper_208_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_209 ( // @[package.scala 93:22:@25652.4]
    .clock(RetimeWrapper_209_clock),
    .reset(RetimeWrapper_209_reset),
    .io_flow(RetimeWrapper_209_io_flow),
    .io_in(RetimeWrapper_209_io_in),
    .io_out(RetimeWrapper_209_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_210 ( // @[package.scala 93:22:@25660.4]
    .clock(RetimeWrapper_210_clock),
    .reset(RetimeWrapper_210_reset),
    .io_flow(RetimeWrapper_210_io_flow),
    .io_in(RetimeWrapper_210_io_in),
    .io_out(RetimeWrapper_210_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_211 ( // @[package.scala 93:22:@25668.4]
    .clock(RetimeWrapper_211_clock),
    .reset(RetimeWrapper_211_reset),
    .io_flow(RetimeWrapper_211_io_flow),
    .io_in(RetimeWrapper_211_io_in),
    .io_out(RetimeWrapper_211_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_212 ( // @[package.scala 93:22:@25676.4]
    .clock(RetimeWrapper_212_clock),
    .reset(RetimeWrapper_212_reset),
    .io_flow(RetimeWrapper_212_io_flow),
    .io_in(RetimeWrapper_212_io_in),
    .io_out(RetimeWrapper_212_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_213 ( // @[package.scala 93:22:@25684.4]
    .clock(RetimeWrapper_213_clock),
    .reset(RetimeWrapper_213_reset),
    .io_flow(RetimeWrapper_213_io_flow),
    .io_in(RetimeWrapper_213_io_in),
    .io_out(RetimeWrapper_213_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_214 ( // @[package.scala 93:22:@25692.4]
    .clock(RetimeWrapper_214_clock),
    .reset(RetimeWrapper_214_reset),
    .io_flow(RetimeWrapper_214_io_flow),
    .io_in(RetimeWrapper_214_io_in),
    .io_out(RetimeWrapper_214_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_215 ( // @[package.scala 93:22:@25700.4]
    .clock(RetimeWrapper_215_clock),
    .reset(RetimeWrapper_215_reset),
    .io_flow(RetimeWrapper_215_io_flow),
    .io_in(RetimeWrapper_215_io_in),
    .io_out(RetimeWrapper_215_io_out)
  );
  assign _T_700 = io_wPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@20535.4]
  assign _T_702 = io_wPort_0_banks_1 == 3'h0; // @[MemPrimitives.scala 82:210:@20536.4]
  assign _T_703 = _T_700 & _T_702; // @[MemPrimitives.scala 82:228:@20537.4]
  assign _T_704 = io_wPort_0_en_0 & _T_703; // @[MemPrimitives.scala 83:102:@20538.4]
  assign _T_706 = io_wPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@20539.4]
  assign _T_708 = io_wPort_2_banks_1 == 3'h0; // @[MemPrimitives.scala 82:210:@20540.4]
  assign _T_709 = _T_706 & _T_708; // @[MemPrimitives.scala 82:228:@20541.4]
  assign _T_710 = io_wPort_2_en_0 & _T_709; // @[MemPrimitives.scala 83:102:@20542.4]
  assign _T_712 = {_T_704,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@20544.4]
  assign _T_714 = {_T_710,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@20546.4]
  assign _T_715 = _T_704 ? _T_712 : _T_714; // @[Mux.scala 31:69:@20547.4]
  assign _T_720 = io_wPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@20554.4]
  assign _T_722 = io_wPort_1_banks_1 == 3'h1; // @[MemPrimitives.scala 82:210:@20555.4]
  assign _T_723 = _T_720 & _T_722; // @[MemPrimitives.scala 82:228:@20556.4]
  assign _T_724 = io_wPort_1_en_0 & _T_723; // @[MemPrimitives.scala 83:102:@20557.4]
  assign _T_726 = io_wPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@20558.4]
  assign _T_728 = io_wPort_3_banks_1 == 3'h1; // @[MemPrimitives.scala 82:210:@20559.4]
  assign _T_729 = _T_726 & _T_728; // @[MemPrimitives.scala 82:228:@20560.4]
  assign _T_730 = io_wPort_3_en_0 & _T_729; // @[MemPrimitives.scala 83:102:@20561.4]
  assign _T_732 = {_T_724,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@20563.4]
  assign _T_734 = {_T_730,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@20565.4]
  assign _T_735 = _T_724 ? _T_732 : _T_734; // @[Mux.scala 31:69:@20566.4]
  assign _T_742 = io_wPort_0_banks_1 == 3'h2; // @[MemPrimitives.scala 82:210:@20574.4]
  assign _T_743 = _T_700 & _T_742; // @[MemPrimitives.scala 82:228:@20575.4]
  assign _T_744 = io_wPort_0_en_0 & _T_743; // @[MemPrimitives.scala 83:102:@20576.4]
  assign _T_748 = io_wPort_2_banks_1 == 3'h2; // @[MemPrimitives.scala 82:210:@20578.4]
  assign _T_749 = _T_706 & _T_748; // @[MemPrimitives.scala 82:228:@20579.4]
  assign _T_750 = io_wPort_2_en_0 & _T_749; // @[MemPrimitives.scala 83:102:@20580.4]
  assign _T_752 = {_T_744,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@20582.4]
  assign _T_754 = {_T_750,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@20584.4]
  assign _T_755 = _T_744 ? _T_752 : _T_754; // @[Mux.scala 31:69:@20585.4]
  assign _T_762 = io_wPort_1_banks_1 == 3'h3; // @[MemPrimitives.scala 82:210:@20593.4]
  assign _T_763 = _T_720 & _T_762; // @[MemPrimitives.scala 82:228:@20594.4]
  assign _T_764 = io_wPort_1_en_0 & _T_763; // @[MemPrimitives.scala 83:102:@20595.4]
  assign _T_768 = io_wPort_3_banks_1 == 3'h3; // @[MemPrimitives.scala 82:210:@20597.4]
  assign _T_769 = _T_726 & _T_768; // @[MemPrimitives.scala 82:228:@20598.4]
  assign _T_770 = io_wPort_3_en_0 & _T_769; // @[MemPrimitives.scala 83:102:@20599.4]
  assign _T_772 = {_T_764,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@20601.4]
  assign _T_774 = {_T_770,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@20603.4]
  assign _T_775 = _T_764 ? _T_772 : _T_774; // @[Mux.scala 31:69:@20604.4]
  assign _T_782 = io_wPort_0_banks_1 == 3'h4; // @[MemPrimitives.scala 82:210:@20612.4]
  assign _T_783 = _T_700 & _T_782; // @[MemPrimitives.scala 82:228:@20613.4]
  assign _T_784 = io_wPort_0_en_0 & _T_783; // @[MemPrimitives.scala 83:102:@20614.4]
  assign _T_788 = io_wPort_2_banks_1 == 3'h4; // @[MemPrimitives.scala 82:210:@20616.4]
  assign _T_789 = _T_706 & _T_788; // @[MemPrimitives.scala 82:228:@20617.4]
  assign _T_790 = io_wPort_2_en_0 & _T_789; // @[MemPrimitives.scala 83:102:@20618.4]
  assign _T_792 = {_T_784,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@20620.4]
  assign _T_794 = {_T_790,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@20622.4]
  assign _T_795 = _T_784 ? _T_792 : _T_794; // @[Mux.scala 31:69:@20623.4]
  assign _T_802 = io_wPort_1_banks_1 == 3'h5; // @[MemPrimitives.scala 82:210:@20631.4]
  assign _T_803 = _T_720 & _T_802; // @[MemPrimitives.scala 82:228:@20632.4]
  assign _T_804 = io_wPort_1_en_0 & _T_803; // @[MemPrimitives.scala 83:102:@20633.4]
  assign _T_808 = io_wPort_3_banks_1 == 3'h5; // @[MemPrimitives.scala 82:210:@20635.4]
  assign _T_809 = _T_726 & _T_808; // @[MemPrimitives.scala 82:228:@20636.4]
  assign _T_810 = io_wPort_3_en_0 & _T_809; // @[MemPrimitives.scala 83:102:@20637.4]
  assign _T_812 = {_T_804,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@20639.4]
  assign _T_814 = {_T_810,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@20641.4]
  assign _T_815 = _T_804 ? _T_812 : _T_814; // @[Mux.scala 31:69:@20642.4]
  assign _T_820 = io_wPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@20649.4]
  assign _T_823 = _T_820 & _T_702; // @[MemPrimitives.scala 82:228:@20651.4]
  assign _T_824 = io_wPort_0_en_0 & _T_823; // @[MemPrimitives.scala 83:102:@20652.4]
  assign _T_826 = io_wPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@20653.4]
  assign _T_829 = _T_826 & _T_708; // @[MemPrimitives.scala 82:228:@20655.4]
  assign _T_830 = io_wPort_2_en_0 & _T_829; // @[MemPrimitives.scala 83:102:@20656.4]
  assign _T_832 = {_T_824,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@20658.4]
  assign _T_834 = {_T_830,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@20660.4]
  assign _T_835 = _T_824 ? _T_832 : _T_834; // @[Mux.scala 31:69:@20661.4]
  assign _T_840 = io_wPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@20668.4]
  assign _T_843 = _T_840 & _T_722; // @[MemPrimitives.scala 82:228:@20670.4]
  assign _T_844 = io_wPort_1_en_0 & _T_843; // @[MemPrimitives.scala 83:102:@20671.4]
  assign _T_846 = io_wPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@20672.4]
  assign _T_849 = _T_846 & _T_728; // @[MemPrimitives.scala 82:228:@20674.4]
  assign _T_850 = io_wPort_3_en_0 & _T_849; // @[MemPrimitives.scala 83:102:@20675.4]
  assign _T_852 = {_T_844,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@20677.4]
  assign _T_854 = {_T_850,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@20679.4]
  assign _T_855 = _T_844 ? _T_852 : _T_854; // @[Mux.scala 31:69:@20680.4]
  assign _T_863 = _T_820 & _T_742; // @[MemPrimitives.scala 82:228:@20689.4]
  assign _T_864 = io_wPort_0_en_0 & _T_863; // @[MemPrimitives.scala 83:102:@20690.4]
  assign _T_869 = _T_826 & _T_748; // @[MemPrimitives.scala 82:228:@20693.4]
  assign _T_870 = io_wPort_2_en_0 & _T_869; // @[MemPrimitives.scala 83:102:@20694.4]
  assign _T_872 = {_T_864,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@20696.4]
  assign _T_874 = {_T_870,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@20698.4]
  assign _T_875 = _T_864 ? _T_872 : _T_874; // @[Mux.scala 31:69:@20699.4]
  assign _T_883 = _T_840 & _T_762; // @[MemPrimitives.scala 82:228:@20708.4]
  assign _T_884 = io_wPort_1_en_0 & _T_883; // @[MemPrimitives.scala 83:102:@20709.4]
  assign _T_889 = _T_846 & _T_768; // @[MemPrimitives.scala 82:228:@20712.4]
  assign _T_890 = io_wPort_3_en_0 & _T_889; // @[MemPrimitives.scala 83:102:@20713.4]
  assign _T_892 = {_T_884,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@20715.4]
  assign _T_894 = {_T_890,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@20717.4]
  assign _T_895 = _T_884 ? _T_892 : _T_894; // @[Mux.scala 31:69:@20718.4]
  assign _T_903 = _T_820 & _T_782; // @[MemPrimitives.scala 82:228:@20727.4]
  assign _T_904 = io_wPort_0_en_0 & _T_903; // @[MemPrimitives.scala 83:102:@20728.4]
  assign _T_909 = _T_826 & _T_788; // @[MemPrimitives.scala 82:228:@20731.4]
  assign _T_910 = io_wPort_2_en_0 & _T_909; // @[MemPrimitives.scala 83:102:@20732.4]
  assign _T_912 = {_T_904,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@20734.4]
  assign _T_914 = {_T_910,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@20736.4]
  assign _T_915 = _T_904 ? _T_912 : _T_914; // @[Mux.scala 31:69:@20737.4]
  assign _T_923 = _T_840 & _T_802; // @[MemPrimitives.scala 82:228:@20746.4]
  assign _T_924 = io_wPort_1_en_0 & _T_923; // @[MemPrimitives.scala 83:102:@20747.4]
  assign _T_929 = _T_846 & _T_808; // @[MemPrimitives.scala 82:228:@20750.4]
  assign _T_930 = io_wPort_3_en_0 & _T_929; // @[MemPrimitives.scala 83:102:@20751.4]
  assign _T_932 = {_T_924,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@20753.4]
  assign _T_934 = {_T_930,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@20755.4]
  assign _T_935 = _T_924 ? _T_932 : _T_934; // @[Mux.scala 31:69:@20756.4]
  assign _T_940 = io_wPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@20763.4]
  assign _T_943 = _T_940 & _T_702; // @[MemPrimitives.scala 82:228:@20765.4]
  assign _T_944 = io_wPort_0_en_0 & _T_943; // @[MemPrimitives.scala 83:102:@20766.4]
  assign _T_946 = io_wPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@20767.4]
  assign _T_949 = _T_946 & _T_708; // @[MemPrimitives.scala 82:228:@20769.4]
  assign _T_950 = io_wPort_2_en_0 & _T_949; // @[MemPrimitives.scala 83:102:@20770.4]
  assign _T_952 = {_T_944,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@20772.4]
  assign _T_954 = {_T_950,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@20774.4]
  assign _T_955 = _T_944 ? _T_952 : _T_954; // @[Mux.scala 31:69:@20775.4]
  assign _T_960 = io_wPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@20782.4]
  assign _T_963 = _T_960 & _T_722; // @[MemPrimitives.scala 82:228:@20784.4]
  assign _T_964 = io_wPort_1_en_0 & _T_963; // @[MemPrimitives.scala 83:102:@20785.4]
  assign _T_966 = io_wPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@20786.4]
  assign _T_969 = _T_966 & _T_728; // @[MemPrimitives.scala 82:228:@20788.4]
  assign _T_970 = io_wPort_3_en_0 & _T_969; // @[MemPrimitives.scala 83:102:@20789.4]
  assign _T_972 = {_T_964,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@20791.4]
  assign _T_974 = {_T_970,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@20793.4]
  assign _T_975 = _T_964 ? _T_972 : _T_974; // @[Mux.scala 31:69:@20794.4]
  assign _T_983 = _T_940 & _T_742; // @[MemPrimitives.scala 82:228:@20803.4]
  assign _T_984 = io_wPort_0_en_0 & _T_983; // @[MemPrimitives.scala 83:102:@20804.4]
  assign _T_989 = _T_946 & _T_748; // @[MemPrimitives.scala 82:228:@20807.4]
  assign _T_990 = io_wPort_2_en_0 & _T_989; // @[MemPrimitives.scala 83:102:@20808.4]
  assign _T_992 = {_T_984,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@20810.4]
  assign _T_994 = {_T_990,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@20812.4]
  assign _T_995 = _T_984 ? _T_992 : _T_994; // @[Mux.scala 31:69:@20813.4]
  assign _T_1003 = _T_960 & _T_762; // @[MemPrimitives.scala 82:228:@20822.4]
  assign _T_1004 = io_wPort_1_en_0 & _T_1003; // @[MemPrimitives.scala 83:102:@20823.4]
  assign _T_1009 = _T_966 & _T_768; // @[MemPrimitives.scala 82:228:@20826.4]
  assign _T_1010 = io_wPort_3_en_0 & _T_1009; // @[MemPrimitives.scala 83:102:@20827.4]
  assign _T_1012 = {_T_1004,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@20829.4]
  assign _T_1014 = {_T_1010,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@20831.4]
  assign _T_1015 = _T_1004 ? _T_1012 : _T_1014; // @[Mux.scala 31:69:@20832.4]
  assign _T_1023 = _T_940 & _T_782; // @[MemPrimitives.scala 82:228:@20841.4]
  assign _T_1024 = io_wPort_0_en_0 & _T_1023; // @[MemPrimitives.scala 83:102:@20842.4]
  assign _T_1029 = _T_946 & _T_788; // @[MemPrimitives.scala 82:228:@20845.4]
  assign _T_1030 = io_wPort_2_en_0 & _T_1029; // @[MemPrimitives.scala 83:102:@20846.4]
  assign _T_1032 = {_T_1024,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@20848.4]
  assign _T_1034 = {_T_1030,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@20850.4]
  assign _T_1035 = _T_1024 ? _T_1032 : _T_1034; // @[Mux.scala 31:69:@20851.4]
  assign _T_1043 = _T_960 & _T_802; // @[MemPrimitives.scala 82:228:@20860.4]
  assign _T_1044 = io_wPort_1_en_0 & _T_1043; // @[MemPrimitives.scala 83:102:@20861.4]
  assign _T_1049 = _T_966 & _T_808; // @[MemPrimitives.scala 82:228:@20864.4]
  assign _T_1050 = io_wPort_3_en_0 & _T_1049; // @[MemPrimitives.scala 83:102:@20865.4]
  assign _T_1052 = {_T_1044,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@20867.4]
  assign _T_1054 = {_T_1050,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@20869.4]
  assign _T_1055 = _T_1044 ? _T_1052 : _T_1054; // @[Mux.scala 31:69:@20870.4]
  assign _T_1060 = io_wPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@20877.4]
  assign _T_1063 = _T_1060 & _T_702; // @[MemPrimitives.scala 82:228:@20879.4]
  assign _T_1064 = io_wPort_0_en_0 & _T_1063; // @[MemPrimitives.scala 83:102:@20880.4]
  assign _T_1066 = io_wPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@20881.4]
  assign _T_1069 = _T_1066 & _T_708; // @[MemPrimitives.scala 82:228:@20883.4]
  assign _T_1070 = io_wPort_2_en_0 & _T_1069; // @[MemPrimitives.scala 83:102:@20884.4]
  assign _T_1072 = {_T_1064,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@20886.4]
  assign _T_1074 = {_T_1070,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@20888.4]
  assign _T_1075 = _T_1064 ? _T_1072 : _T_1074; // @[Mux.scala 31:69:@20889.4]
  assign _T_1080 = io_wPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@20896.4]
  assign _T_1083 = _T_1080 & _T_722; // @[MemPrimitives.scala 82:228:@20898.4]
  assign _T_1084 = io_wPort_1_en_0 & _T_1083; // @[MemPrimitives.scala 83:102:@20899.4]
  assign _T_1086 = io_wPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@20900.4]
  assign _T_1089 = _T_1086 & _T_728; // @[MemPrimitives.scala 82:228:@20902.4]
  assign _T_1090 = io_wPort_3_en_0 & _T_1089; // @[MemPrimitives.scala 83:102:@20903.4]
  assign _T_1092 = {_T_1084,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@20905.4]
  assign _T_1094 = {_T_1090,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@20907.4]
  assign _T_1095 = _T_1084 ? _T_1092 : _T_1094; // @[Mux.scala 31:69:@20908.4]
  assign _T_1103 = _T_1060 & _T_742; // @[MemPrimitives.scala 82:228:@20917.4]
  assign _T_1104 = io_wPort_0_en_0 & _T_1103; // @[MemPrimitives.scala 83:102:@20918.4]
  assign _T_1109 = _T_1066 & _T_748; // @[MemPrimitives.scala 82:228:@20921.4]
  assign _T_1110 = io_wPort_2_en_0 & _T_1109; // @[MemPrimitives.scala 83:102:@20922.4]
  assign _T_1112 = {_T_1104,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@20924.4]
  assign _T_1114 = {_T_1110,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@20926.4]
  assign _T_1115 = _T_1104 ? _T_1112 : _T_1114; // @[Mux.scala 31:69:@20927.4]
  assign _T_1123 = _T_1080 & _T_762; // @[MemPrimitives.scala 82:228:@20936.4]
  assign _T_1124 = io_wPort_1_en_0 & _T_1123; // @[MemPrimitives.scala 83:102:@20937.4]
  assign _T_1129 = _T_1086 & _T_768; // @[MemPrimitives.scala 82:228:@20940.4]
  assign _T_1130 = io_wPort_3_en_0 & _T_1129; // @[MemPrimitives.scala 83:102:@20941.4]
  assign _T_1132 = {_T_1124,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@20943.4]
  assign _T_1134 = {_T_1130,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@20945.4]
  assign _T_1135 = _T_1124 ? _T_1132 : _T_1134; // @[Mux.scala 31:69:@20946.4]
  assign _T_1143 = _T_1060 & _T_782; // @[MemPrimitives.scala 82:228:@20955.4]
  assign _T_1144 = io_wPort_0_en_0 & _T_1143; // @[MemPrimitives.scala 83:102:@20956.4]
  assign _T_1149 = _T_1066 & _T_788; // @[MemPrimitives.scala 82:228:@20959.4]
  assign _T_1150 = io_wPort_2_en_0 & _T_1149; // @[MemPrimitives.scala 83:102:@20960.4]
  assign _T_1152 = {_T_1144,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@20962.4]
  assign _T_1154 = {_T_1150,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@20964.4]
  assign _T_1155 = _T_1144 ? _T_1152 : _T_1154; // @[Mux.scala 31:69:@20965.4]
  assign _T_1163 = _T_1080 & _T_802; // @[MemPrimitives.scala 82:228:@20974.4]
  assign _T_1164 = io_wPort_1_en_0 & _T_1163; // @[MemPrimitives.scala 83:102:@20975.4]
  assign _T_1169 = _T_1086 & _T_808; // @[MemPrimitives.scala 82:228:@20978.4]
  assign _T_1170 = io_wPort_3_en_0 & _T_1169; // @[MemPrimitives.scala 83:102:@20979.4]
  assign _T_1172 = {_T_1164,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@20981.4]
  assign _T_1174 = {_T_1170,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@20983.4]
  assign _T_1175 = _T_1164 ? _T_1172 : _T_1174; // @[Mux.scala 31:69:@20984.4]
  assign _T_1180 = io_rPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@20991.4]
  assign _T_1182 = io_rPort_0_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@20992.4]
  assign _T_1183 = _T_1180 & _T_1182; // @[MemPrimitives.scala 110:228:@20993.4]
  assign _T_1186 = io_rPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@20995.4]
  assign _T_1188 = io_rPort_2_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@20996.4]
  assign _T_1189 = _T_1186 & _T_1188; // @[MemPrimitives.scala 110:228:@20997.4]
  assign _T_1192 = io_rPort_4_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@20999.4]
  assign _T_1194 = io_rPort_4_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@21000.4]
  assign _T_1195 = _T_1192 & _T_1194; // @[MemPrimitives.scala 110:228:@21001.4]
  assign _T_1198 = io_rPort_7_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21003.4]
  assign _T_1200 = io_rPort_7_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@21004.4]
  assign _T_1201 = _T_1198 & _T_1200; // @[MemPrimitives.scala 110:228:@21005.4]
  assign _T_1204 = io_rPort_8_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21007.4]
  assign _T_1206 = io_rPort_8_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@21008.4]
  assign _T_1207 = _T_1204 & _T_1206; // @[MemPrimitives.scala 110:228:@21009.4]
  assign _T_1210 = io_rPort_10_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21011.4]
  assign _T_1212 = io_rPort_10_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@21012.4]
  assign _T_1213 = _T_1210 & _T_1212; // @[MemPrimitives.scala 110:228:@21013.4]
  assign _T_1216 = io_rPort_11_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21015.4]
  assign _T_1218 = io_rPort_11_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@21016.4]
  assign _T_1219 = _T_1216 & _T_1218; // @[MemPrimitives.scala 110:228:@21017.4]
  assign _T_1222 = io_rPort_15_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21019.4]
  assign _T_1224 = io_rPort_15_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@21020.4]
  assign _T_1225 = _T_1222 & _T_1224; // @[MemPrimitives.scala 110:228:@21021.4]
  assign _T_1228 = io_rPort_17_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21023.4]
  assign _T_1230 = io_rPort_17_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@21024.4]
  assign _T_1231 = _T_1228 & _T_1230; // @[MemPrimitives.scala 110:228:@21025.4]
  assign _T_1233 = StickySelects_io_outs_0; // @[MemPrimitives.scala 123:41:@21039.4]
  assign _T_1234 = StickySelects_io_outs_1; // @[MemPrimitives.scala 123:41:@21040.4]
  assign _T_1235 = StickySelects_io_outs_2; // @[MemPrimitives.scala 123:41:@21041.4]
  assign _T_1236 = StickySelects_io_outs_3; // @[MemPrimitives.scala 123:41:@21042.4]
  assign _T_1237 = StickySelects_io_outs_4; // @[MemPrimitives.scala 123:41:@21043.4]
  assign _T_1238 = StickySelects_io_outs_5; // @[MemPrimitives.scala 123:41:@21044.4]
  assign _T_1239 = StickySelects_io_outs_6; // @[MemPrimitives.scala 123:41:@21045.4]
  assign _T_1240 = StickySelects_io_outs_7; // @[MemPrimitives.scala 123:41:@21046.4]
  assign _T_1241 = StickySelects_io_outs_8; // @[MemPrimitives.scala 123:41:@21047.4]
  assign _T_1243 = {_T_1233,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@21049.4]
  assign _T_1245 = {_T_1234,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@21051.4]
  assign _T_1247 = {_T_1235,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@21053.4]
  assign _T_1249 = {_T_1236,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@21055.4]
  assign _T_1251 = {_T_1237,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@21057.4]
  assign _T_1253 = {_T_1238,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@21059.4]
  assign _T_1255 = {_T_1239,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@21061.4]
  assign _T_1257 = {_T_1240,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@21063.4]
  assign _T_1259 = {_T_1241,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@21065.4]
  assign _T_1260 = _T_1240 ? _T_1257 : _T_1259; // @[Mux.scala 31:69:@21066.4]
  assign _T_1261 = _T_1239 ? _T_1255 : _T_1260; // @[Mux.scala 31:69:@21067.4]
  assign _T_1262 = _T_1238 ? _T_1253 : _T_1261; // @[Mux.scala 31:69:@21068.4]
  assign _T_1263 = _T_1237 ? _T_1251 : _T_1262; // @[Mux.scala 31:69:@21069.4]
  assign _T_1264 = _T_1236 ? _T_1249 : _T_1263; // @[Mux.scala 31:69:@21070.4]
  assign _T_1265 = _T_1235 ? _T_1247 : _T_1264; // @[Mux.scala 31:69:@21071.4]
  assign _T_1266 = _T_1234 ? _T_1245 : _T_1265; // @[Mux.scala 31:69:@21072.4]
  assign _T_1267 = _T_1233 ? _T_1243 : _T_1266; // @[Mux.scala 31:69:@21073.4]
  assign _T_1272 = io_rPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21080.4]
  assign _T_1274 = io_rPort_1_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@21081.4]
  assign _T_1275 = _T_1272 & _T_1274; // @[MemPrimitives.scala 110:228:@21082.4]
  assign _T_1278 = io_rPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21084.4]
  assign _T_1280 = io_rPort_3_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@21085.4]
  assign _T_1281 = _T_1278 & _T_1280; // @[MemPrimitives.scala 110:228:@21086.4]
  assign _T_1284 = io_rPort_5_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21088.4]
  assign _T_1286 = io_rPort_5_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@21089.4]
  assign _T_1287 = _T_1284 & _T_1286; // @[MemPrimitives.scala 110:228:@21090.4]
  assign _T_1290 = io_rPort_6_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21092.4]
  assign _T_1292 = io_rPort_6_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@21093.4]
  assign _T_1293 = _T_1290 & _T_1292; // @[MemPrimitives.scala 110:228:@21094.4]
  assign _T_1296 = io_rPort_9_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21096.4]
  assign _T_1298 = io_rPort_9_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@21097.4]
  assign _T_1299 = _T_1296 & _T_1298; // @[MemPrimitives.scala 110:228:@21098.4]
  assign _T_1302 = io_rPort_12_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21100.4]
  assign _T_1304 = io_rPort_12_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@21101.4]
  assign _T_1305 = _T_1302 & _T_1304; // @[MemPrimitives.scala 110:228:@21102.4]
  assign _T_1308 = io_rPort_13_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21104.4]
  assign _T_1310 = io_rPort_13_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@21105.4]
  assign _T_1311 = _T_1308 & _T_1310; // @[MemPrimitives.scala 110:228:@21106.4]
  assign _T_1314 = io_rPort_14_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21108.4]
  assign _T_1316 = io_rPort_14_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@21109.4]
  assign _T_1317 = _T_1314 & _T_1316; // @[MemPrimitives.scala 110:228:@21110.4]
  assign _T_1320 = io_rPort_16_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21112.4]
  assign _T_1322 = io_rPort_16_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@21113.4]
  assign _T_1323 = _T_1320 & _T_1322; // @[MemPrimitives.scala 110:228:@21114.4]
  assign _T_1325 = StickySelects_1_io_outs_0; // @[MemPrimitives.scala 123:41:@21128.4]
  assign _T_1326 = StickySelects_1_io_outs_1; // @[MemPrimitives.scala 123:41:@21129.4]
  assign _T_1327 = StickySelects_1_io_outs_2; // @[MemPrimitives.scala 123:41:@21130.4]
  assign _T_1328 = StickySelects_1_io_outs_3; // @[MemPrimitives.scala 123:41:@21131.4]
  assign _T_1329 = StickySelects_1_io_outs_4; // @[MemPrimitives.scala 123:41:@21132.4]
  assign _T_1330 = StickySelects_1_io_outs_5; // @[MemPrimitives.scala 123:41:@21133.4]
  assign _T_1331 = StickySelects_1_io_outs_6; // @[MemPrimitives.scala 123:41:@21134.4]
  assign _T_1332 = StickySelects_1_io_outs_7; // @[MemPrimitives.scala 123:41:@21135.4]
  assign _T_1333 = StickySelects_1_io_outs_8; // @[MemPrimitives.scala 123:41:@21136.4]
  assign _T_1335 = {_T_1325,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@21138.4]
  assign _T_1337 = {_T_1326,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@21140.4]
  assign _T_1339 = {_T_1327,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@21142.4]
  assign _T_1341 = {_T_1328,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@21144.4]
  assign _T_1343 = {_T_1329,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@21146.4]
  assign _T_1345 = {_T_1330,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@21148.4]
  assign _T_1347 = {_T_1331,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@21150.4]
  assign _T_1349 = {_T_1332,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@21152.4]
  assign _T_1351 = {_T_1333,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@21154.4]
  assign _T_1352 = _T_1332 ? _T_1349 : _T_1351; // @[Mux.scala 31:69:@21155.4]
  assign _T_1353 = _T_1331 ? _T_1347 : _T_1352; // @[Mux.scala 31:69:@21156.4]
  assign _T_1354 = _T_1330 ? _T_1345 : _T_1353; // @[Mux.scala 31:69:@21157.4]
  assign _T_1355 = _T_1329 ? _T_1343 : _T_1354; // @[Mux.scala 31:69:@21158.4]
  assign _T_1356 = _T_1328 ? _T_1341 : _T_1355; // @[Mux.scala 31:69:@21159.4]
  assign _T_1357 = _T_1327 ? _T_1339 : _T_1356; // @[Mux.scala 31:69:@21160.4]
  assign _T_1358 = _T_1326 ? _T_1337 : _T_1357; // @[Mux.scala 31:69:@21161.4]
  assign _T_1359 = _T_1325 ? _T_1335 : _T_1358; // @[Mux.scala 31:69:@21162.4]
  assign _T_1366 = io_rPort_0_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@21170.4]
  assign _T_1367 = _T_1180 & _T_1366; // @[MemPrimitives.scala 110:228:@21171.4]
  assign _T_1372 = io_rPort_2_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@21174.4]
  assign _T_1373 = _T_1186 & _T_1372; // @[MemPrimitives.scala 110:228:@21175.4]
  assign _T_1378 = io_rPort_4_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@21178.4]
  assign _T_1379 = _T_1192 & _T_1378; // @[MemPrimitives.scala 110:228:@21179.4]
  assign _T_1384 = io_rPort_7_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@21182.4]
  assign _T_1385 = _T_1198 & _T_1384; // @[MemPrimitives.scala 110:228:@21183.4]
  assign _T_1390 = io_rPort_8_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@21186.4]
  assign _T_1391 = _T_1204 & _T_1390; // @[MemPrimitives.scala 110:228:@21187.4]
  assign _T_1396 = io_rPort_10_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@21190.4]
  assign _T_1397 = _T_1210 & _T_1396; // @[MemPrimitives.scala 110:228:@21191.4]
  assign _T_1402 = io_rPort_11_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@21194.4]
  assign _T_1403 = _T_1216 & _T_1402; // @[MemPrimitives.scala 110:228:@21195.4]
  assign _T_1408 = io_rPort_15_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@21198.4]
  assign _T_1409 = _T_1222 & _T_1408; // @[MemPrimitives.scala 110:228:@21199.4]
  assign _T_1414 = io_rPort_17_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@21202.4]
  assign _T_1415 = _T_1228 & _T_1414; // @[MemPrimitives.scala 110:228:@21203.4]
  assign _T_1417 = StickySelects_2_io_outs_0; // @[MemPrimitives.scala 123:41:@21217.4]
  assign _T_1418 = StickySelects_2_io_outs_1; // @[MemPrimitives.scala 123:41:@21218.4]
  assign _T_1419 = StickySelects_2_io_outs_2; // @[MemPrimitives.scala 123:41:@21219.4]
  assign _T_1420 = StickySelects_2_io_outs_3; // @[MemPrimitives.scala 123:41:@21220.4]
  assign _T_1421 = StickySelects_2_io_outs_4; // @[MemPrimitives.scala 123:41:@21221.4]
  assign _T_1422 = StickySelects_2_io_outs_5; // @[MemPrimitives.scala 123:41:@21222.4]
  assign _T_1423 = StickySelects_2_io_outs_6; // @[MemPrimitives.scala 123:41:@21223.4]
  assign _T_1424 = StickySelects_2_io_outs_7; // @[MemPrimitives.scala 123:41:@21224.4]
  assign _T_1425 = StickySelects_2_io_outs_8; // @[MemPrimitives.scala 123:41:@21225.4]
  assign _T_1427 = {_T_1417,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@21227.4]
  assign _T_1429 = {_T_1418,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@21229.4]
  assign _T_1431 = {_T_1419,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@21231.4]
  assign _T_1433 = {_T_1420,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@21233.4]
  assign _T_1435 = {_T_1421,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@21235.4]
  assign _T_1437 = {_T_1422,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@21237.4]
  assign _T_1439 = {_T_1423,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@21239.4]
  assign _T_1441 = {_T_1424,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@21241.4]
  assign _T_1443 = {_T_1425,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@21243.4]
  assign _T_1444 = _T_1424 ? _T_1441 : _T_1443; // @[Mux.scala 31:69:@21244.4]
  assign _T_1445 = _T_1423 ? _T_1439 : _T_1444; // @[Mux.scala 31:69:@21245.4]
  assign _T_1446 = _T_1422 ? _T_1437 : _T_1445; // @[Mux.scala 31:69:@21246.4]
  assign _T_1447 = _T_1421 ? _T_1435 : _T_1446; // @[Mux.scala 31:69:@21247.4]
  assign _T_1448 = _T_1420 ? _T_1433 : _T_1447; // @[Mux.scala 31:69:@21248.4]
  assign _T_1449 = _T_1419 ? _T_1431 : _T_1448; // @[Mux.scala 31:69:@21249.4]
  assign _T_1450 = _T_1418 ? _T_1429 : _T_1449; // @[Mux.scala 31:69:@21250.4]
  assign _T_1451 = _T_1417 ? _T_1427 : _T_1450; // @[Mux.scala 31:69:@21251.4]
  assign _T_1458 = io_rPort_1_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@21259.4]
  assign _T_1459 = _T_1272 & _T_1458; // @[MemPrimitives.scala 110:228:@21260.4]
  assign _T_1464 = io_rPort_3_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@21263.4]
  assign _T_1465 = _T_1278 & _T_1464; // @[MemPrimitives.scala 110:228:@21264.4]
  assign _T_1470 = io_rPort_5_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@21267.4]
  assign _T_1471 = _T_1284 & _T_1470; // @[MemPrimitives.scala 110:228:@21268.4]
  assign _T_1476 = io_rPort_6_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@21271.4]
  assign _T_1477 = _T_1290 & _T_1476; // @[MemPrimitives.scala 110:228:@21272.4]
  assign _T_1482 = io_rPort_9_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@21275.4]
  assign _T_1483 = _T_1296 & _T_1482; // @[MemPrimitives.scala 110:228:@21276.4]
  assign _T_1488 = io_rPort_12_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@21279.4]
  assign _T_1489 = _T_1302 & _T_1488; // @[MemPrimitives.scala 110:228:@21280.4]
  assign _T_1494 = io_rPort_13_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@21283.4]
  assign _T_1495 = _T_1308 & _T_1494; // @[MemPrimitives.scala 110:228:@21284.4]
  assign _T_1500 = io_rPort_14_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@21287.4]
  assign _T_1501 = _T_1314 & _T_1500; // @[MemPrimitives.scala 110:228:@21288.4]
  assign _T_1506 = io_rPort_16_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@21291.4]
  assign _T_1507 = _T_1320 & _T_1506; // @[MemPrimitives.scala 110:228:@21292.4]
  assign _T_1509 = StickySelects_3_io_outs_0; // @[MemPrimitives.scala 123:41:@21306.4]
  assign _T_1510 = StickySelects_3_io_outs_1; // @[MemPrimitives.scala 123:41:@21307.4]
  assign _T_1511 = StickySelects_3_io_outs_2; // @[MemPrimitives.scala 123:41:@21308.4]
  assign _T_1512 = StickySelects_3_io_outs_3; // @[MemPrimitives.scala 123:41:@21309.4]
  assign _T_1513 = StickySelects_3_io_outs_4; // @[MemPrimitives.scala 123:41:@21310.4]
  assign _T_1514 = StickySelects_3_io_outs_5; // @[MemPrimitives.scala 123:41:@21311.4]
  assign _T_1515 = StickySelects_3_io_outs_6; // @[MemPrimitives.scala 123:41:@21312.4]
  assign _T_1516 = StickySelects_3_io_outs_7; // @[MemPrimitives.scala 123:41:@21313.4]
  assign _T_1517 = StickySelects_3_io_outs_8; // @[MemPrimitives.scala 123:41:@21314.4]
  assign _T_1519 = {_T_1509,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@21316.4]
  assign _T_1521 = {_T_1510,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@21318.4]
  assign _T_1523 = {_T_1511,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@21320.4]
  assign _T_1525 = {_T_1512,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@21322.4]
  assign _T_1527 = {_T_1513,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@21324.4]
  assign _T_1529 = {_T_1514,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@21326.4]
  assign _T_1531 = {_T_1515,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@21328.4]
  assign _T_1533 = {_T_1516,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@21330.4]
  assign _T_1535 = {_T_1517,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@21332.4]
  assign _T_1536 = _T_1516 ? _T_1533 : _T_1535; // @[Mux.scala 31:69:@21333.4]
  assign _T_1537 = _T_1515 ? _T_1531 : _T_1536; // @[Mux.scala 31:69:@21334.4]
  assign _T_1538 = _T_1514 ? _T_1529 : _T_1537; // @[Mux.scala 31:69:@21335.4]
  assign _T_1539 = _T_1513 ? _T_1527 : _T_1538; // @[Mux.scala 31:69:@21336.4]
  assign _T_1540 = _T_1512 ? _T_1525 : _T_1539; // @[Mux.scala 31:69:@21337.4]
  assign _T_1541 = _T_1511 ? _T_1523 : _T_1540; // @[Mux.scala 31:69:@21338.4]
  assign _T_1542 = _T_1510 ? _T_1521 : _T_1541; // @[Mux.scala 31:69:@21339.4]
  assign _T_1543 = _T_1509 ? _T_1519 : _T_1542; // @[Mux.scala 31:69:@21340.4]
  assign _T_1550 = io_rPort_0_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@21348.4]
  assign _T_1551 = _T_1180 & _T_1550; // @[MemPrimitives.scala 110:228:@21349.4]
  assign _T_1556 = io_rPort_2_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@21352.4]
  assign _T_1557 = _T_1186 & _T_1556; // @[MemPrimitives.scala 110:228:@21353.4]
  assign _T_1562 = io_rPort_4_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@21356.4]
  assign _T_1563 = _T_1192 & _T_1562; // @[MemPrimitives.scala 110:228:@21357.4]
  assign _T_1568 = io_rPort_7_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@21360.4]
  assign _T_1569 = _T_1198 & _T_1568; // @[MemPrimitives.scala 110:228:@21361.4]
  assign _T_1574 = io_rPort_8_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@21364.4]
  assign _T_1575 = _T_1204 & _T_1574; // @[MemPrimitives.scala 110:228:@21365.4]
  assign _T_1580 = io_rPort_10_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@21368.4]
  assign _T_1581 = _T_1210 & _T_1580; // @[MemPrimitives.scala 110:228:@21369.4]
  assign _T_1586 = io_rPort_11_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@21372.4]
  assign _T_1587 = _T_1216 & _T_1586; // @[MemPrimitives.scala 110:228:@21373.4]
  assign _T_1592 = io_rPort_15_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@21376.4]
  assign _T_1593 = _T_1222 & _T_1592; // @[MemPrimitives.scala 110:228:@21377.4]
  assign _T_1598 = io_rPort_17_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@21380.4]
  assign _T_1599 = _T_1228 & _T_1598; // @[MemPrimitives.scala 110:228:@21381.4]
  assign _T_1601 = StickySelects_4_io_outs_0; // @[MemPrimitives.scala 123:41:@21395.4]
  assign _T_1602 = StickySelects_4_io_outs_1; // @[MemPrimitives.scala 123:41:@21396.4]
  assign _T_1603 = StickySelects_4_io_outs_2; // @[MemPrimitives.scala 123:41:@21397.4]
  assign _T_1604 = StickySelects_4_io_outs_3; // @[MemPrimitives.scala 123:41:@21398.4]
  assign _T_1605 = StickySelects_4_io_outs_4; // @[MemPrimitives.scala 123:41:@21399.4]
  assign _T_1606 = StickySelects_4_io_outs_5; // @[MemPrimitives.scala 123:41:@21400.4]
  assign _T_1607 = StickySelects_4_io_outs_6; // @[MemPrimitives.scala 123:41:@21401.4]
  assign _T_1608 = StickySelects_4_io_outs_7; // @[MemPrimitives.scala 123:41:@21402.4]
  assign _T_1609 = StickySelects_4_io_outs_8; // @[MemPrimitives.scala 123:41:@21403.4]
  assign _T_1611 = {_T_1601,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@21405.4]
  assign _T_1613 = {_T_1602,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@21407.4]
  assign _T_1615 = {_T_1603,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@21409.4]
  assign _T_1617 = {_T_1604,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@21411.4]
  assign _T_1619 = {_T_1605,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@21413.4]
  assign _T_1621 = {_T_1606,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@21415.4]
  assign _T_1623 = {_T_1607,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@21417.4]
  assign _T_1625 = {_T_1608,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@21419.4]
  assign _T_1627 = {_T_1609,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@21421.4]
  assign _T_1628 = _T_1608 ? _T_1625 : _T_1627; // @[Mux.scala 31:69:@21422.4]
  assign _T_1629 = _T_1607 ? _T_1623 : _T_1628; // @[Mux.scala 31:69:@21423.4]
  assign _T_1630 = _T_1606 ? _T_1621 : _T_1629; // @[Mux.scala 31:69:@21424.4]
  assign _T_1631 = _T_1605 ? _T_1619 : _T_1630; // @[Mux.scala 31:69:@21425.4]
  assign _T_1632 = _T_1604 ? _T_1617 : _T_1631; // @[Mux.scala 31:69:@21426.4]
  assign _T_1633 = _T_1603 ? _T_1615 : _T_1632; // @[Mux.scala 31:69:@21427.4]
  assign _T_1634 = _T_1602 ? _T_1613 : _T_1633; // @[Mux.scala 31:69:@21428.4]
  assign _T_1635 = _T_1601 ? _T_1611 : _T_1634; // @[Mux.scala 31:69:@21429.4]
  assign _T_1642 = io_rPort_1_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@21437.4]
  assign _T_1643 = _T_1272 & _T_1642; // @[MemPrimitives.scala 110:228:@21438.4]
  assign _T_1648 = io_rPort_3_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@21441.4]
  assign _T_1649 = _T_1278 & _T_1648; // @[MemPrimitives.scala 110:228:@21442.4]
  assign _T_1654 = io_rPort_5_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@21445.4]
  assign _T_1655 = _T_1284 & _T_1654; // @[MemPrimitives.scala 110:228:@21446.4]
  assign _T_1660 = io_rPort_6_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@21449.4]
  assign _T_1661 = _T_1290 & _T_1660; // @[MemPrimitives.scala 110:228:@21450.4]
  assign _T_1666 = io_rPort_9_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@21453.4]
  assign _T_1667 = _T_1296 & _T_1666; // @[MemPrimitives.scala 110:228:@21454.4]
  assign _T_1672 = io_rPort_12_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@21457.4]
  assign _T_1673 = _T_1302 & _T_1672; // @[MemPrimitives.scala 110:228:@21458.4]
  assign _T_1678 = io_rPort_13_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@21461.4]
  assign _T_1679 = _T_1308 & _T_1678; // @[MemPrimitives.scala 110:228:@21462.4]
  assign _T_1684 = io_rPort_14_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@21465.4]
  assign _T_1685 = _T_1314 & _T_1684; // @[MemPrimitives.scala 110:228:@21466.4]
  assign _T_1690 = io_rPort_16_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@21469.4]
  assign _T_1691 = _T_1320 & _T_1690; // @[MemPrimitives.scala 110:228:@21470.4]
  assign _T_1693 = StickySelects_5_io_outs_0; // @[MemPrimitives.scala 123:41:@21484.4]
  assign _T_1694 = StickySelects_5_io_outs_1; // @[MemPrimitives.scala 123:41:@21485.4]
  assign _T_1695 = StickySelects_5_io_outs_2; // @[MemPrimitives.scala 123:41:@21486.4]
  assign _T_1696 = StickySelects_5_io_outs_3; // @[MemPrimitives.scala 123:41:@21487.4]
  assign _T_1697 = StickySelects_5_io_outs_4; // @[MemPrimitives.scala 123:41:@21488.4]
  assign _T_1698 = StickySelects_5_io_outs_5; // @[MemPrimitives.scala 123:41:@21489.4]
  assign _T_1699 = StickySelects_5_io_outs_6; // @[MemPrimitives.scala 123:41:@21490.4]
  assign _T_1700 = StickySelects_5_io_outs_7; // @[MemPrimitives.scala 123:41:@21491.4]
  assign _T_1701 = StickySelects_5_io_outs_8; // @[MemPrimitives.scala 123:41:@21492.4]
  assign _T_1703 = {_T_1693,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@21494.4]
  assign _T_1705 = {_T_1694,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@21496.4]
  assign _T_1707 = {_T_1695,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@21498.4]
  assign _T_1709 = {_T_1696,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@21500.4]
  assign _T_1711 = {_T_1697,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@21502.4]
  assign _T_1713 = {_T_1698,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@21504.4]
  assign _T_1715 = {_T_1699,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@21506.4]
  assign _T_1717 = {_T_1700,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@21508.4]
  assign _T_1719 = {_T_1701,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@21510.4]
  assign _T_1720 = _T_1700 ? _T_1717 : _T_1719; // @[Mux.scala 31:69:@21511.4]
  assign _T_1721 = _T_1699 ? _T_1715 : _T_1720; // @[Mux.scala 31:69:@21512.4]
  assign _T_1722 = _T_1698 ? _T_1713 : _T_1721; // @[Mux.scala 31:69:@21513.4]
  assign _T_1723 = _T_1697 ? _T_1711 : _T_1722; // @[Mux.scala 31:69:@21514.4]
  assign _T_1724 = _T_1696 ? _T_1709 : _T_1723; // @[Mux.scala 31:69:@21515.4]
  assign _T_1725 = _T_1695 ? _T_1707 : _T_1724; // @[Mux.scala 31:69:@21516.4]
  assign _T_1726 = _T_1694 ? _T_1705 : _T_1725; // @[Mux.scala 31:69:@21517.4]
  assign _T_1727 = _T_1693 ? _T_1703 : _T_1726; // @[Mux.scala 31:69:@21518.4]
  assign _T_1732 = io_rPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21525.4]
  assign _T_1735 = _T_1732 & _T_1182; // @[MemPrimitives.scala 110:228:@21527.4]
  assign _T_1738 = io_rPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21529.4]
  assign _T_1741 = _T_1738 & _T_1188; // @[MemPrimitives.scala 110:228:@21531.4]
  assign _T_1744 = io_rPort_4_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21533.4]
  assign _T_1747 = _T_1744 & _T_1194; // @[MemPrimitives.scala 110:228:@21535.4]
  assign _T_1750 = io_rPort_7_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21537.4]
  assign _T_1753 = _T_1750 & _T_1200; // @[MemPrimitives.scala 110:228:@21539.4]
  assign _T_1756 = io_rPort_8_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21541.4]
  assign _T_1759 = _T_1756 & _T_1206; // @[MemPrimitives.scala 110:228:@21543.4]
  assign _T_1762 = io_rPort_10_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21545.4]
  assign _T_1765 = _T_1762 & _T_1212; // @[MemPrimitives.scala 110:228:@21547.4]
  assign _T_1768 = io_rPort_11_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21549.4]
  assign _T_1771 = _T_1768 & _T_1218; // @[MemPrimitives.scala 110:228:@21551.4]
  assign _T_1774 = io_rPort_15_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21553.4]
  assign _T_1777 = _T_1774 & _T_1224; // @[MemPrimitives.scala 110:228:@21555.4]
  assign _T_1780 = io_rPort_17_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21557.4]
  assign _T_1783 = _T_1780 & _T_1230; // @[MemPrimitives.scala 110:228:@21559.4]
  assign _T_1785 = StickySelects_6_io_outs_0; // @[MemPrimitives.scala 123:41:@21573.4]
  assign _T_1786 = StickySelects_6_io_outs_1; // @[MemPrimitives.scala 123:41:@21574.4]
  assign _T_1787 = StickySelects_6_io_outs_2; // @[MemPrimitives.scala 123:41:@21575.4]
  assign _T_1788 = StickySelects_6_io_outs_3; // @[MemPrimitives.scala 123:41:@21576.4]
  assign _T_1789 = StickySelects_6_io_outs_4; // @[MemPrimitives.scala 123:41:@21577.4]
  assign _T_1790 = StickySelects_6_io_outs_5; // @[MemPrimitives.scala 123:41:@21578.4]
  assign _T_1791 = StickySelects_6_io_outs_6; // @[MemPrimitives.scala 123:41:@21579.4]
  assign _T_1792 = StickySelects_6_io_outs_7; // @[MemPrimitives.scala 123:41:@21580.4]
  assign _T_1793 = StickySelects_6_io_outs_8; // @[MemPrimitives.scala 123:41:@21581.4]
  assign _T_1795 = {_T_1785,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@21583.4]
  assign _T_1797 = {_T_1786,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@21585.4]
  assign _T_1799 = {_T_1787,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@21587.4]
  assign _T_1801 = {_T_1788,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@21589.4]
  assign _T_1803 = {_T_1789,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@21591.4]
  assign _T_1805 = {_T_1790,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@21593.4]
  assign _T_1807 = {_T_1791,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@21595.4]
  assign _T_1809 = {_T_1792,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@21597.4]
  assign _T_1811 = {_T_1793,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@21599.4]
  assign _T_1812 = _T_1792 ? _T_1809 : _T_1811; // @[Mux.scala 31:69:@21600.4]
  assign _T_1813 = _T_1791 ? _T_1807 : _T_1812; // @[Mux.scala 31:69:@21601.4]
  assign _T_1814 = _T_1790 ? _T_1805 : _T_1813; // @[Mux.scala 31:69:@21602.4]
  assign _T_1815 = _T_1789 ? _T_1803 : _T_1814; // @[Mux.scala 31:69:@21603.4]
  assign _T_1816 = _T_1788 ? _T_1801 : _T_1815; // @[Mux.scala 31:69:@21604.4]
  assign _T_1817 = _T_1787 ? _T_1799 : _T_1816; // @[Mux.scala 31:69:@21605.4]
  assign _T_1818 = _T_1786 ? _T_1797 : _T_1817; // @[Mux.scala 31:69:@21606.4]
  assign _T_1819 = _T_1785 ? _T_1795 : _T_1818; // @[Mux.scala 31:69:@21607.4]
  assign _T_1824 = io_rPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21614.4]
  assign _T_1827 = _T_1824 & _T_1274; // @[MemPrimitives.scala 110:228:@21616.4]
  assign _T_1830 = io_rPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21618.4]
  assign _T_1833 = _T_1830 & _T_1280; // @[MemPrimitives.scala 110:228:@21620.4]
  assign _T_1836 = io_rPort_5_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21622.4]
  assign _T_1839 = _T_1836 & _T_1286; // @[MemPrimitives.scala 110:228:@21624.4]
  assign _T_1842 = io_rPort_6_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21626.4]
  assign _T_1845 = _T_1842 & _T_1292; // @[MemPrimitives.scala 110:228:@21628.4]
  assign _T_1848 = io_rPort_9_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21630.4]
  assign _T_1851 = _T_1848 & _T_1298; // @[MemPrimitives.scala 110:228:@21632.4]
  assign _T_1854 = io_rPort_12_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21634.4]
  assign _T_1857 = _T_1854 & _T_1304; // @[MemPrimitives.scala 110:228:@21636.4]
  assign _T_1860 = io_rPort_13_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21638.4]
  assign _T_1863 = _T_1860 & _T_1310; // @[MemPrimitives.scala 110:228:@21640.4]
  assign _T_1866 = io_rPort_14_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21642.4]
  assign _T_1869 = _T_1866 & _T_1316; // @[MemPrimitives.scala 110:228:@21644.4]
  assign _T_1872 = io_rPort_16_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21646.4]
  assign _T_1875 = _T_1872 & _T_1322; // @[MemPrimitives.scala 110:228:@21648.4]
  assign _T_1877 = StickySelects_7_io_outs_0; // @[MemPrimitives.scala 123:41:@21662.4]
  assign _T_1878 = StickySelects_7_io_outs_1; // @[MemPrimitives.scala 123:41:@21663.4]
  assign _T_1879 = StickySelects_7_io_outs_2; // @[MemPrimitives.scala 123:41:@21664.4]
  assign _T_1880 = StickySelects_7_io_outs_3; // @[MemPrimitives.scala 123:41:@21665.4]
  assign _T_1881 = StickySelects_7_io_outs_4; // @[MemPrimitives.scala 123:41:@21666.4]
  assign _T_1882 = StickySelects_7_io_outs_5; // @[MemPrimitives.scala 123:41:@21667.4]
  assign _T_1883 = StickySelects_7_io_outs_6; // @[MemPrimitives.scala 123:41:@21668.4]
  assign _T_1884 = StickySelects_7_io_outs_7; // @[MemPrimitives.scala 123:41:@21669.4]
  assign _T_1885 = StickySelects_7_io_outs_8; // @[MemPrimitives.scala 123:41:@21670.4]
  assign _T_1887 = {_T_1877,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@21672.4]
  assign _T_1889 = {_T_1878,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@21674.4]
  assign _T_1891 = {_T_1879,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@21676.4]
  assign _T_1893 = {_T_1880,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@21678.4]
  assign _T_1895 = {_T_1881,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@21680.4]
  assign _T_1897 = {_T_1882,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@21682.4]
  assign _T_1899 = {_T_1883,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@21684.4]
  assign _T_1901 = {_T_1884,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@21686.4]
  assign _T_1903 = {_T_1885,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@21688.4]
  assign _T_1904 = _T_1884 ? _T_1901 : _T_1903; // @[Mux.scala 31:69:@21689.4]
  assign _T_1905 = _T_1883 ? _T_1899 : _T_1904; // @[Mux.scala 31:69:@21690.4]
  assign _T_1906 = _T_1882 ? _T_1897 : _T_1905; // @[Mux.scala 31:69:@21691.4]
  assign _T_1907 = _T_1881 ? _T_1895 : _T_1906; // @[Mux.scala 31:69:@21692.4]
  assign _T_1908 = _T_1880 ? _T_1893 : _T_1907; // @[Mux.scala 31:69:@21693.4]
  assign _T_1909 = _T_1879 ? _T_1891 : _T_1908; // @[Mux.scala 31:69:@21694.4]
  assign _T_1910 = _T_1878 ? _T_1889 : _T_1909; // @[Mux.scala 31:69:@21695.4]
  assign _T_1911 = _T_1877 ? _T_1887 : _T_1910; // @[Mux.scala 31:69:@21696.4]
  assign _T_1919 = _T_1732 & _T_1366; // @[MemPrimitives.scala 110:228:@21705.4]
  assign _T_1925 = _T_1738 & _T_1372; // @[MemPrimitives.scala 110:228:@21709.4]
  assign _T_1931 = _T_1744 & _T_1378; // @[MemPrimitives.scala 110:228:@21713.4]
  assign _T_1937 = _T_1750 & _T_1384; // @[MemPrimitives.scala 110:228:@21717.4]
  assign _T_1943 = _T_1756 & _T_1390; // @[MemPrimitives.scala 110:228:@21721.4]
  assign _T_1949 = _T_1762 & _T_1396; // @[MemPrimitives.scala 110:228:@21725.4]
  assign _T_1955 = _T_1768 & _T_1402; // @[MemPrimitives.scala 110:228:@21729.4]
  assign _T_1961 = _T_1774 & _T_1408; // @[MemPrimitives.scala 110:228:@21733.4]
  assign _T_1967 = _T_1780 & _T_1414; // @[MemPrimitives.scala 110:228:@21737.4]
  assign _T_1969 = StickySelects_8_io_outs_0; // @[MemPrimitives.scala 123:41:@21751.4]
  assign _T_1970 = StickySelects_8_io_outs_1; // @[MemPrimitives.scala 123:41:@21752.4]
  assign _T_1971 = StickySelects_8_io_outs_2; // @[MemPrimitives.scala 123:41:@21753.4]
  assign _T_1972 = StickySelects_8_io_outs_3; // @[MemPrimitives.scala 123:41:@21754.4]
  assign _T_1973 = StickySelects_8_io_outs_4; // @[MemPrimitives.scala 123:41:@21755.4]
  assign _T_1974 = StickySelects_8_io_outs_5; // @[MemPrimitives.scala 123:41:@21756.4]
  assign _T_1975 = StickySelects_8_io_outs_6; // @[MemPrimitives.scala 123:41:@21757.4]
  assign _T_1976 = StickySelects_8_io_outs_7; // @[MemPrimitives.scala 123:41:@21758.4]
  assign _T_1977 = StickySelects_8_io_outs_8; // @[MemPrimitives.scala 123:41:@21759.4]
  assign _T_1979 = {_T_1969,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@21761.4]
  assign _T_1981 = {_T_1970,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@21763.4]
  assign _T_1983 = {_T_1971,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@21765.4]
  assign _T_1985 = {_T_1972,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@21767.4]
  assign _T_1987 = {_T_1973,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@21769.4]
  assign _T_1989 = {_T_1974,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@21771.4]
  assign _T_1991 = {_T_1975,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@21773.4]
  assign _T_1993 = {_T_1976,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@21775.4]
  assign _T_1995 = {_T_1977,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@21777.4]
  assign _T_1996 = _T_1976 ? _T_1993 : _T_1995; // @[Mux.scala 31:69:@21778.4]
  assign _T_1997 = _T_1975 ? _T_1991 : _T_1996; // @[Mux.scala 31:69:@21779.4]
  assign _T_1998 = _T_1974 ? _T_1989 : _T_1997; // @[Mux.scala 31:69:@21780.4]
  assign _T_1999 = _T_1973 ? _T_1987 : _T_1998; // @[Mux.scala 31:69:@21781.4]
  assign _T_2000 = _T_1972 ? _T_1985 : _T_1999; // @[Mux.scala 31:69:@21782.4]
  assign _T_2001 = _T_1971 ? _T_1983 : _T_2000; // @[Mux.scala 31:69:@21783.4]
  assign _T_2002 = _T_1970 ? _T_1981 : _T_2001; // @[Mux.scala 31:69:@21784.4]
  assign _T_2003 = _T_1969 ? _T_1979 : _T_2002; // @[Mux.scala 31:69:@21785.4]
  assign _T_2011 = _T_1824 & _T_1458; // @[MemPrimitives.scala 110:228:@21794.4]
  assign _T_2017 = _T_1830 & _T_1464; // @[MemPrimitives.scala 110:228:@21798.4]
  assign _T_2023 = _T_1836 & _T_1470; // @[MemPrimitives.scala 110:228:@21802.4]
  assign _T_2029 = _T_1842 & _T_1476; // @[MemPrimitives.scala 110:228:@21806.4]
  assign _T_2035 = _T_1848 & _T_1482; // @[MemPrimitives.scala 110:228:@21810.4]
  assign _T_2041 = _T_1854 & _T_1488; // @[MemPrimitives.scala 110:228:@21814.4]
  assign _T_2047 = _T_1860 & _T_1494; // @[MemPrimitives.scala 110:228:@21818.4]
  assign _T_2053 = _T_1866 & _T_1500; // @[MemPrimitives.scala 110:228:@21822.4]
  assign _T_2059 = _T_1872 & _T_1506; // @[MemPrimitives.scala 110:228:@21826.4]
  assign _T_2061 = StickySelects_9_io_outs_0; // @[MemPrimitives.scala 123:41:@21840.4]
  assign _T_2062 = StickySelects_9_io_outs_1; // @[MemPrimitives.scala 123:41:@21841.4]
  assign _T_2063 = StickySelects_9_io_outs_2; // @[MemPrimitives.scala 123:41:@21842.4]
  assign _T_2064 = StickySelects_9_io_outs_3; // @[MemPrimitives.scala 123:41:@21843.4]
  assign _T_2065 = StickySelects_9_io_outs_4; // @[MemPrimitives.scala 123:41:@21844.4]
  assign _T_2066 = StickySelects_9_io_outs_5; // @[MemPrimitives.scala 123:41:@21845.4]
  assign _T_2067 = StickySelects_9_io_outs_6; // @[MemPrimitives.scala 123:41:@21846.4]
  assign _T_2068 = StickySelects_9_io_outs_7; // @[MemPrimitives.scala 123:41:@21847.4]
  assign _T_2069 = StickySelects_9_io_outs_8; // @[MemPrimitives.scala 123:41:@21848.4]
  assign _T_2071 = {_T_2061,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@21850.4]
  assign _T_2073 = {_T_2062,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@21852.4]
  assign _T_2075 = {_T_2063,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@21854.4]
  assign _T_2077 = {_T_2064,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@21856.4]
  assign _T_2079 = {_T_2065,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@21858.4]
  assign _T_2081 = {_T_2066,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@21860.4]
  assign _T_2083 = {_T_2067,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@21862.4]
  assign _T_2085 = {_T_2068,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@21864.4]
  assign _T_2087 = {_T_2069,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@21866.4]
  assign _T_2088 = _T_2068 ? _T_2085 : _T_2087; // @[Mux.scala 31:69:@21867.4]
  assign _T_2089 = _T_2067 ? _T_2083 : _T_2088; // @[Mux.scala 31:69:@21868.4]
  assign _T_2090 = _T_2066 ? _T_2081 : _T_2089; // @[Mux.scala 31:69:@21869.4]
  assign _T_2091 = _T_2065 ? _T_2079 : _T_2090; // @[Mux.scala 31:69:@21870.4]
  assign _T_2092 = _T_2064 ? _T_2077 : _T_2091; // @[Mux.scala 31:69:@21871.4]
  assign _T_2093 = _T_2063 ? _T_2075 : _T_2092; // @[Mux.scala 31:69:@21872.4]
  assign _T_2094 = _T_2062 ? _T_2073 : _T_2093; // @[Mux.scala 31:69:@21873.4]
  assign _T_2095 = _T_2061 ? _T_2071 : _T_2094; // @[Mux.scala 31:69:@21874.4]
  assign _T_2103 = _T_1732 & _T_1550; // @[MemPrimitives.scala 110:228:@21883.4]
  assign _T_2109 = _T_1738 & _T_1556; // @[MemPrimitives.scala 110:228:@21887.4]
  assign _T_2115 = _T_1744 & _T_1562; // @[MemPrimitives.scala 110:228:@21891.4]
  assign _T_2121 = _T_1750 & _T_1568; // @[MemPrimitives.scala 110:228:@21895.4]
  assign _T_2127 = _T_1756 & _T_1574; // @[MemPrimitives.scala 110:228:@21899.4]
  assign _T_2133 = _T_1762 & _T_1580; // @[MemPrimitives.scala 110:228:@21903.4]
  assign _T_2139 = _T_1768 & _T_1586; // @[MemPrimitives.scala 110:228:@21907.4]
  assign _T_2145 = _T_1774 & _T_1592; // @[MemPrimitives.scala 110:228:@21911.4]
  assign _T_2151 = _T_1780 & _T_1598; // @[MemPrimitives.scala 110:228:@21915.4]
  assign _T_2153 = StickySelects_10_io_outs_0; // @[MemPrimitives.scala 123:41:@21929.4]
  assign _T_2154 = StickySelects_10_io_outs_1; // @[MemPrimitives.scala 123:41:@21930.4]
  assign _T_2155 = StickySelects_10_io_outs_2; // @[MemPrimitives.scala 123:41:@21931.4]
  assign _T_2156 = StickySelects_10_io_outs_3; // @[MemPrimitives.scala 123:41:@21932.4]
  assign _T_2157 = StickySelects_10_io_outs_4; // @[MemPrimitives.scala 123:41:@21933.4]
  assign _T_2158 = StickySelects_10_io_outs_5; // @[MemPrimitives.scala 123:41:@21934.4]
  assign _T_2159 = StickySelects_10_io_outs_6; // @[MemPrimitives.scala 123:41:@21935.4]
  assign _T_2160 = StickySelects_10_io_outs_7; // @[MemPrimitives.scala 123:41:@21936.4]
  assign _T_2161 = StickySelects_10_io_outs_8; // @[MemPrimitives.scala 123:41:@21937.4]
  assign _T_2163 = {_T_2153,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@21939.4]
  assign _T_2165 = {_T_2154,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@21941.4]
  assign _T_2167 = {_T_2155,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@21943.4]
  assign _T_2169 = {_T_2156,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@21945.4]
  assign _T_2171 = {_T_2157,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@21947.4]
  assign _T_2173 = {_T_2158,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@21949.4]
  assign _T_2175 = {_T_2159,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@21951.4]
  assign _T_2177 = {_T_2160,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@21953.4]
  assign _T_2179 = {_T_2161,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@21955.4]
  assign _T_2180 = _T_2160 ? _T_2177 : _T_2179; // @[Mux.scala 31:69:@21956.4]
  assign _T_2181 = _T_2159 ? _T_2175 : _T_2180; // @[Mux.scala 31:69:@21957.4]
  assign _T_2182 = _T_2158 ? _T_2173 : _T_2181; // @[Mux.scala 31:69:@21958.4]
  assign _T_2183 = _T_2157 ? _T_2171 : _T_2182; // @[Mux.scala 31:69:@21959.4]
  assign _T_2184 = _T_2156 ? _T_2169 : _T_2183; // @[Mux.scala 31:69:@21960.4]
  assign _T_2185 = _T_2155 ? _T_2167 : _T_2184; // @[Mux.scala 31:69:@21961.4]
  assign _T_2186 = _T_2154 ? _T_2165 : _T_2185; // @[Mux.scala 31:69:@21962.4]
  assign _T_2187 = _T_2153 ? _T_2163 : _T_2186; // @[Mux.scala 31:69:@21963.4]
  assign _T_2195 = _T_1824 & _T_1642; // @[MemPrimitives.scala 110:228:@21972.4]
  assign _T_2201 = _T_1830 & _T_1648; // @[MemPrimitives.scala 110:228:@21976.4]
  assign _T_2207 = _T_1836 & _T_1654; // @[MemPrimitives.scala 110:228:@21980.4]
  assign _T_2213 = _T_1842 & _T_1660; // @[MemPrimitives.scala 110:228:@21984.4]
  assign _T_2219 = _T_1848 & _T_1666; // @[MemPrimitives.scala 110:228:@21988.4]
  assign _T_2225 = _T_1854 & _T_1672; // @[MemPrimitives.scala 110:228:@21992.4]
  assign _T_2231 = _T_1860 & _T_1678; // @[MemPrimitives.scala 110:228:@21996.4]
  assign _T_2237 = _T_1866 & _T_1684; // @[MemPrimitives.scala 110:228:@22000.4]
  assign _T_2243 = _T_1872 & _T_1690; // @[MemPrimitives.scala 110:228:@22004.4]
  assign _T_2245 = StickySelects_11_io_outs_0; // @[MemPrimitives.scala 123:41:@22018.4]
  assign _T_2246 = StickySelects_11_io_outs_1; // @[MemPrimitives.scala 123:41:@22019.4]
  assign _T_2247 = StickySelects_11_io_outs_2; // @[MemPrimitives.scala 123:41:@22020.4]
  assign _T_2248 = StickySelects_11_io_outs_3; // @[MemPrimitives.scala 123:41:@22021.4]
  assign _T_2249 = StickySelects_11_io_outs_4; // @[MemPrimitives.scala 123:41:@22022.4]
  assign _T_2250 = StickySelects_11_io_outs_5; // @[MemPrimitives.scala 123:41:@22023.4]
  assign _T_2251 = StickySelects_11_io_outs_6; // @[MemPrimitives.scala 123:41:@22024.4]
  assign _T_2252 = StickySelects_11_io_outs_7; // @[MemPrimitives.scala 123:41:@22025.4]
  assign _T_2253 = StickySelects_11_io_outs_8; // @[MemPrimitives.scala 123:41:@22026.4]
  assign _T_2255 = {_T_2245,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@22028.4]
  assign _T_2257 = {_T_2246,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@22030.4]
  assign _T_2259 = {_T_2247,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@22032.4]
  assign _T_2261 = {_T_2248,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@22034.4]
  assign _T_2263 = {_T_2249,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@22036.4]
  assign _T_2265 = {_T_2250,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@22038.4]
  assign _T_2267 = {_T_2251,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@22040.4]
  assign _T_2269 = {_T_2252,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@22042.4]
  assign _T_2271 = {_T_2253,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@22044.4]
  assign _T_2272 = _T_2252 ? _T_2269 : _T_2271; // @[Mux.scala 31:69:@22045.4]
  assign _T_2273 = _T_2251 ? _T_2267 : _T_2272; // @[Mux.scala 31:69:@22046.4]
  assign _T_2274 = _T_2250 ? _T_2265 : _T_2273; // @[Mux.scala 31:69:@22047.4]
  assign _T_2275 = _T_2249 ? _T_2263 : _T_2274; // @[Mux.scala 31:69:@22048.4]
  assign _T_2276 = _T_2248 ? _T_2261 : _T_2275; // @[Mux.scala 31:69:@22049.4]
  assign _T_2277 = _T_2247 ? _T_2259 : _T_2276; // @[Mux.scala 31:69:@22050.4]
  assign _T_2278 = _T_2246 ? _T_2257 : _T_2277; // @[Mux.scala 31:69:@22051.4]
  assign _T_2279 = _T_2245 ? _T_2255 : _T_2278; // @[Mux.scala 31:69:@22052.4]
  assign _T_2284 = io_rPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22059.4]
  assign _T_2287 = _T_2284 & _T_1182; // @[MemPrimitives.scala 110:228:@22061.4]
  assign _T_2290 = io_rPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22063.4]
  assign _T_2293 = _T_2290 & _T_1188; // @[MemPrimitives.scala 110:228:@22065.4]
  assign _T_2296 = io_rPort_4_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22067.4]
  assign _T_2299 = _T_2296 & _T_1194; // @[MemPrimitives.scala 110:228:@22069.4]
  assign _T_2302 = io_rPort_7_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22071.4]
  assign _T_2305 = _T_2302 & _T_1200; // @[MemPrimitives.scala 110:228:@22073.4]
  assign _T_2308 = io_rPort_8_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22075.4]
  assign _T_2311 = _T_2308 & _T_1206; // @[MemPrimitives.scala 110:228:@22077.4]
  assign _T_2314 = io_rPort_10_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22079.4]
  assign _T_2317 = _T_2314 & _T_1212; // @[MemPrimitives.scala 110:228:@22081.4]
  assign _T_2320 = io_rPort_11_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22083.4]
  assign _T_2323 = _T_2320 & _T_1218; // @[MemPrimitives.scala 110:228:@22085.4]
  assign _T_2326 = io_rPort_15_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22087.4]
  assign _T_2329 = _T_2326 & _T_1224; // @[MemPrimitives.scala 110:228:@22089.4]
  assign _T_2332 = io_rPort_17_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22091.4]
  assign _T_2335 = _T_2332 & _T_1230; // @[MemPrimitives.scala 110:228:@22093.4]
  assign _T_2337 = StickySelects_12_io_outs_0; // @[MemPrimitives.scala 123:41:@22107.4]
  assign _T_2338 = StickySelects_12_io_outs_1; // @[MemPrimitives.scala 123:41:@22108.4]
  assign _T_2339 = StickySelects_12_io_outs_2; // @[MemPrimitives.scala 123:41:@22109.4]
  assign _T_2340 = StickySelects_12_io_outs_3; // @[MemPrimitives.scala 123:41:@22110.4]
  assign _T_2341 = StickySelects_12_io_outs_4; // @[MemPrimitives.scala 123:41:@22111.4]
  assign _T_2342 = StickySelects_12_io_outs_5; // @[MemPrimitives.scala 123:41:@22112.4]
  assign _T_2343 = StickySelects_12_io_outs_6; // @[MemPrimitives.scala 123:41:@22113.4]
  assign _T_2344 = StickySelects_12_io_outs_7; // @[MemPrimitives.scala 123:41:@22114.4]
  assign _T_2345 = StickySelects_12_io_outs_8; // @[MemPrimitives.scala 123:41:@22115.4]
  assign _T_2347 = {_T_2337,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@22117.4]
  assign _T_2349 = {_T_2338,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@22119.4]
  assign _T_2351 = {_T_2339,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@22121.4]
  assign _T_2353 = {_T_2340,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@22123.4]
  assign _T_2355 = {_T_2341,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@22125.4]
  assign _T_2357 = {_T_2342,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@22127.4]
  assign _T_2359 = {_T_2343,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@22129.4]
  assign _T_2361 = {_T_2344,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@22131.4]
  assign _T_2363 = {_T_2345,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@22133.4]
  assign _T_2364 = _T_2344 ? _T_2361 : _T_2363; // @[Mux.scala 31:69:@22134.4]
  assign _T_2365 = _T_2343 ? _T_2359 : _T_2364; // @[Mux.scala 31:69:@22135.4]
  assign _T_2366 = _T_2342 ? _T_2357 : _T_2365; // @[Mux.scala 31:69:@22136.4]
  assign _T_2367 = _T_2341 ? _T_2355 : _T_2366; // @[Mux.scala 31:69:@22137.4]
  assign _T_2368 = _T_2340 ? _T_2353 : _T_2367; // @[Mux.scala 31:69:@22138.4]
  assign _T_2369 = _T_2339 ? _T_2351 : _T_2368; // @[Mux.scala 31:69:@22139.4]
  assign _T_2370 = _T_2338 ? _T_2349 : _T_2369; // @[Mux.scala 31:69:@22140.4]
  assign _T_2371 = _T_2337 ? _T_2347 : _T_2370; // @[Mux.scala 31:69:@22141.4]
  assign _T_2376 = io_rPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22148.4]
  assign _T_2379 = _T_2376 & _T_1274; // @[MemPrimitives.scala 110:228:@22150.4]
  assign _T_2382 = io_rPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22152.4]
  assign _T_2385 = _T_2382 & _T_1280; // @[MemPrimitives.scala 110:228:@22154.4]
  assign _T_2388 = io_rPort_5_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22156.4]
  assign _T_2391 = _T_2388 & _T_1286; // @[MemPrimitives.scala 110:228:@22158.4]
  assign _T_2394 = io_rPort_6_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22160.4]
  assign _T_2397 = _T_2394 & _T_1292; // @[MemPrimitives.scala 110:228:@22162.4]
  assign _T_2400 = io_rPort_9_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22164.4]
  assign _T_2403 = _T_2400 & _T_1298; // @[MemPrimitives.scala 110:228:@22166.4]
  assign _T_2406 = io_rPort_12_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22168.4]
  assign _T_2409 = _T_2406 & _T_1304; // @[MemPrimitives.scala 110:228:@22170.4]
  assign _T_2412 = io_rPort_13_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22172.4]
  assign _T_2415 = _T_2412 & _T_1310; // @[MemPrimitives.scala 110:228:@22174.4]
  assign _T_2418 = io_rPort_14_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22176.4]
  assign _T_2421 = _T_2418 & _T_1316; // @[MemPrimitives.scala 110:228:@22178.4]
  assign _T_2424 = io_rPort_16_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22180.4]
  assign _T_2427 = _T_2424 & _T_1322; // @[MemPrimitives.scala 110:228:@22182.4]
  assign _T_2429 = StickySelects_13_io_outs_0; // @[MemPrimitives.scala 123:41:@22196.4]
  assign _T_2430 = StickySelects_13_io_outs_1; // @[MemPrimitives.scala 123:41:@22197.4]
  assign _T_2431 = StickySelects_13_io_outs_2; // @[MemPrimitives.scala 123:41:@22198.4]
  assign _T_2432 = StickySelects_13_io_outs_3; // @[MemPrimitives.scala 123:41:@22199.4]
  assign _T_2433 = StickySelects_13_io_outs_4; // @[MemPrimitives.scala 123:41:@22200.4]
  assign _T_2434 = StickySelects_13_io_outs_5; // @[MemPrimitives.scala 123:41:@22201.4]
  assign _T_2435 = StickySelects_13_io_outs_6; // @[MemPrimitives.scala 123:41:@22202.4]
  assign _T_2436 = StickySelects_13_io_outs_7; // @[MemPrimitives.scala 123:41:@22203.4]
  assign _T_2437 = StickySelects_13_io_outs_8; // @[MemPrimitives.scala 123:41:@22204.4]
  assign _T_2439 = {_T_2429,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@22206.4]
  assign _T_2441 = {_T_2430,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@22208.4]
  assign _T_2443 = {_T_2431,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@22210.4]
  assign _T_2445 = {_T_2432,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@22212.4]
  assign _T_2447 = {_T_2433,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@22214.4]
  assign _T_2449 = {_T_2434,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@22216.4]
  assign _T_2451 = {_T_2435,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@22218.4]
  assign _T_2453 = {_T_2436,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@22220.4]
  assign _T_2455 = {_T_2437,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@22222.4]
  assign _T_2456 = _T_2436 ? _T_2453 : _T_2455; // @[Mux.scala 31:69:@22223.4]
  assign _T_2457 = _T_2435 ? _T_2451 : _T_2456; // @[Mux.scala 31:69:@22224.4]
  assign _T_2458 = _T_2434 ? _T_2449 : _T_2457; // @[Mux.scala 31:69:@22225.4]
  assign _T_2459 = _T_2433 ? _T_2447 : _T_2458; // @[Mux.scala 31:69:@22226.4]
  assign _T_2460 = _T_2432 ? _T_2445 : _T_2459; // @[Mux.scala 31:69:@22227.4]
  assign _T_2461 = _T_2431 ? _T_2443 : _T_2460; // @[Mux.scala 31:69:@22228.4]
  assign _T_2462 = _T_2430 ? _T_2441 : _T_2461; // @[Mux.scala 31:69:@22229.4]
  assign _T_2463 = _T_2429 ? _T_2439 : _T_2462; // @[Mux.scala 31:69:@22230.4]
  assign _T_2471 = _T_2284 & _T_1366; // @[MemPrimitives.scala 110:228:@22239.4]
  assign _T_2477 = _T_2290 & _T_1372; // @[MemPrimitives.scala 110:228:@22243.4]
  assign _T_2483 = _T_2296 & _T_1378; // @[MemPrimitives.scala 110:228:@22247.4]
  assign _T_2489 = _T_2302 & _T_1384; // @[MemPrimitives.scala 110:228:@22251.4]
  assign _T_2495 = _T_2308 & _T_1390; // @[MemPrimitives.scala 110:228:@22255.4]
  assign _T_2501 = _T_2314 & _T_1396; // @[MemPrimitives.scala 110:228:@22259.4]
  assign _T_2507 = _T_2320 & _T_1402; // @[MemPrimitives.scala 110:228:@22263.4]
  assign _T_2513 = _T_2326 & _T_1408; // @[MemPrimitives.scala 110:228:@22267.4]
  assign _T_2519 = _T_2332 & _T_1414; // @[MemPrimitives.scala 110:228:@22271.4]
  assign _T_2521 = StickySelects_14_io_outs_0; // @[MemPrimitives.scala 123:41:@22285.4]
  assign _T_2522 = StickySelects_14_io_outs_1; // @[MemPrimitives.scala 123:41:@22286.4]
  assign _T_2523 = StickySelects_14_io_outs_2; // @[MemPrimitives.scala 123:41:@22287.4]
  assign _T_2524 = StickySelects_14_io_outs_3; // @[MemPrimitives.scala 123:41:@22288.4]
  assign _T_2525 = StickySelects_14_io_outs_4; // @[MemPrimitives.scala 123:41:@22289.4]
  assign _T_2526 = StickySelects_14_io_outs_5; // @[MemPrimitives.scala 123:41:@22290.4]
  assign _T_2527 = StickySelects_14_io_outs_6; // @[MemPrimitives.scala 123:41:@22291.4]
  assign _T_2528 = StickySelects_14_io_outs_7; // @[MemPrimitives.scala 123:41:@22292.4]
  assign _T_2529 = StickySelects_14_io_outs_8; // @[MemPrimitives.scala 123:41:@22293.4]
  assign _T_2531 = {_T_2521,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@22295.4]
  assign _T_2533 = {_T_2522,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@22297.4]
  assign _T_2535 = {_T_2523,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@22299.4]
  assign _T_2537 = {_T_2524,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@22301.4]
  assign _T_2539 = {_T_2525,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@22303.4]
  assign _T_2541 = {_T_2526,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@22305.4]
  assign _T_2543 = {_T_2527,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@22307.4]
  assign _T_2545 = {_T_2528,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@22309.4]
  assign _T_2547 = {_T_2529,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@22311.4]
  assign _T_2548 = _T_2528 ? _T_2545 : _T_2547; // @[Mux.scala 31:69:@22312.4]
  assign _T_2549 = _T_2527 ? _T_2543 : _T_2548; // @[Mux.scala 31:69:@22313.4]
  assign _T_2550 = _T_2526 ? _T_2541 : _T_2549; // @[Mux.scala 31:69:@22314.4]
  assign _T_2551 = _T_2525 ? _T_2539 : _T_2550; // @[Mux.scala 31:69:@22315.4]
  assign _T_2552 = _T_2524 ? _T_2537 : _T_2551; // @[Mux.scala 31:69:@22316.4]
  assign _T_2553 = _T_2523 ? _T_2535 : _T_2552; // @[Mux.scala 31:69:@22317.4]
  assign _T_2554 = _T_2522 ? _T_2533 : _T_2553; // @[Mux.scala 31:69:@22318.4]
  assign _T_2555 = _T_2521 ? _T_2531 : _T_2554; // @[Mux.scala 31:69:@22319.4]
  assign _T_2563 = _T_2376 & _T_1458; // @[MemPrimitives.scala 110:228:@22328.4]
  assign _T_2569 = _T_2382 & _T_1464; // @[MemPrimitives.scala 110:228:@22332.4]
  assign _T_2575 = _T_2388 & _T_1470; // @[MemPrimitives.scala 110:228:@22336.4]
  assign _T_2581 = _T_2394 & _T_1476; // @[MemPrimitives.scala 110:228:@22340.4]
  assign _T_2587 = _T_2400 & _T_1482; // @[MemPrimitives.scala 110:228:@22344.4]
  assign _T_2593 = _T_2406 & _T_1488; // @[MemPrimitives.scala 110:228:@22348.4]
  assign _T_2599 = _T_2412 & _T_1494; // @[MemPrimitives.scala 110:228:@22352.4]
  assign _T_2605 = _T_2418 & _T_1500; // @[MemPrimitives.scala 110:228:@22356.4]
  assign _T_2611 = _T_2424 & _T_1506; // @[MemPrimitives.scala 110:228:@22360.4]
  assign _T_2613 = StickySelects_15_io_outs_0; // @[MemPrimitives.scala 123:41:@22374.4]
  assign _T_2614 = StickySelects_15_io_outs_1; // @[MemPrimitives.scala 123:41:@22375.4]
  assign _T_2615 = StickySelects_15_io_outs_2; // @[MemPrimitives.scala 123:41:@22376.4]
  assign _T_2616 = StickySelects_15_io_outs_3; // @[MemPrimitives.scala 123:41:@22377.4]
  assign _T_2617 = StickySelects_15_io_outs_4; // @[MemPrimitives.scala 123:41:@22378.4]
  assign _T_2618 = StickySelects_15_io_outs_5; // @[MemPrimitives.scala 123:41:@22379.4]
  assign _T_2619 = StickySelects_15_io_outs_6; // @[MemPrimitives.scala 123:41:@22380.4]
  assign _T_2620 = StickySelects_15_io_outs_7; // @[MemPrimitives.scala 123:41:@22381.4]
  assign _T_2621 = StickySelects_15_io_outs_8; // @[MemPrimitives.scala 123:41:@22382.4]
  assign _T_2623 = {_T_2613,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@22384.4]
  assign _T_2625 = {_T_2614,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@22386.4]
  assign _T_2627 = {_T_2615,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@22388.4]
  assign _T_2629 = {_T_2616,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@22390.4]
  assign _T_2631 = {_T_2617,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@22392.4]
  assign _T_2633 = {_T_2618,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@22394.4]
  assign _T_2635 = {_T_2619,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@22396.4]
  assign _T_2637 = {_T_2620,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@22398.4]
  assign _T_2639 = {_T_2621,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@22400.4]
  assign _T_2640 = _T_2620 ? _T_2637 : _T_2639; // @[Mux.scala 31:69:@22401.4]
  assign _T_2641 = _T_2619 ? _T_2635 : _T_2640; // @[Mux.scala 31:69:@22402.4]
  assign _T_2642 = _T_2618 ? _T_2633 : _T_2641; // @[Mux.scala 31:69:@22403.4]
  assign _T_2643 = _T_2617 ? _T_2631 : _T_2642; // @[Mux.scala 31:69:@22404.4]
  assign _T_2644 = _T_2616 ? _T_2629 : _T_2643; // @[Mux.scala 31:69:@22405.4]
  assign _T_2645 = _T_2615 ? _T_2627 : _T_2644; // @[Mux.scala 31:69:@22406.4]
  assign _T_2646 = _T_2614 ? _T_2625 : _T_2645; // @[Mux.scala 31:69:@22407.4]
  assign _T_2647 = _T_2613 ? _T_2623 : _T_2646; // @[Mux.scala 31:69:@22408.4]
  assign _T_2655 = _T_2284 & _T_1550; // @[MemPrimitives.scala 110:228:@22417.4]
  assign _T_2661 = _T_2290 & _T_1556; // @[MemPrimitives.scala 110:228:@22421.4]
  assign _T_2667 = _T_2296 & _T_1562; // @[MemPrimitives.scala 110:228:@22425.4]
  assign _T_2673 = _T_2302 & _T_1568; // @[MemPrimitives.scala 110:228:@22429.4]
  assign _T_2679 = _T_2308 & _T_1574; // @[MemPrimitives.scala 110:228:@22433.4]
  assign _T_2685 = _T_2314 & _T_1580; // @[MemPrimitives.scala 110:228:@22437.4]
  assign _T_2691 = _T_2320 & _T_1586; // @[MemPrimitives.scala 110:228:@22441.4]
  assign _T_2697 = _T_2326 & _T_1592; // @[MemPrimitives.scala 110:228:@22445.4]
  assign _T_2703 = _T_2332 & _T_1598; // @[MemPrimitives.scala 110:228:@22449.4]
  assign _T_2705 = StickySelects_16_io_outs_0; // @[MemPrimitives.scala 123:41:@22463.4]
  assign _T_2706 = StickySelects_16_io_outs_1; // @[MemPrimitives.scala 123:41:@22464.4]
  assign _T_2707 = StickySelects_16_io_outs_2; // @[MemPrimitives.scala 123:41:@22465.4]
  assign _T_2708 = StickySelects_16_io_outs_3; // @[MemPrimitives.scala 123:41:@22466.4]
  assign _T_2709 = StickySelects_16_io_outs_4; // @[MemPrimitives.scala 123:41:@22467.4]
  assign _T_2710 = StickySelects_16_io_outs_5; // @[MemPrimitives.scala 123:41:@22468.4]
  assign _T_2711 = StickySelects_16_io_outs_6; // @[MemPrimitives.scala 123:41:@22469.4]
  assign _T_2712 = StickySelects_16_io_outs_7; // @[MemPrimitives.scala 123:41:@22470.4]
  assign _T_2713 = StickySelects_16_io_outs_8; // @[MemPrimitives.scala 123:41:@22471.4]
  assign _T_2715 = {_T_2705,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@22473.4]
  assign _T_2717 = {_T_2706,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@22475.4]
  assign _T_2719 = {_T_2707,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@22477.4]
  assign _T_2721 = {_T_2708,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@22479.4]
  assign _T_2723 = {_T_2709,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@22481.4]
  assign _T_2725 = {_T_2710,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@22483.4]
  assign _T_2727 = {_T_2711,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@22485.4]
  assign _T_2729 = {_T_2712,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@22487.4]
  assign _T_2731 = {_T_2713,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@22489.4]
  assign _T_2732 = _T_2712 ? _T_2729 : _T_2731; // @[Mux.scala 31:69:@22490.4]
  assign _T_2733 = _T_2711 ? _T_2727 : _T_2732; // @[Mux.scala 31:69:@22491.4]
  assign _T_2734 = _T_2710 ? _T_2725 : _T_2733; // @[Mux.scala 31:69:@22492.4]
  assign _T_2735 = _T_2709 ? _T_2723 : _T_2734; // @[Mux.scala 31:69:@22493.4]
  assign _T_2736 = _T_2708 ? _T_2721 : _T_2735; // @[Mux.scala 31:69:@22494.4]
  assign _T_2737 = _T_2707 ? _T_2719 : _T_2736; // @[Mux.scala 31:69:@22495.4]
  assign _T_2738 = _T_2706 ? _T_2717 : _T_2737; // @[Mux.scala 31:69:@22496.4]
  assign _T_2739 = _T_2705 ? _T_2715 : _T_2738; // @[Mux.scala 31:69:@22497.4]
  assign _T_2747 = _T_2376 & _T_1642; // @[MemPrimitives.scala 110:228:@22506.4]
  assign _T_2753 = _T_2382 & _T_1648; // @[MemPrimitives.scala 110:228:@22510.4]
  assign _T_2759 = _T_2388 & _T_1654; // @[MemPrimitives.scala 110:228:@22514.4]
  assign _T_2765 = _T_2394 & _T_1660; // @[MemPrimitives.scala 110:228:@22518.4]
  assign _T_2771 = _T_2400 & _T_1666; // @[MemPrimitives.scala 110:228:@22522.4]
  assign _T_2777 = _T_2406 & _T_1672; // @[MemPrimitives.scala 110:228:@22526.4]
  assign _T_2783 = _T_2412 & _T_1678; // @[MemPrimitives.scala 110:228:@22530.4]
  assign _T_2789 = _T_2418 & _T_1684; // @[MemPrimitives.scala 110:228:@22534.4]
  assign _T_2795 = _T_2424 & _T_1690; // @[MemPrimitives.scala 110:228:@22538.4]
  assign _T_2797 = StickySelects_17_io_outs_0; // @[MemPrimitives.scala 123:41:@22552.4]
  assign _T_2798 = StickySelects_17_io_outs_1; // @[MemPrimitives.scala 123:41:@22553.4]
  assign _T_2799 = StickySelects_17_io_outs_2; // @[MemPrimitives.scala 123:41:@22554.4]
  assign _T_2800 = StickySelects_17_io_outs_3; // @[MemPrimitives.scala 123:41:@22555.4]
  assign _T_2801 = StickySelects_17_io_outs_4; // @[MemPrimitives.scala 123:41:@22556.4]
  assign _T_2802 = StickySelects_17_io_outs_5; // @[MemPrimitives.scala 123:41:@22557.4]
  assign _T_2803 = StickySelects_17_io_outs_6; // @[MemPrimitives.scala 123:41:@22558.4]
  assign _T_2804 = StickySelects_17_io_outs_7; // @[MemPrimitives.scala 123:41:@22559.4]
  assign _T_2805 = StickySelects_17_io_outs_8; // @[MemPrimitives.scala 123:41:@22560.4]
  assign _T_2807 = {_T_2797,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@22562.4]
  assign _T_2809 = {_T_2798,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@22564.4]
  assign _T_2811 = {_T_2799,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@22566.4]
  assign _T_2813 = {_T_2800,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@22568.4]
  assign _T_2815 = {_T_2801,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@22570.4]
  assign _T_2817 = {_T_2802,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@22572.4]
  assign _T_2819 = {_T_2803,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@22574.4]
  assign _T_2821 = {_T_2804,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@22576.4]
  assign _T_2823 = {_T_2805,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@22578.4]
  assign _T_2824 = _T_2804 ? _T_2821 : _T_2823; // @[Mux.scala 31:69:@22579.4]
  assign _T_2825 = _T_2803 ? _T_2819 : _T_2824; // @[Mux.scala 31:69:@22580.4]
  assign _T_2826 = _T_2802 ? _T_2817 : _T_2825; // @[Mux.scala 31:69:@22581.4]
  assign _T_2827 = _T_2801 ? _T_2815 : _T_2826; // @[Mux.scala 31:69:@22582.4]
  assign _T_2828 = _T_2800 ? _T_2813 : _T_2827; // @[Mux.scala 31:69:@22583.4]
  assign _T_2829 = _T_2799 ? _T_2811 : _T_2828; // @[Mux.scala 31:69:@22584.4]
  assign _T_2830 = _T_2798 ? _T_2809 : _T_2829; // @[Mux.scala 31:69:@22585.4]
  assign _T_2831 = _T_2797 ? _T_2807 : _T_2830; // @[Mux.scala 31:69:@22586.4]
  assign _T_2836 = io_rPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22593.4]
  assign _T_2839 = _T_2836 & _T_1182; // @[MemPrimitives.scala 110:228:@22595.4]
  assign _T_2842 = io_rPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22597.4]
  assign _T_2845 = _T_2842 & _T_1188; // @[MemPrimitives.scala 110:228:@22599.4]
  assign _T_2848 = io_rPort_4_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22601.4]
  assign _T_2851 = _T_2848 & _T_1194; // @[MemPrimitives.scala 110:228:@22603.4]
  assign _T_2854 = io_rPort_7_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22605.4]
  assign _T_2857 = _T_2854 & _T_1200; // @[MemPrimitives.scala 110:228:@22607.4]
  assign _T_2860 = io_rPort_8_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22609.4]
  assign _T_2863 = _T_2860 & _T_1206; // @[MemPrimitives.scala 110:228:@22611.4]
  assign _T_2866 = io_rPort_10_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22613.4]
  assign _T_2869 = _T_2866 & _T_1212; // @[MemPrimitives.scala 110:228:@22615.4]
  assign _T_2872 = io_rPort_11_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22617.4]
  assign _T_2875 = _T_2872 & _T_1218; // @[MemPrimitives.scala 110:228:@22619.4]
  assign _T_2878 = io_rPort_15_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22621.4]
  assign _T_2881 = _T_2878 & _T_1224; // @[MemPrimitives.scala 110:228:@22623.4]
  assign _T_2884 = io_rPort_17_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22625.4]
  assign _T_2887 = _T_2884 & _T_1230; // @[MemPrimitives.scala 110:228:@22627.4]
  assign _T_2889 = StickySelects_18_io_outs_0; // @[MemPrimitives.scala 123:41:@22641.4]
  assign _T_2890 = StickySelects_18_io_outs_1; // @[MemPrimitives.scala 123:41:@22642.4]
  assign _T_2891 = StickySelects_18_io_outs_2; // @[MemPrimitives.scala 123:41:@22643.4]
  assign _T_2892 = StickySelects_18_io_outs_3; // @[MemPrimitives.scala 123:41:@22644.4]
  assign _T_2893 = StickySelects_18_io_outs_4; // @[MemPrimitives.scala 123:41:@22645.4]
  assign _T_2894 = StickySelects_18_io_outs_5; // @[MemPrimitives.scala 123:41:@22646.4]
  assign _T_2895 = StickySelects_18_io_outs_6; // @[MemPrimitives.scala 123:41:@22647.4]
  assign _T_2896 = StickySelects_18_io_outs_7; // @[MemPrimitives.scala 123:41:@22648.4]
  assign _T_2897 = StickySelects_18_io_outs_8; // @[MemPrimitives.scala 123:41:@22649.4]
  assign _T_2899 = {_T_2889,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@22651.4]
  assign _T_2901 = {_T_2890,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@22653.4]
  assign _T_2903 = {_T_2891,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@22655.4]
  assign _T_2905 = {_T_2892,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@22657.4]
  assign _T_2907 = {_T_2893,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@22659.4]
  assign _T_2909 = {_T_2894,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@22661.4]
  assign _T_2911 = {_T_2895,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@22663.4]
  assign _T_2913 = {_T_2896,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@22665.4]
  assign _T_2915 = {_T_2897,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@22667.4]
  assign _T_2916 = _T_2896 ? _T_2913 : _T_2915; // @[Mux.scala 31:69:@22668.4]
  assign _T_2917 = _T_2895 ? _T_2911 : _T_2916; // @[Mux.scala 31:69:@22669.4]
  assign _T_2918 = _T_2894 ? _T_2909 : _T_2917; // @[Mux.scala 31:69:@22670.4]
  assign _T_2919 = _T_2893 ? _T_2907 : _T_2918; // @[Mux.scala 31:69:@22671.4]
  assign _T_2920 = _T_2892 ? _T_2905 : _T_2919; // @[Mux.scala 31:69:@22672.4]
  assign _T_2921 = _T_2891 ? _T_2903 : _T_2920; // @[Mux.scala 31:69:@22673.4]
  assign _T_2922 = _T_2890 ? _T_2901 : _T_2921; // @[Mux.scala 31:69:@22674.4]
  assign _T_2923 = _T_2889 ? _T_2899 : _T_2922; // @[Mux.scala 31:69:@22675.4]
  assign _T_2928 = io_rPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22682.4]
  assign _T_2931 = _T_2928 & _T_1274; // @[MemPrimitives.scala 110:228:@22684.4]
  assign _T_2934 = io_rPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22686.4]
  assign _T_2937 = _T_2934 & _T_1280; // @[MemPrimitives.scala 110:228:@22688.4]
  assign _T_2940 = io_rPort_5_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22690.4]
  assign _T_2943 = _T_2940 & _T_1286; // @[MemPrimitives.scala 110:228:@22692.4]
  assign _T_2946 = io_rPort_6_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22694.4]
  assign _T_2949 = _T_2946 & _T_1292; // @[MemPrimitives.scala 110:228:@22696.4]
  assign _T_2952 = io_rPort_9_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22698.4]
  assign _T_2955 = _T_2952 & _T_1298; // @[MemPrimitives.scala 110:228:@22700.4]
  assign _T_2958 = io_rPort_12_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22702.4]
  assign _T_2961 = _T_2958 & _T_1304; // @[MemPrimitives.scala 110:228:@22704.4]
  assign _T_2964 = io_rPort_13_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22706.4]
  assign _T_2967 = _T_2964 & _T_1310; // @[MemPrimitives.scala 110:228:@22708.4]
  assign _T_2970 = io_rPort_14_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22710.4]
  assign _T_2973 = _T_2970 & _T_1316; // @[MemPrimitives.scala 110:228:@22712.4]
  assign _T_2976 = io_rPort_16_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22714.4]
  assign _T_2979 = _T_2976 & _T_1322; // @[MemPrimitives.scala 110:228:@22716.4]
  assign _T_2981 = StickySelects_19_io_outs_0; // @[MemPrimitives.scala 123:41:@22730.4]
  assign _T_2982 = StickySelects_19_io_outs_1; // @[MemPrimitives.scala 123:41:@22731.4]
  assign _T_2983 = StickySelects_19_io_outs_2; // @[MemPrimitives.scala 123:41:@22732.4]
  assign _T_2984 = StickySelects_19_io_outs_3; // @[MemPrimitives.scala 123:41:@22733.4]
  assign _T_2985 = StickySelects_19_io_outs_4; // @[MemPrimitives.scala 123:41:@22734.4]
  assign _T_2986 = StickySelects_19_io_outs_5; // @[MemPrimitives.scala 123:41:@22735.4]
  assign _T_2987 = StickySelects_19_io_outs_6; // @[MemPrimitives.scala 123:41:@22736.4]
  assign _T_2988 = StickySelects_19_io_outs_7; // @[MemPrimitives.scala 123:41:@22737.4]
  assign _T_2989 = StickySelects_19_io_outs_8; // @[MemPrimitives.scala 123:41:@22738.4]
  assign _T_2991 = {_T_2981,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@22740.4]
  assign _T_2993 = {_T_2982,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@22742.4]
  assign _T_2995 = {_T_2983,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@22744.4]
  assign _T_2997 = {_T_2984,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@22746.4]
  assign _T_2999 = {_T_2985,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@22748.4]
  assign _T_3001 = {_T_2986,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@22750.4]
  assign _T_3003 = {_T_2987,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@22752.4]
  assign _T_3005 = {_T_2988,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@22754.4]
  assign _T_3007 = {_T_2989,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@22756.4]
  assign _T_3008 = _T_2988 ? _T_3005 : _T_3007; // @[Mux.scala 31:69:@22757.4]
  assign _T_3009 = _T_2987 ? _T_3003 : _T_3008; // @[Mux.scala 31:69:@22758.4]
  assign _T_3010 = _T_2986 ? _T_3001 : _T_3009; // @[Mux.scala 31:69:@22759.4]
  assign _T_3011 = _T_2985 ? _T_2999 : _T_3010; // @[Mux.scala 31:69:@22760.4]
  assign _T_3012 = _T_2984 ? _T_2997 : _T_3011; // @[Mux.scala 31:69:@22761.4]
  assign _T_3013 = _T_2983 ? _T_2995 : _T_3012; // @[Mux.scala 31:69:@22762.4]
  assign _T_3014 = _T_2982 ? _T_2993 : _T_3013; // @[Mux.scala 31:69:@22763.4]
  assign _T_3015 = _T_2981 ? _T_2991 : _T_3014; // @[Mux.scala 31:69:@22764.4]
  assign _T_3023 = _T_2836 & _T_1366; // @[MemPrimitives.scala 110:228:@22773.4]
  assign _T_3029 = _T_2842 & _T_1372; // @[MemPrimitives.scala 110:228:@22777.4]
  assign _T_3035 = _T_2848 & _T_1378; // @[MemPrimitives.scala 110:228:@22781.4]
  assign _T_3041 = _T_2854 & _T_1384; // @[MemPrimitives.scala 110:228:@22785.4]
  assign _T_3047 = _T_2860 & _T_1390; // @[MemPrimitives.scala 110:228:@22789.4]
  assign _T_3053 = _T_2866 & _T_1396; // @[MemPrimitives.scala 110:228:@22793.4]
  assign _T_3059 = _T_2872 & _T_1402; // @[MemPrimitives.scala 110:228:@22797.4]
  assign _T_3065 = _T_2878 & _T_1408; // @[MemPrimitives.scala 110:228:@22801.4]
  assign _T_3071 = _T_2884 & _T_1414; // @[MemPrimitives.scala 110:228:@22805.4]
  assign _T_3073 = StickySelects_20_io_outs_0; // @[MemPrimitives.scala 123:41:@22819.4]
  assign _T_3074 = StickySelects_20_io_outs_1; // @[MemPrimitives.scala 123:41:@22820.4]
  assign _T_3075 = StickySelects_20_io_outs_2; // @[MemPrimitives.scala 123:41:@22821.4]
  assign _T_3076 = StickySelects_20_io_outs_3; // @[MemPrimitives.scala 123:41:@22822.4]
  assign _T_3077 = StickySelects_20_io_outs_4; // @[MemPrimitives.scala 123:41:@22823.4]
  assign _T_3078 = StickySelects_20_io_outs_5; // @[MemPrimitives.scala 123:41:@22824.4]
  assign _T_3079 = StickySelects_20_io_outs_6; // @[MemPrimitives.scala 123:41:@22825.4]
  assign _T_3080 = StickySelects_20_io_outs_7; // @[MemPrimitives.scala 123:41:@22826.4]
  assign _T_3081 = StickySelects_20_io_outs_8; // @[MemPrimitives.scala 123:41:@22827.4]
  assign _T_3083 = {_T_3073,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@22829.4]
  assign _T_3085 = {_T_3074,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@22831.4]
  assign _T_3087 = {_T_3075,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@22833.4]
  assign _T_3089 = {_T_3076,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@22835.4]
  assign _T_3091 = {_T_3077,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@22837.4]
  assign _T_3093 = {_T_3078,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@22839.4]
  assign _T_3095 = {_T_3079,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@22841.4]
  assign _T_3097 = {_T_3080,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@22843.4]
  assign _T_3099 = {_T_3081,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@22845.4]
  assign _T_3100 = _T_3080 ? _T_3097 : _T_3099; // @[Mux.scala 31:69:@22846.4]
  assign _T_3101 = _T_3079 ? _T_3095 : _T_3100; // @[Mux.scala 31:69:@22847.4]
  assign _T_3102 = _T_3078 ? _T_3093 : _T_3101; // @[Mux.scala 31:69:@22848.4]
  assign _T_3103 = _T_3077 ? _T_3091 : _T_3102; // @[Mux.scala 31:69:@22849.4]
  assign _T_3104 = _T_3076 ? _T_3089 : _T_3103; // @[Mux.scala 31:69:@22850.4]
  assign _T_3105 = _T_3075 ? _T_3087 : _T_3104; // @[Mux.scala 31:69:@22851.4]
  assign _T_3106 = _T_3074 ? _T_3085 : _T_3105; // @[Mux.scala 31:69:@22852.4]
  assign _T_3107 = _T_3073 ? _T_3083 : _T_3106; // @[Mux.scala 31:69:@22853.4]
  assign _T_3115 = _T_2928 & _T_1458; // @[MemPrimitives.scala 110:228:@22862.4]
  assign _T_3121 = _T_2934 & _T_1464; // @[MemPrimitives.scala 110:228:@22866.4]
  assign _T_3127 = _T_2940 & _T_1470; // @[MemPrimitives.scala 110:228:@22870.4]
  assign _T_3133 = _T_2946 & _T_1476; // @[MemPrimitives.scala 110:228:@22874.4]
  assign _T_3139 = _T_2952 & _T_1482; // @[MemPrimitives.scala 110:228:@22878.4]
  assign _T_3145 = _T_2958 & _T_1488; // @[MemPrimitives.scala 110:228:@22882.4]
  assign _T_3151 = _T_2964 & _T_1494; // @[MemPrimitives.scala 110:228:@22886.4]
  assign _T_3157 = _T_2970 & _T_1500; // @[MemPrimitives.scala 110:228:@22890.4]
  assign _T_3163 = _T_2976 & _T_1506; // @[MemPrimitives.scala 110:228:@22894.4]
  assign _T_3165 = StickySelects_21_io_outs_0; // @[MemPrimitives.scala 123:41:@22908.4]
  assign _T_3166 = StickySelects_21_io_outs_1; // @[MemPrimitives.scala 123:41:@22909.4]
  assign _T_3167 = StickySelects_21_io_outs_2; // @[MemPrimitives.scala 123:41:@22910.4]
  assign _T_3168 = StickySelects_21_io_outs_3; // @[MemPrimitives.scala 123:41:@22911.4]
  assign _T_3169 = StickySelects_21_io_outs_4; // @[MemPrimitives.scala 123:41:@22912.4]
  assign _T_3170 = StickySelects_21_io_outs_5; // @[MemPrimitives.scala 123:41:@22913.4]
  assign _T_3171 = StickySelects_21_io_outs_6; // @[MemPrimitives.scala 123:41:@22914.4]
  assign _T_3172 = StickySelects_21_io_outs_7; // @[MemPrimitives.scala 123:41:@22915.4]
  assign _T_3173 = StickySelects_21_io_outs_8; // @[MemPrimitives.scala 123:41:@22916.4]
  assign _T_3175 = {_T_3165,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@22918.4]
  assign _T_3177 = {_T_3166,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@22920.4]
  assign _T_3179 = {_T_3167,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@22922.4]
  assign _T_3181 = {_T_3168,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@22924.4]
  assign _T_3183 = {_T_3169,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@22926.4]
  assign _T_3185 = {_T_3170,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@22928.4]
  assign _T_3187 = {_T_3171,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@22930.4]
  assign _T_3189 = {_T_3172,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@22932.4]
  assign _T_3191 = {_T_3173,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@22934.4]
  assign _T_3192 = _T_3172 ? _T_3189 : _T_3191; // @[Mux.scala 31:69:@22935.4]
  assign _T_3193 = _T_3171 ? _T_3187 : _T_3192; // @[Mux.scala 31:69:@22936.4]
  assign _T_3194 = _T_3170 ? _T_3185 : _T_3193; // @[Mux.scala 31:69:@22937.4]
  assign _T_3195 = _T_3169 ? _T_3183 : _T_3194; // @[Mux.scala 31:69:@22938.4]
  assign _T_3196 = _T_3168 ? _T_3181 : _T_3195; // @[Mux.scala 31:69:@22939.4]
  assign _T_3197 = _T_3167 ? _T_3179 : _T_3196; // @[Mux.scala 31:69:@22940.4]
  assign _T_3198 = _T_3166 ? _T_3177 : _T_3197; // @[Mux.scala 31:69:@22941.4]
  assign _T_3199 = _T_3165 ? _T_3175 : _T_3198; // @[Mux.scala 31:69:@22942.4]
  assign _T_3207 = _T_2836 & _T_1550; // @[MemPrimitives.scala 110:228:@22951.4]
  assign _T_3213 = _T_2842 & _T_1556; // @[MemPrimitives.scala 110:228:@22955.4]
  assign _T_3219 = _T_2848 & _T_1562; // @[MemPrimitives.scala 110:228:@22959.4]
  assign _T_3225 = _T_2854 & _T_1568; // @[MemPrimitives.scala 110:228:@22963.4]
  assign _T_3231 = _T_2860 & _T_1574; // @[MemPrimitives.scala 110:228:@22967.4]
  assign _T_3237 = _T_2866 & _T_1580; // @[MemPrimitives.scala 110:228:@22971.4]
  assign _T_3243 = _T_2872 & _T_1586; // @[MemPrimitives.scala 110:228:@22975.4]
  assign _T_3249 = _T_2878 & _T_1592; // @[MemPrimitives.scala 110:228:@22979.4]
  assign _T_3255 = _T_2884 & _T_1598; // @[MemPrimitives.scala 110:228:@22983.4]
  assign _T_3257 = StickySelects_22_io_outs_0; // @[MemPrimitives.scala 123:41:@22997.4]
  assign _T_3258 = StickySelects_22_io_outs_1; // @[MemPrimitives.scala 123:41:@22998.4]
  assign _T_3259 = StickySelects_22_io_outs_2; // @[MemPrimitives.scala 123:41:@22999.4]
  assign _T_3260 = StickySelects_22_io_outs_3; // @[MemPrimitives.scala 123:41:@23000.4]
  assign _T_3261 = StickySelects_22_io_outs_4; // @[MemPrimitives.scala 123:41:@23001.4]
  assign _T_3262 = StickySelects_22_io_outs_5; // @[MemPrimitives.scala 123:41:@23002.4]
  assign _T_3263 = StickySelects_22_io_outs_6; // @[MemPrimitives.scala 123:41:@23003.4]
  assign _T_3264 = StickySelects_22_io_outs_7; // @[MemPrimitives.scala 123:41:@23004.4]
  assign _T_3265 = StickySelects_22_io_outs_8; // @[MemPrimitives.scala 123:41:@23005.4]
  assign _T_3267 = {_T_3257,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@23007.4]
  assign _T_3269 = {_T_3258,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@23009.4]
  assign _T_3271 = {_T_3259,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@23011.4]
  assign _T_3273 = {_T_3260,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@23013.4]
  assign _T_3275 = {_T_3261,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@23015.4]
  assign _T_3277 = {_T_3262,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@23017.4]
  assign _T_3279 = {_T_3263,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@23019.4]
  assign _T_3281 = {_T_3264,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@23021.4]
  assign _T_3283 = {_T_3265,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@23023.4]
  assign _T_3284 = _T_3264 ? _T_3281 : _T_3283; // @[Mux.scala 31:69:@23024.4]
  assign _T_3285 = _T_3263 ? _T_3279 : _T_3284; // @[Mux.scala 31:69:@23025.4]
  assign _T_3286 = _T_3262 ? _T_3277 : _T_3285; // @[Mux.scala 31:69:@23026.4]
  assign _T_3287 = _T_3261 ? _T_3275 : _T_3286; // @[Mux.scala 31:69:@23027.4]
  assign _T_3288 = _T_3260 ? _T_3273 : _T_3287; // @[Mux.scala 31:69:@23028.4]
  assign _T_3289 = _T_3259 ? _T_3271 : _T_3288; // @[Mux.scala 31:69:@23029.4]
  assign _T_3290 = _T_3258 ? _T_3269 : _T_3289; // @[Mux.scala 31:69:@23030.4]
  assign _T_3291 = _T_3257 ? _T_3267 : _T_3290; // @[Mux.scala 31:69:@23031.4]
  assign _T_3299 = _T_2928 & _T_1642; // @[MemPrimitives.scala 110:228:@23040.4]
  assign _T_3305 = _T_2934 & _T_1648; // @[MemPrimitives.scala 110:228:@23044.4]
  assign _T_3311 = _T_2940 & _T_1654; // @[MemPrimitives.scala 110:228:@23048.4]
  assign _T_3317 = _T_2946 & _T_1660; // @[MemPrimitives.scala 110:228:@23052.4]
  assign _T_3323 = _T_2952 & _T_1666; // @[MemPrimitives.scala 110:228:@23056.4]
  assign _T_3329 = _T_2958 & _T_1672; // @[MemPrimitives.scala 110:228:@23060.4]
  assign _T_3335 = _T_2964 & _T_1678; // @[MemPrimitives.scala 110:228:@23064.4]
  assign _T_3341 = _T_2970 & _T_1684; // @[MemPrimitives.scala 110:228:@23068.4]
  assign _T_3347 = _T_2976 & _T_1690; // @[MemPrimitives.scala 110:228:@23072.4]
  assign _T_3349 = StickySelects_23_io_outs_0; // @[MemPrimitives.scala 123:41:@23086.4]
  assign _T_3350 = StickySelects_23_io_outs_1; // @[MemPrimitives.scala 123:41:@23087.4]
  assign _T_3351 = StickySelects_23_io_outs_2; // @[MemPrimitives.scala 123:41:@23088.4]
  assign _T_3352 = StickySelects_23_io_outs_3; // @[MemPrimitives.scala 123:41:@23089.4]
  assign _T_3353 = StickySelects_23_io_outs_4; // @[MemPrimitives.scala 123:41:@23090.4]
  assign _T_3354 = StickySelects_23_io_outs_5; // @[MemPrimitives.scala 123:41:@23091.4]
  assign _T_3355 = StickySelects_23_io_outs_6; // @[MemPrimitives.scala 123:41:@23092.4]
  assign _T_3356 = StickySelects_23_io_outs_7; // @[MemPrimitives.scala 123:41:@23093.4]
  assign _T_3357 = StickySelects_23_io_outs_8; // @[MemPrimitives.scala 123:41:@23094.4]
  assign _T_3359 = {_T_3349,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@23096.4]
  assign _T_3361 = {_T_3350,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@23098.4]
  assign _T_3363 = {_T_3351,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@23100.4]
  assign _T_3365 = {_T_3352,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@23102.4]
  assign _T_3367 = {_T_3353,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@23104.4]
  assign _T_3369 = {_T_3354,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@23106.4]
  assign _T_3371 = {_T_3355,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@23108.4]
  assign _T_3373 = {_T_3356,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@23110.4]
  assign _T_3375 = {_T_3357,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@23112.4]
  assign _T_3376 = _T_3356 ? _T_3373 : _T_3375; // @[Mux.scala 31:69:@23113.4]
  assign _T_3377 = _T_3355 ? _T_3371 : _T_3376; // @[Mux.scala 31:69:@23114.4]
  assign _T_3378 = _T_3354 ? _T_3369 : _T_3377; // @[Mux.scala 31:69:@23115.4]
  assign _T_3379 = _T_3353 ? _T_3367 : _T_3378; // @[Mux.scala 31:69:@23116.4]
  assign _T_3380 = _T_3352 ? _T_3365 : _T_3379; // @[Mux.scala 31:69:@23117.4]
  assign _T_3381 = _T_3351 ? _T_3363 : _T_3380; // @[Mux.scala 31:69:@23118.4]
  assign _T_3382 = _T_3350 ? _T_3361 : _T_3381; // @[Mux.scala 31:69:@23119.4]
  assign _T_3383 = _T_3349 ? _T_3359 : _T_3382; // @[Mux.scala 31:69:@23120.4]
  assign _T_3479 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@23249.4 package.scala 96:25:@23250.4]
  assign _T_3483 = _T_3479 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@23259.4]
  assign _T_3476 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@23241.4 package.scala 96:25:@23242.4]
  assign _T_3484 = _T_3476 ? Mem1D_18_io_output : _T_3483; // @[Mux.scala 31:69:@23260.4]
  assign _T_3473 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@23233.4 package.scala 96:25:@23234.4]
  assign _T_3485 = _T_3473 ? Mem1D_16_io_output : _T_3484; // @[Mux.scala 31:69:@23261.4]
  assign _T_3470 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@23225.4 package.scala 96:25:@23226.4]
  assign _T_3486 = _T_3470 ? Mem1D_14_io_output : _T_3485; // @[Mux.scala 31:69:@23262.4]
  assign _T_3467 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@23217.4 package.scala 96:25:@23218.4]
  assign _T_3487 = _T_3467 ? Mem1D_12_io_output : _T_3486; // @[Mux.scala 31:69:@23263.4]
  assign _T_3464 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@23209.4 package.scala 96:25:@23210.4]
  assign _T_3488 = _T_3464 ? Mem1D_10_io_output : _T_3487; // @[Mux.scala 31:69:@23264.4]
  assign _T_3461 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@23201.4 package.scala 96:25:@23202.4]
  assign _T_3489 = _T_3461 ? Mem1D_8_io_output : _T_3488; // @[Mux.scala 31:69:@23265.4]
  assign _T_3458 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@23193.4 package.scala 96:25:@23194.4]
  assign _T_3490 = _T_3458 ? Mem1D_6_io_output : _T_3489; // @[Mux.scala 31:69:@23266.4]
  assign _T_3455 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@23185.4 package.scala 96:25:@23186.4]
  assign _T_3491 = _T_3455 ? Mem1D_4_io_output : _T_3490; // @[Mux.scala 31:69:@23267.4]
  assign _T_3452 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@23177.4 package.scala 96:25:@23178.4]
  assign _T_3492 = _T_3452 ? Mem1D_2_io_output : _T_3491; // @[Mux.scala 31:69:@23268.4]
  assign _T_3449 = RetimeWrapper_io_out; // @[package.scala 96:25:@23169.4 package.scala 96:25:@23170.4]
  assign _T_3586 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@23393.4 package.scala 96:25:@23394.4]
  assign _T_3590 = _T_3586 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@23403.4]
  assign _T_3583 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@23385.4 package.scala 96:25:@23386.4]
  assign _T_3591 = _T_3583 ? Mem1D_19_io_output : _T_3590; // @[Mux.scala 31:69:@23404.4]
  assign _T_3580 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@23377.4 package.scala 96:25:@23378.4]
  assign _T_3592 = _T_3580 ? Mem1D_17_io_output : _T_3591; // @[Mux.scala 31:69:@23405.4]
  assign _T_3577 = RetimeWrapper_19_io_out; // @[package.scala 96:25:@23369.4 package.scala 96:25:@23370.4]
  assign _T_3593 = _T_3577 ? Mem1D_15_io_output : _T_3592; // @[Mux.scala 31:69:@23406.4]
  assign _T_3574 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@23361.4 package.scala 96:25:@23362.4]
  assign _T_3594 = _T_3574 ? Mem1D_13_io_output : _T_3593; // @[Mux.scala 31:69:@23407.4]
  assign _T_3571 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@23353.4 package.scala 96:25:@23354.4]
  assign _T_3595 = _T_3571 ? Mem1D_11_io_output : _T_3594; // @[Mux.scala 31:69:@23408.4]
  assign _T_3568 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@23345.4 package.scala 96:25:@23346.4]
  assign _T_3596 = _T_3568 ? Mem1D_9_io_output : _T_3595; // @[Mux.scala 31:69:@23409.4]
  assign _T_3565 = RetimeWrapper_15_io_out; // @[package.scala 96:25:@23337.4 package.scala 96:25:@23338.4]
  assign _T_3597 = _T_3565 ? Mem1D_7_io_output : _T_3596; // @[Mux.scala 31:69:@23410.4]
  assign _T_3562 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@23329.4 package.scala 96:25:@23330.4]
  assign _T_3598 = _T_3562 ? Mem1D_5_io_output : _T_3597; // @[Mux.scala 31:69:@23411.4]
  assign _T_3559 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@23321.4 package.scala 96:25:@23322.4]
  assign _T_3599 = _T_3559 ? Mem1D_3_io_output : _T_3598; // @[Mux.scala 31:69:@23412.4]
  assign _T_3556 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@23313.4 package.scala 96:25:@23314.4]
  assign _T_3693 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@23537.4 package.scala 96:25:@23538.4]
  assign _T_3697 = _T_3693 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@23547.4]
  assign _T_3690 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@23529.4 package.scala 96:25:@23530.4]
  assign _T_3698 = _T_3690 ? Mem1D_18_io_output : _T_3697; // @[Mux.scala 31:69:@23548.4]
  assign _T_3687 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@23521.4 package.scala 96:25:@23522.4]
  assign _T_3699 = _T_3687 ? Mem1D_16_io_output : _T_3698; // @[Mux.scala 31:69:@23549.4]
  assign _T_3684 = RetimeWrapper_31_io_out; // @[package.scala 96:25:@23513.4 package.scala 96:25:@23514.4]
  assign _T_3700 = _T_3684 ? Mem1D_14_io_output : _T_3699; // @[Mux.scala 31:69:@23550.4]
  assign _T_3681 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@23505.4 package.scala 96:25:@23506.4]
  assign _T_3701 = _T_3681 ? Mem1D_12_io_output : _T_3700; // @[Mux.scala 31:69:@23551.4]
  assign _T_3678 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@23497.4 package.scala 96:25:@23498.4]
  assign _T_3702 = _T_3678 ? Mem1D_10_io_output : _T_3701; // @[Mux.scala 31:69:@23552.4]
  assign _T_3675 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@23489.4 package.scala 96:25:@23490.4]
  assign _T_3703 = _T_3675 ? Mem1D_8_io_output : _T_3702; // @[Mux.scala 31:69:@23553.4]
  assign _T_3672 = RetimeWrapper_27_io_out; // @[package.scala 96:25:@23481.4 package.scala 96:25:@23482.4]
  assign _T_3704 = _T_3672 ? Mem1D_6_io_output : _T_3703; // @[Mux.scala 31:69:@23554.4]
  assign _T_3669 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@23473.4 package.scala 96:25:@23474.4]
  assign _T_3705 = _T_3669 ? Mem1D_4_io_output : _T_3704; // @[Mux.scala 31:69:@23555.4]
  assign _T_3666 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@23465.4 package.scala 96:25:@23466.4]
  assign _T_3706 = _T_3666 ? Mem1D_2_io_output : _T_3705; // @[Mux.scala 31:69:@23556.4]
  assign _T_3663 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@23457.4 package.scala 96:25:@23458.4]
  assign _T_3800 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@23681.4 package.scala 96:25:@23682.4]
  assign _T_3804 = _T_3800 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@23691.4]
  assign _T_3797 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@23673.4 package.scala 96:25:@23674.4]
  assign _T_3805 = _T_3797 ? Mem1D_19_io_output : _T_3804; // @[Mux.scala 31:69:@23692.4]
  assign _T_3794 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@23665.4 package.scala 96:25:@23666.4]
  assign _T_3806 = _T_3794 ? Mem1D_17_io_output : _T_3805; // @[Mux.scala 31:69:@23693.4]
  assign _T_3791 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@23657.4 package.scala 96:25:@23658.4]
  assign _T_3807 = _T_3791 ? Mem1D_15_io_output : _T_3806; // @[Mux.scala 31:69:@23694.4]
  assign _T_3788 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@23649.4 package.scala 96:25:@23650.4]
  assign _T_3808 = _T_3788 ? Mem1D_13_io_output : _T_3807; // @[Mux.scala 31:69:@23695.4]
  assign _T_3785 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@23641.4 package.scala 96:25:@23642.4]
  assign _T_3809 = _T_3785 ? Mem1D_11_io_output : _T_3808; // @[Mux.scala 31:69:@23696.4]
  assign _T_3782 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@23633.4 package.scala 96:25:@23634.4]
  assign _T_3810 = _T_3782 ? Mem1D_9_io_output : _T_3809; // @[Mux.scala 31:69:@23697.4]
  assign _T_3779 = RetimeWrapper_39_io_out; // @[package.scala 96:25:@23625.4 package.scala 96:25:@23626.4]
  assign _T_3811 = _T_3779 ? Mem1D_7_io_output : _T_3810; // @[Mux.scala 31:69:@23698.4]
  assign _T_3776 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@23617.4 package.scala 96:25:@23618.4]
  assign _T_3812 = _T_3776 ? Mem1D_5_io_output : _T_3811; // @[Mux.scala 31:69:@23699.4]
  assign _T_3773 = RetimeWrapper_37_io_out; // @[package.scala 96:25:@23609.4 package.scala 96:25:@23610.4]
  assign _T_3813 = _T_3773 ? Mem1D_3_io_output : _T_3812; // @[Mux.scala 31:69:@23700.4]
  assign _T_3770 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@23601.4 package.scala 96:25:@23602.4]
  assign _T_3907 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@23825.4 package.scala 96:25:@23826.4]
  assign _T_3911 = _T_3907 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@23835.4]
  assign _T_3904 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@23817.4 package.scala 96:25:@23818.4]
  assign _T_3912 = _T_3904 ? Mem1D_18_io_output : _T_3911; // @[Mux.scala 31:69:@23836.4]
  assign _T_3901 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@23809.4 package.scala 96:25:@23810.4]
  assign _T_3913 = _T_3901 ? Mem1D_16_io_output : _T_3912; // @[Mux.scala 31:69:@23837.4]
  assign _T_3898 = RetimeWrapper_55_io_out; // @[package.scala 96:25:@23801.4 package.scala 96:25:@23802.4]
  assign _T_3914 = _T_3898 ? Mem1D_14_io_output : _T_3913; // @[Mux.scala 31:69:@23838.4]
  assign _T_3895 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@23793.4 package.scala 96:25:@23794.4]
  assign _T_3915 = _T_3895 ? Mem1D_12_io_output : _T_3914; // @[Mux.scala 31:69:@23839.4]
  assign _T_3892 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@23785.4 package.scala 96:25:@23786.4]
  assign _T_3916 = _T_3892 ? Mem1D_10_io_output : _T_3915; // @[Mux.scala 31:69:@23840.4]
  assign _T_3889 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@23777.4 package.scala 96:25:@23778.4]
  assign _T_3917 = _T_3889 ? Mem1D_8_io_output : _T_3916; // @[Mux.scala 31:69:@23841.4]
  assign _T_3886 = RetimeWrapper_51_io_out; // @[package.scala 96:25:@23769.4 package.scala 96:25:@23770.4]
  assign _T_3918 = _T_3886 ? Mem1D_6_io_output : _T_3917; // @[Mux.scala 31:69:@23842.4]
  assign _T_3883 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@23761.4 package.scala 96:25:@23762.4]
  assign _T_3919 = _T_3883 ? Mem1D_4_io_output : _T_3918; // @[Mux.scala 31:69:@23843.4]
  assign _T_3880 = RetimeWrapper_49_io_out; // @[package.scala 96:25:@23753.4 package.scala 96:25:@23754.4]
  assign _T_3920 = _T_3880 ? Mem1D_2_io_output : _T_3919; // @[Mux.scala 31:69:@23844.4]
  assign _T_3877 = RetimeWrapper_48_io_out; // @[package.scala 96:25:@23745.4 package.scala 96:25:@23746.4]
  assign _T_4014 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@23969.4 package.scala 96:25:@23970.4]
  assign _T_4018 = _T_4014 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@23979.4]
  assign _T_4011 = RetimeWrapper_69_io_out; // @[package.scala 96:25:@23961.4 package.scala 96:25:@23962.4]
  assign _T_4019 = _T_4011 ? Mem1D_19_io_output : _T_4018; // @[Mux.scala 31:69:@23980.4]
  assign _T_4008 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@23953.4 package.scala 96:25:@23954.4]
  assign _T_4020 = _T_4008 ? Mem1D_17_io_output : _T_4019; // @[Mux.scala 31:69:@23981.4]
  assign _T_4005 = RetimeWrapper_67_io_out; // @[package.scala 96:25:@23945.4 package.scala 96:25:@23946.4]
  assign _T_4021 = _T_4005 ? Mem1D_15_io_output : _T_4020; // @[Mux.scala 31:69:@23982.4]
  assign _T_4002 = RetimeWrapper_66_io_out; // @[package.scala 96:25:@23937.4 package.scala 96:25:@23938.4]
  assign _T_4022 = _T_4002 ? Mem1D_13_io_output : _T_4021; // @[Mux.scala 31:69:@23983.4]
  assign _T_3999 = RetimeWrapper_65_io_out; // @[package.scala 96:25:@23929.4 package.scala 96:25:@23930.4]
  assign _T_4023 = _T_3999 ? Mem1D_11_io_output : _T_4022; // @[Mux.scala 31:69:@23984.4]
  assign _T_3996 = RetimeWrapper_64_io_out; // @[package.scala 96:25:@23921.4 package.scala 96:25:@23922.4]
  assign _T_4024 = _T_3996 ? Mem1D_9_io_output : _T_4023; // @[Mux.scala 31:69:@23985.4]
  assign _T_3993 = RetimeWrapper_63_io_out; // @[package.scala 96:25:@23913.4 package.scala 96:25:@23914.4]
  assign _T_4025 = _T_3993 ? Mem1D_7_io_output : _T_4024; // @[Mux.scala 31:69:@23986.4]
  assign _T_3990 = RetimeWrapper_62_io_out; // @[package.scala 96:25:@23905.4 package.scala 96:25:@23906.4]
  assign _T_4026 = _T_3990 ? Mem1D_5_io_output : _T_4025; // @[Mux.scala 31:69:@23987.4]
  assign _T_3987 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@23897.4 package.scala 96:25:@23898.4]
  assign _T_4027 = _T_3987 ? Mem1D_3_io_output : _T_4026; // @[Mux.scala 31:69:@23988.4]
  assign _T_3984 = RetimeWrapper_60_io_out; // @[package.scala 96:25:@23889.4 package.scala 96:25:@23890.4]
  assign _T_4121 = RetimeWrapper_82_io_out; // @[package.scala 96:25:@24113.4 package.scala 96:25:@24114.4]
  assign _T_4125 = _T_4121 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@24123.4]
  assign _T_4118 = RetimeWrapper_81_io_out; // @[package.scala 96:25:@24105.4 package.scala 96:25:@24106.4]
  assign _T_4126 = _T_4118 ? Mem1D_19_io_output : _T_4125; // @[Mux.scala 31:69:@24124.4]
  assign _T_4115 = RetimeWrapper_80_io_out; // @[package.scala 96:25:@24097.4 package.scala 96:25:@24098.4]
  assign _T_4127 = _T_4115 ? Mem1D_17_io_output : _T_4126; // @[Mux.scala 31:69:@24125.4]
  assign _T_4112 = RetimeWrapper_79_io_out; // @[package.scala 96:25:@24089.4 package.scala 96:25:@24090.4]
  assign _T_4128 = _T_4112 ? Mem1D_15_io_output : _T_4127; // @[Mux.scala 31:69:@24126.4]
  assign _T_4109 = RetimeWrapper_78_io_out; // @[package.scala 96:25:@24081.4 package.scala 96:25:@24082.4]
  assign _T_4129 = _T_4109 ? Mem1D_13_io_output : _T_4128; // @[Mux.scala 31:69:@24127.4]
  assign _T_4106 = RetimeWrapper_77_io_out; // @[package.scala 96:25:@24073.4 package.scala 96:25:@24074.4]
  assign _T_4130 = _T_4106 ? Mem1D_11_io_output : _T_4129; // @[Mux.scala 31:69:@24128.4]
  assign _T_4103 = RetimeWrapper_76_io_out; // @[package.scala 96:25:@24065.4 package.scala 96:25:@24066.4]
  assign _T_4131 = _T_4103 ? Mem1D_9_io_output : _T_4130; // @[Mux.scala 31:69:@24129.4]
  assign _T_4100 = RetimeWrapper_75_io_out; // @[package.scala 96:25:@24057.4 package.scala 96:25:@24058.4]
  assign _T_4132 = _T_4100 ? Mem1D_7_io_output : _T_4131; // @[Mux.scala 31:69:@24130.4]
  assign _T_4097 = RetimeWrapper_74_io_out; // @[package.scala 96:25:@24049.4 package.scala 96:25:@24050.4]
  assign _T_4133 = _T_4097 ? Mem1D_5_io_output : _T_4132; // @[Mux.scala 31:69:@24131.4]
  assign _T_4094 = RetimeWrapper_73_io_out; // @[package.scala 96:25:@24041.4 package.scala 96:25:@24042.4]
  assign _T_4134 = _T_4094 ? Mem1D_3_io_output : _T_4133; // @[Mux.scala 31:69:@24132.4]
  assign _T_4091 = RetimeWrapper_72_io_out; // @[package.scala 96:25:@24033.4 package.scala 96:25:@24034.4]
  assign _T_4228 = RetimeWrapper_94_io_out; // @[package.scala 96:25:@24257.4 package.scala 96:25:@24258.4]
  assign _T_4232 = _T_4228 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@24267.4]
  assign _T_4225 = RetimeWrapper_93_io_out; // @[package.scala 96:25:@24249.4 package.scala 96:25:@24250.4]
  assign _T_4233 = _T_4225 ? Mem1D_18_io_output : _T_4232; // @[Mux.scala 31:69:@24268.4]
  assign _T_4222 = RetimeWrapper_92_io_out; // @[package.scala 96:25:@24241.4 package.scala 96:25:@24242.4]
  assign _T_4234 = _T_4222 ? Mem1D_16_io_output : _T_4233; // @[Mux.scala 31:69:@24269.4]
  assign _T_4219 = RetimeWrapper_91_io_out; // @[package.scala 96:25:@24233.4 package.scala 96:25:@24234.4]
  assign _T_4235 = _T_4219 ? Mem1D_14_io_output : _T_4234; // @[Mux.scala 31:69:@24270.4]
  assign _T_4216 = RetimeWrapper_90_io_out; // @[package.scala 96:25:@24225.4 package.scala 96:25:@24226.4]
  assign _T_4236 = _T_4216 ? Mem1D_12_io_output : _T_4235; // @[Mux.scala 31:69:@24271.4]
  assign _T_4213 = RetimeWrapper_89_io_out; // @[package.scala 96:25:@24217.4 package.scala 96:25:@24218.4]
  assign _T_4237 = _T_4213 ? Mem1D_10_io_output : _T_4236; // @[Mux.scala 31:69:@24272.4]
  assign _T_4210 = RetimeWrapper_88_io_out; // @[package.scala 96:25:@24209.4 package.scala 96:25:@24210.4]
  assign _T_4238 = _T_4210 ? Mem1D_8_io_output : _T_4237; // @[Mux.scala 31:69:@24273.4]
  assign _T_4207 = RetimeWrapper_87_io_out; // @[package.scala 96:25:@24201.4 package.scala 96:25:@24202.4]
  assign _T_4239 = _T_4207 ? Mem1D_6_io_output : _T_4238; // @[Mux.scala 31:69:@24274.4]
  assign _T_4204 = RetimeWrapper_86_io_out; // @[package.scala 96:25:@24193.4 package.scala 96:25:@24194.4]
  assign _T_4240 = _T_4204 ? Mem1D_4_io_output : _T_4239; // @[Mux.scala 31:69:@24275.4]
  assign _T_4201 = RetimeWrapper_85_io_out; // @[package.scala 96:25:@24185.4 package.scala 96:25:@24186.4]
  assign _T_4241 = _T_4201 ? Mem1D_2_io_output : _T_4240; // @[Mux.scala 31:69:@24276.4]
  assign _T_4198 = RetimeWrapper_84_io_out; // @[package.scala 96:25:@24177.4 package.scala 96:25:@24178.4]
  assign _T_4335 = RetimeWrapper_106_io_out; // @[package.scala 96:25:@24401.4 package.scala 96:25:@24402.4]
  assign _T_4339 = _T_4335 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@24411.4]
  assign _T_4332 = RetimeWrapper_105_io_out; // @[package.scala 96:25:@24393.4 package.scala 96:25:@24394.4]
  assign _T_4340 = _T_4332 ? Mem1D_18_io_output : _T_4339; // @[Mux.scala 31:69:@24412.4]
  assign _T_4329 = RetimeWrapper_104_io_out; // @[package.scala 96:25:@24385.4 package.scala 96:25:@24386.4]
  assign _T_4341 = _T_4329 ? Mem1D_16_io_output : _T_4340; // @[Mux.scala 31:69:@24413.4]
  assign _T_4326 = RetimeWrapper_103_io_out; // @[package.scala 96:25:@24377.4 package.scala 96:25:@24378.4]
  assign _T_4342 = _T_4326 ? Mem1D_14_io_output : _T_4341; // @[Mux.scala 31:69:@24414.4]
  assign _T_4323 = RetimeWrapper_102_io_out; // @[package.scala 96:25:@24369.4 package.scala 96:25:@24370.4]
  assign _T_4343 = _T_4323 ? Mem1D_12_io_output : _T_4342; // @[Mux.scala 31:69:@24415.4]
  assign _T_4320 = RetimeWrapper_101_io_out; // @[package.scala 96:25:@24361.4 package.scala 96:25:@24362.4]
  assign _T_4344 = _T_4320 ? Mem1D_10_io_output : _T_4343; // @[Mux.scala 31:69:@24416.4]
  assign _T_4317 = RetimeWrapper_100_io_out; // @[package.scala 96:25:@24353.4 package.scala 96:25:@24354.4]
  assign _T_4345 = _T_4317 ? Mem1D_8_io_output : _T_4344; // @[Mux.scala 31:69:@24417.4]
  assign _T_4314 = RetimeWrapper_99_io_out; // @[package.scala 96:25:@24345.4 package.scala 96:25:@24346.4]
  assign _T_4346 = _T_4314 ? Mem1D_6_io_output : _T_4345; // @[Mux.scala 31:69:@24418.4]
  assign _T_4311 = RetimeWrapper_98_io_out; // @[package.scala 96:25:@24337.4 package.scala 96:25:@24338.4]
  assign _T_4347 = _T_4311 ? Mem1D_4_io_output : _T_4346; // @[Mux.scala 31:69:@24419.4]
  assign _T_4308 = RetimeWrapper_97_io_out; // @[package.scala 96:25:@24329.4 package.scala 96:25:@24330.4]
  assign _T_4348 = _T_4308 ? Mem1D_2_io_output : _T_4347; // @[Mux.scala 31:69:@24420.4]
  assign _T_4305 = RetimeWrapper_96_io_out; // @[package.scala 96:25:@24321.4 package.scala 96:25:@24322.4]
  assign _T_4442 = RetimeWrapper_118_io_out; // @[package.scala 96:25:@24545.4 package.scala 96:25:@24546.4]
  assign _T_4446 = _T_4442 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@24555.4]
  assign _T_4439 = RetimeWrapper_117_io_out; // @[package.scala 96:25:@24537.4 package.scala 96:25:@24538.4]
  assign _T_4447 = _T_4439 ? Mem1D_19_io_output : _T_4446; // @[Mux.scala 31:69:@24556.4]
  assign _T_4436 = RetimeWrapper_116_io_out; // @[package.scala 96:25:@24529.4 package.scala 96:25:@24530.4]
  assign _T_4448 = _T_4436 ? Mem1D_17_io_output : _T_4447; // @[Mux.scala 31:69:@24557.4]
  assign _T_4433 = RetimeWrapper_115_io_out; // @[package.scala 96:25:@24521.4 package.scala 96:25:@24522.4]
  assign _T_4449 = _T_4433 ? Mem1D_15_io_output : _T_4448; // @[Mux.scala 31:69:@24558.4]
  assign _T_4430 = RetimeWrapper_114_io_out; // @[package.scala 96:25:@24513.4 package.scala 96:25:@24514.4]
  assign _T_4450 = _T_4430 ? Mem1D_13_io_output : _T_4449; // @[Mux.scala 31:69:@24559.4]
  assign _T_4427 = RetimeWrapper_113_io_out; // @[package.scala 96:25:@24505.4 package.scala 96:25:@24506.4]
  assign _T_4451 = _T_4427 ? Mem1D_11_io_output : _T_4450; // @[Mux.scala 31:69:@24560.4]
  assign _T_4424 = RetimeWrapper_112_io_out; // @[package.scala 96:25:@24497.4 package.scala 96:25:@24498.4]
  assign _T_4452 = _T_4424 ? Mem1D_9_io_output : _T_4451; // @[Mux.scala 31:69:@24561.4]
  assign _T_4421 = RetimeWrapper_111_io_out; // @[package.scala 96:25:@24489.4 package.scala 96:25:@24490.4]
  assign _T_4453 = _T_4421 ? Mem1D_7_io_output : _T_4452; // @[Mux.scala 31:69:@24562.4]
  assign _T_4418 = RetimeWrapper_110_io_out; // @[package.scala 96:25:@24481.4 package.scala 96:25:@24482.4]
  assign _T_4454 = _T_4418 ? Mem1D_5_io_output : _T_4453; // @[Mux.scala 31:69:@24563.4]
  assign _T_4415 = RetimeWrapper_109_io_out; // @[package.scala 96:25:@24473.4 package.scala 96:25:@24474.4]
  assign _T_4455 = _T_4415 ? Mem1D_3_io_output : _T_4454; // @[Mux.scala 31:69:@24564.4]
  assign _T_4412 = RetimeWrapper_108_io_out; // @[package.scala 96:25:@24465.4 package.scala 96:25:@24466.4]
  assign _T_4549 = RetimeWrapper_130_io_out; // @[package.scala 96:25:@24689.4 package.scala 96:25:@24690.4]
  assign _T_4553 = _T_4549 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@24699.4]
  assign _T_4546 = RetimeWrapper_129_io_out; // @[package.scala 96:25:@24681.4 package.scala 96:25:@24682.4]
  assign _T_4554 = _T_4546 ? Mem1D_18_io_output : _T_4553; // @[Mux.scala 31:69:@24700.4]
  assign _T_4543 = RetimeWrapper_128_io_out; // @[package.scala 96:25:@24673.4 package.scala 96:25:@24674.4]
  assign _T_4555 = _T_4543 ? Mem1D_16_io_output : _T_4554; // @[Mux.scala 31:69:@24701.4]
  assign _T_4540 = RetimeWrapper_127_io_out; // @[package.scala 96:25:@24665.4 package.scala 96:25:@24666.4]
  assign _T_4556 = _T_4540 ? Mem1D_14_io_output : _T_4555; // @[Mux.scala 31:69:@24702.4]
  assign _T_4537 = RetimeWrapper_126_io_out; // @[package.scala 96:25:@24657.4 package.scala 96:25:@24658.4]
  assign _T_4557 = _T_4537 ? Mem1D_12_io_output : _T_4556; // @[Mux.scala 31:69:@24703.4]
  assign _T_4534 = RetimeWrapper_125_io_out; // @[package.scala 96:25:@24649.4 package.scala 96:25:@24650.4]
  assign _T_4558 = _T_4534 ? Mem1D_10_io_output : _T_4557; // @[Mux.scala 31:69:@24704.4]
  assign _T_4531 = RetimeWrapper_124_io_out; // @[package.scala 96:25:@24641.4 package.scala 96:25:@24642.4]
  assign _T_4559 = _T_4531 ? Mem1D_8_io_output : _T_4558; // @[Mux.scala 31:69:@24705.4]
  assign _T_4528 = RetimeWrapper_123_io_out; // @[package.scala 96:25:@24633.4 package.scala 96:25:@24634.4]
  assign _T_4560 = _T_4528 ? Mem1D_6_io_output : _T_4559; // @[Mux.scala 31:69:@24706.4]
  assign _T_4525 = RetimeWrapper_122_io_out; // @[package.scala 96:25:@24625.4 package.scala 96:25:@24626.4]
  assign _T_4561 = _T_4525 ? Mem1D_4_io_output : _T_4560; // @[Mux.scala 31:69:@24707.4]
  assign _T_4522 = RetimeWrapper_121_io_out; // @[package.scala 96:25:@24617.4 package.scala 96:25:@24618.4]
  assign _T_4562 = _T_4522 ? Mem1D_2_io_output : _T_4561; // @[Mux.scala 31:69:@24708.4]
  assign _T_4519 = RetimeWrapper_120_io_out; // @[package.scala 96:25:@24609.4 package.scala 96:25:@24610.4]
  assign _T_4656 = RetimeWrapper_142_io_out; // @[package.scala 96:25:@24833.4 package.scala 96:25:@24834.4]
  assign _T_4660 = _T_4656 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@24843.4]
  assign _T_4653 = RetimeWrapper_141_io_out; // @[package.scala 96:25:@24825.4 package.scala 96:25:@24826.4]
  assign _T_4661 = _T_4653 ? Mem1D_18_io_output : _T_4660; // @[Mux.scala 31:69:@24844.4]
  assign _T_4650 = RetimeWrapper_140_io_out; // @[package.scala 96:25:@24817.4 package.scala 96:25:@24818.4]
  assign _T_4662 = _T_4650 ? Mem1D_16_io_output : _T_4661; // @[Mux.scala 31:69:@24845.4]
  assign _T_4647 = RetimeWrapper_139_io_out; // @[package.scala 96:25:@24809.4 package.scala 96:25:@24810.4]
  assign _T_4663 = _T_4647 ? Mem1D_14_io_output : _T_4662; // @[Mux.scala 31:69:@24846.4]
  assign _T_4644 = RetimeWrapper_138_io_out; // @[package.scala 96:25:@24801.4 package.scala 96:25:@24802.4]
  assign _T_4664 = _T_4644 ? Mem1D_12_io_output : _T_4663; // @[Mux.scala 31:69:@24847.4]
  assign _T_4641 = RetimeWrapper_137_io_out; // @[package.scala 96:25:@24793.4 package.scala 96:25:@24794.4]
  assign _T_4665 = _T_4641 ? Mem1D_10_io_output : _T_4664; // @[Mux.scala 31:69:@24848.4]
  assign _T_4638 = RetimeWrapper_136_io_out; // @[package.scala 96:25:@24785.4 package.scala 96:25:@24786.4]
  assign _T_4666 = _T_4638 ? Mem1D_8_io_output : _T_4665; // @[Mux.scala 31:69:@24849.4]
  assign _T_4635 = RetimeWrapper_135_io_out; // @[package.scala 96:25:@24777.4 package.scala 96:25:@24778.4]
  assign _T_4667 = _T_4635 ? Mem1D_6_io_output : _T_4666; // @[Mux.scala 31:69:@24850.4]
  assign _T_4632 = RetimeWrapper_134_io_out; // @[package.scala 96:25:@24769.4 package.scala 96:25:@24770.4]
  assign _T_4668 = _T_4632 ? Mem1D_4_io_output : _T_4667; // @[Mux.scala 31:69:@24851.4]
  assign _T_4629 = RetimeWrapper_133_io_out; // @[package.scala 96:25:@24761.4 package.scala 96:25:@24762.4]
  assign _T_4669 = _T_4629 ? Mem1D_2_io_output : _T_4668; // @[Mux.scala 31:69:@24852.4]
  assign _T_4626 = RetimeWrapper_132_io_out; // @[package.scala 96:25:@24753.4 package.scala 96:25:@24754.4]
  assign _T_4763 = RetimeWrapper_154_io_out; // @[package.scala 96:25:@24977.4 package.scala 96:25:@24978.4]
  assign _T_4767 = _T_4763 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@24987.4]
  assign _T_4760 = RetimeWrapper_153_io_out; // @[package.scala 96:25:@24969.4 package.scala 96:25:@24970.4]
  assign _T_4768 = _T_4760 ? Mem1D_19_io_output : _T_4767; // @[Mux.scala 31:69:@24988.4]
  assign _T_4757 = RetimeWrapper_152_io_out; // @[package.scala 96:25:@24961.4 package.scala 96:25:@24962.4]
  assign _T_4769 = _T_4757 ? Mem1D_17_io_output : _T_4768; // @[Mux.scala 31:69:@24989.4]
  assign _T_4754 = RetimeWrapper_151_io_out; // @[package.scala 96:25:@24953.4 package.scala 96:25:@24954.4]
  assign _T_4770 = _T_4754 ? Mem1D_15_io_output : _T_4769; // @[Mux.scala 31:69:@24990.4]
  assign _T_4751 = RetimeWrapper_150_io_out; // @[package.scala 96:25:@24945.4 package.scala 96:25:@24946.4]
  assign _T_4771 = _T_4751 ? Mem1D_13_io_output : _T_4770; // @[Mux.scala 31:69:@24991.4]
  assign _T_4748 = RetimeWrapper_149_io_out; // @[package.scala 96:25:@24937.4 package.scala 96:25:@24938.4]
  assign _T_4772 = _T_4748 ? Mem1D_11_io_output : _T_4771; // @[Mux.scala 31:69:@24992.4]
  assign _T_4745 = RetimeWrapper_148_io_out; // @[package.scala 96:25:@24929.4 package.scala 96:25:@24930.4]
  assign _T_4773 = _T_4745 ? Mem1D_9_io_output : _T_4772; // @[Mux.scala 31:69:@24993.4]
  assign _T_4742 = RetimeWrapper_147_io_out; // @[package.scala 96:25:@24921.4 package.scala 96:25:@24922.4]
  assign _T_4774 = _T_4742 ? Mem1D_7_io_output : _T_4773; // @[Mux.scala 31:69:@24994.4]
  assign _T_4739 = RetimeWrapper_146_io_out; // @[package.scala 96:25:@24913.4 package.scala 96:25:@24914.4]
  assign _T_4775 = _T_4739 ? Mem1D_5_io_output : _T_4774; // @[Mux.scala 31:69:@24995.4]
  assign _T_4736 = RetimeWrapper_145_io_out; // @[package.scala 96:25:@24905.4 package.scala 96:25:@24906.4]
  assign _T_4776 = _T_4736 ? Mem1D_3_io_output : _T_4775; // @[Mux.scala 31:69:@24996.4]
  assign _T_4733 = RetimeWrapper_144_io_out; // @[package.scala 96:25:@24897.4 package.scala 96:25:@24898.4]
  assign _T_4870 = RetimeWrapper_166_io_out; // @[package.scala 96:25:@25121.4 package.scala 96:25:@25122.4]
  assign _T_4874 = _T_4870 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@25131.4]
  assign _T_4867 = RetimeWrapper_165_io_out; // @[package.scala 96:25:@25113.4 package.scala 96:25:@25114.4]
  assign _T_4875 = _T_4867 ? Mem1D_19_io_output : _T_4874; // @[Mux.scala 31:69:@25132.4]
  assign _T_4864 = RetimeWrapper_164_io_out; // @[package.scala 96:25:@25105.4 package.scala 96:25:@25106.4]
  assign _T_4876 = _T_4864 ? Mem1D_17_io_output : _T_4875; // @[Mux.scala 31:69:@25133.4]
  assign _T_4861 = RetimeWrapper_163_io_out; // @[package.scala 96:25:@25097.4 package.scala 96:25:@25098.4]
  assign _T_4877 = _T_4861 ? Mem1D_15_io_output : _T_4876; // @[Mux.scala 31:69:@25134.4]
  assign _T_4858 = RetimeWrapper_162_io_out; // @[package.scala 96:25:@25089.4 package.scala 96:25:@25090.4]
  assign _T_4878 = _T_4858 ? Mem1D_13_io_output : _T_4877; // @[Mux.scala 31:69:@25135.4]
  assign _T_4855 = RetimeWrapper_161_io_out; // @[package.scala 96:25:@25081.4 package.scala 96:25:@25082.4]
  assign _T_4879 = _T_4855 ? Mem1D_11_io_output : _T_4878; // @[Mux.scala 31:69:@25136.4]
  assign _T_4852 = RetimeWrapper_160_io_out; // @[package.scala 96:25:@25073.4 package.scala 96:25:@25074.4]
  assign _T_4880 = _T_4852 ? Mem1D_9_io_output : _T_4879; // @[Mux.scala 31:69:@25137.4]
  assign _T_4849 = RetimeWrapper_159_io_out; // @[package.scala 96:25:@25065.4 package.scala 96:25:@25066.4]
  assign _T_4881 = _T_4849 ? Mem1D_7_io_output : _T_4880; // @[Mux.scala 31:69:@25138.4]
  assign _T_4846 = RetimeWrapper_158_io_out; // @[package.scala 96:25:@25057.4 package.scala 96:25:@25058.4]
  assign _T_4882 = _T_4846 ? Mem1D_5_io_output : _T_4881; // @[Mux.scala 31:69:@25139.4]
  assign _T_4843 = RetimeWrapper_157_io_out; // @[package.scala 96:25:@25049.4 package.scala 96:25:@25050.4]
  assign _T_4883 = _T_4843 ? Mem1D_3_io_output : _T_4882; // @[Mux.scala 31:69:@25140.4]
  assign _T_4840 = RetimeWrapper_156_io_out; // @[package.scala 96:25:@25041.4 package.scala 96:25:@25042.4]
  assign _T_4977 = RetimeWrapper_178_io_out; // @[package.scala 96:25:@25265.4 package.scala 96:25:@25266.4]
  assign _T_4981 = _T_4977 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@25275.4]
  assign _T_4974 = RetimeWrapper_177_io_out; // @[package.scala 96:25:@25257.4 package.scala 96:25:@25258.4]
  assign _T_4982 = _T_4974 ? Mem1D_19_io_output : _T_4981; // @[Mux.scala 31:69:@25276.4]
  assign _T_4971 = RetimeWrapper_176_io_out; // @[package.scala 96:25:@25249.4 package.scala 96:25:@25250.4]
  assign _T_4983 = _T_4971 ? Mem1D_17_io_output : _T_4982; // @[Mux.scala 31:69:@25277.4]
  assign _T_4968 = RetimeWrapper_175_io_out; // @[package.scala 96:25:@25241.4 package.scala 96:25:@25242.4]
  assign _T_4984 = _T_4968 ? Mem1D_15_io_output : _T_4983; // @[Mux.scala 31:69:@25278.4]
  assign _T_4965 = RetimeWrapper_174_io_out; // @[package.scala 96:25:@25233.4 package.scala 96:25:@25234.4]
  assign _T_4985 = _T_4965 ? Mem1D_13_io_output : _T_4984; // @[Mux.scala 31:69:@25279.4]
  assign _T_4962 = RetimeWrapper_173_io_out; // @[package.scala 96:25:@25225.4 package.scala 96:25:@25226.4]
  assign _T_4986 = _T_4962 ? Mem1D_11_io_output : _T_4985; // @[Mux.scala 31:69:@25280.4]
  assign _T_4959 = RetimeWrapper_172_io_out; // @[package.scala 96:25:@25217.4 package.scala 96:25:@25218.4]
  assign _T_4987 = _T_4959 ? Mem1D_9_io_output : _T_4986; // @[Mux.scala 31:69:@25281.4]
  assign _T_4956 = RetimeWrapper_171_io_out; // @[package.scala 96:25:@25209.4 package.scala 96:25:@25210.4]
  assign _T_4988 = _T_4956 ? Mem1D_7_io_output : _T_4987; // @[Mux.scala 31:69:@25282.4]
  assign _T_4953 = RetimeWrapper_170_io_out; // @[package.scala 96:25:@25201.4 package.scala 96:25:@25202.4]
  assign _T_4989 = _T_4953 ? Mem1D_5_io_output : _T_4988; // @[Mux.scala 31:69:@25283.4]
  assign _T_4950 = RetimeWrapper_169_io_out; // @[package.scala 96:25:@25193.4 package.scala 96:25:@25194.4]
  assign _T_4990 = _T_4950 ? Mem1D_3_io_output : _T_4989; // @[Mux.scala 31:69:@25284.4]
  assign _T_4947 = RetimeWrapper_168_io_out; // @[package.scala 96:25:@25185.4 package.scala 96:25:@25186.4]
  assign _T_5084 = RetimeWrapper_190_io_out; // @[package.scala 96:25:@25409.4 package.scala 96:25:@25410.4]
  assign _T_5088 = _T_5084 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@25419.4]
  assign _T_5081 = RetimeWrapper_189_io_out; // @[package.scala 96:25:@25401.4 package.scala 96:25:@25402.4]
  assign _T_5089 = _T_5081 ? Mem1D_18_io_output : _T_5088; // @[Mux.scala 31:69:@25420.4]
  assign _T_5078 = RetimeWrapper_188_io_out; // @[package.scala 96:25:@25393.4 package.scala 96:25:@25394.4]
  assign _T_5090 = _T_5078 ? Mem1D_16_io_output : _T_5089; // @[Mux.scala 31:69:@25421.4]
  assign _T_5075 = RetimeWrapper_187_io_out; // @[package.scala 96:25:@25385.4 package.scala 96:25:@25386.4]
  assign _T_5091 = _T_5075 ? Mem1D_14_io_output : _T_5090; // @[Mux.scala 31:69:@25422.4]
  assign _T_5072 = RetimeWrapper_186_io_out; // @[package.scala 96:25:@25377.4 package.scala 96:25:@25378.4]
  assign _T_5092 = _T_5072 ? Mem1D_12_io_output : _T_5091; // @[Mux.scala 31:69:@25423.4]
  assign _T_5069 = RetimeWrapper_185_io_out; // @[package.scala 96:25:@25369.4 package.scala 96:25:@25370.4]
  assign _T_5093 = _T_5069 ? Mem1D_10_io_output : _T_5092; // @[Mux.scala 31:69:@25424.4]
  assign _T_5066 = RetimeWrapper_184_io_out; // @[package.scala 96:25:@25361.4 package.scala 96:25:@25362.4]
  assign _T_5094 = _T_5066 ? Mem1D_8_io_output : _T_5093; // @[Mux.scala 31:69:@25425.4]
  assign _T_5063 = RetimeWrapper_183_io_out; // @[package.scala 96:25:@25353.4 package.scala 96:25:@25354.4]
  assign _T_5095 = _T_5063 ? Mem1D_6_io_output : _T_5094; // @[Mux.scala 31:69:@25426.4]
  assign _T_5060 = RetimeWrapper_182_io_out; // @[package.scala 96:25:@25345.4 package.scala 96:25:@25346.4]
  assign _T_5096 = _T_5060 ? Mem1D_4_io_output : _T_5095; // @[Mux.scala 31:69:@25427.4]
  assign _T_5057 = RetimeWrapper_181_io_out; // @[package.scala 96:25:@25337.4 package.scala 96:25:@25338.4]
  assign _T_5097 = _T_5057 ? Mem1D_2_io_output : _T_5096; // @[Mux.scala 31:69:@25428.4]
  assign _T_5054 = RetimeWrapper_180_io_out; // @[package.scala 96:25:@25329.4 package.scala 96:25:@25330.4]
  assign _T_5191 = RetimeWrapper_202_io_out; // @[package.scala 96:25:@25553.4 package.scala 96:25:@25554.4]
  assign _T_5195 = _T_5191 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@25563.4]
  assign _T_5188 = RetimeWrapper_201_io_out; // @[package.scala 96:25:@25545.4 package.scala 96:25:@25546.4]
  assign _T_5196 = _T_5188 ? Mem1D_19_io_output : _T_5195; // @[Mux.scala 31:69:@25564.4]
  assign _T_5185 = RetimeWrapper_200_io_out; // @[package.scala 96:25:@25537.4 package.scala 96:25:@25538.4]
  assign _T_5197 = _T_5185 ? Mem1D_17_io_output : _T_5196; // @[Mux.scala 31:69:@25565.4]
  assign _T_5182 = RetimeWrapper_199_io_out; // @[package.scala 96:25:@25529.4 package.scala 96:25:@25530.4]
  assign _T_5198 = _T_5182 ? Mem1D_15_io_output : _T_5197; // @[Mux.scala 31:69:@25566.4]
  assign _T_5179 = RetimeWrapper_198_io_out; // @[package.scala 96:25:@25521.4 package.scala 96:25:@25522.4]
  assign _T_5199 = _T_5179 ? Mem1D_13_io_output : _T_5198; // @[Mux.scala 31:69:@25567.4]
  assign _T_5176 = RetimeWrapper_197_io_out; // @[package.scala 96:25:@25513.4 package.scala 96:25:@25514.4]
  assign _T_5200 = _T_5176 ? Mem1D_11_io_output : _T_5199; // @[Mux.scala 31:69:@25568.4]
  assign _T_5173 = RetimeWrapper_196_io_out; // @[package.scala 96:25:@25505.4 package.scala 96:25:@25506.4]
  assign _T_5201 = _T_5173 ? Mem1D_9_io_output : _T_5200; // @[Mux.scala 31:69:@25569.4]
  assign _T_5170 = RetimeWrapper_195_io_out; // @[package.scala 96:25:@25497.4 package.scala 96:25:@25498.4]
  assign _T_5202 = _T_5170 ? Mem1D_7_io_output : _T_5201; // @[Mux.scala 31:69:@25570.4]
  assign _T_5167 = RetimeWrapper_194_io_out; // @[package.scala 96:25:@25489.4 package.scala 96:25:@25490.4]
  assign _T_5203 = _T_5167 ? Mem1D_5_io_output : _T_5202; // @[Mux.scala 31:69:@25571.4]
  assign _T_5164 = RetimeWrapper_193_io_out; // @[package.scala 96:25:@25481.4 package.scala 96:25:@25482.4]
  assign _T_5204 = _T_5164 ? Mem1D_3_io_output : _T_5203; // @[Mux.scala 31:69:@25572.4]
  assign _T_5161 = RetimeWrapper_192_io_out; // @[package.scala 96:25:@25473.4 package.scala 96:25:@25474.4]
  assign _T_5298 = RetimeWrapper_214_io_out; // @[package.scala 96:25:@25697.4 package.scala 96:25:@25698.4]
  assign _T_5302 = _T_5298 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@25707.4]
  assign _T_5295 = RetimeWrapper_213_io_out; // @[package.scala 96:25:@25689.4 package.scala 96:25:@25690.4]
  assign _T_5303 = _T_5295 ? Mem1D_18_io_output : _T_5302; // @[Mux.scala 31:69:@25708.4]
  assign _T_5292 = RetimeWrapper_212_io_out; // @[package.scala 96:25:@25681.4 package.scala 96:25:@25682.4]
  assign _T_5304 = _T_5292 ? Mem1D_16_io_output : _T_5303; // @[Mux.scala 31:69:@25709.4]
  assign _T_5289 = RetimeWrapper_211_io_out; // @[package.scala 96:25:@25673.4 package.scala 96:25:@25674.4]
  assign _T_5305 = _T_5289 ? Mem1D_14_io_output : _T_5304; // @[Mux.scala 31:69:@25710.4]
  assign _T_5286 = RetimeWrapper_210_io_out; // @[package.scala 96:25:@25665.4 package.scala 96:25:@25666.4]
  assign _T_5306 = _T_5286 ? Mem1D_12_io_output : _T_5305; // @[Mux.scala 31:69:@25711.4]
  assign _T_5283 = RetimeWrapper_209_io_out; // @[package.scala 96:25:@25657.4 package.scala 96:25:@25658.4]
  assign _T_5307 = _T_5283 ? Mem1D_10_io_output : _T_5306; // @[Mux.scala 31:69:@25712.4]
  assign _T_5280 = RetimeWrapper_208_io_out; // @[package.scala 96:25:@25649.4 package.scala 96:25:@25650.4]
  assign _T_5308 = _T_5280 ? Mem1D_8_io_output : _T_5307; // @[Mux.scala 31:69:@25713.4]
  assign _T_5277 = RetimeWrapper_207_io_out; // @[package.scala 96:25:@25641.4 package.scala 96:25:@25642.4]
  assign _T_5309 = _T_5277 ? Mem1D_6_io_output : _T_5308; // @[Mux.scala 31:69:@25714.4]
  assign _T_5274 = RetimeWrapper_206_io_out; // @[package.scala 96:25:@25633.4 package.scala 96:25:@25634.4]
  assign _T_5310 = _T_5274 ? Mem1D_4_io_output : _T_5309; // @[Mux.scala 31:69:@25715.4]
  assign _T_5271 = RetimeWrapper_205_io_out; // @[package.scala 96:25:@25625.4 package.scala 96:25:@25626.4]
  assign _T_5311 = _T_5271 ? Mem1D_2_io_output : _T_5310; // @[Mux.scala 31:69:@25716.4]
  assign _T_5268 = RetimeWrapper_204_io_out; // @[package.scala 96:25:@25617.4 package.scala 96:25:@25618.4]
  assign io_rPort_17_output_0 = _T_5268 ? Mem1D_io_output : _T_5311; // @[MemPrimitives.scala 148:13:@25718.4]
  assign io_rPort_16_output_0 = _T_5161 ? Mem1D_1_io_output : _T_5204; // @[MemPrimitives.scala 148:13:@25574.4]
  assign io_rPort_15_output_0 = _T_5054 ? Mem1D_io_output : _T_5097; // @[MemPrimitives.scala 148:13:@25430.4]
  assign io_rPort_14_output_0 = _T_4947 ? Mem1D_1_io_output : _T_4990; // @[MemPrimitives.scala 148:13:@25286.4]
  assign io_rPort_13_output_0 = _T_4840 ? Mem1D_1_io_output : _T_4883; // @[MemPrimitives.scala 148:13:@25142.4]
  assign io_rPort_12_output_0 = _T_4733 ? Mem1D_1_io_output : _T_4776; // @[MemPrimitives.scala 148:13:@24998.4]
  assign io_rPort_11_output_0 = _T_4626 ? Mem1D_io_output : _T_4669; // @[MemPrimitives.scala 148:13:@24854.4]
  assign io_rPort_10_output_0 = _T_4519 ? Mem1D_io_output : _T_4562; // @[MemPrimitives.scala 148:13:@24710.4]
  assign io_rPort_9_output_0 = _T_4412 ? Mem1D_1_io_output : _T_4455; // @[MemPrimitives.scala 148:13:@24566.4]
  assign io_rPort_8_output_0 = _T_4305 ? Mem1D_io_output : _T_4348; // @[MemPrimitives.scala 148:13:@24422.4]
  assign io_rPort_7_output_0 = _T_4198 ? Mem1D_io_output : _T_4241; // @[MemPrimitives.scala 148:13:@24278.4]
  assign io_rPort_6_output_0 = _T_4091 ? Mem1D_1_io_output : _T_4134; // @[MemPrimitives.scala 148:13:@24134.4]
  assign io_rPort_5_output_0 = _T_3984 ? Mem1D_1_io_output : _T_4027; // @[MemPrimitives.scala 148:13:@23990.4]
  assign io_rPort_4_output_0 = _T_3877 ? Mem1D_io_output : _T_3920; // @[MemPrimitives.scala 148:13:@23846.4]
  assign io_rPort_3_output_0 = _T_3770 ? Mem1D_1_io_output : _T_3813; // @[MemPrimitives.scala 148:13:@23702.4]
  assign io_rPort_2_output_0 = _T_3663 ? Mem1D_io_output : _T_3706; // @[MemPrimitives.scala 148:13:@23558.4]
  assign io_rPort_1_output_0 = _T_3556 ? Mem1D_1_io_output : _T_3599; // @[MemPrimitives.scala 148:13:@23414.4]
  assign io_rPort_0_output_0 = _T_3449 ? Mem1D_io_output : _T_3492; // @[MemPrimitives.scala 148:13:@23270.4]
  assign Mem1D_clock = clock; // @[:@20152.4]
  assign Mem1D_reset = reset; // @[:@20153.4]
  assign Mem1D_io_r_ofs_0 = _T_1267[8:0]; // @[MemPrimitives.scala 127:28:@21077.4]
  assign Mem1D_io_r_backpressure = _T_1267[9]; // @[MemPrimitives.scala 128:32:@21078.4]
  assign Mem1D_io_w_ofs_0 = _T_715[8:0]; // @[MemPrimitives.scala 94:28:@20551.4]
  assign Mem1D_io_w_data_0 = _T_715[16:9]; // @[MemPrimitives.scala 95:29:@20552.4]
  assign Mem1D_io_w_en_0 = _T_715[17]; // @[MemPrimitives.scala 96:27:@20553.4]
  assign Mem1D_1_clock = clock; // @[:@20168.4]
  assign Mem1D_1_reset = reset; // @[:@20169.4]
  assign Mem1D_1_io_r_ofs_0 = _T_1359[8:0]; // @[MemPrimitives.scala 127:28:@21166.4]
  assign Mem1D_1_io_r_backpressure = _T_1359[9]; // @[MemPrimitives.scala 128:32:@21167.4]
  assign Mem1D_1_io_w_ofs_0 = _T_735[8:0]; // @[MemPrimitives.scala 94:28:@20570.4]
  assign Mem1D_1_io_w_data_0 = _T_735[16:9]; // @[MemPrimitives.scala 95:29:@20571.4]
  assign Mem1D_1_io_w_en_0 = _T_735[17]; // @[MemPrimitives.scala 96:27:@20572.4]
  assign Mem1D_2_clock = clock; // @[:@20184.4]
  assign Mem1D_2_reset = reset; // @[:@20185.4]
  assign Mem1D_2_io_r_ofs_0 = _T_1451[8:0]; // @[MemPrimitives.scala 127:28:@21255.4]
  assign Mem1D_2_io_r_backpressure = _T_1451[9]; // @[MemPrimitives.scala 128:32:@21256.4]
  assign Mem1D_2_io_w_ofs_0 = _T_755[8:0]; // @[MemPrimitives.scala 94:28:@20589.4]
  assign Mem1D_2_io_w_data_0 = _T_755[16:9]; // @[MemPrimitives.scala 95:29:@20590.4]
  assign Mem1D_2_io_w_en_0 = _T_755[17]; // @[MemPrimitives.scala 96:27:@20591.4]
  assign Mem1D_3_clock = clock; // @[:@20200.4]
  assign Mem1D_3_reset = reset; // @[:@20201.4]
  assign Mem1D_3_io_r_ofs_0 = _T_1543[8:0]; // @[MemPrimitives.scala 127:28:@21344.4]
  assign Mem1D_3_io_r_backpressure = _T_1543[9]; // @[MemPrimitives.scala 128:32:@21345.4]
  assign Mem1D_3_io_w_ofs_0 = _T_775[8:0]; // @[MemPrimitives.scala 94:28:@20608.4]
  assign Mem1D_3_io_w_data_0 = _T_775[16:9]; // @[MemPrimitives.scala 95:29:@20609.4]
  assign Mem1D_3_io_w_en_0 = _T_775[17]; // @[MemPrimitives.scala 96:27:@20610.4]
  assign Mem1D_4_clock = clock; // @[:@20216.4]
  assign Mem1D_4_reset = reset; // @[:@20217.4]
  assign Mem1D_4_io_r_ofs_0 = _T_1635[8:0]; // @[MemPrimitives.scala 127:28:@21433.4]
  assign Mem1D_4_io_r_backpressure = _T_1635[9]; // @[MemPrimitives.scala 128:32:@21434.4]
  assign Mem1D_4_io_w_ofs_0 = _T_795[8:0]; // @[MemPrimitives.scala 94:28:@20627.4]
  assign Mem1D_4_io_w_data_0 = _T_795[16:9]; // @[MemPrimitives.scala 95:29:@20628.4]
  assign Mem1D_4_io_w_en_0 = _T_795[17]; // @[MemPrimitives.scala 96:27:@20629.4]
  assign Mem1D_5_clock = clock; // @[:@20232.4]
  assign Mem1D_5_reset = reset; // @[:@20233.4]
  assign Mem1D_5_io_r_ofs_0 = _T_1727[8:0]; // @[MemPrimitives.scala 127:28:@21522.4]
  assign Mem1D_5_io_r_backpressure = _T_1727[9]; // @[MemPrimitives.scala 128:32:@21523.4]
  assign Mem1D_5_io_w_ofs_0 = _T_815[8:0]; // @[MemPrimitives.scala 94:28:@20646.4]
  assign Mem1D_5_io_w_data_0 = _T_815[16:9]; // @[MemPrimitives.scala 95:29:@20647.4]
  assign Mem1D_5_io_w_en_0 = _T_815[17]; // @[MemPrimitives.scala 96:27:@20648.4]
  assign Mem1D_6_clock = clock; // @[:@20248.4]
  assign Mem1D_6_reset = reset; // @[:@20249.4]
  assign Mem1D_6_io_r_ofs_0 = _T_1819[8:0]; // @[MemPrimitives.scala 127:28:@21611.4]
  assign Mem1D_6_io_r_backpressure = _T_1819[9]; // @[MemPrimitives.scala 128:32:@21612.4]
  assign Mem1D_6_io_w_ofs_0 = _T_835[8:0]; // @[MemPrimitives.scala 94:28:@20665.4]
  assign Mem1D_6_io_w_data_0 = _T_835[16:9]; // @[MemPrimitives.scala 95:29:@20666.4]
  assign Mem1D_6_io_w_en_0 = _T_835[17]; // @[MemPrimitives.scala 96:27:@20667.4]
  assign Mem1D_7_clock = clock; // @[:@20264.4]
  assign Mem1D_7_reset = reset; // @[:@20265.4]
  assign Mem1D_7_io_r_ofs_0 = _T_1911[8:0]; // @[MemPrimitives.scala 127:28:@21700.4]
  assign Mem1D_7_io_r_backpressure = _T_1911[9]; // @[MemPrimitives.scala 128:32:@21701.4]
  assign Mem1D_7_io_w_ofs_0 = _T_855[8:0]; // @[MemPrimitives.scala 94:28:@20684.4]
  assign Mem1D_7_io_w_data_0 = _T_855[16:9]; // @[MemPrimitives.scala 95:29:@20685.4]
  assign Mem1D_7_io_w_en_0 = _T_855[17]; // @[MemPrimitives.scala 96:27:@20686.4]
  assign Mem1D_8_clock = clock; // @[:@20280.4]
  assign Mem1D_8_reset = reset; // @[:@20281.4]
  assign Mem1D_8_io_r_ofs_0 = _T_2003[8:0]; // @[MemPrimitives.scala 127:28:@21789.4]
  assign Mem1D_8_io_r_backpressure = _T_2003[9]; // @[MemPrimitives.scala 128:32:@21790.4]
  assign Mem1D_8_io_w_ofs_0 = _T_875[8:0]; // @[MemPrimitives.scala 94:28:@20703.4]
  assign Mem1D_8_io_w_data_0 = _T_875[16:9]; // @[MemPrimitives.scala 95:29:@20704.4]
  assign Mem1D_8_io_w_en_0 = _T_875[17]; // @[MemPrimitives.scala 96:27:@20705.4]
  assign Mem1D_9_clock = clock; // @[:@20296.4]
  assign Mem1D_9_reset = reset; // @[:@20297.4]
  assign Mem1D_9_io_r_ofs_0 = _T_2095[8:0]; // @[MemPrimitives.scala 127:28:@21878.4]
  assign Mem1D_9_io_r_backpressure = _T_2095[9]; // @[MemPrimitives.scala 128:32:@21879.4]
  assign Mem1D_9_io_w_ofs_0 = _T_895[8:0]; // @[MemPrimitives.scala 94:28:@20722.4]
  assign Mem1D_9_io_w_data_0 = _T_895[16:9]; // @[MemPrimitives.scala 95:29:@20723.4]
  assign Mem1D_9_io_w_en_0 = _T_895[17]; // @[MemPrimitives.scala 96:27:@20724.4]
  assign Mem1D_10_clock = clock; // @[:@20312.4]
  assign Mem1D_10_reset = reset; // @[:@20313.4]
  assign Mem1D_10_io_r_ofs_0 = _T_2187[8:0]; // @[MemPrimitives.scala 127:28:@21967.4]
  assign Mem1D_10_io_r_backpressure = _T_2187[9]; // @[MemPrimitives.scala 128:32:@21968.4]
  assign Mem1D_10_io_w_ofs_0 = _T_915[8:0]; // @[MemPrimitives.scala 94:28:@20741.4]
  assign Mem1D_10_io_w_data_0 = _T_915[16:9]; // @[MemPrimitives.scala 95:29:@20742.4]
  assign Mem1D_10_io_w_en_0 = _T_915[17]; // @[MemPrimitives.scala 96:27:@20743.4]
  assign Mem1D_11_clock = clock; // @[:@20328.4]
  assign Mem1D_11_reset = reset; // @[:@20329.4]
  assign Mem1D_11_io_r_ofs_0 = _T_2279[8:0]; // @[MemPrimitives.scala 127:28:@22056.4]
  assign Mem1D_11_io_r_backpressure = _T_2279[9]; // @[MemPrimitives.scala 128:32:@22057.4]
  assign Mem1D_11_io_w_ofs_0 = _T_935[8:0]; // @[MemPrimitives.scala 94:28:@20760.4]
  assign Mem1D_11_io_w_data_0 = _T_935[16:9]; // @[MemPrimitives.scala 95:29:@20761.4]
  assign Mem1D_11_io_w_en_0 = _T_935[17]; // @[MemPrimitives.scala 96:27:@20762.4]
  assign Mem1D_12_clock = clock; // @[:@20344.4]
  assign Mem1D_12_reset = reset; // @[:@20345.4]
  assign Mem1D_12_io_r_ofs_0 = _T_2371[8:0]; // @[MemPrimitives.scala 127:28:@22145.4]
  assign Mem1D_12_io_r_backpressure = _T_2371[9]; // @[MemPrimitives.scala 128:32:@22146.4]
  assign Mem1D_12_io_w_ofs_0 = _T_955[8:0]; // @[MemPrimitives.scala 94:28:@20779.4]
  assign Mem1D_12_io_w_data_0 = _T_955[16:9]; // @[MemPrimitives.scala 95:29:@20780.4]
  assign Mem1D_12_io_w_en_0 = _T_955[17]; // @[MemPrimitives.scala 96:27:@20781.4]
  assign Mem1D_13_clock = clock; // @[:@20360.4]
  assign Mem1D_13_reset = reset; // @[:@20361.4]
  assign Mem1D_13_io_r_ofs_0 = _T_2463[8:0]; // @[MemPrimitives.scala 127:28:@22234.4]
  assign Mem1D_13_io_r_backpressure = _T_2463[9]; // @[MemPrimitives.scala 128:32:@22235.4]
  assign Mem1D_13_io_w_ofs_0 = _T_975[8:0]; // @[MemPrimitives.scala 94:28:@20798.4]
  assign Mem1D_13_io_w_data_0 = _T_975[16:9]; // @[MemPrimitives.scala 95:29:@20799.4]
  assign Mem1D_13_io_w_en_0 = _T_975[17]; // @[MemPrimitives.scala 96:27:@20800.4]
  assign Mem1D_14_clock = clock; // @[:@20376.4]
  assign Mem1D_14_reset = reset; // @[:@20377.4]
  assign Mem1D_14_io_r_ofs_0 = _T_2555[8:0]; // @[MemPrimitives.scala 127:28:@22323.4]
  assign Mem1D_14_io_r_backpressure = _T_2555[9]; // @[MemPrimitives.scala 128:32:@22324.4]
  assign Mem1D_14_io_w_ofs_0 = _T_995[8:0]; // @[MemPrimitives.scala 94:28:@20817.4]
  assign Mem1D_14_io_w_data_0 = _T_995[16:9]; // @[MemPrimitives.scala 95:29:@20818.4]
  assign Mem1D_14_io_w_en_0 = _T_995[17]; // @[MemPrimitives.scala 96:27:@20819.4]
  assign Mem1D_15_clock = clock; // @[:@20392.4]
  assign Mem1D_15_reset = reset; // @[:@20393.4]
  assign Mem1D_15_io_r_ofs_0 = _T_2647[8:0]; // @[MemPrimitives.scala 127:28:@22412.4]
  assign Mem1D_15_io_r_backpressure = _T_2647[9]; // @[MemPrimitives.scala 128:32:@22413.4]
  assign Mem1D_15_io_w_ofs_0 = _T_1015[8:0]; // @[MemPrimitives.scala 94:28:@20836.4]
  assign Mem1D_15_io_w_data_0 = _T_1015[16:9]; // @[MemPrimitives.scala 95:29:@20837.4]
  assign Mem1D_15_io_w_en_0 = _T_1015[17]; // @[MemPrimitives.scala 96:27:@20838.4]
  assign Mem1D_16_clock = clock; // @[:@20408.4]
  assign Mem1D_16_reset = reset; // @[:@20409.4]
  assign Mem1D_16_io_r_ofs_0 = _T_2739[8:0]; // @[MemPrimitives.scala 127:28:@22501.4]
  assign Mem1D_16_io_r_backpressure = _T_2739[9]; // @[MemPrimitives.scala 128:32:@22502.4]
  assign Mem1D_16_io_w_ofs_0 = _T_1035[8:0]; // @[MemPrimitives.scala 94:28:@20855.4]
  assign Mem1D_16_io_w_data_0 = _T_1035[16:9]; // @[MemPrimitives.scala 95:29:@20856.4]
  assign Mem1D_16_io_w_en_0 = _T_1035[17]; // @[MemPrimitives.scala 96:27:@20857.4]
  assign Mem1D_17_clock = clock; // @[:@20424.4]
  assign Mem1D_17_reset = reset; // @[:@20425.4]
  assign Mem1D_17_io_r_ofs_0 = _T_2831[8:0]; // @[MemPrimitives.scala 127:28:@22590.4]
  assign Mem1D_17_io_r_backpressure = _T_2831[9]; // @[MemPrimitives.scala 128:32:@22591.4]
  assign Mem1D_17_io_w_ofs_0 = _T_1055[8:0]; // @[MemPrimitives.scala 94:28:@20874.4]
  assign Mem1D_17_io_w_data_0 = _T_1055[16:9]; // @[MemPrimitives.scala 95:29:@20875.4]
  assign Mem1D_17_io_w_en_0 = _T_1055[17]; // @[MemPrimitives.scala 96:27:@20876.4]
  assign Mem1D_18_clock = clock; // @[:@20440.4]
  assign Mem1D_18_reset = reset; // @[:@20441.4]
  assign Mem1D_18_io_r_ofs_0 = _T_2923[8:0]; // @[MemPrimitives.scala 127:28:@22679.4]
  assign Mem1D_18_io_r_backpressure = _T_2923[9]; // @[MemPrimitives.scala 128:32:@22680.4]
  assign Mem1D_18_io_w_ofs_0 = _T_1075[8:0]; // @[MemPrimitives.scala 94:28:@20893.4]
  assign Mem1D_18_io_w_data_0 = _T_1075[16:9]; // @[MemPrimitives.scala 95:29:@20894.4]
  assign Mem1D_18_io_w_en_0 = _T_1075[17]; // @[MemPrimitives.scala 96:27:@20895.4]
  assign Mem1D_19_clock = clock; // @[:@20456.4]
  assign Mem1D_19_reset = reset; // @[:@20457.4]
  assign Mem1D_19_io_r_ofs_0 = _T_3015[8:0]; // @[MemPrimitives.scala 127:28:@22768.4]
  assign Mem1D_19_io_r_backpressure = _T_3015[9]; // @[MemPrimitives.scala 128:32:@22769.4]
  assign Mem1D_19_io_w_ofs_0 = _T_1095[8:0]; // @[MemPrimitives.scala 94:28:@20912.4]
  assign Mem1D_19_io_w_data_0 = _T_1095[16:9]; // @[MemPrimitives.scala 95:29:@20913.4]
  assign Mem1D_19_io_w_en_0 = _T_1095[17]; // @[MemPrimitives.scala 96:27:@20914.4]
  assign Mem1D_20_clock = clock; // @[:@20472.4]
  assign Mem1D_20_reset = reset; // @[:@20473.4]
  assign Mem1D_20_io_r_ofs_0 = _T_3107[8:0]; // @[MemPrimitives.scala 127:28:@22857.4]
  assign Mem1D_20_io_r_backpressure = _T_3107[9]; // @[MemPrimitives.scala 128:32:@22858.4]
  assign Mem1D_20_io_w_ofs_0 = _T_1115[8:0]; // @[MemPrimitives.scala 94:28:@20931.4]
  assign Mem1D_20_io_w_data_0 = _T_1115[16:9]; // @[MemPrimitives.scala 95:29:@20932.4]
  assign Mem1D_20_io_w_en_0 = _T_1115[17]; // @[MemPrimitives.scala 96:27:@20933.4]
  assign Mem1D_21_clock = clock; // @[:@20488.4]
  assign Mem1D_21_reset = reset; // @[:@20489.4]
  assign Mem1D_21_io_r_ofs_0 = _T_3199[8:0]; // @[MemPrimitives.scala 127:28:@22946.4]
  assign Mem1D_21_io_r_backpressure = _T_3199[9]; // @[MemPrimitives.scala 128:32:@22947.4]
  assign Mem1D_21_io_w_ofs_0 = _T_1135[8:0]; // @[MemPrimitives.scala 94:28:@20950.4]
  assign Mem1D_21_io_w_data_0 = _T_1135[16:9]; // @[MemPrimitives.scala 95:29:@20951.4]
  assign Mem1D_21_io_w_en_0 = _T_1135[17]; // @[MemPrimitives.scala 96:27:@20952.4]
  assign Mem1D_22_clock = clock; // @[:@20504.4]
  assign Mem1D_22_reset = reset; // @[:@20505.4]
  assign Mem1D_22_io_r_ofs_0 = _T_3291[8:0]; // @[MemPrimitives.scala 127:28:@23035.4]
  assign Mem1D_22_io_r_backpressure = _T_3291[9]; // @[MemPrimitives.scala 128:32:@23036.4]
  assign Mem1D_22_io_w_ofs_0 = _T_1155[8:0]; // @[MemPrimitives.scala 94:28:@20969.4]
  assign Mem1D_22_io_w_data_0 = _T_1155[16:9]; // @[MemPrimitives.scala 95:29:@20970.4]
  assign Mem1D_22_io_w_en_0 = _T_1155[17]; // @[MemPrimitives.scala 96:27:@20971.4]
  assign Mem1D_23_clock = clock; // @[:@20520.4]
  assign Mem1D_23_reset = reset; // @[:@20521.4]
  assign Mem1D_23_io_r_ofs_0 = _T_3383[8:0]; // @[MemPrimitives.scala 127:28:@23124.4]
  assign Mem1D_23_io_r_backpressure = _T_3383[9]; // @[MemPrimitives.scala 128:32:@23125.4]
  assign Mem1D_23_io_w_ofs_0 = _T_1175[8:0]; // @[MemPrimitives.scala 94:28:@20988.4]
  assign Mem1D_23_io_w_data_0 = _T_1175[16:9]; // @[MemPrimitives.scala 95:29:@20989.4]
  assign Mem1D_23_io_w_en_0 = _T_1175[17]; // @[MemPrimitives.scala 96:27:@20990.4]
  assign StickySelects_clock = clock; // @[:@21028.4]
  assign StickySelects_reset = reset; // @[:@21029.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0 & _T_1183; // @[MemPrimitives.scala 122:60:@21030.4]
  assign StickySelects_io_ins_1 = io_rPort_2_en_0 & _T_1189; // @[MemPrimitives.scala 122:60:@21031.4]
  assign StickySelects_io_ins_2 = io_rPort_4_en_0 & _T_1195; // @[MemPrimitives.scala 122:60:@21032.4]
  assign StickySelects_io_ins_3 = io_rPort_7_en_0 & _T_1201; // @[MemPrimitives.scala 122:60:@21033.4]
  assign StickySelects_io_ins_4 = io_rPort_8_en_0 & _T_1207; // @[MemPrimitives.scala 122:60:@21034.4]
  assign StickySelects_io_ins_5 = io_rPort_10_en_0 & _T_1213; // @[MemPrimitives.scala 122:60:@21035.4]
  assign StickySelects_io_ins_6 = io_rPort_11_en_0 & _T_1219; // @[MemPrimitives.scala 122:60:@21036.4]
  assign StickySelects_io_ins_7 = io_rPort_15_en_0 & _T_1225; // @[MemPrimitives.scala 122:60:@21037.4]
  assign StickySelects_io_ins_8 = io_rPort_17_en_0 & _T_1231; // @[MemPrimitives.scala 122:60:@21038.4]
  assign StickySelects_1_clock = clock; // @[:@21117.4]
  assign StickySelects_1_reset = reset; // @[:@21118.4]
  assign StickySelects_1_io_ins_0 = io_rPort_1_en_0 & _T_1275; // @[MemPrimitives.scala 122:60:@21119.4]
  assign StickySelects_1_io_ins_1 = io_rPort_3_en_0 & _T_1281; // @[MemPrimitives.scala 122:60:@21120.4]
  assign StickySelects_1_io_ins_2 = io_rPort_5_en_0 & _T_1287; // @[MemPrimitives.scala 122:60:@21121.4]
  assign StickySelects_1_io_ins_3 = io_rPort_6_en_0 & _T_1293; // @[MemPrimitives.scala 122:60:@21122.4]
  assign StickySelects_1_io_ins_4 = io_rPort_9_en_0 & _T_1299; // @[MemPrimitives.scala 122:60:@21123.4]
  assign StickySelects_1_io_ins_5 = io_rPort_12_en_0 & _T_1305; // @[MemPrimitives.scala 122:60:@21124.4]
  assign StickySelects_1_io_ins_6 = io_rPort_13_en_0 & _T_1311; // @[MemPrimitives.scala 122:60:@21125.4]
  assign StickySelects_1_io_ins_7 = io_rPort_14_en_0 & _T_1317; // @[MemPrimitives.scala 122:60:@21126.4]
  assign StickySelects_1_io_ins_8 = io_rPort_16_en_0 & _T_1323; // @[MemPrimitives.scala 122:60:@21127.4]
  assign StickySelects_2_clock = clock; // @[:@21206.4]
  assign StickySelects_2_reset = reset; // @[:@21207.4]
  assign StickySelects_2_io_ins_0 = io_rPort_0_en_0 & _T_1367; // @[MemPrimitives.scala 122:60:@21208.4]
  assign StickySelects_2_io_ins_1 = io_rPort_2_en_0 & _T_1373; // @[MemPrimitives.scala 122:60:@21209.4]
  assign StickySelects_2_io_ins_2 = io_rPort_4_en_0 & _T_1379; // @[MemPrimitives.scala 122:60:@21210.4]
  assign StickySelects_2_io_ins_3 = io_rPort_7_en_0 & _T_1385; // @[MemPrimitives.scala 122:60:@21211.4]
  assign StickySelects_2_io_ins_4 = io_rPort_8_en_0 & _T_1391; // @[MemPrimitives.scala 122:60:@21212.4]
  assign StickySelects_2_io_ins_5 = io_rPort_10_en_0 & _T_1397; // @[MemPrimitives.scala 122:60:@21213.4]
  assign StickySelects_2_io_ins_6 = io_rPort_11_en_0 & _T_1403; // @[MemPrimitives.scala 122:60:@21214.4]
  assign StickySelects_2_io_ins_7 = io_rPort_15_en_0 & _T_1409; // @[MemPrimitives.scala 122:60:@21215.4]
  assign StickySelects_2_io_ins_8 = io_rPort_17_en_0 & _T_1415; // @[MemPrimitives.scala 122:60:@21216.4]
  assign StickySelects_3_clock = clock; // @[:@21295.4]
  assign StickySelects_3_reset = reset; // @[:@21296.4]
  assign StickySelects_3_io_ins_0 = io_rPort_1_en_0 & _T_1459; // @[MemPrimitives.scala 122:60:@21297.4]
  assign StickySelects_3_io_ins_1 = io_rPort_3_en_0 & _T_1465; // @[MemPrimitives.scala 122:60:@21298.4]
  assign StickySelects_3_io_ins_2 = io_rPort_5_en_0 & _T_1471; // @[MemPrimitives.scala 122:60:@21299.4]
  assign StickySelects_3_io_ins_3 = io_rPort_6_en_0 & _T_1477; // @[MemPrimitives.scala 122:60:@21300.4]
  assign StickySelects_3_io_ins_4 = io_rPort_9_en_0 & _T_1483; // @[MemPrimitives.scala 122:60:@21301.4]
  assign StickySelects_3_io_ins_5 = io_rPort_12_en_0 & _T_1489; // @[MemPrimitives.scala 122:60:@21302.4]
  assign StickySelects_3_io_ins_6 = io_rPort_13_en_0 & _T_1495; // @[MemPrimitives.scala 122:60:@21303.4]
  assign StickySelects_3_io_ins_7 = io_rPort_14_en_0 & _T_1501; // @[MemPrimitives.scala 122:60:@21304.4]
  assign StickySelects_3_io_ins_8 = io_rPort_16_en_0 & _T_1507; // @[MemPrimitives.scala 122:60:@21305.4]
  assign StickySelects_4_clock = clock; // @[:@21384.4]
  assign StickySelects_4_reset = reset; // @[:@21385.4]
  assign StickySelects_4_io_ins_0 = io_rPort_0_en_0 & _T_1551; // @[MemPrimitives.scala 122:60:@21386.4]
  assign StickySelects_4_io_ins_1 = io_rPort_2_en_0 & _T_1557; // @[MemPrimitives.scala 122:60:@21387.4]
  assign StickySelects_4_io_ins_2 = io_rPort_4_en_0 & _T_1563; // @[MemPrimitives.scala 122:60:@21388.4]
  assign StickySelects_4_io_ins_3 = io_rPort_7_en_0 & _T_1569; // @[MemPrimitives.scala 122:60:@21389.4]
  assign StickySelects_4_io_ins_4 = io_rPort_8_en_0 & _T_1575; // @[MemPrimitives.scala 122:60:@21390.4]
  assign StickySelects_4_io_ins_5 = io_rPort_10_en_0 & _T_1581; // @[MemPrimitives.scala 122:60:@21391.4]
  assign StickySelects_4_io_ins_6 = io_rPort_11_en_0 & _T_1587; // @[MemPrimitives.scala 122:60:@21392.4]
  assign StickySelects_4_io_ins_7 = io_rPort_15_en_0 & _T_1593; // @[MemPrimitives.scala 122:60:@21393.4]
  assign StickySelects_4_io_ins_8 = io_rPort_17_en_0 & _T_1599; // @[MemPrimitives.scala 122:60:@21394.4]
  assign StickySelects_5_clock = clock; // @[:@21473.4]
  assign StickySelects_5_reset = reset; // @[:@21474.4]
  assign StickySelects_5_io_ins_0 = io_rPort_1_en_0 & _T_1643; // @[MemPrimitives.scala 122:60:@21475.4]
  assign StickySelects_5_io_ins_1 = io_rPort_3_en_0 & _T_1649; // @[MemPrimitives.scala 122:60:@21476.4]
  assign StickySelects_5_io_ins_2 = io_rPort_5_en_0 & _T_1655; // @[MemPrimitives.scala 122:60:@21477.4]
  assign StickySelects_5_io_ins_3 = io_rPort_6_en_0 & _T_1661; // @[MemPrimitives.scala 122:60:@21478.4]
  assign StickySelects_5_io_ins_4 = io_rPort_9_en_0 & _T_1667; // @[MemPrimitives.scala 122:60:@21479.4]
  assign StickySelects_5_io_ins_5 = io_rPort_12_en_0 & _T_1673; // @[MemPrimitives.scala 122:60:@21480.4]
  assign StickySelects_5_io_ins_6 = io_rPort_13_en_0 & _T_1679; // @[MemPrimitives.scala 122:60:@21481.4]
  assign StickySelects_5_io_ins_7 = io_rPort_14_en_0 & _T_1685; // @[MemPrimitives.scala 122:60:@21482.4]
  assign StickySelects_5_io_ins_8 = io_rPort_16_en_0 & _T_1691; // @[MemPrimitives.scala 122:60:@21483.4]
  assign StickySelects_6_clock = clock; // @[:@21562.4]
  assign StickySelects_6_reset = reset; // @[:@21563.4]
  assign StickySelects_6_io_ins_0 = io_rPort_0_en_0 & _T_1735; // @[MemPrimitives.scala 122:60:@21564.4]
  assign StickySelects_6_io_ins_1 = io_rPort_2_en_0 & _T_1741; // @[MemPrimitives.scala 122:60:@21565.4]
  assign StickySelects_6_io_ins_2 = io_rPort_4_en_0 & _T_1747; // @[MemPrimitives.scala 122:60:@21566.4]
  assign StickySelects_6_io_ins_3 = io_rPort_7_en_0 & _T_1753; // @[MemPrimitives.scala 122:60:@21567.4]
  assign StickySelects_6_io_ins_4 = io_rPort_8_en_0 & _T_1759; // @[MemPrimitives.scala 122:60:@21568.4]
  assign StickySelects_6_io_ins_5 = io_rPort_10_en_0 & _T_1765; // @[MemPrimitives.scala 122:60:@21569.4]
  assign StickySelects_6_io_ins_6 = io_rPort_11_en_0 & _T_1771; // @[MemPrimitives.scala 122:60:@21570.4]
  assign StickySelects_6_io_ins_7 = io_rPort_15_en_0 & _T_1777; // @[MemPrimitives.scala 122:60:@21571.4]
  assign StickySelects_6_io_ins_8 = io_rPort_17_en_0 & _T_1783; // @[MemPrimitives.scala 122:60:@21572.4]
  assign StickySelects_7_clock = clock; // @[:@21651.4]
  assign StickySelects_7_reset = reset; // @[:@21652.4]
  assign StickySelects_7_io_ins_0 = io_rPort_1_en_0 & _T_1827; // @[MemPrimitives.scala 122:60:@21653.4]
  assign StickySelects_7_io_ins_1 = io_rPort_3_en_0 & _T_1833; // @[MemPrimitives.scala 122:60:@21654.4]
  assign StickySelects_7_io_ins_2 = io_rPort_5_en_0 & _T_1839; // @[MemPrimitives.scala 122:60:@21655.4]
  assign StickySelects_7_io_ins_3 = io_rPort_6_en_0 & _T_1845; // @[MemPrimitives.scala 122:60:@21656.4]
  assign StickySelects_7_io_ins_4 = io_rPort_9_en_0 & _T_1851; // @[MemPrimitives.scala 122:60:@21657.4]
  assign StickySelects_7_io_ins_5 = io_rPort_12_en_0 & _T_1857; // @[MemPrimitives.scala 122:60:@21658.4]
  assign StickySelects_7_io_ins_6 = io_rPort_13_en_0 & _T_1863; // @[MemPrimitives.scala 122:60:@21659.4]
  assign StickySelects_7_io_ins_7 = io_rPort_14_en_0 & _T_1869; // @[MemPrimitives.scala 122:60:@21660.4]
  assign StickySelects_7_io_ins_8 = io_rPort_16_en_0 & _T_1875; // @[MemPrimitives.scala 122:60:@21661.4]
  assign StickySelects_8_clock = clock; // @[:@21740.4]
  assign StickySelects_8_reset = reset; // @[:@21741.4]
  assign StickySelects_8_io_ins_0 = io_rPort_0_en_0 & _T_1919; // @[MemPrimitives.scala 122:60:@21742.4]
  assign StickySelects_8_io_ins_1 = io_rPort_2_en_0 & _T_1925; // @[MemPrimitives.scala 122:60:@21743.4]
  assign StickySelects_8_io_ins_2 = io_rPort_4_en_0 & _T_1931; // @[MemPrimitives.scala 122:60:@21744.4]
  assign StickySelects_8_io_ins_3 = io_rPort_7_en_0 & _T_1937; // @[MemPrimitives.scala 122:60:@21745.4]
  assign StickySelects_8_io_ins_4 = io_rPort_8_en_0 & _T_1943; // @[MemPrimitives.scala 122:60:@21746.4]
  assign StickySelects_8_io_ins_5 = io_rPort_10_en_0 & _T_1949; // @[MemPrimitives.scala 122:60:@21747.4]
  assign StickySelects_8_io_ins_6 = io_rPort_11_en_0 & _T_1955; // @[MemPrimitives.scala 122:60:@21748.4]
  assign StickySelects_8_io_ins_7 = io_rPort_15_en_0 & _T_1961; // @[MemPrimitives.scala 122:60:@21749.4]
  assign StickySelects_8_io_ins_8 = io_rPort_17_en_0 & _T_1967; // @[MemPrimitives.scala 122:60:@21750.4]
  assign StickySelects_9_clock = clock; // @[:@21829.4]
  assign StickySelects_9_reset = reset; // @[:@21830.4]
  assign StickySelects_9_io_ins_0 = io_rPort_1_en_0 & _T_2011; // @[MemPrimitives.scala 122:60:@21831.4]
  assign StickySelects_9_io_ins_1 = io_rPort_3_en_0 & _T_2017; // @[MemPrimitives.scala 122:60:@21832.4]
  assign StickySelects_9_io_ins_2 = io_rPort_5_en_0 & _T_2023; // @[MemPrimitives.scala 122:60:@21833.4]
  assign StickySelects_9_io_ins_3 = io_rPort_6_en_0 & _T_2029; // @[MemPrimitives.scala 122:60:@21834.4]
  assign StickySelects_9_io_ins_4 = io_rPort_9_en_0 & _T_2035; // @[MemPrimitives.scala 122:60:@21835.4]
  assign StickySelects_9_io_ins_5 = io_rPort_12_en_0 & _T_2041; // @[MemPrimitives.scala 122:60:@21836.4]
  assign StickySelects_9_io_ins_6 = io_rPort_13_en_0 & _T_2047; // @[MemPrimitives.scala 122:60:@21837.4]
  assign StickySelects_9_io_ins_7 = io_rPort_14_en_0 & _T_2053; // @[MemPrimitives.scala 122:60:@21838.4]
  assign StickySelects_9_io_ins_8 = io_rPort_16_en_0 & _T_2059; // @[MemPrimitives.scala 122:60:@21839.4]
  assign StickySelects_10_clock = clock; // @[:@21918.4]
  assign StickySelects_10_reset = reset; // @[:@21919.4]
  assign StickySelects_10_io_ins_0 = io_rPort_0_en_0 & _T_2103; // @[MemPrimitives.scala 122:60:@21920.4]
  assign StickySelects_10_io_ins_1 = io_rPort_2_en_0 & _T_2109; // @[MemPrimitives.scala 122:60:@21921.4]
  assign StickySelects_10_io_ins_2 = io_rPort_4_en_0 & _T_2115; // @[MemPrimitives.scala 122:60:@21922.4]
  assign StickySelects_10_io_ins_3 = io_rPort_7_en_0 & _T_2121; // @[MemPrimitives.scala 122:60:@21923.4]
  assign StickySelects_10_io_ins_4 = io_rPort_8_en_0 & _T_2127; // @[MemPrimitives.scala 122:60:@21924.4]
  assign StickySelects_10_io_ins_5 = io_rPort_10_en_0 & _T_2133; // @[MemPrimitives.scala 122:60:@21925.4]
  assign StickySelects_10_io_ins_6 = io_rPort_11_en_0 & _T_2139; // @[MemPrimitives.scala 122:60:@21926.4]
  assign StickySelects_10_io_ins_7 = io_rPort_15_en_0 & _T_2145; // @[MemPrimitives.scala 122:60:@21927.4]
  assign StickySelects_10_io_ins_8 = io_rPort_17_en_0 & _T_2151; // @[MemPrimitives.scala 122:60:@21928.4]
  assign StickySelects_11_clock = clock; // @[:@22007.4]
  assign StickySelects_11_reset = reset; // @[:@22008.4]
  assign StickySelects_11_io_ins_0 = io_rPort_1_en_0 & _T_2195; // @[MemPrimitives.scala 122:60:@22009.4]
  assign StickySelects_11_io_ins_1 = io_rPort_3_en_0 & _T_2201; // @[MemPrimitives.scala 122:60:@22010.4]
  assign StickySelects_11_io_ins_2 = io_rPort_5_en_0 & _T_2207; // @[MemPrimitives.scala 122:60:@22011.4]
  assign StickySelects_11_io_ins_3 = io_rPort_6_en_0 & _T_2213; // @[MemPrimitives.scala 122:60:@22012.4]
  assign StickySelects_11_io_ins_4 = io_rPort_9_en_0 & _T_2219; // @[MemPrimitives.scala 122:60:@22013.4]
  assign StickySelects_11_io_ins_5 = io_rPort_12_en_0 & _T_2225; // @[MemPrimitives.scala 122:60:@22014.4]
  assign StickySelects_11_io_ins_6 = io_rPort_13_en_0 & _T_2231; // @[MemPrimitives.scala 122:60:@22015.4]
  assign StickySelects_11_io_ins_7 = io_rPort_14_en_0 & _T_2237; // @[MemPrimitives.scala 122:60:@22016.4]
  assign StickySelects_11_io_ins_8 = io_rPort_16_en_0 & _T_2243; // @[MemPrimitives.scala 122:60:@22017.4]
  assign StickySelects_12_clock = clock; // @[:@22096.4]
  assign StickySelects_12_reset = reset; // @[:@22097.4]
  assign StickySelects_12_io_ins_0 = io_rPort_0_en_0 & _T_2287; // @[MemPrimitives.scala 122:60:@22098.4]
  assign StickySelects_12_io_ins_1 = io_rPort_2_en_0 & _T_2293; // @[MemPrimitives.scala 122:60:@22099.4]
  assign StickySelects_12_io_ins_2 = io_rPort_4_en_0 & _T_2299; // @[MemPrimitives.scala 122:60:@22100.4]
  assign StickySelects_12_io_ins_3 = io_rPort_7_en_0 & _T_2305; // @[MemPrimitives.scala 122:60:@22101.4]
  assign StickySelects_12_io_ins_4 = io_rPort_8_en_0 & _T_2311; // @[MemPrimitives.scala 122:60:@22102.4]
  assign StickySelects_12_io_ins_5 = io_rPort_10_en_0 & _T_2317; // @[MemPrimitives.scala 122:60:@22103.4]
  assign StickySelects_12_io_ins_6 = io_rPort_11_en_0 & _T_2323; // @[MemPrimitives.scala 122:60:@22104.4]
  assign StickySelects_12_io_ins_7 = io_rPort_15_en_0 & _T_2329; // @[MemPrimitives.scala 122:60:@22105.4]
  assign StickySelects_12_io_ins_8 = io_rPort_17_en_0 & _T_2335; // @[MemPrimitives.scala 122:60:@22106.4]
  assign StickySelects_13_clock = clock; // @[:@22185.4]
  assign StickySelects_13_reset = reset; // @[:@22186.4]
  assign StickySelects_13_io_ins_0 = io_rPort_1_en_0 & _T_2379; // @[MemPrimitives.scala 122:60:@22187.4]
  assign StickySelects_13_io_ins_1 = io_rPort_3_en_0 & _T_2385; // @[MemPrimitives.scala 122:60:@22188.4]
  assign StickySelects_13_io_ins_2 = io_rPort_5_en_0 & _T_2391; // @[MemPrimitives.scala 122:60:@22189.4]
  assign StickySelects_13_io_ins_3 = io_rPort_6_en_0 & _T_2397; // @[MemPrimitives.scala 122:60:@22190.4]
  assign StickySelects_13_io_ins_4 = io_rPort_9_en_0 & _T_2403; // @[MemPrimitives.scala 122:60:@22191.4]
  assign StickySelects_13_io_ins_5 = io_rPort_12_en_0 & _T_2409; // @[MemPrimitives.scala 122:60:@22192.4]
  assign StickySelects_13_io_ins_6 = io_rPort_13_en_0 & _T_2415; // @[MemPrimitives.scala 122:60:@22193.4]
  assign StickySelects_13_io_ins_7 = io_rPort_14_en_0 & _T_2421; // @[MemPrimitives.scala 122:60:@22194.4]
  assign StickySelects_13_io_ins_8 = io_rPort_16_en_0 & _T_2427; // @[MemPrimitives.scala 122:60:@22195.4]
  assign StickySelects_14_clock = clock; // @[:@22274.4]
  assign StickySelects_14_reset = reset; // @[:@22275.4]
  assign StickySelects_14_io_ins_0 = io_rPort_0_en_0 & _T_2471; // @[MemPrimitives.scala 122:60:@22276.4]
  assign StickySelects_14_io_ins_1 = io_rPort_2_en_0 & _T_2477; // @[MemPrimitives.scala 122:60:@22277.4]
  assign StickySelects_14_io_ins_2 = io_rPort_4_en_0 & _T_2483; // @[MemPrimitives.scala 122:60:@22278.4]
  assign StickySelects_14_io_ins_3 = io_rPort_7_en_0 & _T_2489; // @[MemPrimitives.scala 122:60:@22279.4]
  assign StickySelects_14_io_ins_4 = io_rPort_8_en_0 & _T_2495; // @[MemPrimitives.scala 122:60:@22280.4]
  assign StickySelects_14_io_ins_5 = io_rPort_10_en_0 & _T_2501; // @[MemPrimitives.scala 122:60:@22281.4]
  assign StickySelects_14_io_ins_6 = io_rPort_11_en_0 & _T_2507; // @[MemPrimitives.scala 122:60:@22282.4]
  assign StickySelects_14_io_ins_7 = io_rPort_15_en_0 & _T_2513; // @[MemPrimitives.scala 122:60:@22283.4]
  assign StickySelects_14_io_ins_8 = io_rPort_17_en_0 & _T_2519; // @[MemPrimitives.scala 122:60:@22284.4]
  assign StickySelects_15_clock = clock; // @[:@22363.4]
  assign StickySelects_15_reset = reset; // @[:@22364.4]
  assign StickySelects_15_io_ins_0 = io_rPort_1_en_0 & _T_2563; // @[MemPrimitives.scala 122:60:@22365.4]
  assign StickySelects_15_io_ins_1 = io_rPort_3_en_0 & _T_2569; // @[MemPrimitives.scala 122:60:@22366.4]
  assign StickySelects_15_io_ins_2 = io_rPort_5_en_0 & _T_2575; // @[MemPrimitives.scala 122:60:@22367.4]
  assign StickySelects_15_io_ins_3 = io_rPort_6_en_0 & _T_2581; // @[MemPrimitives.scala 122:60:@22368.4]
  assign StickySelects_15_io_ins_4 = io_rPort_9_en_0 & _T_2587; // @[MemPrimitives.scala 122:60:@22369.4]
  assign StickySelects_15_io_ins_5 = io_rPort_12_en_0 & _T_2593; // @[MemPrimitives.scala 122:60:@22370.4]
  assign StickySelects_15_io_ins_6 = io_rPort_13_en_0 & _T_2599; // @[MemPrimitives.scala 122:60:@22371.4]
  assign StickySelects_15_io_ins_7 = io_rPort_14_en_0 & _T_2605; // @[MemPrimitives.scala 122:60:@22372.4]
  assign StickySelects_15_io_ins_8 = io_rPort_16_en_0 & _T_2611; // @[MemPrimitives.scala 122:60:@22373.4]
  assign StickySelects_16_clock = clock; // @[:@22452.4]
  assign StickySelects_16_reset = reset; // @[:@22453.4]
  assign StickySelects_16_io_ins_0 = io_rPort_0_en_0 & _T_2655; // @[MemPrimitives.scala 122:60:@22454.4]
  assign StickySelects_16_io_ins_1 = io_rPort_2_en_0 & _T_2661; // @[MemPrimitives.scala 122:60:@22455.4]
  assign StickySelects_16_io_ins_2 = io_rPort_4_en_0 & _T_2667; // @[MemPrimitives.scala 122:60:@22456.4]
  assign StickySelects_16_io_ins_3 = io_rPort_7_en_0 & _T_2673; // @[MemPrimitives.scala 122:60:@22457.4]
  assign StickySelects_16_io_ins_4 = io_rPort_8_en_0 & _T_2679; // @[MemPrimitives.scala 122:60:@22458.4]
  assign StickySelects_16_io_ins_5 = io_rPort_10_en_0 & _T_2685; // @[MemPrimitives.scala 122:60:@22459.4]
  assign StickySelects_16_io_ins_6 = io_rPort_11_en_0 & _T_2691; // @[MemPrimitives.scala 122:60:@22460.4]
  assign StickySelects_16_io_ins_7 = io_rPort_15_en_0 & _T_2697; // @[MemPrimitives.scala 122:60:@22461.4]
  assign StickySelects_16_io_ins_8 = io_rPort_17_en_0 & _T_2703; // @[MemPrimitives.scala 122:60:@22462.4]
  assign StickySelects_17_clock = clock; // @[:@22541.4]
  assign StickySelects_17_reset = reset; // @[:@22542.4]
  assign StickySelects_17_io_ins_0 = io_rPort_1_en_0 & _T_2747; // @[MemPrimitives.scala 122:60:@22543.4]
  assign StickySelects_17_io_ins_1 = io_rPort_3_en_0 & _T_2753; // @[MemPrimitives.scala 122:60:@22544.4]
  assign StickySelects_17_io_ins_2 = io_rPort_5_en_0 & _T_2759; // @[MemPrimitives.scala 122:60:@22545.4]
  assign StickySelects_17_io_ins_3 = io_rPort_6_en_0 & _T_2765; // @[MemPrimitives.scala 122:60:@22546.4]
  assign StickySelects_17_io_ins_4 = io_rPort_9_en_0 & _T_2771; // @[MemPrimitives.scala 122:60:@22547.4]
  assign StickySelects_17_io_ins_5 = io_rPort_12_en_0 & _T_2777; // @[MemPrimitives.scala 122:60:@22548.4]
  assign StickySelects_17_io_ins_6 = io_rPort_13_en_0 & _T_2783; // @[MemPrimitives.scala 122:60:@22549.4]
  assign StickySelects_17_io_ins_7 = io_rPort_14_en_0 & _T_2789; // @[MemPrimitives.scala 122:60:@22550.4]
  assign StickySelects_17_io_ins_8 = io_rPort_16_en_0 & _T_2795; // @[MemPrimitives.scala 122:60:@22551.4]
  assign StickySelects_18_clock = clock; // @[:@22630.4]
  assign StickySelects_18_reset = reset; // @[:@22631.4]
  assign StickySelects_18_io_ins_0 = io_rPort_0_en_0 & _T_2839; // @[MemPrimitives.scala 122:60:@22632.4]
  assign StickySelects_18_io_ins_1 = io_rPort_2_en_0 & _T_2845; // @[MemPrimitives.scala 122:60:@22633.4]
  assign StickySelects_18_io_ins_2 = io_rPort_4_en_0 & _T_2851; // @[MemPrimitives.scala 122:60:@22634.4]
  assign StickySelects_18_io_ins_3 = io_rPort_7_en_0 & _T_2857; // @[MemPrimitives.scala 122:60:@22635.4]
  assign StickySelects_18_io_ins_4 = io_rPort_8_en_0 & _T_2863; // @[MemPrimitives.scala 122:60:@22636.4]
  assign StickySelects_18_io_ins_5 = io_rPort_10_en_0 & _T_2869; // @[MemPrimitives.scala 122:60:@22637.4]
  assign StickySelects_18_io_ins_6 = io_rPort_11_en_0 & _T_2875; // @[MemPrimitives.scala 122:60:@22638.4]
  assign StickySelects_18_io_ins_7 = io_rPort_15_en_0 & _T_2881; // @[MemPrimitives.scala 122:60:@22639.4]
  assign StickySelects_18_io_ins_8 = io_rPort_17_en_0 & _T_2887; // @[MemPrimitives.scala 122:60:@22640.4]
  assign StickySelects_19_clock = clock; // @[:@22719.4]
  assign StickySelects_19_reset = reset; // @[:@22720.4]
  assign StickySelects_19_io_ins_0 = io_rPort_1_en_0 & _T_2931; // @[MemPrimitives.scala 122:60:@22721.4]
  assign StickySelects_19_io_ins_1 = io_rPort_3_en_0 & _T_2937; // @[MemPrimitives.scala 122:60:@22722.4]
  assign StickySelects_19_io_ins_2 = io_rPort_5_en_0 & _T_2943; // @[MemPrimitives.scala 122:60:@22723.4]
  assign StickySelects_19_io_ins_3 = io_rPort_6_en_0 & _T_2949; // @[MemPrimitives.scala 122:60:@22724.4]
  assign StickySelects_19_io_ins_4 = io_rPort_9_en_0 & _T_2955; // @[MemPrimitives.scala 122:60:@22725.4]
  assign StickySelects_19_io_ins_5 = io_rPort_12_en_0 & _T_2961; // @[MemPrimitives.scala 122:60:@22726.4]
  assign StickySelects_19_io_ins_6 = io_rPort_13_en_0 & _T_2967; // @[MemPrimitives.scala 122:60:@22727.4]
  assign StickySelects_19_io_ins_7 = io_rPort_14_en_0 & _T_2973; // @[MemPrimitives.scala 122:60:@22728.4]
  assign StickySelects_19_io_ins_8 = io_rPort_16_en_0 & _T_2979; // @[MemPrimitives.scala 122:60:@22729.4]
  assign StickySelects_20_clock = clock; // @[:@22808.4]
  assign StickySelects_20_reset = reset; // @[:@22809.4]
  assign StickySelects_20_io_ins_0 = io_rPort_0_en_0 & _T_3023; // @[MemPrimitives.scala 122:60:@22810.4]
  assign StickySelects_20_io_ins_1 = io_rPort_2_en_0 & _T_3029; // @[MemPrimitives.scala 122:60:@22811.4]
  assign StickySelects_20_io_ins_2 = io_rPort_4_en_0 & _T_3035; // @[MemPrimitives.scala 122:60:@22812.4]
  assign StickySelects_20_io_ins_3 = io_rPort_7_en_0 & _T_3041; // @[MemPrimitives.scala 122:60:@22813.4]
  assign StickySelects_20_io_ins_4 = io_rPort_8_en_0 & _T_3047; // @[MemPrimitives.scala 122:60:@22814.4]
  assign StickySelects_20_io_ins_5 = io_rPort_10_en_0 & _T_3053; // @[MemPrimitives.scala 122:60:@22815.4]
  assign StickySelects_20_io_ins_6 = io_rPort_11_en_0 & _T_3059; // @[MemPrimitives.scala 122:60:@22816.4]
  assign StickySelects_20_io_ins_7 = io_rPort_15_en_0 & _T_3065; // @[MemPrimitives.scala 122:60:@22817.4]
  assign StickySelects_20_io_ins_8 = io_rPort_17_en_0 & _T_3071; // @[MemPrimitives.scala 122:60:@22818.4]
  assign StickySelects_21_clock = clock; // @[:@22897.4]
  assign StickySelects_21_reset = reset; // @[:@22898.4]
  assign StickySelects_21_io_ins_0 = io_rPort_1_en_0 & _T_3115; // @[MemPrimitives.scala 122:60:@22899.4]
  assign StickySelects_21_io_ins_1 = io_rPort_3_en_0 & _T_3121; // @[MemPrimitives.scala 122:60:@22900.4]
  assign StickySelects_21_io_ins_2 = io_rPort_5_en_0 & _T_3127; // @[MemPrimitives.scala 122:60:@22901.4]
  assign StickySelects_21_io_ins_3 = io_rPort_6_en_0 & _T_3133; // @[MemPrimitives.scala 122:60:@22902.4]
  assign StickySelects_21_io_ins_4 = io_rPort_9_en_0 & _T_3139; // @[MemPrimitives.scala 122:60:@22903.4]
  assign StickySelects_21_io_ins_5 = io_rPort_12_en_0 & _T_3145; // @[MemPrimitives.scala 122:60:@22904.4]
  assign StickySelects_21_io_ins_6 = io_rPort_13_en_0 & _T_3151; // @[MemPrimitives.scala 122:60:@22905.4]
  assign StickySelects_21_io_ins_7 = io_rPort_14_en_0 & _T_3157; // @[MemPrimitives.scala 122:60:@22906.4]
  assign StickySelects_21_io_ins_8 = io_rPort_16_en_0 & _T_3163; // @[MemPrimitives.scala 122:60:@22907.4]
  assign StickySelects_22_clock = clock; // @[:@22986.4]
  assign StickySelects_22_reset = reset; // @[:@22987.4]
  assign StickySelects_22_io_ins_0 = io_rPort_0_en_0 & _T_3207; // @[MemPrimitives.scala 122:60:@22988.4]
  assign StickySelects_22_io_ins_1 = io_rPort_2_en_0 & _T_3213; // @[MemPrimitives.scala 122:60:@22989.4]
  assign StickySelects_22_io_ins_2 = io_rPort_4_en_0 & _T_3219; // @[MemPrimitives.scala 122:60:@22990.4]
  assign StickySelects_22_io_ins_3 = io_rPort_7_en_0 & _T_3225; // @[MemPrimitives.scala 122:60:@22991.4]
  assign StickySelects_22_io_ins_4 = io_rPort_8_en_0 & _T_3231; // @[MemPrimitives.scala 122:60:@22992.4]
  assign StickySelects_22_io_ins_5 = io_rPort_10_en_0 & _T_3237; // @[MemPrimitives.scala 122:60:@22993.4]
  assign StickySelects_22_io_ins_6 = io_rPort_11_en_0 & _T_3243; // @[MemPrimitives.scala 122:60:@22994.4]
  assign StickySelects_22_io_ins_7 = io_rPort_15_en_0 & _T_3249; // @[MemPrimitives.scala 122:60:@22995.4]
  assign StickySelects_22_io_ins_8 = io_rPort_17_en_0 & _T_3255; // @[MemPrimitives.scala 122:60:@22996.4]
  assign StickySelects_23_clock = clock; // @[:@23075.4]
  assign StickySelects_23_reset = reset; // @[:@23076.4]
  assign StickySelects_23_io_ins_0 = io_rPort_1_en_0 & _T_3299; // @[MemPrimitives.scala 122:60:@23077.4]
  assign StickySelects_23_io_ins_1 = io_rPort_3_en_0 & _T_3305; // @[MemPrimitives.scala 122:60:@23078.4]
  assign StickySelects_23_io_ins_2 = io_rPort_5_en_0 & _T_3311; // @[MemPrimitives.scala 122:60:@23079.4]
  assign StickySelects_23_io_ins_3 = io_rPort_6_en_0 & _T_3317; // @[MemPrimitives.scala 122:60:@23080.4]
  assign StickySelects_23_io_ins_4 = io_rPort_9_en_0 & _T_3323; // @[MemPrimitives.scala 122:60:@23081.4]
  assign StickySelects_23_io_ins_5 = io_rPort_12_en_0 & _T_3329; // @[MemPrimitives.scala 122:60:@23082.4]
  assign StickySelects_23_io_ins_6 = io_rPort_13_en_0 & _T_3335; // @[MemPrimitives.scala 122:60:@23083.4]
  assign StickySelects_23_io_ins_7 = io_rPort_14_en_0 & _T_3341; // @[MemPrimitives.scala 122:60:@23084.4]
  assign StickySelects_23_io_ins_8 = io_rPort_16_en_0 & _T_3347; // @[MemPrimitives.scala 122:60:@23085.4]
  assign RetimeWrapper_clock = clock; // @[:@23165.4]
  assign RetimeWrapper_reset = reset; // @[:@23166.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@23168.4]
  assign RetimeWrapper_io_in = _T_1183 & io_rPort_0_en_0; // @[package.scala 94:16:@23167.4]
  assign RetimeWrapper_1_clock = clock; // @[:@23173.4]
  assign RetimeWrapper_1_reset = reset; // @[:@23174.4]
  assign RetimeWrapper_1_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@23176.4]
  assign RetimeWrapper_1_io_in = _T_1367 & io_rPort_0_en_0; // @[package.scala 94:16:@23175.4]
  assign RetimeWrapper_2_clock = clock; // @[:@23181.4]
  assign RetimeWrapper_2_reset = reset; // @[:@23182.4]
  assign RetimeWrapper_2_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@23184.4]
  assign RetimeWrapper_2_io_in = _T_1551 & io_rPort_0_en_0; // @[package.scala 94:16:@23183.4]
  assign RetimeWrapper_3_clock = clock; // @[:@23189.4]
  assign RetimeWrapper_3_reset = reset; // @[:@23190.4]
  assign RetimeWrapper_3_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@23192.4]
  assign RetimeWrapper_3_io_in = _T_1735 & io_rPort_0_en_0; // @[package.scala 94:16:@23191.4]
  assign RetimeWrapper_4_clock = clock; // @[:@23197.4]
  assign RetimeWrapper_4_reset = reset; // @[:@23198.4]
  assign RetimeWrapper_4_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@23200.4]
  assign RetimeWrapper_4_io_in = _T_1919 & io_rPort_0_en_0; // @[package.scala 94:16:@23199.4]
  assign RetimeWrapper_5_clock = clock; // @[:@23205.4]
  assign RetimeWrapper_5_reset = reset; // @[:@23206.4]
  assign RetimeWrapper_5_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@23208.4]
  assign RetimeWrapper_5_io_in = _T_2103 & io_rPort_0_en_0; // @[package.scala 94:16:@23207.4]
  assign RetimeWrapper_6_clock = clock; // @[:@23213.4]
  assign RetimeWrapper_6_reset = reset; // @[:@23214.4]
  assign RetimeWrapper_6_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@23216.4]
  assign RetimeWrapper_6_io_in = _T_2287 & io_rPort_0_en_0; // @[package.scala 94:16:@23215.4]
  assign RetimeWrapper_7_clock = clock; // @[:@23221.4]
  assign RetimeWrapper_7_reset = reset; // @[:@23222.4]
  assign RetimeWrapper_7_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@23224.4]
  assign RetimeWrapper_7_io_in = _T_2471 & io_rPort_0_en_0; // @[package.scala 94:16:@23223.4]
  assign RetimeWrapper_8_clock = clock; // @[:@23229.4]
  assign RetimeWrapper_8_reset = reset; // @[:@23230.4]
  assign RetimeWrapper_8_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@23232.4]
  assign RetimeWrapper_8_io_in = _T_2655 & io_rPort_0_en_0; // @[package.scala 94:16:@23231.4]
  assign RetimeWrapper_9_clock = clock; // @[:@23237.4]
  assign RetimeWrapper_9_reset = reset; // @[:@23238.4]
  assign RetimeWrapper_9_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@23240.4]
  assign RetimeWrapper_9_io_in = _T_2839 & io_rPort_0_en_0; // @[package.scala 94:16:@23239.4]
  assign RetimeWrapper_10_clock = clock; // @[:@23245.4]
  assign RetimeWrapper_10_reset = reset; // @[:@23246.4]
  assign RetimeWrapper_10_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@23248.4]
  assign RetimeWrapper_10_io_in = _T_3023 & io_rPort_0_en_0; // @[package.scala 94:16:@23247.4]
  assign RetimeWrapper_11_clock = clock; // @[:@23253.4]
  assign RetimeWrapper_11_reset = reset; // @[:@23254.4]
  assign RetimeWrapper_11_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@23256.4]
  assign RetimeWrapper_11_io_in = _T_3207 & io_rPort_0_en_0; // @[package.scala 94:16:@23255.4]
  assign RetimeWrapper_12_clock = clock; // @[:@23309.4]
  assign RetimeWrapper_12_reset = reset; // @[:@23310.4]
  assign RetimeWrapper_12_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@23312.4]
  assign RetimeWrapper_12_io_in = _T_1275 & io_rPort_1_en_0; // @[package.scala 94:16:@23311.4]
  assign RetimeWrapper_13_clock = clock; // @[:@23317.4]
  assign RetimeWrapper_13_reset = reset; // @[:@23318.4]
  assign RetimeWrapper_13_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@23320.4]
  assign RetimeWrapper_13_io_in = _T_1459 & io_rPort_1_en_0; // @[package.scala 94:16:@23319.4]
  assign RetimeWrapper_14_clock = clock; // @[:@23325.4]
  assign RetimeWrapper_14_reset = reset; // @[:@23326.4]
  assign RetimeWrapper_14_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@23328.4]
  assign RetimeWrapper_14_io_in = _T_1643 & io_rPort_1_en_0; // @[package.scala 94:16:@23327.4]
  assign RetimeWrapper_15_clock = clock; // @[:@23333.4]
  assign RetimeWrapper_15_reset = reset; // @[:@23334.4]
  assign RetimeWrapper_15_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@23336.4]
  assign RetimeWrapper_15_io_in = _T_1827 & io_rPort_1_en_0; // @[package.scala 94:16:@23335.4]
  assign RetimeWrapper_16_clock = clock; // @[:@23341.4]
  assign RetimeWrapper_16_reset = reset; // @[:@23342.4]
  assign RetimeWrapper_16_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@23344.4]
  assign RetimeWrapper_16_io_in = _T_2011 & io_rPort_1_en_0; // @[package.scala 94:16:@23343.4]
  assign RetimeWrapper_17_clock = clock; // @[:@23349.4]
  assign RetimeWrapper_17_reset = reset; // @[:@23350.4]
  assign RetimeWrapper_17_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@23352.4]
  assign RetimeWrapper_17_io_in = _T_2195 & io_rPort_1_en_0; // @[package.scala 94:16:@23351.4]
  assign RetimeWrapper_18_clock = clock; // @[:@23357.4]
  assign RetimeWrapper_18_reset = reset; // @[:@23358.4]
  assign RetimeWrapper_18_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@23360.4]
  assign RetimeWrapper_18_io_in = _T_2379 & io_rPort_1_en_0; // @[package.scala 94:16:@23359.4]
  assign RetimeWrapper_19_clock = clock; // @[:@23365.4]
  assign RetimeWrapper_19_reset = reset; // @[:@23366.4]
  assign RetimeWrapper_19_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@23368.4]
  assign RetimeWrapper_19_io_in = _T_2563 & io_rPort_1_en_0; // @[package.scala 94:16:@23367.4]
  assign RetimeWrapper_20_clock = clock; // @[:@23373.4]
  assign RetimeWrapper_20_reset = reset; // @[:@23374.4]
  assign RetimeWrapper_20_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@23376.4]
  assign RetimeWrapper_20_io_in = _T_2747 & io_rPort_1_en_0; // @[package.scala 94:16:@23375.4]
  assign RetimeWrapper_21_clock = clock; // @[:@23381.4]
  assign RetimeWrapper_21_reset = reset; // @[:@23382.4]
  assign RetimeWrapper_21_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@23384.4]
  assign RetimeWrapper_21_io_in = _T_2931 & io_rPort_1_en_0; // @[package.scala 94:16:@23383.4]
  assign RetimeWrapper_22_clock = clock; // @[:@23389.4]
  assign RetimeWrapper_22_reset = reset; // @[:@23390.4]
  assign RetimeWrapper_22_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@23392.4]
  assign RetimeWrapper_22_io_in = _T_3115 & io_rPort_1_en_0; // @[package.scala 94:16:@23391.4]
  assign RetimeWrapper_23_clock = clock; // @[:@23397.4]
  assign RetimeWrapper_23_reset = reset; // @[:@23398.4]
  assign RetimeWrapper_23_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@23400.4]
  assign RetimeWrapper_23_io_in = _T_3299 & io_rPort_1_en_0; // @[package.scala 94:16:@23399.4]
  assign RetimeWrapper_24_clock = clock; // @[:@23453.4]
  assign RetimeWrapper_24_reset = reset; // @[:@23454.4]
  assign RetimeWrapper_24_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@23456.4]
  assign RetimeWrapper_24_io_in = _T_1189 & io_rPort_2_en_0; // @[package.scala 94:16:@23455.4]
  assign RetimeWrapper_25_clock = clock; // @[:@23461.4]
  assign RetimeWrapper_25_reset = reset; // @[:@23462.4]
  assign RetimeWrapper_25_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@23464.4]
  assign RetimeWrapper_25_io_in = _T_1373 & io_rPort_2_en_0; // @[package.scala 94:16:@23463.4]
  assign RetimeWrapper_26_clock = clock; // @[:@23469.4]
  assign RetimeWrapper_26_reset = reset; // @[:@23470.4]
  assign RetimeWrapper_26_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@23472.4]
  assign RetimeWrapper_26_io_in = _T_1557 & io_rPort_2_en_0; // @[package.scala 94:16:@23471.4]
  assign RetimeWrapper_27_clock = clock; // @[:@23477.4]
  assign RetimeWrapper_27_reset = reset; // @[:@23478.4]
  assign RetimeWrapper_27_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@23480.4]
  assign RetimeWrapper_27_io_in = _T_1741 & io_rPort_2_en_0; // @[package.scala 94:16:@23479.4]
  assign RetimeWrapper_28_clock = clock; // @[:@23485.4]
  assign RetimeWrapper_28_reset = reset; // @[:@23486.4]
  assign RetimeWrapper_28_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@23488.4]
  assign RetimeWrapper_28_io_in = _T_1925 & io_rPort_2_en_0; // @[package.scala 94:16:@23487.4]
  assign RetimeWrapper_29_clock = clock; // @[:@23493.4]
  assign RetimeWrapper_29_reset = reset; // @[:@23494.4]
  assign RetimeWrapper_29_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@23496.4]
  assign RetimeWrapper_29_io_in = _T_2109 & io_rPort_2_en_0; // @[package.scala 94:16:@23495.4]
  assign RetimeWrapper_30_clock = clock; // @[:@23501.4]
  assign RetimeWrapper_30_reset = reset; // @[:@23502.4]
  assign RetimeWrapper_30_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@23504.4]
  assign RetimeWrapper_30_io_in = _T_2293 & io_rPort_2_en_0; // @[package.scala 94:16:@23503.4]
  assign RetimeWrapper_31_clock = clock; // @[:@23509.4]
  assign RetimeWrapper_31_reset = reset; // @[:@23510.4]
  assign RetimeWrapper_31_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@23512.4]
  assign RetimeWrapper_31_io_in = _T_2477 & io_rPort_2_en_0; // @[package.scala 94:16:@23511.4]
  assign RetimeWrapper_32_clock = clock; // @[:@23517.4]
  assign RetimeWrapper_32_reset = reset; // @[:@23518.4]
  assign RetimeWrapper_32_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@23520.4]
  assign RetimeWrapper_32_io_in = _T_2661 & io_rPort_2_en_0; // @[package.scala 94:16:@23519.4]
  assign RetimeWrapper_33_clock = clock; // @[:@23525.4]
  assign RetimeWrapper_33_reset = reset; // @[:@23526.4]
  assign RetimeWrapper_33_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@23528.4]
  assign RetimeWrapper_33_io_in = _T_2845 & io_rPort_2_en_0; // @[package.scala 94:16:@23527.4]
  assign RetimeWrapper_34_clock = clock; // @[:@23533.4]
  assign RetimeWrapper_34_reset = reset; // @[:@23534.4]
  assign RetimeWrapper_34_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@23536.4]
  assign RetimeWrapper_34_io_in = _T_3029 & io_rPort_2_en_0; // @[package.scala 94:16:@23535.4]
  assign RetimeWrapper_35_clock = clock; // @[:@23541.4]
  assign RetimeWrapper_35_reset = reset; // @[:@23542.4]
  assign RetimeWrapper_35_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@23544.4]
  assign RetimeWrapper_35_io_in = _T_3213 & io_rPort_2_en_0; // @[package.scala 94:16:@23543.4]
  assign RetimeWrapper_36_clock = clock; // @[:@23597.4]
  assign RetimeWrapper_36_reset = reset; // @[:@23598.4]
  assign RetimeWrapper_36_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@23600.4]
  assign RetimeWrapper_36_io_in = _T_1281 & io_rPort_3_en_0; // @[package.scala 94:16:@23599.4]
  assign RetimeWrapper_37_clock = clock; // @[:@23605.4]
  assign RetimeWrapper_37_reset = reset; // @[:@23606.4]
  assign RetimeWrapper_37_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@23608.4]
  assign RetimeWrapper_37_io_in = _T_1465 & io_rPort_3_en_0; // @[package.scala 94:16:@23607.4]
  assign RetimeWrapper_38_clock = clock; // @[:@23613.4]
  assign RetimeWrapper_38_reset = reset; // @[:@23614.4]
  assign RetimeWrapper_38_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@23616.4]
  assign RetimeWrapper_38_io_in = _T_1649 & io_rPort_3_en_0; // @[package.scala 94:16:@23615.4]
  assign RetimeWrapper_39_clock = clock; // @[:@23621.4]
  assign RetimeWrapper_39_reset = reset; // @[:@23622.4]
  assign RetimeWrapper_39_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@23624.4]
  assign RetimeWrapper_39_io_in = _T_1833 & io_rPort_3_en_0; // @[package.scala 94:16:@23623.4]
  assign RetimeWrapper_40_clock = clock; // @[:@23629.4]
  assign RetimeWrapper_40_reset = reset; // @[:@23630.4]
  assign RetimeWrapper_40_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@23632.4]
  assign RetimeWrapper_40_io_in = _T_2017 & io_rPort_3_en_0; // @[package.scala 94:16:@23631.4]
  assign RetimeWrapper_41_clock = clock; // @[:@23637.4]
  assign RetimeWrapper_41_reset = reset; // @[:@23638.4]
  assign RetimeWrapper_41_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@23640.4]
  assign RetimeWrapper_41_io_in = _T_2201 & io_rPort_3_en_0; // @[package.scala 94:16:@23639.4]
  assign RetimeWrapper_42_clock = clock; // @[:@23645.4]
  assign RetimeWrapper_42_reset = reset; // @[:@23646.4]
  assign RetimeWrapper_42_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@23648.4]
  assign RetimeWrapper_42_io_in = _T_2385 & io_rPort_3_en_0; // @[package.scala 94:16:@23647.4]
  assign RetimeWrapper_43_clock = clock; // @[:@23653.4]
  assign RetimeWrapper_43_reset = reset; // @[:@23654.4]
  assign RetimeWrapper_43_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@23656.4]
  assign RetimeWrapper_43_io_in = _T_2569 & io_rPort_3_en_0; // @[package.scala 94:16:@23655.4]
  assign RetimeWrapper_44_clock = clock; // @[:@23661.4]
  assign RetimeWrapper_44_reset = reset; // @[:@23662.4]
  assign RetimeWrapper_44_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@23664.4]
  assign RetimeWrapper_44_io_in = _T_2753 & io_rPort_3_en_0; // @[package.scala 94:16:@23663.4]
  assign RetimeWrapper_45_clock = clock; // @[:@23669.4]
  assign RetimeWrapper_45_reset = reset; // @[:@23670.4]
  assign RetimeWrapper_45_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@23672.4]
  assign RetimeWrapper_45_io_in = _T_2937 & io_rPort_3_en_0; // @[package.scala 94:16:@23671.4]
  assign RetimeWrapper_46_clock = clock; // @[:@23677.4]
  assign RetimeWrapper_46_reset = reset; // @[:@23678.4]
  assign RetimeWrapper_46_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@23680.4]
  assign RetimeWrapper_46_io_in = _T_3121 & io_rPort_3_en_0; // @[package.scala 94:16:@23679.4]
  assign RetimeWrapper_47_clock = clock; // @[:@23685.4]
  assign RetimeWrapper_47_reset = reset; // @[:@23686.4]
  assign RetimeWrapper_47_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@23688.4]
  assign RetimeWrapper_47_io_in = _T_3305 & io_rPort_3_en_0; // @[package.scala 94:16:@23687.4]
  assign RetimeWrapper_48_clock = clock; // @[:@23741.4]
  assign RetimeWrapper_48_reset = reset; // @[:@23742.4]
  assign RetimeWrapper_48_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23744.4]
  assign RetimeWrapper_48_io_in = _T_1195 & io_rPort_4_en_0; // @[package.scala 94:16:@23743.4]
  assign RetimeWrapper_49_clock = clock; // @[:@23749.4]
  assign RetimeWrapper_49_reset = reset; // @[:@23750.4]
  assign RetimeWrapper_49_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23752.4]
  assign RetimeWrapper_49_io_in = _T_1379 & io_rPort_4_en_0; // @[package.scala 94:16:@23751.4]
  assign RetimeWrapper_50_clock = clock; // @[:@23757.4]
  assign RetimeWrapper_50_reset = reset; // @[:@23758.4]
  assign RetimeWrapper_50_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23760.4]
  assign RetimeWrapper_50_io_in = _T_1563 & io_rPort_4_en_0; // @[package.scala 94:16:@23759.4]
  assign RetimeWrapper_51_clock = clock; // @[:@23765.4]
  assign RetimeWrapper_51_reset = reset; // @[:@23766.4]
  assign RetimeWrapper_51_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23768.4]
  assign RetimeWrapper_51_io_in = _T_1747 & io_rPort_4_en_0; // @[package.scala 94:16:@23767.4]
  assign RetimeWrapper_52_clock = clock; // @[:@23773.4]
  assign RetimeWrapper_52_reset = reset; // @[:@23774.4]
  assign RetimeWrapper_52_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23776.4]
  assign RetimeWrapper_52_io_in = _T_1931 & io_rPort_4_en_0; // @[package.scala 94:16:@23775.4]
  assign RetimeWrapper_53_clock = clock; // @[:@23781.4]
  assign RetimeWrapper_53_reset = reset; // @[:@23782.4]
  assign RetimeWrapper_53_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23784.4]
  assign RetimeWrapper_53_io_in = _T_2115 & io_rPort_4_en_0; // @[package.scala 94:16:@23783.4]
  assign RetimeWrapper_54_clock = clock; // @[:@23789.4]
  assign RetimeWrapper_54_reset = reset; // @[:@23790.4]
  assign RetimeWrapper_54_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23792.4]
  assign RetimeWrapper_54_io_in = _T_2299 & io_rPort_4_en_0; // @[package.scala 94:16:@23791.4]
  assign RetimeWrapper_55_clock = clock; // @[:@23797.4]
  assign RetimeWrapper_55_reset = reset; // @[:@23798.4]
  assign RetimeWrapper_55_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23800.4]
  assign RetimeWrapper_55_io_in = _T_2483 & io_rPort_4_en_0; // @[package.scala 94:16:@23799.4]
  assign RetimeWrapper_56_clock = clock; // @[:@23805.4]
  assign RetimeWrapper_56_reset = reset; // @[:@23806.4]
  assign RetimeWrapper_56_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23808.4]
  assign RetimeWrapper_56_io_in = _T_2667 & io_rPort_4_en_0; // @[package.scala 94:16:@23807.4]
  assign RetimeWrapper_57_clock = clock; // @[:@23813.4]
  assign RetimeWrapper_57_reset = reset; // @[:@23814.4]
  assign RetimeWrapper_57_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23816.4]
  assign RetimeWrapper_57_io_in = _T_2851 & io_rPort_4_en_0; // @[package.scala 94:16:@23815.4]
  assign RetimeWrapper_58_clock = clock; // @[:@23821.4]
  assign RetimeWrapper_58_reset = reset; // @[:@23822.4]
  assign RetimeWrapper_58_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23824.4]
  assign RetimeWrapper_58_io_in = _T_3035 & io_rPort_4_en_0; // @[package.scala 94:16:@23823.4]
  assign RetimeWrapper_59_clock = clock; // @[:@23829.4]
  assign RetimeWrapper_59_reset = reset; // @[:@23830.4]
  assign RetimeWrapper_59_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23832.4]
  assign RetimeWrapper_59_io_in = _T_3219 & io_rPort_4_en_0; // @[package.scala 94:16:@23831.4]
  assign RetimeWrapper_60_clock = clock; // @[:@23885.4]
  assign RetimeWrapper_60_reset = reset; // @[:@23886.4]
  assign RetimeWrapper_60_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23888.4]
  assign RetimeWrapper_60_io_in = _T_1287 & io_rPort_5_en_0; // @[package.scala 94:16:@23887.4]
  assign RetimeWrapper_61_clock = clock; // @[:@23893.4]
  assign RetimeWrapper_61_reset = reset; // @[:@23894.4]
  assign RetimeWrapper_61_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23896.4]
  assign RetimeWrapper_61_io_in = _T_1471 & io_rPort_5_en_0; // @[package.scala 94:16:@23895.4]
  assign RetimeWrapper_62_clock = clock; // @[:@23901.4]
  assign RetimeWrapper_62_reset = reset; // @[:@23902.4]
  assign RetimeWrapper_62_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23904.4]
  assign RetimeWrapper_62_io_in = _T_1655 & io_rPort_5_en_0; // @[package.scala 94:16:@23903.4]
  assign RetimeWrapper_63_clock = clock; // @[:@23909.4]
  assign RetimeWrapper_63_reset = reset; // @[:@23910.4]
  assign RetimeWrapper_63_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23912.4]
  assign RetimeWrapper_63_io_in = _T_1839 & io_rPort_5_en_0; // @[package.scala 94:16:@23911.4]
  assign RetimeWrapper_64_clock = clock; // @[:@23917.4]
  assign RetimeWrapper_64_reset = reset; // @[:@23918.4]
  assign RetimeWrapper_64_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23920.4]
  assign RetimeWrapper_64_io_in = _T_2023 & io_rPort_5_en_0; // @[package.scala 94:16:@23919.4]
  assign RetimeWrapper_65_clock = clock; // @[:@23925.4]
  assign RetimeWrapper_65_reset = reset; // @[:@23926.4]
  assign RetimeWrapper_65_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23928.4]
  assign RetimeWrapper_65_io_in = _T_2207 & io_rPort_5_en_0; // @[package.scala 94:16:@23927.4]
  assign RetimeWrapper_66_clock = clock; // @[:@23933.4]
  assign RetimeWrapper_66_reset = reset; // @[:@23934.4]
  assign RetimeWrapper_66_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23936.4]
  assign RetimeWrapper_66_io_in = _T_2391 & io_rPort_5_en_0; // @[package.scala 94:16:@23935.4]
  assign RetimeWrapper_67_clock = clock; // @[:@23941.4]
  assign RetimeWrapper_67_reset = reset; // @[:@23942.4]
  assign RetimeWrapper_67_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23944.4]
  assign RetimeWrapper_67_io_in = _T_2575 & io_rPort_5_en_0; // @[package.scala 94:16:@23943.4]
  assign RetimeWrapper_68_clock = clock; // @[:@23949.4]
  assign RetimeWrapper_68_reset = reset; // @[:@23950.4]
  assign RetimeWrapper_68_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23952.4]
  assign RetimeWrapper_68_io_in = _T_2759 & io_rPort_5_en_0; // @[package.scala 94:16:@23951.4]
  assign RetimeWrapper_69_clock = clock; // @[:@23957.4]
  assign RetimeWrapper_69_reset = reset; // @[:@23958.4]
  assign RetimeWrapper_69_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23960.4]
  assign RetimeWrapper_69_io_in = _T_2943 & io_rPort_5_en_0; // @[package.scala 94:16:@23959.4]
  assign RetimeWrapper_70_clock = clock; // @[:@23965.4]
  assign RetimeWrapper_70_reset = reset; // @[:@23966.4]
  assign RetimeWrapper_70_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23968.4]
  assign RetimeWrapper_70_io_in = _T_3127 & io_rPort_5_en_0; // @[package.scala 94:16:@23967.4]
  assign RetimeWrapper_71_clock = clock; // @[:@23973.4]
  assign RetimeWrapper_71_reset = reset; // @[:@23974.4]
  assign RetimeWrapper_71_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23976.4]
  assign RetimeWrapper_71_io_in = _T_3311 & io_rPort_5_en_0; // @[package.scala 94:16:@23975.4]
  assign RetimeWrapper_72_clock = clock; // @[:@24029.4]
  assign RetimeWrapper_72_reset = reset; // @[:@24030.4]
  assign RetimeWrapper_72_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@24032.4]
  assign RetimeWrapper_72_io_in = _T_1293 & io_rPort_6_en_0; // @[package.scala 94:16:@24031.4]
  assign RetimeWrapper_73_clock = clock; // @[:@24037.4]
  assign RetimeWrapper_73_reset = reset; // @[:@24038.4]
  assign RetimeWrapper_73_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@24040.4]
  assign RetimeWrapper_73_io_in = _T_1477 & io_rPort_6_en_0; // @[package.scala 94:16:@24039.4]
  assign RetimeWrapper_74_clock = clock; // @[:@24045.4]
  assign RetimeWrapper_74_reset = reset; // @[:@24046.4]
  assign RetimeWrapper_74_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@24048.4]
  assign RetimeWrapper_74_io_in = _T_1661 & io_rPort_6_en_0; // @[package.scala 94:16:@24047.4]
  assign RetimeWrapper_75_clock = clock; // @[:@24053.4]
  assign RetimeWrapper_75_reset = reset; // @[:@24054.4]
  assign RetimeWrapper_75_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@24056.4]
  assign RetimeWrapper_75_io_in = _T_1845 & io_rPort_6_en_0; // @[package.scala 94:16:@24055.4]
  assign RetimeWrapper_76_clock = clock; // @[:@24061.4]
  assign RetimeWrapper_76_reset = reset; // @[:@24062.4]
  assign RetimeWrapper_76_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@24064.4]
  assign RetimeWrapper_76_io_in = _T_2029 & io_rPort_6_en_0; // @[package.scala 94:16:@24063.4]
  assign RetimeWrapper_77_clock = clock; // @[:@24069.4]
  assign RetimeWrapper_77_reset = reset; // @[:@24070.4]
  assign RetimeWrapper_77_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@24072.4]
  assign RetimeWrapper_77_io_in = _T_2213 & io_rPort_6_en_0; // @[package.scala 94:16:@24071.4]
  assign RetimeWrapper_78_clock = clock; // @[:@24077.4]
  assign RetimeWrapper_78_reset = reset; // @[:@24078.4]
  assign RetimeWrapper_78_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@24080.4]
  assign RetimeWrapper_78_io_in = _T_2397 & io_rPort_6_en_0; // @[package.scala 94:16:@24079.4]
  assign RetimeWrapper_79_clock = clock; // @[:@24085.4]
  assign RetimeWrapper_79_reset = reset; // @[:@24086.4]
  assign RetimeWrapper_79_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@24088.4]
  assign RetimeWrapper_79_io_in = _T_2581 & io_rPort_6_en_0; // @[package.scala 94:16:@24087.4]
  assign RetimeWrapper_80_clock = clock; // @[:@24093.4]
  assign RetimeWrapper_80_reset = reset; // @[:@24094.4]
  assign RetimeWrapper_80_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@24096.4]
  assign RetimeWrapper_80_io_in = _T_2765 & io_rPort_6_en_0; // @[package.scala 94:16:@24095.4]
  assign RetimeWrapper_81_clock = clock; // @[:@24101.4]
  assign RetimeWrapper_81_reset = reset; // @[:@24102.4]
  assign RetimeWrapper_81_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@24104.4]
  assign RetimeWrapper_81_io_in = _T_2949 & io_rPort_6_en_0; // @[package.scala 94:16:@24103.4]
  assign RetimeWrapper_82_clock = clock; // @[:@24109.4]
  assign RetimeWrapper_82_reset = reset; // @[:@24110.4]
  assign RetimeWrapper_82_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@24112.4]
  assign RetimeWrapper_82_io_in = _T_3133 & io_rPort_6_en_0; // @[package.scala 94:16:@24111.4]
  assign RetimeWrapper_83_clock = clock; // @[:@24117.4]
  assign RetimeWrapper_83_reset = reset; // @[:@24118.4]
  assign RetimeWrapper_83_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@24120.4]
  assign RetimeWrapper_83_io_in = _T_3317 & io_rPort_6_en_0; // @[package.scala 94:16:@24119.4]
  assign RetimeWrapper_84_clock = clock; // @[:@24173.4]
  assign RetimeWrapper_84_reset = reset; // @[:@24174.4]
  assign RetimeWrapper_84_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@24176.4]
  assign RetimeWrapper_84_io_in = _T_1201 & io_rPort_7_en_0; // @[package.scala 94:16:@24175.4]
  assign RetimeWrapper_85_clock = clock; // @[:@24181.4]
  assign RetimeWrapper_85_reset = reset; // @[:@24182.4]
  assign RetimeWrapper_85_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@24184.4]
  assign RetimeWrapper_85_io_in = _T_1385 & io_rPort_7_en_0; // @[package.scala 94:16:@24183.4]
  assign RetimeWrapper_86_clock = clock; // @[:@24189.4]
  assign RetimeWrapper_86_reset = reset; // @[:@24190.4]
  assign RetimeWrapper_86_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@24192.4]
  assign RetimeWrapper_86_io_in = _T_1569 & io_rPort_7_en_0; // @[package.scala 94:16:@24191.4]
  assign RetimeWrapper_87_clock = clock; // @[:@24197.4]
  assign RetimeWrapper_87_reset = reset; // @[:@24198.4]
  assign RetimeWrapper_87_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@24200.4]
  assign RetimeWrapper_87_io_in = _T_1753 & io_rPort_7_en_0; // @[package.scala 94:16:@24199.4]
  assign RetimeWrapper_88_clock = clock; // @[:@24205.4]
  assign RetimeWrapper_88_reset = reset; // @[:@24206.4]
  assign RetimeWrapper_88_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@24208.4]
  assign RetimeWrapper_88_io_in = _T_1937 & io_rPort_7_en_0; // @[package.scala 94:16:@24207.4]
  assign RetimeWrapper_89_clock = clock; // @[:@24213.4]
  assign RetimeWrapper_89_reset = reset; // @[:@24214.4]
  assign RetimeWrapper_89_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@24216.4]
  assign RetimeWrapper_89_io_in = _T_2121 & io_rPort_7_en_0; // @[package.scala 94:16:@24215.4]
  assign RetimeWrapper_90_clock = clock; // @[:@24221.4]
  assign RetimeWrapper_90_reset = reset; // @[:@24222.4]
  assign RetimeWrapper_90_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@24224.4]
  assign RetimeWrapper_90_io_in = _T_2305 & io_rPort_7_en_0; // @[package.scala 94:16:@24223.4]
  assign RetimeWrapper_91_clock = clock; // @[:@24229.4]
  assign RetimeWrapper_91_reset = reset; // @[:@24230.4]
  assign RetimeWrapper_91_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@24232.4]
  assign RetimeWrapper_91_io_in = _T_2489 & io_rPort_7_en_0; // @[package.scala 94:16:@24231.4]
  assign RetimeWrapper_92_clock = clock; // @[:@24237.4]
  assign RetimeWrapper_92_reset = reset; // @[:@24238.4]
  assign RetimeWrapper_92_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@24240.4]
  assign RetimeWrapper_92_io_in = _T_2673 & io_rPort_7_en_0; // @[package.scala 94:16:@24239.4]
  assign RetimeWrapper_93_clock = clock; // @[:@24245.4]
  assign RetimeWrapper_93_reset = reset; // @[:@24246.4]
  assign RetimeWrapper_93_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@24248.4]
  assign RetimeWrapper_93_io_in = _T_2857 & io_rPort_7_en_0; // @[package.scala 94:16:@24247.4]
  assign RetimeWrapper_94_clock = clock; // @[:@24253.4]
  assign RetimeWrapper_94_reset = reset; // @[:@24254.4]
  assign RetimeWrapper_94_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@24256.4]
  assign RetimeWrapper_94_io_in = _T_3041 & io_rPort_7_en_0; // @[package.scala 94:16:@24255.4]
  assign RetimeWrapper_95_clock = clock; // @[:@24261.4]
  assign RetimeWrapper_95_reset = reset; // @[:@24262.4]
  assign RetimeWrapper_95_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@24264.4]
  assign RetimeWrapper_95_io_in = _T_3225 & io_rPort_7_en_0; // @[package.scala 94:16:@24263.4]
  assign RetimeWrapper_96_clock = clock; // @[:@24317.4]
  assign RetimeWrapper_96_reset = reset; // @[:@24318.4]
  assign RetimeWrapper_96_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@24320.4]
  assign RetimeWrapper_96_io_in = _T_1207 & io_rPort_8_en_0; // @[package.scala 94:16:@24319.4]
  assign RetimeWrapper_97_clock = clock; // @[:@24325.4]
  assign RetimeWrapper_97_reset = reset; // @[:@24326.4]
  assign RetimeWrapper_97_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@24328.4]
  assign RetimeWrapper_97_io_in = _T_1391 & io_rPort_8_en_0; // @[package.scala 94:16:@24327.4]
  assign RetimeWrapper_98_clock = clock; // @[:@24333.4]
  assign RetimeWrapper_98_reset = reset; // @[:@24334.4]
  assign RetimeWrapper_98_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@24336.4]
  assign RetimeWrapper_98_io_in = _T_1575 & io_rPort_8_en_0; // @[package.scala 94:16:@24335.4]
  assign RetimeWrapper_99_clock = clock; // @[:@24341.4]
  assign RetimeWrapper_99_reset = reset; // @[:@24342.4]
  assign RetimeWrapper_99_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@24344.4]
  assign RetimeWrapper_99_io_in = _T_1759 & io_rPort_8_en_0; // @[package.scala 94:16:@24343.4]
  assign RetimeWrapper_100_clock = clock; // @[:@24349.4]
  assign RetimeWrapper_100_reset = reset; // @[:@24350.4]
  assign RetimeWrapper_100_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@24352.4]
  assign RetimeWrapper_100_io_in = _T_1943 & io_rPort_8_en_0; // @[package.scala 94:16:@24351.4]
  assign RetimeWrapper_101_clock = clock; // @[:@24357.4]
  assign RetimeWrapper_101_reset = reset; // @[:@24358.4]
  assign RetimeWrapper_101_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@24360.4]
  assign RetimeWrapper_101_io_in = _T_2127 & io_rPort_8_en_0; // @[package.scala 94:16:@24359.4]
  assign RetimeWrapper_102_clock = clock; // @[:@24365.4]
  assign RetimeWrapper_102_reset = reset; // @[:@24366.4]
  assign RetimeWrapper_102_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@24368.4]
  assign RetimeWrapper_102_io_in = _T_2311 & io_rPort_8_en_0; // @[package.scala 94:16:@24367.4]
  assign RetimeWrapper_103_clock = clock; // @[:@24373.4]
  assign RetimeWrapper_103_reset = reset; // @[:@24374.4]
  assign RetimeWrapper_103_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@24376.4]
  assign RetimeWrapper_103_io_in = _T_2495 & io_rPort_8_en_0; // @[package.scala 94:16:@24375.4]
  assign RetimeWrapper_104_clock = clock; // @[:@24381.4]
  assign RetimeWrapper_104_reset = reset; // @[:@24382.4]
  assign RetimeWrapper_104_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@24384.4]
  assign RetimeWrapper_104_io_in = _T_2679 & io_rPort_8_en_0; // @[package.scala 94:16:@24383.4]
  assign RetimeWrapper_105_clock = clock; // @[:@24389.4]
  assign RetimeWrapper_105_reset = reset; // @[:@24390.4]
  assign RetimeWrapper_105_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@24392.4]
  assign RetimeWrapper_105_io_in = _T_2863 & io_rPort_8_en_0; // @[package.scala 94:16:@24391.4]
  assign RetimeWrapper_106_clock = clock; // @[:@24397.4]
  assign RetimeWrapper_106_reset = reset; // @[:@24398.4]
  assign RetimeWrapper_106_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@24400.4]
  assign RetimeWrapper_106_io_in = _T_3047 & io_rPort_8_en_0; // @[package.scala 94:16:@24399.4]
  assign RetimeWrapper_107_clock = clock; // @[:@24405.4]
  assign RetimeWrapper_107_reset = reset; // @[:@24406.4]
  assign RetimeWrapper_107_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@24408.4]
  assign RetimeWrapper_107_io_in = _T_3231 & io_rPort_8_en_0; // @[package.scala 94:16:@24407.4]
  assign RetimeWrapper_108_clock = clock; // @[:@24461.4]
  assign RetimeWrapper_108_reset = reset; // @[:@24462.4]
  assign RetimeWrapper_108_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@24464.4]
  assign RetimeWrapper_108_io_in = _T_1299 & io_rPort_9_en_0; // @[package.scala 94:16:@24463.4]
  assign RetimeWrapper_109_clock = clock; // @[:@24469.4]
  assign RetimeWrapper_109_reset = reset; // @[:@24470.4]
  assign RetimeWrapper_109_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@24472.4]
  assign RetimeWrapper_109_io_in = _T_1483 & io_rPort_9_en_0; // @[package.scala 94:16:@24471.4]
  assign RetimeWrapper_110_clock = clock; // @[:@24477.4]
  assign RetimeWrapper_110_reset = reset; // @[:@24478.4]
  assign RetimeWrapper_110_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@24480.4]
  assign RetimeWrapper_110_io_in = _T_1667 & io_rPort_9_en_0; // @[package.scala 94:16:@24479.4]
  assign RetimeWrapper_111_clock = clock; // @[:@24485.4]
  assign RetimeWrapper_111_reset = reset; // @[:@24486.4]
  assign RetimeWrapper_111_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@24488.4]
  assign RetimeWrapper_111_io_in = _T_1851 & io_rPort_9_en_0; // @[package.scala 94:16:@24487.4]
  assign RetimeWrapper_112_clock = clock; // @[:@24493.4]
  assign RetimeWrapper_112_reset = reset; // @[:@24494.4]
  assign RetimeWrapper_112_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@24496.4]
  assign RetimeWrapper_112_io_in = _T_2035 & io_rPort_9_en_0; // @[package.scala 94:16:@24495.4]
  assign RetimeWrapper_113_clock = clock; // @[:@24501.4]
  assign RetimeWrapper_113_reset = reset; // @[:@24502.4]
  assign RetimeWrapper_113_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@24504.4]
  assign RetimeWrapper_113_io_in = _T_2219 & io_rPort_9_en_0; // @[package.scala 94:16:@24503.4]
  assign RetimeWrapper_114_clock = clock; // @[:@24509.4]
  assign RetimeWrapper_114_reset = reset; // @[:@24510.4]
  assign RetimeWrapper_114_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@24512.4]
  assign RetimeWrapper_114_io_in = _T_2403 & io_rPort_9_en_0; // @[package.scala 94:16:@24511.4]
  assign RetimeWrapper_115_clock = clock; // @[:@24517.4]
  assign RetimeWrapper_115_reset = reset; // @[:@24518.4]
  assign RetimeWrapper_115_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@24520.4]
  assign RetimeWrapper_115_io_in = _T_2587 & io_rPort_9_en_0; // @[package.scala 94:16:@24519.4]
  assign RetimeWrapper_116_clock = clock; // @[:@24525.4]
  assign RetimeWrapper_116_reset = reset; // @[:@24526.4]
  assign RetimeWrapper_116_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@24528.4]
  assign RetimeWrapper_116_io_in = _T_2771 & io_rPort_9_en_0; // @[package.scala 94:16:@24527.4]
  assign RetimeWrapper_117_clock = clock; // @[:@24533.4]
  assign RetimeWrapper_117_reset = reset; // @[:@24534.4]
  assign RetimeWrapper_117_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@24536.4]
  assign RetimeWrapper_117_io_in = _T_2955 & io_rPort_9_en_0; // @[package.scala 94:16:@24535.4]
  assign RetimeWrapper_118_clock = clock; // @[:@24541.4]
  assign RetimeWrapper_118_reset = reset; // @[:@24542.4]
  assign RetimeWrapper_118_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@24544.4]
  assign RetimeWrapper_118_io_in = _T_3139 & io_rPort_9_en_0; // @[package.scala 94:16:@24543.4]
  assign RetimeWrapper_119_clock = clock; // @[:@24549.4]
  assign RetimeWrapper_119_reset = reset; // @[:@24550.4]
  assign RetimeWrapper_119_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@24552.4]
  assign RetimeWrapper_119_io_in = _T_3323 & io_rPort_9_en_0; // @[package.scala 94:16:@24551.4]
  assign RetimeWrapper_120_clock = clock; // @[:@24605.4]
  assign RetimeWrapper_120_reset = reset; // @[:@24606.4]
  assign RetimeWrapper_120_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@24608.4]
  assign RetimeWrapper_120_io_in = _T_1213 & io_rPort_10_en_0; // @[package.scala 94:16:@24607.4]
  assign RetimeWrapper_121_clock = clock; // @[:@24613.4]
  assign RetimeWrapper_121_reset = reset; // @[:@24614.4]
  assign RetimeWrapper_121_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@24616.4]
  assign RetimeWrapper_121_io_in = _T_1397 & io_rPort_10_en_0; // @[package.scala 94:16:@24615.4]
  assign RetimeWrapper_122_clock = clock; // @[:@24621.4]
  assign RetimeWrapper_122_reset = reset; // @[:@24622.4]
  assign RetimeWrapper_122_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@24624.4]
  assign RetimeWrapper_122_io_in = _T_1581 & io_rPort_10_en_0; // @[package.scala 94:16:@24623.4]
  assign RetimeWrapper_123_clock = clock; // @[:@24629.4]
  assign RetimeWrapper_123_reset = reset; // @[:@24630.4]
  assign RetimeWrapper_123_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@24632.4]
  assign RetimeWrapper_123_io_in = _T_1765 & io_rPort_10_en_0; // @[package.scala 94:16:@24631.4]
  assign RetimeWrapper_124_clock = clock; // @[:@24637.4]
  assign RetimeWrapper_124_reset = reset; // @[:@24638.4]
  assign RetimeWrapper_124_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@24640.4]
  assign RetimeWrapper_124_io_in = _T_1949 & io_rPort_10_en_0; // @[package.scala 94:16:@24639.4]
  assign RetimeWrapper_125_clock = clock; // @[:@24645.4]
  assign RetimeWrapper_125_reset = reset; // @[:@24646.4]
  assign RetimeWrapper_125_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@24648.4]
  assign RetimeWrapper_125_io_in = _T_2133 & io_rPort_10_en_0; // @[package.scala 94:16:@24647.4]
  assign RetimeWrapper_126_clock = clock; // @[:@24653.4]
  assign RetimeWrapper_126_reset = reset; // @[:@24654.4]
  assign RetimeWrapper_126_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@24656.4]
  assign RetimeWrapper_126_io_in = _T_2317 & io_rPort_10_en_0; // @[package.scala 94:16:@24655.4]
  assign RetimeWrapper_127_clock = clock; // @[:@24661.4]
  assign RetimeWrapper_127_reset = reset; // @[:@24662.4]
  assign RetimeWrapper_127_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@24664.4]
  assign RetimeWrapper_127_io_in = _T_2501 & io_rPort_10_en_0; // @[package.scala 94:16:@24663.4]
  assign RetimeWrapper_128_clock = clock; // @[:@24669.4]
  assign RetimeWrapper_128_reset = reset; // @[:@24670.4]
  assign RetimeWrapper_128_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@24672.4]
  assign RetimeWrapper_128_io_in = _T_2685 & io_rPort_10_en_0; // @[package.scala 94:16:@24671.4]
  assign RetimeWrapper_129_clock = clock; // @[:@24677.4]
  assign RetimeWrapper_129_reset = reset; // @[:@24678.4]
  assign RetimeWrapper_129_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@24680.4]
  assign RetimeWrapper_129_io_in = _T_2869 & io_rPort_10_en_0; // @[package.scala 94:16:@24679.4]
  assign RetimeWrapper_130_clock = clock; // @[:@24685.4]
  assign RetimeWrapper_130_reset = reset; // @[:@24686.4]
  assign RetimeWrapper_130_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@24688.4]
  assign RetimeWrapper_130_io_in = _T_3053 & io_rPort_10_en_0; // @[package.scala 94:16:@24687.4]
  assign RetimeWrapper_131_clock = clock; // @[:@24693.4]
  assign RetimeWrapper_131_reset = reset; // @[:@24694.4]
  assign RetimeWrapper_131_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@24696.4]
  assign RetimeWrapper_131_io_in = _T_3237 & io_rPort_10_en_0; // @[package.scala 94:16:@24695.4]
  assign RetimeWrapper_132_clock = clock; // @[:@24749.4]
  assign RetimeWrapper_132_reset = reset; // @[:@24750.4]
  assign RetimeWrapper_132_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24752.4]
  assign RetimeWrapper_132_io_in = _T_1219 & io_rPort_11_en_0; // @[package.scala 94:16:@24751.4]
  assign RetimeWrapper_133_clock = clock; // @[:@24757.4]
  assign RetimeWrapper_133_reset = reset; // @[:@24758.4]
  assign RetimeWrapper_133_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24760.4]
  assign RetimeWrapper_133_io_in = _T_1403 & io_rPort_11_en_0; // @[package.scala 94:16:@24759.4]
  assign RetimeWrapper_134_clock = clock; // @[:@24765.4]
  assign RetimeWrapper_134_reset = reset; // @[:@24766.4]
  assign RetimeWrapper_134_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24768.4]
  assign RetimeWrapper_134_io_in = _T_1587 & io_rPort_11_en_0; // @[package.scala 94:16:@24767.4]
  assign RetimeWrapper_135_clock = clock; // @[:@24773.4]
  assign RetimeWrapper_135_reset = reset; // @[:@24774.4]
  assign RetimeWrapper_135_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24776.4]
  assign RetimeWrapper_135_io_in = _T_1771 & io_rPort_11_en_0; // @[package.scala 94:16:@24775.4]
  assign RetimeWrapper_136_clock = clock; // @[:@24781.4]
  assign RetimeWrapper_136_reset = reset; // @[:@24782.4]
  assign RetimeWrapper_136_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24784.4]
  assign RetimeWrapper_136_io_in = _T_1955 & io_rPort_11_en_0; // @[package.scala 94:16:@24783.4]
  assign RetimeWrapper_137_clock = clock; // @[:@24789.4]
  assign RetimeWrapper_137_reset = reset; // @[:@24790.4]
  assign RetimeWrapper_137_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24792.4]
  assign RetimeWrapper_137_io_in = _T_2139 & io_rPort_11_en_0; // @[package.scala 94:16:@24791.4]
  assign RetimeWrapper_138_clock = clock; // @[:@24797.4]
  assign RetimeWrapper_138_reset = reset; // @[:@24798.4]
  assign RetimeWrapper_138_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24800.4]
  assign RetimeWrapper_138_io_in = _T_2323 & io_rPort_11_en_0; // @[package.scala 94:16:@24799.4]
  assign RetimeWrapper_139_clock = clock; // @[:@24805.4]
  assign RetimeWrapper_139_reset = reset; // @[:@24806.4]
  assign RetimeWrapper_139_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24808.4]
  assign RetimeWrapper_139_io_in = _T_2507 & io_rPort_11_en_0; // @[package.scala 94:16:@24807.4]
  assign RetimeWrapper_140_clock = clock; // @[:@24813.4]
  assign RetimeWrapper_140_reset = reset; // @[:@24814.4]
  assign RetimeWrapper_140_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24816.4]
  assign RetimeWrapper_140_io_in = _T_2691 & io_rPort_11_en_0; // @[package.scala 94:16:@24815.4]
  assign RetimeWrapper_141_clock = clock; // @[:@24821.4]
  assign RetimeWrapper_141_reset = reset; // @[:@24822.4]
  assign RetimeWrapper_141_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24824.4]
  assign RetimeWrapper_141_io_in = _T_2875 & io_rPort_11_en_0; // @[package.scala 94:16:@24823.4]
  assign RetimeWrapper_142_clock = clock; // @[:@24829.4]
  assign RetimeWrapper_142_reset = reset; // @[:@24830.4]
  assign RetimeWrapper_142_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24832.4]
  assign RetimeWrapper_142_io_in = _T_3059 & io_rPort_11_en_0; // @[package.scala 94:16:@24831.4]
  assign RetimeWrapper_143_clock = clock; // @[:@24837.4]
  assign RetimeWrapper_143_reset = reset; // @[:@24838.4]
  assign RetimeWrapper_143_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24840.4]
  assign RetimeWrapper_143_io_in = _T_3243 & io_rPort_11_en_0; // @[package.scala 94:16:@24839.4]
  assign RetimeWrapper_144_clock = clock; // @[:@24893.4]
  assign RetimeWrapper_144_reset = reset; // @[:@24894.4]
  assign RetimeWrapper_144_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@24896.4]
  assign RetimeWrapper_144_io_in = _T_1305 & io_rPort_12_en_0; // @[package.scala 94:16:@24895.4]
  assign RetimeWrapper_145_clock = clock; // @[:@24901.4]
  assign RetimeWrapper_145_reset = reset; // @[:@24902.4]
  assign RetimeWrapper_145_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@24904.4]
  assign RetimeWrapper_145_io_in = _T_1489 & io_rPort_12_en_0; // @[package.scala 94:16:@24903.4]
  assign RetimeWrapper_146_clock = clock; // @[:@24909.4]
  assign RetimeWrapper_146_reset = reset; // @[:@24910.4]
  assign RetimeWrapper_146_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@24912.4]
  assign RetimeWrapper_146_io_in = _T_1673 & io_rPort_12_en_0; // @[package.scala 94:16:@24911.4]
  assign RetimeWrapper_147_clock = clock; // @[:@24917.4]
  assign RetimeWrapper_147_reset = reset; // @[:@24918.4]
  assign RetimeWrapper_147_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@24920.4]
  assign RetimeWrapper_147_io_in = _T_1857 & io_rPort_12_en_0; // @[package.scala 94:16:@24919.4]
  assign RetimeWrapper_148_clock = clock; // @[:@24925.4]
  assign RetimeWrapper_148_reset = reset; // @[:@24926.4]
  assign RetimeWrapper_148_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@24928.4]
  assign RetimeWrapper_148_io_in = _T_2041 & io_rPort_12_en_0; // @[package.scala 94:16:@24927.4]
  assign RetimeWrapper_149_clock = clock; // @[:@24933.4]
  assign RetimeWrapper_149_reset = reset; // @[:@24934.4]
  assign RetimeWrapper_149_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@24936.4]
  assign RetimeWrapper_149_io_in = _T_2225 & io_rPort_12_en_0; // @[package.scala 94:16:@24935.4]
  assign RetimeWrapper_150_clock = clock; // @[:@24941.4]
  assign RetimeWrapper_150_reset = reset; // @[:@24942.4]
  assign RetimeWrapper_150_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@24944.4]
  assign RetimeWrapper_150_io_in = _T_2409 & io_rPort_12_en_0; // @[package.scala 94:16:@24943.4]
  assign RetimeWrapper_151_clock = clock; // @[:@24949.4]
  assign RetimeWrapper_151_reset = reset; // @[:@24950.4]
  assign RetimeWrapper_151_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@24952.4]
  assign RetimeWrapper_151_io_in = _T_2593 & io_rPort_12_en_0; // @[package.scala 94:16:@24951.4]
  assign RetimeWrapper_152_clock = clock; // @[:@24957.4]
  assign RetimeWrapper_152_reset = reset; // @[:@24958.4]
  assign RetimeWrapper_152_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@24960.4]
  assign RetimeWrapper_152_io_in = _T_2777 & io_rPort_12_en_0; // @[package.scala 94:16:@24959.4]
  assign RetimeWrapper_153_clock = clock; // @[:@24965.4]
  assign RetimeWrapper_153_reset = reset; // @[:@24966.4]
  assign RetimeWrapper_153_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@24968.4]
  assign RetimeWrapper_153_io_in = _T_2961 & io_rPort_12_en_0; // @[package.scala 94:16:@24967.4]
  assign RetimeWrapper_154_clock = clock; // @[:@24973.4]
  assign RetimeWrapper_154_reset = reset; // @[:@24974.4]
  assign RetimeWrapper_154_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@24976.4]
  assign RetimeWrapper_154_io_in = _T_3145 & io_rPort_12_en_0; // @[package.scala 94:16:@24975.4]
  assign RetimeWrapper_155_clock = clock; // @[:@24981.4]
  assign RetimeWrapper_155_reset = reset; // @[:@24982.4]
  assign RetimeWrapper_155_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@24984.4]
  assign RetimeWrapper_155_io_in = _T_3329 & io_rPort_12_en_0; // @[package.scala 94:16:@24983.4]
  assign RetimeWrapper_156_clock = clock; // @[:@25037.4]
  assign RetimeWrapper_156_reset = reset; // @[:@25038.4]
  assign RetimeWrapper_156_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@25040.4]
  assign RetimeWrapper_156_io_in = _T_1311 & io_rPort_13_en_0; // @[package.scala 94:16:@25039.4]
  assign RetimeWrapper_157_clock = clock; // @[:@25045.4]
  assign RetimeWrapper_157_reset = reset; // @[:@25046.4]
  assign RetimeWrapper_157_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@25048.4]
  assign RetimeWrapper_157_io_in = _T_1495 & io_rPort_13_en_0; // @[package.scala 94:16:@25047.4]
  assign RetimeWrapper_158_clock = clock; // @[:@25053.4]
  assign RetimeWrapper_158_reset = reset; // @[:@25054.4]
  assign RetimeWrapper_158_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@25056.4]
  assign RetimeWrapper_158_io_in = _T_1679 & io_rPort_13_en_0; // @[package.scala 94:16:@25055.4]
  assign RetimeWrapper_159_clock = clock; // @[:@25061.4]
  assign RetimeWrapper_159_reset = reset; // @[:@25062.4]
  assign RetimeWrapper_159_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@25064.4]
  assign RetimeWrapper_159_io_in = _T_1863 & io_rPort_13_en_0; // @[package.scala 94:16:@25063.4]
  assign RetimeWrapper_160_clock = clock; // @[:@25069.4]
  assign RetimeWrapper_160_reset = reset; // @[:@25070.4]
  assign RetimeWrapper_160_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@25072.4]
  assign RetimeWrapper_160_io_in = _T_2047 & io_rPort_13_en_0; // @[package.scala 94:16:@25071.4]
  assign RetimeWrapper_161_clock = clock; // @[:@25077.4]
  assign RetimeWrapper_161_reset = reset; // @[:@25078.4]
  assign RetimeWrapper_161_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@25080.4]
  assign RetimeWrapper_161_io_in = _T_2231 & io_rPort_13_en_0; // @[package.scala 94:16:@25079.4]
  assign RetimeWrapper_162_clock = clock; // @[:@25085.4]
  assign RetimeWrapper_162_reset = reset; // @[:@25086.4]
  assign RetimeWrapper_162_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@25088.4]
  assign RetimeWrapper_162_io_in = _T_2415 & io_rPort_13_en_0; // @[package.scala 94:16:@25087.4]
  assign RetimeWrapper_163_clock = clock; // @[:@25093.4]
  assign RetimeWrapper_163_reset = reset; // @[:@25094.4]
  assign RetimeWrapper_163_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@25096.4]
  assign RetimeWrapper_163_io_in = _T_2599 & io_rPort_13_en_0; // @[package.scala 94:16:@25095.4]
  assign RetimeWrapper_164_clock = clock; // @[:@25101.4]
  assign RetimeWrapper_164_reset = reset; // @[:@25102.4]
  assign RetimeWrapper_164_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@25104.4]
  assign RetimeWrapper_164_io_in = _T_2783 & io_rPort_13_en_0; // @[package.scala 94:16:@25103.4]
  assign RetimeWrapper_165_clock = clock; // @[:@25109.4]
  assign RetimeWrapper_165_reset = reset; // @[:@25110.4]
  assign RetimeWrapper_165_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@25112.4]
  assign RetimeWrapper_165_io_in = _T_2967 & io_rPort_13_en_0; // @[package.scala 94:16:@25111.4]
  assign RetimeWrapper_166_clock = clock; // @[:@25117.4]
  assign RetimeWrapper_166_reset = reset; // @[:@25118.4]
  assign RetimeWrapper_166_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@25120.4]
  assign RetimeWrapper_166_io_in = _T_3151 & io_rPort_13_en_0; // @[package.scala 94:16:@25119.4]
  assign RetimeWrapper_167_clock = clock; // @[:@25125.4]
  assign RetimeWrapper_167_reset = reset; // @[:@25126.4]
  assign RetimeWrapper_167_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@25128.4]
  assign RetimeWrapper_167_io_in = _T_3335 & io_rPort_13_en_0; // @[package.scala 94:16:@25127.4]
  assign RetimeWrapper_168_clock = clock; // @[:@25181.4]
  assign RetimeWrapper_168_reset = reset; // @[:@25182.4]
  assign RetimeWrapper_168_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@25184.4]
  assign RetimeWrapper_168_io_in = _T_1317 & io_rPort_14_en_0; // @[package.scala 94:16:@25183.4]
  assign RetimeWrapper_169_clock = clock; // @[:@25189.4]
  assign RetimeWrapper_169_reset = reset; // @[:@25190.4]
  assign RetimeWrapper_169_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@25192.4]
  assign RetimeWrapper_169_io_in = _T_1501 & io_rPort_14_en_0; // @[package.scala 94:16:@25191.4]
  assign RetimeWrapper_170_clock = clock; // @[:@25197.4]
  assign RetimeWrapper_170_reset = reset; // @[:@25198.4]
  assign RetimeWrapper_170_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@25200.4]
  assign RetimeWrapper_170_io_in = _T_1685 & io_rPort_14_en_0; // @[package.scala 94:16:@25199.4]
  assign RetimeWrapper_171_clock = clock; // @[:@25205.4]
  assign RetimeWrapper_171_reset = reset; // @[:@25206.4]
  assign RetimeWrapper_171_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@25208.4]
  assign RetimeWrapper_171_io_in = _T_1869 & io_rPort_14_en_0; // @[package.scala 94:16:@25207.4]
  assign RetimeWrapper_172_clock = clock; // @[:@25213.4]
  assign RetimeWrapper_172_reset = reset; // @[:@25214.4]
  assign RetimeWrapper_172_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@25216.4]
  assign RetimeWrapper_172_io_in = _T_2053 & io_rPort_14_en_0; // @[package.scala 94:16:@25215.4]
  assign RetimeWrapper_173_clock = clock; // @[:@25221.4]
  assign RetimeWrapper_173_reset = reset; // @[:@25222.4]
  assign RetimeWrapper_173_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@25224.4]
  assign RetimeWrapper_173_io_in = _T_2237 & io_rPort_14_en_0; // @[package.scala 94:16:@25223.4]
  assign RetimeWrapper_174_clock = clock; // @[:@25229.4]
  assign RetimeWrapper_174_reset = reset; // @[:@25230.4]
  assign RetimeWrapper_174_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@25232.4]
  assign RetimeWrapper_174_io_in = _T_2421 & io_rPort_14_en_0; // @[package.scala 94:16:@25231.4]
  assign RetimeWrapper_175_clock = clock; // @[:@25237.4]
  assign RetimeWrapper_175_reset = reset; // @[:@25238.4]
  assign RetimeWrapper_175_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@25240.4]
  assign RetimeWrapper_175_io_in = _T_2605 & io_rPort_14_en_0; // @[package.scala 94:16:@25239.4]
  assign RetimeWrapper_176_clock = clock; // @[:@25245.4]
  assign RetimeWrapper_176_reset = reset; // @[:@25246.4]
  assign RetimeWrapper_176_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@25248.4]
  assign RetimeWrapper_176_io_in = _T_2789 & io_rPort_14_en_0; // @[package.scala 94:16:@25247.4]
  assign RetimeWrapper_177_clock = clock; // @[:@25253.4]
  assign RetimeWrapper_177_reset = reset; // @[:@25254.4]
  assign RetimeWrapper_177_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@25256.4]
  assign RetimeWrapper_177_io_in = _T_2973 & io_rPort_14_en_0; // @[package.scala 94:16:@25255.4]
  assign RetimeWrapper_178_clock = clock; // @[:@25261.4]
  assign RetimeWrapper_178_reset = reset; // @[:@25262.4]
  assign RetimeWrapper_178_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@25264.4]
  assign RetimeWrapper_178_io_in = _T_3157 & io_rPort_14_en_0; // @[package.scala 94:16:@25263.4]
  assign RetimeWrapper_179_clock = clock; // @[:@25269.4]
  assign RetimeWrapper_179_reset = reset; // @[:@25270.4]
  assign RetimeWrapper_179_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@25272.4]
  assign RetimeWrapper_179_io_in = _T_3341 & io_rPort_14_en_0; // @[package.scala 94:16:@25271.4]
  assign RetimeWrapper_180_clock = clock; // @[:@25325.4]
  assign RetimeWrapper_180_reset = reset; // @[:@25326.4]
  assign RetimeWrapper_180_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@25328.4]
  assign RetimeWrapper_180_io_in = _T_1225 & io_rPort_15_en_0; // @[package.scala 94:16:@25327.4]
  assign RetimeWrapper_181_clock = clock; // @[:@25333.4]
  assign RetimeWrapper_181_reset = reset; // @[:@25334.4]
  assign RetimeWrapper_181_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@25336.4]
  assign RetimeWrapper_181_io_in = _T_1409 & io_rPort_15_en_0; // @[package.scala 94:16:@25335.4]
  assign RetimeWrapper_182_clock = clock; // @[:@25341.4]
  assign RetimeWrapper_182_reset = reset; // @[:@25342.4]
  assign RetimeWrapper_182_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@25344.4]
  assign RetimeWrapper_182_io_in = _T_1593 & io_rPort_15_en_0; // @[package.scala 94:16:@25343.4]
  assign RetimeWrapper_183_clock = clock; // @[:@25349.4]
  assign RetimeWrapper_183_reset = reset; // @[:@25350.4]
  assign RetimeWrapper_183_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@25352.4]
  assign RetimeWrapper_183_io_in = _T_1777 & io_rPort_15_en_0; // @[package.scala 94:16:@25351.4]
  assign RetimeWrapper_184_clock = clock; // @[:@25357.4]
  assign RetimeWrapper_184_reset = reset; // @[:@25358.4]
  assign RetimeWrapper_184_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@25360.4]
  assign RetimeWrapper_184_io_in = _T_1961 & io_rPort_15_en_0; // @[package.scala 94:16:@25359.4]
  assign RetimeWrapper_185_clock = clock; // @[:@25365.4]
  assign RetimeWrapper_185_reset = reset; // @[:@25366.4]
  assign RetimeWrapper_185_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@25368.4]
  assign RetimeWrapper_185_io_in = _T_2145 & io_rPort_15_en_0; // @[package.scala 94:16:@25367.4]
  assign RetimeWrapper_186_clock = clock; // @[:@25373.4]
  assign RetimeWrapper_186_reset = reset; // @[:@25374.4]
  assign RetimeWrapper_186_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@25376.4]
  assign RetimeWrapper_186_io_in = _T_2329 & io_rPort_15_en_0; // @[package.scala 94:16:@25375.4]
  assign RetimeWrapper_187_clock = clock; // @[:@25381.4]
  assign RetimeWrapper_187_reset = reset; // @[:@25382.4]
  assign RetimeWrapper_187_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@25384.4]
  assign RetimeWrapper_187_io_in = _T_2513 & io_rPort_15_en_0; // @[package.scala 94:16:@25383.4]
  assign RetimeWrapper_188_clock = clock; // @[:@25389.4]
  assign RetimeWrapper_188_reset = reset; // @[:@25390.4]
  assign RetimeWrapper_188_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@25392.4]
  assign RetimeWrapper_188_io_in = _T_2697 & io_rPort_15_en_0; // @[package.scala 94:16:@25391.4]
  assign RetimeWrapper_189_clock = clock; // @[:@25397.4]
  assign RetimeWrapper_189_reset = reset; // @[:@25398.4]
  assign RetimeWrapper_189_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@25400.4]
  assign RetimeWrapper_189_io_in = _T_2881 & io_rPort_15_en_0; // @[package.scala 94:16:@25399.4]
  assign RetimeWrapper_190_clock = clock; // @[:@25405.4]
  assign RetimeWrapper_190_reset = reset; // @[:@25406.4]
  assign RetimeWrapper_190_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@25408.4]
  assign RetimeWrapper_190_io_in = _T_3065 & io_rPort_15_en_0; // @[package.scala 94:16:@25407.4]
  assign RetimeWrapper_191_clock = clock; // @[:@25413.4]
  assign RetimeWrapper_191_reset = reset; // @[:@25414.4]
  assign RetimeWrapper_191_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@25416.4]
  assign RetimeWrapper_191_io_in = _T_3249 & io_rPort_15_en_0; // @[package.scala 94:16:@25415.4]
  assign RetimeWrapper_192_clock = clock; // @[:@25469.4]
  assign RetimeWrapper_192_reset = reset; // @[:@25470.4]
  assign RetimeWrapper_192_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@25472.4]
  assign RetimeWrapper_192_io_in = _T_1323 & io_rPort_16_en_0; // @[package.scala 94:16:@25471.4]
  assign RetimeWrapper_193_clock = clock; // @[:@25477.4]
  assign RetimeWrapper_193_reset = reset; // @[:@25478.4]
  assign RetimeWrapper_193_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@25480.4]
  assign RetimeWrapper_193_io_in = _T_1507 & io_rPort_16_en_0; // @[package.scala 94:16:@25479.4]
  assign RetimeWrapper_194_clock = clock; // @[:@25485.4]
  assign RetimeWrapper_194_reset = reset; // @[:@25486.4]
  assign RetimeWrapper_194_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@25488.4]
  assign RetimeWrapper_194_io_in = _T_1691 & io_rPort_16_en_0; // @[package.scala 94:16:@25487.4]
  assign RetimeWrapper_195_clock = clock; // @[:@25493.4]
  assign RetimeWrapper_195_reset = reset; // @[:@25494.4]
  assign RetimeWrapper_195_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@25496.4]
  assign RetimeWrapper_195_io_in = _T_1875 & io_rPort_16_en_0; // @[package.scala 94:16:@25495.4]
  assign RetimeWrapper_196_clock = clock; // @[:@25501.4]
  assign RetimeWrapper_196_reset = reset; // @[:@25502.4]
  assign RetimeWrapper_196_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@25504.4]
  assign RetimeWrapper_196_io_in = _T_2059 & io_rPort_16_en_0; // @[package.scala 94:16:@25503.4]
  assign RetimeWrapper_197_clock = clock; // @[:@25509.4]
  assign RetimeWrapper_197_reset = reset; // @[:@25510.4]
  assign RetimeWrapper_197_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@25512.4]
  assign RetimeWrapper_197_io_in = _T_2243 & io_rPort_16_en_0; // @[package.scala 94:16:@25511.4]
  assign RetimeWrapper_198_clock = clock; // @[:@25517.4]
  assign RetimeWrapper_198_reset = reset; // @[:@25518.4]
  assign RetimeWrapper_198_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@25520.4]
  assign RetimeWrapper_198_io_in = _T_2427 & io_rPort_16_en_0; // @[package.scala 94:16:@25519.4]
  assign RetimeWrapper_199_clock = clock; // @[:@25525.4]
  assign RetimeWrapper_199_reset = reset; // @[:@25526.4]
  assign RetimeWrapper_199_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@25528.4]
  assign RetimeWrapper_199_io_in = _T_2611 & io_rPort_16_en_0; // @[package.scala 94:16:@25527.4]
  assign RetimeWrapper_200_clock = clock; // @[:@25533.4]
  assign RetimeWrapper_200_reset = reset; // @[:@25534.4]
  assign RetimeWrapper_200_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@25536.4]
  assign RetimeWrapper_200_io_in = _T_2795 & io_rPort_16_en_0; // @[package.scala 94:16:@25535.4]
  assign RetimeWrapper_201_clock = clock; // @[:@25541.4]
  assign RetimeWrapper_201_reset = reset; // @[:@25542.4]
  assign RetimeWrapper_201_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@25544.4]
  assign RetimeWrapper_201_io_in = _T_2979 & io_rPort_16_en_0; // @[package.scala 94:16:@25543.4]
  assign RetimeWrapper_202_clock = clock; // @[:@25549.4]
  assign RetimeWrapper_202_reset = reset; // @[:@25550.4]
  assign RetimeWrapper_202_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@25552.4]
  assign RetimeWrapper_202_io_in = _T_3163 & io_rPort_16_en_0; // @[package.scala 94:16:@25551.4]
  assign RetimeWrapper_203_clock = clock; // @[:@25557.4]
  assign RetimeWrapper_203_reset = reset; // @[:@25558.4]
  assign RetimeWrapper_203_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@25560.4]
  assign RetimeWrapper_203_io_in = _T_3347 & io_rPort_16_en_0; // @[package.scala 94:16:@25559.4]
  assign RetimeWrapper_204_clock = clock; // @[:@25613.4]
  assign RetimeWrapper_204_reset = reset; // @[:@25614.4]
  assign RetimeWrapper_204_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@25616.4]
  assign RetimeWrapper_204_io_in = _T_1231 & io_rPort_17_en_0; // @[package.scala 94:16:@25615.4]
  assign RetimeWrapper_205_clock = clock; // @[:@25621.4]
  assign RetimeWrapper_205_reset = reset; // @[:@25622.4]
  assign RetimeWrapper_205_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@25624.4]
  assign RetimeWrapper_205_io_in = _T_1415 & io_rPort_17_en_0; // @[package.scala 94:16:@25623.4]
  assign RetimeWrapper_206_clock = clock; // @[:@25629.4]
  assign RetimeWrapper_206_reset = reset; // @[:@25630.4]
  assign RetimeWrapper_206_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@25632.4]
  assign RetimeWrapper_206_io_in = _T_1599 & io_rPort_17_en_0; // @[package.scala 94:16:@25631.4]
  assign RetimeWrapper_207_clock = clock; // @[:@25637.4]
  assign RetimeWrapper_207_reset = reset; // @[:@25638.4]
  assign RetimeWrapper_207_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@25640.4]
  assign RetimeWrapper_207_io_in = _T_1783 & io_rPort_17_en_0; // @[package.scala 94:16:@25639.4]
  assign RetimeWrapper_208_clock = clock; // @[:@25645.4]
  assign RetimeWrapper_208_reset = reset; // @[:@25646.4]
  assign RetimeWrapper_208_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@25648.4]
  assign RetimeWrapper_208_io_in = _T_1967 & io_rPort_17_en_0; // @[package.scala 94:16:@25647.4]
  assign RetimeWrapper_209_clock = clock; // @[:@25653.4]
  assign RetimeWrapper_209_reset = reset; // @[:@25654.4]
  assign RetimeWrapper_209_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@25656.4]
  assign RetimeWrapper_209_io_in = _T_2151 & io_rPort_17_en_0; // @[package.scala 94:16:@25655.4]
  assign RetimeWrapper_210_clock = clock; // @[:@25661.4]
  assign RetimeWrapper_210_reset = reset; // @[:@25662.4]
  assign RetimeWrapper_210_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@25664.4]
  assign RetimeWrapper_210_io_in = _T_2335 & io_rPort_17_en_0; // @[package.scala 94:16:@25663.4]
  assign RetimeWrapper_211_clock = clock; // @[:@25669.4]
  assign RetimeWrapper_211_reset = reset; // @[:@25670.4]
  assign RetimeWrapper_211_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@25672.4]
  assign RetimeWrapper_211_io_in = _T_2519 & io_rPort_17_en_0; // @[package.scala 94:16:@25671.4]
  assign RetimeWrapper_212_clock = clock; // @[:@25677.4]
  assign RetimeWrapper_212_reset = reset; // @[:@25678.4]
  assign RetimeWrapper_212_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@25680.4]
  assign RetimeWrapper_212_io_in = _T_2703 & io_rPort_17_en_0; // @[package.scala 94:16:@25679.4]
  assign RetimeWrapper_213_clock = clock; // @[:@25685.4]
  assign RetimeWrapper_213_reset = reset; // @[:@25686.4]
  assign RetimeWrapper_213_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@25688.4]
  assign RetimeWrapper_213_io_in = _T_2887 & io_rPort_17_en_0; // @[package.scala 94:16:@25687.4]
  assign RetimeWrapper_214_clock = clock; // @[:@25693.4]
  assign RetimeWrapper_214_reset = reset; // @[:@25694.4]
  assign RetimeWrapper_214_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@25696.4]
  assign RetimeWrapper_214_io_in = _T_3071 & io_rPort_17_en_0; // @[package.scala 94:16:@25695.4]
  assign RetimeWrapper_215_clock = clock; // @[:@25701.4]
  assign RetimeWrapper_215_reset = reset; // @[:@25702.4]
  assign RetimeWrapper_215_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@25704.4]
  assign RetimeWrapper_215_io_in = _T_3255 & io_rPort_17_en_0; // @[package.scala 94:16:@25703.4]
endmodule
module RetimeWrapper_297( // @[:@25732.2]
  input         clock, // @[:@25733.4]
  input         reset, // @[:@25734.4]
  input         io_flow, // @[:@25735.4]
  input  [31:0] io_in, // @[:@25735.4]
  output [31:0] io_out // @[:@25735.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@25737.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@25737.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@25737.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@25737.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@25737.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@25737.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@25737.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@25750.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@25749.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@25748.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@25747.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@25746.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@25744.4]
endmodule
module RetimeWrapper_298( // @[:@25764.2]
  input         clock, // @[:@25765.4]
  input         reset, // @[:@25766.4]
  input         io_flow, // @[:@25767.4]
  input  [31:0] io_in, // @[:@25767.4]
  output [31:0] io_out // @[:@25767.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@25769.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@25769.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@25769.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@25769.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@25769.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@25769.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(16)) sr ( // @[RetimeShiftRegister.scala 15:20:@25769.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@25782.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@25781.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@25780.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@25779.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@25778.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@25776.4]
endmodule
module fix2fixBox_10( // @[:@25784.2]
  input  [63:0] io_a, // @[:@25787.4]
  output [31:0] io_b // @[:@25787.4]
);
  assign io_b = io_a[31:0]; // @[Converter.scala 95:38:@25800.4]
endmodule
module x534( // @[:@25802.2]
  input         clock, // @[:@25803.4]
  input         reset, // @[:@25804.4]
  input  [31:0] io_a, // @[:@25805.4]
  input         io_flow, // @[:@25805.4]
  output [31:0] io_result // @[:@25805.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@25814.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@25814.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@25814.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@25814.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@25814.4]
  wire [63:0] fix2fixBox_io_a; // @[Math.scala 357:30:@25822.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 357:30:@25822.4]
  wire [31:0] _T_19; // @[package.scala 96:25:@25819.4 package.scala 96:25:@25820.4]
  wire [31:0] _GEN_0; // @[package.scala 94:16:@25817.4]
  RetimeWrapper_298 RetimeWrapper ( // @[package.scala 93:22:@25814.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  fix2fixBox_10 fix2fixBox ( // @[Math.scala 357:30:@25822.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign _T_19 = RetimeWrapper_io_out; // @[package.scala 96:25:@25819.4 package.scala 96:25:@25820.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 363:17:@25830.4]
  assign RetimeWrapper_clock = clock; // @[:@25815.4]
  assign RetimeWrapper_reset = reset; // @[:@25816.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@25818.4]
  assign _GEN_0 = io_a % 32'h6; // @[package.scala 94:16:@25817.4]
  assign RetimeWrapper_io_in = _GEN_0[31:0]; // @[package.scala 94:16:@25817.4]
  assign fix2fixBox_io_a = {{32'd0}, _T_19}; // @[Math.scala 358:23:@25825.4]
endmodule
module RetimeWrapper_300( // @[:@26033.2]
  input         clock, // @[:@26034.4]
  input         reset, // @[:@26035.4]
  input         io_flow, // @[:@26036.4]
  input  [31:0] io_in, // @[:@26036.4]
  output [31:0] io_out // @[:@26036.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@26038.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@26038.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@26038.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@26038.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@26038.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@26038.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(20)) sr ( // @[RetimeShiftRegister.scala 15:20:@26038.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@26051.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@26050.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@26049.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@26048.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@26047.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@26045.4]
endmodule
module x537_div( // @[:@26094.2]
  input         clock, // @[:@26095.4]
  input         reset, // @[:@26096.4]
  input  [31:0] io_a, // @[:@26097.4]
  input         io_flow, // @[:@26097.4]
  output [31:0] io_result // @[:@26097.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@26106.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@26106.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@26106.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@26106.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@26106.4]
  wire [31:0] __io_b; // @[Math.scala 709:24:@26119.4]
  wire [31:0] __io_result; // @[Math.scala 709:24:@26119.4]
  wire [31:0] _T_15; // @[FixedPoint.scala 24:59:@26103.4]
  wire [32:0] _T_17; // @[BigIPSim.scala 23:39:@26105.4]
  wire [32:0] _T_18; // @[package.scala 94:23:@26109.4]
  wire [31:0] _T_21; // @[package.scala 96:25:@26113.4]
  RetimeWrapper_300 RetimeWrapper ( // @[package.scala 93:22:@26106.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  _ _ ( // @[Math.scala 709:24:@26119.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  assign _T_15 = $signed(io_a); // @[FixedPoint.scala 24:59:@26103.4]
  assign _T_17 = $signed(_T_15) / $signed(32'sh6); // @[BigIPSim.scala 23:39:@26105.4]
  assign _T_18 = $unsigned(_T_17); // @[package.scala 94:23:@26109.4]
  assign _T_21 = $signed(RetimeWrapper_io_out); // @[package.scala 96:25:@26113.4]
  assign io_result = __io_result; // @[Math.scala 290:34:@26127.4]
  assign RetimeWrapper_clock = clock; // @[:@26107.4]
  assign RetimeWrapper_reset = reset; // @[:@26108.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@26111.4]
  assign RetimeWrapper_io_in = _T_18[31:0]; // @[package.scala 94:16:@26110.4]
  assign __io_b = $unsigned(_T_21); // @[Math.scala 710:17:@26122.4]
endmodule
module RetimeWrapper_301( // @[:@26141.2]
  input         clock, // @[:@26142.4]
  input         reset, // @[:@26143.4]
  input         io_flow, // @[:@26144.4]
  input  [31:0] io_in, // @[:@26144.4]
  output [31:0] io_out // @[:@26144.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@26146.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@26146.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@26146.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@26146.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@26146.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@26146.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(17)) sr ( // @[RetimeShiftRegister.scala 15:20:@26146.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@26159.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@26158.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@26157.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@26156.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@26155.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@26153.4]
endmodule
module RetimeWrapper_303( // @[:@26362.2]
  input         clock, // @[:@26363.4]
  input         reset, // @[:@26364.4]
  input         io_flow, // @[:@26365.4]
  input  [31:0] io_in, // @[:@26365.4]
  output [31:0] io_out // @[:@26365.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@26367.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@26367.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@26367.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@26367.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@26367.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@26367.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@26367.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@26380.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@26379.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@26378.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@26377.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@26376.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@26374.4]
endmodule
module RetimeWrapper_304( // @[:@26394.2]
  input         clock, // @[:@26395.4]
  input         reset, // @[:@26396.4]
  input         io_flow, // @[:@26397.4]
  input  [31:0] io_in, // @[:@26397.4]
  output [31:0] io_out // @[:@26397.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@26399.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@26399.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@26399.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@26399.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@26399.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@26399.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(8)) sr ( // @[RetimeShiftRegister.scala 15:20:@26399.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@26412.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@26411.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@26410.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@26409.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@26408.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@26406.4]
endmodule
module RetimeWrapper_305( // @[:@26426.2]
  input   clock, // @[:@26427.4]
  input   reset, // @[:@26428.4]
  input   io_flow, // @[:@26429.4]
  input   io_in, // @[:@26429.4]
  output  io_out // @[:@26429.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@26431.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@26431.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@26431.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@26431.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@26431.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@26431.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(24)) sr ( // @[RetimeShiftRegister.scala 15:20:@26431.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@26444.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@26443.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@26442.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@26441.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@26440.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@26438.4]
endmodule
module RetimeWrapper_307( // @[:@26490.2]
  input         clock, // @[:@26491.4]
  input         reset, // @[:@26492.4]
  input         io_flow, // @[:@26493.4]
  input  [31:0] io_in, // @[:@26493.4]
  output [31:0] io_out // @[:@26493.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@26495.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@26495.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@26495.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@26495.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@26495.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@26495.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(22)) sr ( // @[RetimeShiftRegister.scala 15:20:@26495.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@26508.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@26507.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@26506.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@26505.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@26504.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@26502.4]
endmodule
module RetimeWrapper_308( // @[:@26522.2]
  input        clock, // @[:@26523.4]
  input        reset, // @[:@26524.4]
  input        io_flow, // @[:@26525.4]
  input  [7:0] io_in, // @[:@26525.4]
  output [7:0] io_out // @[:@26525.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@26527.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@26527.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@26527.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@26527.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@26527.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@26527.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(23)) sr ( // @[RetimeShiftRegister.scala 15:20:@26527.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@26540.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@26539.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@26538.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@26537.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@26536.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@26534.4]
endmodule
module RetimeWrapper_313( // @[:@26963.2]
  input         clock, // @[:@26964.4]
  input         reset, // @[:@26965.4]
  input         io_flow, // @[:@26966.4]
  input  [31:0] io_in, // @[:@26966.4]
  output [31:0] io_out // @[:@26966.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@26968.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@26968.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@26968.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@26968.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@26968.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@26968.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(18)) sr ( // @[RetimeShiftRegister.scala 15:20:@26968.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@26981.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@26980.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@26979.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@26978.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@26977.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@26975.4]
endmodule
module RetimeWrapper_315( // @[:@27184.2]
  input         clock, // @[:@27185.4]
  input         reset, // @[:@27186.4]
  input         io_flow, // @[:@27187.4]
  input  [31:0] io_in, // @[:@27187.4]
  output [31:0] io_out // @[:@27187.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@27189.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@27189.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@27189.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@27189.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@27189.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@27189.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(7)) sr ( // @[RetimeShiftRegister.scala 15:20:@27189.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@27202.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@27201.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@27200.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@27199.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@27198.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@27196.4]
endmodule
module RetimeWrapper_335( // @[:@28700.2]
  input         clock, // @[:@28701.4]
  input         reset, // @[:@28702.4]
  input         io_flow, // @[:@28703.4]
  input  [31:0] io_in, // @[:@28703.4]
  output [31:0] io_out // @[:@28703.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@28705.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@28705.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@28705.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@28705.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@28705.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@28705.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(26)) sr ( // @[RetimeShiftRegister.scala 15:20:@28705.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@28718.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@28717.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@28716.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@28715.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@28714.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@28712.4]
endmodule
module RetimeWrapper_342( // @[:@29081.2]
  input         clock, // @[:@29082.4]
  input         reset, // @[:@29083.4]
  input         io_flow, // @[:@29084.4]
  input  [31:0] io_in, // @[:@29084.4]
  output [31:0] io_out // @[:@29084.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@29086.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@29086.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@29086.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@29086.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@29086.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@29086.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(19)) sr ( // @[RetimeShiftRegister.scala 15:20:@29086.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@29099.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@29098.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@29097.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@29096.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@29095.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@29093.4]
endmodule
module RetimeWrapper_345( // @[:@29334.2]
  input   clock, // @[:@29335.4]
  input   reset, // @[:@29336.4]
  input   io_flow, // @[:@29337.4]
  input   io_in, // @[:@29337.4]
  output  io_out // @[:@29337.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@29339.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@29339.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@29339.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@29339.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@29339.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@29339.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(48)) sr ( // @[RetimeShiftRegister.scala 15:20:@29339.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@29352.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@29351.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@29350.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@29349.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@29348.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@29346.4]
endmodule
module RetimeWrapper_346( // @[:@29366.2]
  input         clock, // @[:@29367.4]
  input         reset, // @[:@29368.4]
  input         io_flow, // @[:@29369.4]
  input  [31:0] io_in, // @[:@29369.4]
  output [31:0] io_out // @[:@29369.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@29371.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@29371.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@29371.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@29371.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@29371.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@29371.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(31)) sr ( // @[RetimeShiftRegister.scala 15:20:@29371.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@29384.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@29383.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@29382.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@29381.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@29380.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@29378.4]
endmodule
module RetimeWrapper_347( // @[:@29398.2]
  input         clock, // @[:@29399.4]
  input         reset, // @[:@29400.4]
  input         io_flow, // @[:@29401.4]
  input  [31:0] io_in, // @[:@29401.4]
  output [31:0] io_out // @[:@29401.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@29403.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@29403.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@29403.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@29403.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@29403.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@29403.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(21)) sr ( // @[RetimeShiftRegister.scala 15:20:@29403.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@29416.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@29415.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@29414.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@29413.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@29412.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@29410.4]
endmodule
module RetimeWrapper_349( // @[:@29462.2]
  input   clock, // @[:@29463.4]
  input   reset, // @[:@29464.4]
  input   io_flow, // @[:@29465.4]
  input   io_in, // @[:@29465.4]
  output  io_out // @[:@29465.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@29467.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@29467.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@29467.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@29467.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@29467.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@29467.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(20)) sr ( // @[RetimeShiftRegister.scala 15:20:@29467.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@29480.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@29479.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@29478.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@29477.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@29476.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@29474.4]
endmodule
module RetimeWrapper_370( // @[:@30605.2]
  input         clock, // @[:@30606.4]
  input         reset, // @[:@30607.4]
  input         io_flow, // @[:@30608.4]
  input  [31:0] io_in, // @[:@30608.4]
  output [31:0] io_out // @[:@30608.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@30610.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@30610.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@30610.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@30610.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@30610.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@30610.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(32)) sr ( // @[RetimeShiftRegister.scala 15:20:@30610.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@30623.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@30622.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@30621.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@30620.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@30619.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@30617.4]
endmodule
module RetimeWrapper_371( // @[:@30637.2]
  input   clock, // @[:@30638.4]
  input   reset, // @[:@30639.4]
  input   io_flow, // @[:@30640.4]
  input   io_in, // @[:@30640.4]
  output  io_out // @[:@30640.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@30642.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@30642.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@30642.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@30642.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@30642.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@30642.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(21)) sr ( // @[RetimeShiftRegister.scala 15:20:@30642.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@30655.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@30654.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@30653.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@30652.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@30651.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@30649.4]
endmodule
module RetimeWrapper_380( // @[:@31363.2]
  input         clock, // @[:@31364.4]
  input         reset, // @[:@31365.4]
  input         io_flow, // @[:@31366.4]
  input  [31:0] io_in, // @[:@31366.4]
  output [31:0] io_out // @[:@31366.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@31368.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@31368.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@31368.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@31368.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@31368.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@31368.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(5)) sr ( // @[RetimeShiftRegister.scala 15:20:@31368.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@31381.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@31380.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@31379.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@31378.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@31377.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@31375.4]
endmodule
module RetimeWrapper_445( // @[:@36395.2]
  input        clock, // @[:@36396.4]
  input        reset, // @[:@36397.4]
  input        io_flow, // @[:@36398.4]
  input  [9:0] io_in, // @[:@36398.4]
  output [9:0] io_out // @[:@36398.4]
);
  wire [9:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@36400.4]
  wire [9:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@36400.4]
  wire [9:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@36400.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@36400.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@36400.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@36400.4]
  RetimeShiftRegister #(.WIDTH(10), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@36400.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@36413.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@36412.4]
  assign sr_init = 10'h0; // @[RetimeShiftRegister.scala 19:16:@36411.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@36410.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@36409.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@36407.4]
endmodule
module RetimeWrapper_448( // @[:@36491.2]
  input        clock, // @[:@36492.4]
  input        reset, // @[:@36493.4]
  input        io_flow, // @[:@36494.4]
  input  [7:0] io_in, // @[:@36494.4]
  output [7:0] io_out // @[:@36494.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@36496.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@36496.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@36496.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@36496.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@36496.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@36496.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@36496.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@36509.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@36508.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@36507.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@36506.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@36505.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@36503.4]
endmodule
module SimBlackBoxesfix2fixBox_100( // @[:@36511.2]
  input  [7:0] io_a, // @[:@36514.4]
  output [8:0] io_b // @[:@36514.4]
);
  assign io_b = {1'h0,io_a}; // @[SimBlackBoxes.scala 99:40:@36528.4]
endmodule
module __96( // @[:@36530.2]
  input  [7:0] io_b, // @[:@36533.4]
  output [8:0] io_result // @[:@36533.4]
);
  wire [7:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@36538.4]
  wire [8:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@36538.4]
  SimBlackBoxesfix2fixBox_100 SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@36538.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@36551.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@36546.4]
endmodule
module fix2fixBox_49( // @[:@36595.2]
  input  [8:0] io_a, // @[:@36598.4]
  output [7:0] io_b // @[:@36598.4]
);
  assign io_b = io_a[7:0]; // @[Converter.scala 95:38:@36611.4]
endmodule
module x683_x15( // @[:@36613.2]
  input  [7:0] io_a, // @[:@36616.4]
  input  [7:0] io_b, // @[:@36616.4]
  output [7:0] io_result // @[:@36616.4]
);
  wire [7:0] __io_b; // @[Math.scala 709:24:@36624.4]
  wire [8:0] __io_result; // @[Math.scala 709:24:@36624.4]
  wire [7:0] __1_io_b; // @[Math.scala 709:24:@36631.4]
  wire [8:0] __1_io_result; // @[Math.scala 709:24:@36631.4]
  wire [8:0] fix2fixBox_io_a; // @[Math.scala 141:30:@36641.4]
  wire [7:0] fix2fixBox_io_b; // @[Math.scala 141:30:@36641.4]
  wire [8:0] a_upcast_number; // @[Math.scala 712:22:@36629.4 Math.scala 713:14:@36630.4]
  wire [8:0] b_upcast_number; // @[Math.scala 712:22:@36636.4 Math.scala 713:14:@36637.4]
  wire [9:0] _T_21; // @[Math.scala 136:37:@36638.4]
  __96 _ ( // @[Math.scala 709:24:@36624.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __96 __1 ( // @[Math.scala 709:24:@36631.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_49 fix2fixBox ( // @[Math.scala 141:30:@36641.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@36629.4 Math.scala 713:14:@36630.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@36636.4 Math.scala 713:14:@36637.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@36638.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@36649.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@36627.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@36634.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@36644.4]
endmodule
module fix2fixBox_56( // @[:@37703.2]
  input        clock, // @[:@37704.4]
  input        reset, // @[:@37705.4]
  input  [8:0] io_a, // @[:@37706.4]
  input        io_flow, // @[:@37706.4]
  output [7:0] io_b // @[:@37706.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@37719.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@37719.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@37719.4]
  wire [7:0] RetimeWrapper_io_in; // @[package.scala 93:22:@37719.4]
  wire [7:0] RetimeWrapper_io_out; // @[package.scala 93:22:@37719.4]
  RetimeWrapper_448 RetimeWrapper ( // @[package.scala 93:22:@37719.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@37726.4]
  assign RetimeWrapper_clock = clock; // @[:@37720.4]
  assign RetimeWrapper_reset = reset; // @[:@37721.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@37723.4]
  assign RetimeWrapper_io_in = io_a[7:0]; // @[package.scala 94:16:@37722.4]
endmodule
module x690_sum( // @[:@37728.2]
  input        clock, // @[:@37729.4]
  input        reset, // @[:@37730.4]
  input  [7:0] io_a, // @[:@37731.4]
  input  [7:0] io_b, // @[:@37731.4]
  input        io_flow, // @[:@37731.4]
  output [7:0] io_result // @[:@37731.4]
);
  wire [7:0] __io_b; // @[Math.scala 709:24:@37739.4]
  wire [8:0] __io_result; // @[Math.scala 709:24:@37739.4]
  wire [7:0] __1_io_b; // @[Math.scala 709:24:@37746.4]
  wire [8:0] __1_io_result; // @[Math.scala 709:24:@37746.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@37756.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@37756.4]
  wire [8:0] fix2fixBox_io_a; // @[Math.scala 141:30:@37756.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@37756.4]
  wire [7:0] fix2fixBox_io_b; // @[Math.scala 141:30:@37756.4]
  wire [8:0] a_upcast_number; // @[Math.scala 712:22:@37744.4 Math.scala 713:14:@37745.4]
  wire [8:0] b_upcast_number; // @[Math.scala 712:22:@37751.4 Math.scala 713:14:@37752.4]
  wire [9:0] _T_21; // @[Math.scala 136:37:@37753.4]
  __96 _ ( // @[Math.scala 709:24:@37739.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __96 __1 ( // @[Math.scala 709:24:@37746.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_56 fix2fixBox ( // @[Math.scala 141:30:@37756.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@37744.4 Math.scala 713:14:@37745.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@37751.4 Math.scala 713:14:@37752.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@37753.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@37764.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@37742.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@37749.4]
  assign fix2fixBox_clock = clock; // @[:@37757.4]
  assign fix2fixBox_reset = reset; // @[:@37758.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@37759.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@37762.4]
endmodule
module x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1( // @[:@42043.2]
  input          clock, // @[:@42044.4]
  input          reset, // @[:@42045.4]
  output         io_in_x481_TVALID, // @[:@42046.4]
  input          io_in_x481_TREADY, // @[:@42046.4]
  output [255:0] io_in_x481_TDATA, // @[:@42046.4]
  output         io_in_x480_TREADY, // @[:@42046.4]
  input  [255:0] io_in_x480_TDATA, // @[:@42046.4]
  input  [7:0]   io_in_x480_TID, // @[:@42046.4]
  input  [7:0]   io_in_x480_TDEST, // @[:@42046.4]
  input          io_sigsIn_backpressure, // @[:@42046.4]
  input          io_sigsIn_datapathEn, // @[:@42046.4]
  input          io_sigsIn_break, // @[:@42046.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_1, // @[:@42046.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_0, // @[:@42046.4]
  input          io_sigsIn_cchainOutputs_0_oobs_0, // @[:@42046.4]
  input          io_sigsIn_cchainOutputs_0_oobs_1, // @[:@42046.4]
  input          io_rr // @[:@42046.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@42060.4]
  wire [31:0] __io_result; // @[Math.scala 709:24:@42060.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@42072.4]
  wire [31:0] __1_io_result; // @[Math.scala 709:24:@42072.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@42095.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@42095.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@42095.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@42095.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@42095.4]
  wire  x525_lb_0_clock; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire  x525_lb_0_reset; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_rPort_17_banks_1; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_rPort_17_banks_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [8:0] x525_lb_0_io_rPort_17_ofs_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire  x525_lb_0_io_rPort_17_en_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire  x525_lb_0_io_rPort_17_backpressure; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [7:0] x525_lb_0_io_rPort_17_output_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_rPort_16_banks_1; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_rPort_16_banks_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [8:0] x525_lb_0_io_rPort_16_ofs_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire  x525_lb_0_io_rPort_16_en_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire  x525_lb_0_io_rPort_16_backpressure; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [7:0] x525_lb_0_io_rPort_16_output_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_rPort_15_banks_1; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_rPort_15_banks_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [8:0] x525_lb_0_io_rPort_15_ofs_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire  x525_lb_0_io_rPort_15_en_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire  x525_lb_0_io_rPort_15_backpressure; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [7:0] x525_lb_0_io_rPort_15_output_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_rPort_14_banks_1; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_rPort_14_banks_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [8:0] x525_lb_0_io_rPort_14_ofs_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire  x525_lb_0_io_rPort_14_en_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire  x525_lb_0_io_rPort_14_backpressure; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [7:0] x525_lb_0_io_rPort_14_output_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_rPort_13_banks_1; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_rPort_13_banks_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [8:0] x525_lb_0_io_rPort_13_ofs_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire  x525_lb_0_io_rPort_13_en_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire  x525_lb_0_io_rPort_13_backpressure; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [7:0] x525_lb_0_io_rPort_13_output_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_rPort_12_banks_1; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_rPort_12_banks_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [8:0] x525_lb_0_io_rPort_12_ofs_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire  x525_lb_0_io_rPort_12_en_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire  x525_lb_0_io_rPort_12_backpressure; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [7:0] x525_lb_0_io_rPort_12_output_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_rPort_11_banks_1; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_rPort_11_banks_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [8:0] x525_lb_0_io_rPort_11_ofs_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire  x525_lb_0_io_rPort_11_en_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire  x525_lb_0_io_rPort_11_backpressure; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [7:0] x525_lb_0_io_rPort_11_output_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_rPort_10_banks_1; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_rPort_10_banks_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [8:0] x525_lb_0_io_rPort_10_ofs_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire  x525_lb_0_io_rPort_10_en_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire  x525_lb_0_io_rPort_10_backpressure; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [7:0] x525_lb_0_io_rPort_10_output_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_rPort_9_banks_1; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_rPort_9_banks_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [8:0] x525_lb_0_io_rPort_9_ofs_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire  x525_lb_0_io_rPort_9_en_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire  x525_lb_0_io_rPort_9_backpressure; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [7:0] x525_lb_0_io_rPort_9_output_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_rPort_8_banks_1; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_rPort_8_banks_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [8:0] x525_lb_0_io_rPort_8_ofs_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire  x525_lb_0_io_rPort_8_en_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire  x525_lb_0_io_rPort_8_backpressure; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [7:0] x525_lb_0_io_rPort_8_output_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_rPort_7_banks_1; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_rPort_7_banks_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [8:0] x525_lb_0_io_rPort_7_ofs_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire  x525_lb_0_io_rPort_7_en_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire  x525_lb_0_io_rPort_7_backpressure; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [7:0] x525_lb_0_io_rPort_7_output_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_rPort_6_banks_1; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_rPort_6_banks_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [8:0] x525_lb_0_io_rPort_6_ofs_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire  x525_lb_0_io_rPort_6_en_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire  x525_lb_0_io_rPort_6_backpressure; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [7:0] x525_lb_0_io_rPort_6_output_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_rPort_5_banks_1; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_rPort_5_banks_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [8:0] x525_lb_0_io_rPort_5_ofs_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire  x525_lb_0_io_rPort_5_en_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire  x525_lb_0_io_rPort_5_backpressure; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [7:0] x525_lb_0_io_rPort_5_output_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_rPort_4_banks_1; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_rPort_4_banks_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [8:0] x525_lb_0_io_rPort_4_ofs_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire  x525_lb_0_io_rPort_4_en_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire  x525_lb_0_io_rPort_4_backpressure; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [7:0] x525_lb_0_io_rPort_4_output_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_rPort_3_banks_1; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_rPort_3_banks_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [8:0] x525_lb_0_io_rPort_3_ofs_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire  x525_lb_0_io_rPort_3_en_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire  x525_lb_0_io_rPort_3_backpressure; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [7:0] x525_lb_0_io_rPort_3_output_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_rPort_2_banks_1; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_rPort_2_banks_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [8:0] x525_lb_0_io_rPort_2_ofs_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire  x525_lb_0_io_rPort_2_en_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire  x525_lb_0_io_rPort_2_backpressure; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [7:0] x525_lb_0_io_rPort_2_output_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_rPort_1_banks_1; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_rPort_1_banks_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [8:0] x525_lb_0_io_rPort_1_ofs_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire  x525_lb_0_io_rPort_1_en_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire  x525_lb_0_io_rPort_1_backpressure; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [7:0] x525_lb_0_io_rPort_1_output_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_rPort_0_banks_1; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_rPort_0_banks_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [8:0] x525_lb_0_io_rPort_0_ofs_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire  x525_lb_0_io_rPort_0_en_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire  x525_lb_0_io_rPort_0_backpressure; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [7:0] x525_lb_0_io_rPort_0_output_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_wPort_3_banks_1; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_wPort_3_banks_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [8:0] x525_lb_0_io_wPort_3_ofs_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [7:0] x525_lb_0_io_wPort_3_data_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire  x525_lb_0_io_wPort_3_en_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_wPort_2_banks_1; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_wPort_2_banks_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [8:0] x525_lb_0_io_wPort_2_ofs_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [7:0] x525_lb_0_io_wPort_2_data_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire  x525_lb_0_io_wPort_2_en_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_wPort_1_banks_1; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_wPort_1_banks_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [8:0] x525_lb_0_io_wPort_1_ofs_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [7:0] x525_lb_0_io_wPort_1_data_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire  x525_lb_0_io_wPort_1_en_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_wPort_0_banks_1; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [2:0] x525_lb_0_io_wPort_0_banks_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [8:0] x525_lb_0_io_wPort_0_ofs_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire [7:0] x525_lb_0_io_wPort_0_data_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire  x525_lb_0_io_wPort_0_en_0; // @[m_x525_lb_0.scala 47:17:@42105.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@42311.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@42311.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@42311.4]
  wire [31:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@42311.4]
  wire [31:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@42311.4]
  wire  x534_1_clock; // @[Math.scala 366:24:@42333.4]
  wire  x534_1_reset; // @[Math.scala 366:24:@42333.4]
  wire [31:0] x534_1_io_a; // @[Math.scala 366:24:@42333.4]
  wire  x534_1_io_flow; // @[Math.scala 366:24:@42333.4]
  wire [31:0] x534_1_io_result; // @[Math.scala 366:24:@42333.4]
  wire  x803_sum_1_clock; // @[Math.scala 150:24:@42362.4]
  wire  x803_sum_1_reset; // @[Math.scala 150:24:@42362.4]
  wire [31:0] x803_sum_1_io_a; // @[Math.scala 150:24:@42362.4]
  wire [31:0] x803_sum_1_io_b; // @[Math.scala 150:24:@42362.4]
  wire  x803_sum_1_io_flow; // @[Math.scala 150:24:@42362.4]
  wire [31:0] x803_sum_1_io_result; // @[Math.scala 150:24:@42362.4]
  wire  x537_div_1_clock; // @[Math.scala 327:24:@42374.4]
  wire  x537_div_1_reset; // @[Math.scala 327:24:@42374.4]
  wire [31:0] x537_div_1_io_a; // @[Math.scala 327:24:@42374.4]
  wire  x537_div_1_io_flow; // @[Math.scala 327:24:@42374.4]
  wire [31:0] x537_div_1_io_result; // @[Math.scala 327:24:@42374.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@42384.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@42384.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@42384.4]
  wire [31:0] RetimeWrapper_2_io_in; // @[package.scala 93:22:@42384.4]
  wire [31:0] RetimeWrapper_2_io_out; // @[package.scala 93:22:@42384.4]
  wire  x538_sum_1_clock; // @[Math.scala 150:24:@42393.4]
  wire  x538_sum_1_reset; // @[Math.scala 150:24:@42393.4]
  wire [31:0] x538_sum_1_io_a; // @[Math.scala 150:24:@42393.4]
  wire [31:0] x538_sum_1_io_b; // @[Math.scala 150:24:@42393.4]
  wire  x538_sum_1_io_flow; // @[Math.scala 150:24:@42393.4]
  wire [31:0] x538_sum_1_io_result; // @[Math.scala 150:24:@42393.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@42403.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@42403.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@42403.4]
  wire [31:0] RetimeWrapper_3_io_in; // @[package.scala 93:22:@42403.4]
  wire [31:0] RetimeWrapper_3_io_out; // @[package.scala 93:22:@42403.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@42412.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@42412.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@42412.4]
  wire [31:0] RetimeWrapper_4_io_in; // @[package.scala 93:22:@42412.4]
  wire [31:0] RetimeWrapper_4_io_out; // @[package.scala 93:22:@42412.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@42421.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@42421.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@42421.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@42421.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@42421.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@42430.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@42430.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@42430.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@42430.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@42430.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@42439.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@42439.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@42439.4]
  wire [31:0] RetimeWrapper_7_io_in; // @[package.scala 93:22:@42439.4]
  wire [31:0] RetimeWrapper_7_io_out; // @[package.scala 93:22:@42439.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@42448.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@42448.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@42448.4]
  wire [7:0] RetimeWrapper_8_io_in; // @[package.scala 93:22:@42448.4]
  wire [7:0] RetimeWrapper_8_io_out; // @[package.scala 93:22:@42448.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@42459.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@42459.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@42459.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@42459.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@42459.4]
  wire  x540_rdcol_1_clock; // @[Math.scala 150:24:@42482.4]
  wire  x540_rdcol_1_reset; // @[Math.scala 150:24:@42482.4]
  wire [31:0] x540_rdcol_1_io_a; // @[Math.scala 150:24:@42482.4]
  wire [31:0] x540_rdcol_1_io_b; // @[Math.scala 150:24:@42482.4]
  wire  x540_rdcol_1_io_flow; // @[Math.scala 150:24:@42482.4]
  wire [31:0] x540_rdcol_1_io_result; // @[Math.scala 150:24:@42482.4]
  wire  x542_1_clock; // @[Math.scala 366:24:@42496.4]
  wire  x542_1_reset; // @[Math.scala 366:24:@42496.4]
  wire [31:0] x542_1_io_a; // @[Math.scala 366:24:@42496.4]
  wire  x542_1_io_flow; // @[Math.scala 366:24:@42496.4]
  wire [31:0] x542_1_io_result; // @[Math.scala 366:24:@42496.4]
  wire  x543_div_1_clock; // @[Math.scala 327:24:@42508.4]
  wire  x543_div_1_reset; // @[Math.scala 327:24:@42508.4]
  wire [31:0] x543_div_1_io_a; // @[Math.scala 327:24:@42508.4]
  wire  x543_div_1_io_flow; // @[Math.scala 327:24:@42508.4]
  wire [31:0] x543_div_1_io_result; // @[Math.scala 327:24:@42508.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@42518.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@42518.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@42518.4]
  wire [31:0] RetimeWrapper_10_io_in; // @[package.scala 93:22:@42518.4]
  wire [31:0] RetimeWrapper_10_io_out; // @[package.scala 93:22:@42518.4]
  wire  x544_sum_1_clock; // @[Math.scala 150:24:@42527.4]
  wire  x544_sum_1_reset; // @[Math.scala 150:24:@42527.4]
  wire [31:0] x544_sum_1_io_a; // @[Math.scala 150:24:@42527.4]
  wire [31:0] x544_sum_1_io_b; // @[Math.scala 150:24:@42527.4]
  wire  x544_sum_1_io_flow; // @[Math.scala 150:24:@42527.4]
  wire [31:0] x544_sum_1_io_result; // @[Math.scala 150:24:@42527.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@42537.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@42537.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@42537.4]
  wire [31:0] RetimeWrapper_11_io_in; // @[package.scala 93:22:@42537.4]
  wire [31:0] RetimeWrapper_11_io_out; // @[package.scala 93:22:@42537.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@42546.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@42546.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@42546.4]
  wire [7:0] RetimeWrapper_12_io_in; // @[package.scala 93:22:@42546.4]
  wire [7:0] RetimeWrapper_12_io_out; // @[package.scala 93:22:@42546.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@42555.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@42555.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@42555.4]
  wire [31:0] RetimeWrapper_13_io_in; // @[package.scala 93:22:@42555.4]
  wire [31:0] RetimeWrapper_13_io_out; // @[package.scala 93:22:@42555.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@42566.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@42566.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@42566.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@42566.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@42566.4]
  wire  x546_rdcol_1_clock; // @[Math.scala 150:24:@42589.4]
  wire  x546_rdcol_1_reset; // @[Math.scala 150:24:@42589.4]
  wire [31:0] x546_rdcol_1_io_a; // @[Math.scala 150:24:@42589.4]
  wire [31:0] x546_rdcol_1_io_b; // @[Math.scala 150:24:@42589.4]
  wire  x546_rdcol_1_io_flow; // @[Math.scala 150:24:@42589.4]
  wire [31:0] x546_rdcol_1_io_result; // @[Math.scala 150:24:@42589.4]
  wire  x548_1_clock; // @[Math.scala 366:24:@42603.4]
  wire  x548_1_reset; // @[Math.scala 366:24:@42603.4]
  wire [31:0] x548_1_io_a; // @[Math.scala 366:24:@42603.4]
  wire  x548_1_io_flow; // @[Math.scala 366:24:@42603.4]
  wire [31:0] x548_1_io_result; // @[Math.scala 366:24:@42603.4]
  wire  x549_div_1_clock; // @[Math.scala 327:24:@42615.4]
  wire  x549_div_1_reset; // @[Math.scala 327:24:@42615.4]
  wire [31:0] x549_div_1_io_a; // @[Math.scala 327:24:@42615.4]
  wire  x549_div_1_io_flow; // @[Math.scala 327:24:@42615.4]
  wire [31:0] x549_div_1_io_result; // @[Math.scala 327:24:@42615.4]
  wire  x550_sum_1_clock; // @[Math.scala 150:24:@42625.4]
  wire  x550_sum_1_reset; // @[Math.scala 150:24:@42625.4]
  wire [31:0] x550_sum_1_io_a; // @[Math.scala 150:24:@42625.4]
  wire [31:0] x550_sum_1_io_b; // @[Math.scala 150:24:@42625.4]
  wire  x550_sum_1_io_flow; // @[Math.scala 150:24:@42625.4]
  wire [31:0] x550_sum_1_io_result; // @[Math.scala 150:24:@42625.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@42635.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@42635.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@42635.4]
  wire [31:0] RetimeWrapper_15_io_in; // @[package.scala 93:22:@42635.4]
  wire [31:0] RetimeWrapper_15_io_out; // @[package.scala 93:22:@42635.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@42644.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@42644.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@42644.4]
  wire [7:0] RetimeWrapper_16_io_in; // @[package.scala 93:22:@42644.4]
  wire [7:0] RetimeWrapper_16_io_out; // @[package.scala 93:22:@42644.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@42653.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@42653.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@42653.4]
  wire [31:0] RetimeWrapper_17_io_in; // @[package.scala 93:22:@42653.4]
  wire [31:0] RetimeWrapper_17_io_out; // @[package.scala 93:22:@42653.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@42664.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@42664.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@42664.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@42664.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@42664.4]
  wire  x552_rdcol_1_clock; // @[Math.scala 150:24:@42687.4]
  wire  x552_rdcol_1_reset; // @[Math.scala 150:24:@42687.4]
  wire [31:0] x552_rdcol_1_io_a; // @[Math.scala 150:24:@42687.4]
  wire [31:0] x552_rdcol_1_io_b; // @[Math.scala 150:24:@42687.4]
  wire  x552_rdcol_1_io_flow; // @[Math.scala 150:24:@42687.4]
  wire [31:0] x552_rdcol_1_io_result; // @[Math.scala 150:24:@42687.4]
  wire  x554_1_clock; // @[Math.scala 366:24:@42703.4]
  wire  x554_1_reset; // @[Math.scala 366:24:@42703.4]
  wire [31:0] x554_1_io_a; // @[Math.scala 366:24:@42703.4]
  wire  x554_1_io_flow; // @[Math.scala 366:24:@42703.4]
  wire [31:0] x554_1_io_result; // @[Math.scala 366:24:@42703.4]
  wire  x555_div_1_clock; // @[Math.scala 327:24:@42715.4]
  wire  x555_div_1_reset; // @[Math.scala 327:24:@42715.4]
  wire [31:0] x555_div_1_io_a; // @[Math.scala 327:24:@42715.4]
  wire  x555_div_1_io_flow; // @[Math.scala 327:24:@42715.4]
  wire [31:0] x555_div_1_io_result; // @[Math.scala 327:24:@42715.4]
  wire  x556_sum_1_clock; // @[Math.scala 150:24:@42725.4]
  wire  x556_sum_1_reset; // @[Math.scala 150:24:@42725.4]
  wire [31:0] x556_sum_1_io_a; // @[Math.scala 150:24:@42725.4]
  wire [31:0] x556_sum_1_io_b; // @[Math.scala 150:24:@42725.4]
  wire  x556_sum_1_io_flow; // @[Math.scala 150:24:@42725.4]
  wire [31:0] x556_sum_1_io_result; // @[Math.scala 150:24:@42725.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@42735.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@42735.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@42735.4]
  wire [31:0] RetimeWrapper_19_io_in; // @[package.scala 93:22:@42735.4]
  wire [31:0] RetimeWrapper_19_io_out; // @[package.scala 93:22:@42735.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@42744.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@42744.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@42744.4]
  wire [7:0] RetimeWrapper_20_io_in; // @[package.scala 93:22:@42744.4]
  wire [7:0] RetimeWrapper_20_io_out; // @[package.scala 93:22:@42744.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@42753.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@42753.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@42753.4]
  wire [31:0] RetimeWrapper_21_io_in; // @[package.scala 93:22:@42753.4]
  wire [31:0] RetimeWrapper_21_io_out; // @[package.scala 93:22:@42753.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@42764.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@42764.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@42764.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@42764.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@42764.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@42785.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@42785.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@42785.4]
  wire [31:0] RetimeWrapper_23_io_in; // @[package.scala 93:22:@42785.4]
  wire [31:0] RetimeWrapper_23_io_out; // @[package.scala 93:22:@42785.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@42801.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@42801.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@42801.4]
  wire [31:0] RetimeWrapper_24_io_in; // @[package.scala 93:22:@42801.4]
  wire [31:0] RetimeWrapper_24_io_out; // @[package.scala 93:22:@42801.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@42819.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@42819.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@42819.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@42819.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@42819.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@42828.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@42828.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@42828.4]
  wire [31:0] RetimeWrapper_26_io_in; // @[package.scala 93:22:@42828.4]
  wire [31:0] RetimeWrapper_26_io_out; // @[package.scala 93:22:@42828.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@42842.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@42842.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@42842.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@42842.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@42842.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@42851.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@42851.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@42851.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@42851.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@42851.4]
  wire  x808_sum_1_clock; // @[Math.scala 150:24:@42896.4]
  wire  x808_sum_1_reset; // @[Math.scala 150:24:@42896.4]
  wire [31:0] x808_sum_1_io_a; // @[Math.scala 150:24:@42896.4]
  wire [31:0] x808_sum_1_io_b; // @[Math.scala 150:24:@42896.4]
  wire  x808_sum_1_io_flow; // @[Math.scala 150:24:@42896.4]
  wire [31:0] x808_sum_1_io_result; // @[Math.scala 150:24:@42896.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@42906.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@42906.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@42906.4]
  wire [31:0] RetimeWrapper_29_io_in; // @[package.scala 93:22:@42906.4]
  wire [31:0] RetimeWrapper_29_io_out; // @[package.scala 93:22:@42906.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@42915.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@42915.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@42915.4]
  wire [31:0] RetimeWrapper_30_io_in; // @[package.scala 93:22:@42915.4]
  wire [31:0] RetimeWrapper_30_io_out; // @[package.scala 93:22:@42915.4]
  wire  x567_sum_1_clock; // @[Math.scala 150:24:@42924.4]
  wire  x567_sum_1_reset; // @[Math.scala 150:24:@42924.4]
  wire [31:0] x567_sum_1_io_a; // @[Math.scala 150:24:@42924.4]
  wire [31:0] x567_sum_1_io_b; // @[Math.scala 150:24:@42924.4]
  wire  x567_sum_1_io_flow; // @[Math.scala 150:24:@42924.4]
  wire [31:0] x567_sum_1_io_result; // @[Math.scala 150:24:@42924.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@42934.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@42934.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@42934.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@42934.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@42934.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@42943.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@42943.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@42943.4]
  wire [31:0] RetimeWrapper_32_io_in; // @[package.scala 93:22:@42943.4]
  wire [31:0] RetimeWrapper_32_io_out; // @[package.scala 93:22:@42943.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@42952.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@42952.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@42952.4]
  wire [31:0] RetimeWrapper_33_io_in; // @[package.scala 93:22:@42952.4]
  wire [31:0] RetimeWrapper_33_io_out; // @[package.scala 93:22:@42952.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@42961.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@42961.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@42961.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@42961.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@42961.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@42970.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@42970.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@42970.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@42970.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@42970.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@42982.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@42982.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@42982.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@42982.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@42982.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@43003.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@43003.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@43003.4]
  wire [31:0] RetimeWrapper_37_io_in; // @[package.scala 93:22:@43003.4]
  wire [31:0] RetimeWrapper_37_io_out; // @[package.scala 93:22:@43003.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@43017.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@43017.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@43017.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@43017.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@43017.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@43032.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@43032.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@43032.4]
  wire [31:0] RetimeWrapper_39_io_in; // @[package.scala 93:22:@43032.4]
  wire [31:0] RetimeWrapper_39_io_out; // @[package.scala 93:22:@43032.4]
  wire  x573_sum_1_clock; // @[Math.scala 150:24:@43041.4]
  wire  x573_sum_1_reset; // @[Math.scala 150:24:@43041.4]
  wire [31:0] x573_sum_1_io_a; // @[Math.scala 150:24:@43041.4]
  wire [31:0] x573_sum_1_io_b; // @[Math.scala 150:24:@43041.4]
  wire  x573_sum_1_io_flow; // @[Math.scala 150:24:@43041.4]
  wire [31:0] x573_sum_1_io_result; // @[Math.scala 150:24:@43041.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@43051.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@43051.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@43051.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@43051.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@43051.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@43060.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@43060.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@43060.4]
  wire [31:0] RetimeWrapper_41_io_in; // @[package.scala 93:22:@43060.4]
  wire [31:0] RetimeWrapper_41_io_out; // @[package.scala 93:22:@43060.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@43072.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@43072.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@43072.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@43072.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@43072.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@43093.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@43093.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@43093.4]
  wire [31:0] RetimeWrapper_43_io_in; // @[package.scala 93:22:@43093.4]
  wire [31:0] RetimeWrapper_43_io_out; // @[package.scala 93:22:@43093.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@43107.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@43107.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@43107.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@43107.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@43107.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@43122.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@43122.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@43122.4]
  wire [31:0] RetimeWrapper_45_io_in; // @[package.scala 93:22:@43122.4]
  wire [31:0] RetimeWrapper_45_io_out; // @[package.scala 93:22:@43122.4]
  wire  x579_sum_1_clock; // @[Math.scala 150:24:@43131.4]
  wire  x579_sum_1_reset; // @[Math.scala 150:24:@43131.4]
  wire [31:0] x579_sum_1_io_a; // @[Math.scala 150:24:@43131.4]
  wire [31:0] x579_sum_1_io_b; // @[Math.scala 150:24:@43131.4]
  wire  x579_sum_1_io_flow; // @[Math.scala 150:24:@43131.4]
  wire [31:0] x579_sum_1_io_result; // @[Math.scala 150:24:@43131.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@43141.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@43141.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@43141.4]
  wire [31:0] RetimeWrapper_46_io_in; // @[package.scala 93:22:@43141.4]
  wire [31:0] RetimeWrapper_46_io_out; // @[package.scala 93:22:@43141.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@43150.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@43150.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@43150.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@43150.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@43150.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@43162.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@43162.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@43162.4]
  wire  RetimeWrapper_48_io_in; // @[package.scala 93:22:@43162.4]
  wire  RetimeWrapper_48_io_out; // @[package.scala 93:22:@43162.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@43183.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@43183.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@43183.4]
  wire [31:0] RetimeWrapper_49_io_in; // @[package.scala 93:22:@43183.4]
  wire [31:0] RetimeWrapper_49_io_out; // @[package.scala 93:22:@43183.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@43199.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@43199.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@43199.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@43199.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@43199.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@43214.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@43214.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@43214.4]
  wire [31:0] RetimeWrapper_51_io_in; // @[package.scala 93:22:@43214.4]
  wire [31:0] RetimeWrapper_51_io_out; // @[package.scala 93:22:@43214.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@43223.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@43223.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@43223.4]
  wire [31:0] RetimeWrapper_52_io_in; // @[package.scala 93:22:@43223.4]
  wire [31:0] RetimeWrapper_52_io_out; // @[package.scala 93:22:@43223.4]
  wire  x585_sum_1_clock; // @[Math.scala 150:24:@43232.4]
  wire  x585_sum_1_reset; // @[Math.scala 150:24:@43232.4]
  wire [31:0] x585_sum_1_io_a; // @[Math.scala 150:24:@43232.4]
  wire [31:0] x585_sum_1_io_b; // @[Math.scala 150:24:@43232.4]
  wire  x585_sum_1_io_flow; // @[Math.scala 150:24:@43232.4]
  wire [31:0] x585_sum_1_io_result; // @[Math.scala 150:24:@43232.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@43242.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@43242.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@43242.4]
  wire [31:0] RetimeWrapper_53_io_in; // @[package.scala 93:22:@43242.4]
  wire [31:0] RetimeWrapper_53_io_out; // @[package.scala 93:22:@43242.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@43251.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@43251.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@43251.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@43251.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@43251.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@43260.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@43260.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@43260.4]
  wire [31:0] RetimeWrapper_55_io_in; // @[package.scala 93:22:@43260.4]
  wire [31:0] RetimeWrapper_55_io_out; // @[package.scala 93:22:@43260.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@43272.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@43272.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@43272.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@43272.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@43272.4]
  wire  x588_rdcol_1_clock; // @[Math.scala 150:24:@43295.4]
  wire  x588_rdcol_1_reset; // @[Math.scala 150:24:@43295.4]
  wire [31:0] x588_rdcol_1_io_a; // @[Math.scala 150:24:@43295.4]
  wire [31:0] x588_rdcol_1_io_b; // @[Math.scala 150:24:@43295.4]
  wire  x588_rdcol_1_io_flow; // @[Math.scala 150:24:@43295.4]
  wire [31:0] x588_rdcol_1_io_result; // @[Math.scala 150:24:@43295.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@43310.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@43310.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@43310.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@43310.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@43310.4]
  wire  x592_1_clock; // @[Math.scala 366:24:@43327.4]
  wire  x592_1_reset; // @[Math.scala 366:24:@43327.4]
  wire [31:0] x592_1_io_a; // @[Math.scala 366:24:@43327.4]
  wire  x592_1_io_flow; // @[Math.scala 366:24:@43327.4]
  wire [31:0] x592_1_io_result; // @[Math.scala 366:24:@43327.4]
  wire  x593_div_1_clock; // @[Math.scala 327:24:@43339.4]
  wire  x593_div_1_reset; // @[Math.scala 327:24:@43339.4]
  wire [31:0] x593_div_1_io_a; // @[Math.scala 327:24:@43339.4]
  wire  x593_div_1_io_flow; // @[Math.scala 327:24:@43339.4]
  wire [31:0] x593_div_1_io_result; // @[Math.scala 327:24:@43339.4]
  wire  x594_sum_1_clock; // @[Math.scala 150:24:@43349.4]
  wire  x594_sum_1_reset; // @[Math.scala 150:24:@43349.4]
  wire [31:0] x594_sum_1_io_a; // @[Math.scala 150:24:@43349.4]
  wire [31:0] x594_sum_1_io_b; // @[Math.scala 150:24:@43349.4]
  wire  x594_sum_1_io_flow; // @[Math.scala 150:24:@43349.4]
  wire [31:0] x594_sum_1_io_result; // @[Math.scala 150:24:@43349.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@43359.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@43359.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@43359.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@43359.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@43359.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@43368.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@43368.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@43368.4]
  wire [31:0] RetimeWrapper_59_io_in; // @[package.scala 93:22:@43368.4]
  wire [31:0] RetimeWrapper_59_io_out; // @[package.scala 93:22:@43368.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@43380.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@43380.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@43380.4]
  wire  RetimeWrapper_60_io_in; // @[package.scala 93:22:@43380.4]
  wire  RetimeWrapper_60_io_out; // @[package.scala 93:22:@43380.4]
  wire  x597_rdcol_1_clock; // @[Math.scala 150:24:@43403.4]
  wire  x597_rdcol_1_reset; // @[Math.scala 150:24:@43403.4]
  wire [31:0] x597_rdcol_1_io_a; // @[Math.scala 150:24:@43403.4]
  wire [31:0] x597_rdcol_1_io_b; // @[Math.scala 150:24:@43403.4]
  wire  x597_rdcol_1_io_flow; // @[Math.scala 150:24:@43403.4]
  wire [31:0] x597_rdcol_1_io_result; // @[Math.scala 150:24:@43403.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@43418.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@43418.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@43418.4]
  wire  RetimeWrapper_61_io_in; // @[package.scala 93:22:@43418.4]
  wire  RetimeWrapper_61_io_out; // @[package.scala 93:22:@43418.4]
  wire  x601_1_clock; // @[Math.scala 366:24:@43435.4]
  wire  x601_1_reset; // @[Math.scala 366:24:@43435.4]
  wire [31:0] x601_1_io_a; // @[Math.scala 366:24:@43435.4]
  wire  x601_1_io_flow; // @[Math.scala 366:24:@43435.4]
  wire [31:0] x601_1_io_result; // @[Math.scala 366:24:@43435.4]
  wire  x602_div_1_clock; // @[Math.scala 327:24:@43447.4]
  wire  x602_div_1_reset; // @[Math.scala 327:24:@43447.4]
  wire [31:0] x602_div_1_io_a; // @[Math.scala 327:24:@43447.4]
  wire  x602_div_1_io_flow; // @[Math.scala 327:24:@43447.4]
  wire [31:0] x602_div_1_io_result; // @[Math.scala 327:24:@43447.4]
  wire  x603_sum_1_clock; // @[Math.scala 150:24:@43457.4]
  wire  x603_sum_1_reset; // @[Math.scala 150:24:@43457.4]
  wire [31:0] x603_sum_1_io_a; // @[Math.scala 150:24:@43457.4]
  wire [31:0] x603_sum_1_io_b; // @[Math.scala 150:24:@43457.4]
  wire  x603_sum_1_io_flow; // @[Math.scala 150:24:@43457.4]
  wire [31:0] x603_sum_1_io_result; // @[Math.scala 150:24:@43457.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@43467.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@43467.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@43467.4]
  wire [31:0] RetimeWrapper_62_io_in; // @[package.scala 93:22:@43467.4]
  wire [31:0] RetimeWrapper_62_io_out; // @[package.scala 93:22:@43467.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@43476.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@43476.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@43476.4]
  wire  RetimeWrapper_63_io_in; // @[package.scala 93:22:@43476.4]
  wire  RetimeWrapper_63_io_out; // @[package.scala 93:22:@43476.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@43488.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@43488.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@43488.4]
  wire  RetimeWrapper_64_io_in; // @[package.scala 93:22:@43488.4]
  wire  RetimeWrapper_64_io_out; // @[package.scala 93:22:@43488.4]
  wire  x606_rdrow_1_clock; // @[Math.scala 191:24:@43511.4]
  wire  x606_rdrow_1_reset; // @[Math.scala 191:24:@43511.4]
  wire [31:0] x606_rdrow_1_io_a; // @[Math.scala 191:24:@43511.4]
  wire [31:0] x606_rdrow_1_io_b; // @[Math.scala 191:24:@43511.4]
  wire  x606_rdrow_1_io_flow; // @[Math.scala 191:24:@43511.4]
  wire [31:0] x606_rdrow_1_io_result; // @[Math.scala 191:24:@43511.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@43528.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@43528.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@43528.4]
  wire [31:0] RetimeWrapper_65_io_in; // @[package.scala 93:22:@43528.4]
  wire [31:0] RetimeWrapper_65_io_out; // @[package.scala 93:22:@43528.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@43546.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@43546.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@43546.4]
  wire  RetimeWrapper_66_io_in; // @[package.scala 93:22:@43546.4]
  wire  RetimeWrapper_66_io_out; // @[package.scala 93:22:@43546.4]
  wire  x813_sum_1_clock; // @[Math.scala 150:24:@43591.4]
  wire  x813_sum_1_reset; // @[Math.scala 150:24:@43591.4]
  wire [31:0] x813_sum_1_io_a; // @[Math.scala 150:24:@43591.4]
  wire [31:0] x813_sum_1_io_b; // @[Math.scala 150:24:@43591.4]
  wire  x813_sum_1_io_flow; // @[Math.scala 150:24:@43591.4]
  wire [31:0] x813_sum_1_io_result; // @[Math.scala 150:24:@43591.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@43601.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@43601.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@43601.4]
  wire [31:0] RetimeWrapper_67_io_in; // @[package.scala 93:22:@43601.4]
  wire [31:0] RetimeWrapper_67_io_out; // @[package.scala 93:22:@43601.4]
  wire  x614_sum_1_clock; // @[Math.scala 150:24:@43610.4]
  wire  x614_sum_1_reset; // @[Math.scala 150:24:@43610.4]
  wire [31:0] x614_sum_1_io_a; // @[Math.scala 150:24:@43610.4]
  wire [31:0] x614_sum_1_io_b; // @[Math.scala 150:24:@43610.4]
  wire  x614_sum_1_io_flow; // @[Math.scala 150:24:@43610.4]
  wire [31:0] x614_sum_1_io_result; // @[Math.scala 150:24:@43610.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@43620.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@43620.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@43620.4]
  wire [31:0] RetimeWrapper_68_io_in; // @[package.scala 93:22:@43620.4]
  wire [31:0] RetimeWrapper_68_io_out; // @[package.scala 93:22:@43620.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@43629.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@43629.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@43629.4]
  wire  RetimeWrapper_69_io_in; // @[package.scala 93:22:@43629.4]
  wire  RetimeWrapper_69_io_out; // @[package.scala 93:22:@43629.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@43641.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@43641.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@43641.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@43641.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@43641.4]
  wire  x619_sum_1_clock; // @[Math.scala 150:24:@43670.4]
  wire  x619_sum_1_reset; // @[Math.scala 150:24:@43670.4]
  wire [31:0] x619_sum_1_io_a; // @[Math.scala 150:24:@43670.4]
  wire [31:0] x619_sum_1_io_b; // @[Math.scala 150:24:@43670.4]
  wire  x619_sum_1_io_flow; // @[Math.scala 150:24:@43670.4]
  wire [31:0] x619_sum_1_io_result; // @[Math.scala 150:24:@43670.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@43680.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@43680.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@43680.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@43680.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@43680.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@43692.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@43692.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@43692.4]
  wire  RetimeWrapper_72_io_in; // @[package.scala 93:22:@43692.4]
  wire  RetimeWrapper_72_io_out; // @[package.scala 93:22:@43692.4]
  wire  x624_sum_1_clock; // @[Math.scala 150:24:@43719.4]
  wire  x624_sum_1_reset; // @[Math.scala 150:24:@43719.4]
  wire [31:0] x624_sum_1_io_a; // @[Math.scala 150:24:@43719.4]
  wire [31:0] x624_sum_1_io_b; // @[Math.scala 150:24:@43719.4]
  wire  x624_sum_1_io_flow; // @[Math.scala 150:24:@43719.4]
  wire [31:0] x624_sum_1_io_result; // @[Math.scala 150:24:@43719.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@43729.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@43729.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@43729.4]
  wire  RetimeWrapper_73_io_in; // @[package.scala 93:22:@43729.4]
  wire  RetimeWrapper_73_io_out; // @[package.scala 93:22:@43729.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@43741.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@43741.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@43741.4]
  wire  RetimeWrapper_74_io_in; // @[package.scala 93:22:@43741.4]
  wire  RetimeWrapper_74_io_out; // @[package.scala 93:22:@43741.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@43762.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@43762.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@43762.4]
  wire  RetimeWrapper_75_io_in; // @[package.scala 93:22:@43762.4]
  wire  RetimeWrapper_75_io_out; // @[package.scala 93:22:@43762.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@43777.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@43777.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@43777.4]
  wire [31:0] RetimeWrapper_76_io_in; // @[package.scala 93:22:@43777.4]
  wire [31:0] RetimeWrapper_76_io_out; // @[package.scala 93:22:@43777.4]
  wire  x629_sum_1_clock; // @[Math.scala 150:24:@43786.4]
  wire  x629_sum_1_reset; // @[Math.scala 150:24:@43786.4]
  wire [31:0] x629_sum_1_io_a; // @[Math.scala 150:24:@43786.4]
  wire [31:0] x629_sum_1_io_b; // @[Math.scala 150:24:@43786.4]
  wire  x629_sum_1_io_flow; // @[Math.scala 150:24:@43786.4]
  wire [31:0] x629_sum_1_io_result; // @[Math.scala 150:24:@43786.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@43796.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@43796.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@43796.4]
  wire [31:0] RetimeWrapper_77_io_in; // @[package.scala 93:22:@43796.4]
  wire [31:0] RetimeWrapper_77_io_out; // @[package.scala 93:22:@43796.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@43805.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@43805.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@43805.4]
  wire  RetimeWrapper_78_io_in; // @[package.scala 93:22:@43805.4]
  wire  RetimeWrapper_78_io_out; // @[package.scala 93:22:@43805.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@43817.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@43817.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@43817.4]
  wire  RetimeWrapper_79_io_in; // @[package.scala 93:22:@43817.4]
  wire  RetimeWrapper_79_io_out; // @[package.scala 93:22:@43817.4]
  wire  x634_sum_1_clock; // @[Math.scala 150:24:@43844.4]
  wire  x634_sum_1_reset; // @[Math.scala 150:24:@43844.4]
  wire [31:0] x634_sum_1_io_a; // @[Math.scala 150:24:@43844.4]
  wire [31:0] x634_sum_1_io_b; // @[Math.scala 150:24:@43844.4]
  wire  x634_sum_1_io_flow; // @[Math.scala 150:24:@43844.4]
  wire [31:0] x634_sum_1_io_result; // @[Math.scala 150:24:@43844.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@43854.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@43854.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@43854.4]
  wire  RetimeWrapper_80_io_in; // @[package.scala 93:22:@43854.4]
  wire  RetimeWrapper_80_io_out; // @[package.scala 93:22:@43854.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@43866.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@43866.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@43866.4]
  wire  RetimeWrapper_81_io_in; // @[package.scala 93:22:@43866.4]
  wire  RetimeWrapper_81_io_out; // @[package.scala 93:22:@43866.4]
  wire  x639_sum_1_clock; // @[Math.scala 150:24:@43893.4]
  wire  x639_sum_1_reset; // @[Math.scala 150:24:@43893.4]
  wire [31:0] x639_sum_1_io_a; // @[Math.scala 150:24:@43893.4]
  wire [31:0] x639_sum_1_io_b; // @[Math.scala 150:24:@43893.4]
  wire  x639_sum_1_io_flow; // @[Math.scala 150:24:@43893.4]
  wire [31:0] x639_sum_1_io_result; // @[Math.scala 150:24:@43893.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@43903.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@43903.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@43903.4]
  wire  RetimeWrapper_82_io_in; // @[package.scala 93:22:@43903.4]
  wire  RetimeWrapper_82_io_out; // @[package.scala 93:22:@43903.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@43915.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@43915.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@43915.4]
  wire  RetimeWrapper_83_io_in; // @[package.scala 93:22:@43915.4]
  wire  RetimeWrapper_83_io_out; // @[package.scala 93:22:@43915.4]
  wire  x642_rdrow_1_clock; // @[Math.scala 191:24:@43938.4]
  wire  x642_rdrow_1_reset; // @[Math.scala 191:24:@43938.4]
  wire [31:0] x642_rdrow_1_io_a; // @[Math.scala 191:24:@43938.4]
  wire [31:0] x642_rdrow_1_io_b; // @[Math.scala 191:24:@43938.4]
  wire  x642_rdrow_1_io_flow; // @[Math.scala 191:24:@43938.4]
  wire [31:0] x642_rdrow_1_io_result; // @[Math.scala 191:24:@43938.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@43955.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@43955.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@43955.4]
  wire [31:0] RetimeWrapper_84_io_in; // @[package.scala 93:22:@43955.4]
  wire [31:0] RetimeWrapper_84_io_out; // @[package.scala 93:22:@43955.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@43973.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@43973.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@43973.4]
  wire  RetimeWrapper_85_io_in; // @[package.scala 93:22:@43973.4]
  wire  RetimeWrapper_85_io_out; // @[package.scala 93:22:@43973.4]
  wire  x818_sum_1_clock; // @[Math.scala 150:24:@44018.4]
  wire  x818_sum_1_reset; // @[Math.scala 150:24:@44018.4]
  wire [31:0] x818_sum_1_io_a; // @[Math.scala 150:24:@44018.4]
  wire [31:0] x818_sum_1_io_b; // @[Math.scala 150:24:@44018.4]
  wire  x818_sum_1_io_flow; // @[Math.scala 150:24:@44018.4]
  wire [31:0] x818_sum_1_io_result; // @[Math.scala 150:24:@44018.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@44028.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@44028.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@44028.4]
  wire [31:0] RetimeWrapper_86_io_in; // @[package.scala 93:22:@44028.4]
  wire [31:0] RetimeWrapper_86_io_out; // @[package.scala 93:22:@44028.4]
  wire  x650_sum_1_clock; // @[Math.scala 150:24:@44037.4]
  wire  x650_sum_1_reset; // @[Math.scala 150:24:@44037.4]
  wire [31:0] x650_sum_1_io_a; // @[Math.scala 150:24:@44037.4]
  wire [31:0] x650_sum_1_io_b; // @[Math.scala 150:24:@44037.4]
  wire  x650_sum_1_io_flow; // @[Math.scala 150:24:@44037.4]
  wire [31:0] x650_sum_1_io_result; // @[Math.scala 150:24:@44037.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@44047.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@44047.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@44047.4]
  wire  RetimeWrapper_87_io_in; // @[package.scala 93:22:@44047.4]
  wire  RetimeWrapper_87_io_out; // @[package.scala 93:22:@44047.4]
  wire  RetimeWrapper_88_clock; // @[package.scala 93:22:@44056.4]
  wire  RetimeWrapper_88_reset; // @[package.scala 93:22:@44056.4]
  wire  RetimeWrapper_88_io_flow; // @[package.scala 93:22:@44056.4]
  wire [31:0] RetimeWrapper_88_io_in; // @[package.scala 93:22:@44056.4]
  wire [31:0] RetimeWrapper_88_io_out; // @[package.scala 93:22:@44056.4]
  wire  RetimeWrapper_89_clock; // @[package.scala 93:22:@44068.4]
  wire  RetimeWrapper_89_reset; // @[package.scala 93:22:@44068.4]
  wire  RetimeWrapper_89_io_flow; // @[package.scala 93:22:@44068.4]
  wire  RetimeWrapper_89_io_in; // @[package.scala 93:22:@44068.4]
  wire  RetimeWrapper_89_io_out; // @[package.scala 93:22:@44068.4]
  wire  x655_sum_1_clock; // @[Math.scala 150:24:@44097.4]
  wire  x655_sum_1_reset; // @[Math.scala 150:24:@44097.4]
  wire [31:0] x655_sum_1_io_a; // @[Math.scala 150:24:@44097.4]
  wire [31:0] x655_sum_1_io_b; // @[Math.scala 150:24:@44097.4]
  wire  x655_sum_1_io_flow; // @[Math.scala 150:24:@44097.4]
  wire [31:0] x655_sum_1_io_result; // @[Math.scala 150:24:@44097.4]
  wire  RetimeWrapper_90_clock; // @[package.scala 93:22:@44107.4]
  wire  RetimeWrapper_90_reset; // @[package.scala 93:22:@44107.4]
  wire  RetimeWrapper_90_io_flow; // @[package.scala 93:22:@44107.4]
  wire  RetimeWrapper_90_io_in; // @[package.scala 93:22:@44107.4]
  wire  RetimeWrapper_90_io_out; // @[package.scala 93:22:@44107.4]
  wire  RetimeWrapper_91_clock; // @[package.scala 93:22:@44119.4]
  wire  RetimeWrapper_91_reset; // @[package.scala 93:22:@44119.4]
  wire  RetimeWrapper_91_io_flow; // @[package.scala 93:22:@44119.4]
  wire  RetimeWrapper_91_io_in; // @[package.scala 93:22:@44119.4]
  wire  RetimeWrapper_91_io_out; // @[package.scala 93:22:@44119.4]
  wire  x660_sum_1_clock; // @[Math.scala 150:24:@44146.4]
  wire  x660_sum_1_reset; // @[Math.scala 150:24:@44146.4]
  wire [31:0] x660_sum_1_io_a; // @[Math.scala 150:24:@44146.4]
  wire [31:0] x660_sum_1_io_b; // @[Math.scala 150:24:@44146.4]
  wire  x660_sum_1_io_flow; // @[Math.scala 150:24:@44146.4]
  wire [31:0] x660_sum_1_io_result; // @[Math.scala 150:24:@44146.4]
  wire  RetimeWrapper_92_clock; // @[package.scala 93:22:@44156.4]
  wire  RetimeWrapper_92_reset; // @[package.scala 93:22:@44156.4]
  wire  RetimeWrapper_92_io_flow; // @[package.scala 93:22:@44156.4]
  wire  RetimeWrapper_92_io_in; // @[package.scala 93:22:@44156.4]
  wire  RetimeWrapper_92_io_out; // @[package.scala 93:22:@44156.4]
  wire  RetimeWrapper_93_clock; // @[package.scala 93:22:@44168.4]
  wire  RetimeWrapper_93_reset; // @[package.scala 93:22:@44168.4]
  wire  RetimeWrapper_93_io_flow; // @[package.scala 93:22:@44168.4]
  wire  RetimeWrapper_93_io_in; // @[package.scala 93:22:@44168.4]
  wire  RetimeWrapper_93_io_out; // @[package.scala 93:22:@44168.4]
  wire  RetimeWrapper_94_clock; // @[package.scala 93:22:@44195.4]
  wire  RetimeWrapper_94_reset; // @[package.scala 93:22:@44195.4]
  wire  RetimeWrapper_94_io_flow; // @[package.scala 93:22:@44195.4]
  wire [31:0] RetimeWrapper_94_io_in; // @[package.scala 93:22:@44195.4]
  wire [31:0] RetimeWrapper_94_io_out; // @[package.scala 93:22:@44195.4]
  wire  x665_sum_1_clock; // @[Math.scala 150:24:@44204.4]
  wire  x665_sum_1_reset; // @[Math.scala 150:24:@44204.4]
  wire [31:0] x665_sum_1_io_a; // @[Math.scala 150:24:@44204.4]
  wire [31:0] x665_sum_1_io_b; // @[Math.scala 150:24:@44204.4]
  wire  x665_sum_1_io_flow; // @[Math.scala 150:24:@44204.4]
  wire [31:0] x665_sum_1_io_result; // @[Math.scala 150:24:@44204.4]
  wire  RetimeWrapper_95_clock; // @[package.scala 93:22:@44214.4]
  wire  RetimeWrapper_95_reset; // @[package.scala 93:22:@44214.4]
  wire  RetimeWrapper_95_io_flow; // @[package.scala 93:22:@44214.4]
  wire [31:0] RetimeWrapper_95_io_in; // @[package.scala 93:22:@44214.4]
  wire [31:0] RetimeWrapper_95_io_out; // @[package.scala 93:22:@44214.4]
  wire  RetimeWrapper_96_clock; // @[package.scala 93:22:@44223.4]
  wire  RetimeWrapper_96_reset; // @[package.scala 93:22:@44223.4]
  wire  RetimeWrapper_96_io_flow; // @[package.scala 93:22:@44223.4]
  wire  RetimeWrapper_96_io_in; // @[package.scala 93:22:@44223.4]
  wire  RetimeWrapper_96_io_out; // @[package.scala 93:22:@44223.4]
  wire  RetimeWrapper_97_clock; // @[package.scala 93:22:@44235.4]
  wire  RetimeWrapper_97_reset; // @[package.scala 93:22:@44235.4]
  wire  RetimeWrapper_97_io_flow; // @[package.scala 93:22:@44235.4]
  wire  RetimeWrapper_97_io_in; // @[package.scala 93:22:@44235.4]
  wire  RetimeWrapper_97_io_out; // @[package.scala 93:22:@44235.4]
  wire  x670_sum_1_clock; // @[Math.scala 150:24:@44262.4]
  wire  x670_sum_1_reset; // @[Math.scala 150:24:@44262.4]
  wire [31:0] x670_sum_1_io_a; // @[Math.scala 150:24:@44262.4]
  wire [31:0] x670_sum_1_io_b; // @[Math.scala 150:24:@44262.4]
  wire  x670_sum_1_io_flow; // @[Math.scala 150:24:@44262.4]
  wire [31:0] x670_sum_1_io_result; // @[Math.scala 150:24:@44262.4]
  wire  RetimeWrapper_98_clock; // @[package.scala 93:22:@44272.4]
  wire  RetimeWrapper_98_reset; // @[package.scala 93:22:@44272.4]
  wire  RetimeWrapper_98_io_flow; // @[package.scala 93:22:@44272.4]
  wire  RetimeWrapper_98_io_in; // @[package.scala 93:22:@44272.4]
  wire  RetimeWrapper_98_io_out; // @[package.scala 93:22:@44272.4]
  wire  RetimeWrapper_99_clock; // @[package.scala 93:22:@44284.4]
  wire  RetimeWrapper_99_reset; // @[package.scala 93:22:@44284.4]
  wire  RetimeWrapper_99_io_flow; // @[package.scala 93:22:@44284.4]
  wire  RetimeWrapper_99_io_in; // @[package.scala 93:22:@44284.4]
  wire  RetimeWrapper_99_io_out; // @[package.scala 93:22:@44284.4]
  wire  x675_sum_1_clock; // @[Math.scala 150:24:@44311.4]
  wire  x675_sum_1_reset; // @[Math.scala 150:24:@44311.4]
  wire [31:0] x675_sum_1_io_a; // @[Math.scala 150:24:@44311.4]
  wire [31:0] x675_sum_1_io_b; // @[Math.scala 150:24:@44311.4]
  wire  x675_sum_1_io_flow; // @[Math.scala 150:24:@44311.4]
  wire [31:0] x675_sum_1_io_result; // @[Math.scala 150:24:@44311.4]
  wire  RetimeWrapper_100_clock; // @[package.scala 93:22:@44321.4]
  wire  RetimeWrapper_100_reset; // @[package.scala 93:22:@44321.4]
  wire  RetimeWrapper_100_io_flow; // @[package.scala 93:22:@44321.4]
  wire  RetimeWrapper_100_io_in; // @[package.scala 93:22:@44321.4]
  wire  RetimeWrapper_100_io_out; // @[package.scala 93:22:@44321.4]
  wire  RetimeWrapper_101_clock; // @[package.scala 93:22:@44333.4]
  wire  RetimeWrapper_101_reset; // @[package.scala 93:22:@44333.4]
  wire  RetimeWrapper_101_io_flow; // @[package.scala 93:22:@44333.4]
  wire  RetimeWrapper_101_io_in; // @[package.scala 93:22:@44333.4]
  wire  RetimeWrapper_101_io_out; // @[package.scala 93:22:@44333.4]
  wire  RetimeWrapper_102_clock; // @[package.scala 93:22:@44356.4]
  wire  RetimeWrapper_102_reset; // @[package.scala 93:22:@44356.4]
  wire  RetimeWrapper_102_io_flow; // @[package.scala 93:22:@44356.4]
  wire [8:0] RetimeWrapper_102_io_in; // @[package.scala 93:22:@44356.4]
  wire [8:0] RetimeWrapper_102_io_out; // @[package.scala 93:22:@44356.4]
  wire  RetimeWrapper_103_clock; // @[package.scala 93:22:@44368.4]
  wire  RetimeWrapper_103_reset; // @[package.scala 93:22:@44368.4]
  wire  RetimeWrapper_103_io_flow; // @[package.scala 93:22:@44368.4]
  wire [8:0] RetimeWrapper_103_io_in; // @[package.scala 93:22:@44368.4]
  wire [8:0] RetimeWrapper_103_io_out; // @[package.scala 93:22:@44368.4]
  wire  RetimeWrapper_104_clock; // @[package.scala 93:22:@44380.4]
  wire  RetimeWrapper_104_reset; // @[package.scala 93:22:@44380.4]
  wire  RetimeWrapper_104_io_flow; // @[package.scala 93:22:@44380.4]
  wire [9:0] RetimeWrapper_104_io_in; // @[package.scala 93:22:@44380.4]
  wire [9:0] RetimeWrapper_104_io_out; // @[package.scala 93:22:@44380.4]
  wire  RetimeWrapper_105_clock; // @[package.scala 93:22:@44392.4]
  wire  RetimeWrapper_105_reset; // @[package.scala 93:22:@44392.4]
  wire  RetimeWrapper_105_io_flow; // @[package.scala 93:22:@44392.4]
  wire [8:0] RetimeWrapper_105_io_in; // @[package.scala 93:22:@44392.4]
  wire [8:0] RetimeWrapper_105_io_out; // @[package.scala 93:22:@44392.4]
  wire  RetimeWrapper_106_clock; // @[package.scala 93:22:@44404.4]
  wire  RetimeWrapper_106_reset; // @[package.scala 93:22:@44404.4]
  wire  RetimeWrapper_106_io_flow; // @[package.scala 93:22:@44404.4]
  wire [8:0] RetimeWrapper_106_io_in; // @[package.scala 93:22:@44404.4]
  wire [8:0] RetimeWrapper_106_io_out; // @[package.scala 93:22:@44404.4]
  wire  RetimeWrapper_107_clock; // @[package.scala 93:22:@44414.4]
  wire  RetimeWrapper_107_reset; // @[package.scala 93:22:@44414.4]
  wire  RetimeWrapper_107_io_flow; // @[package.scala 93:22:@44414.4]
  wire [7:0] RetimeWrapper_107_io_in; // @[package.scala 93:22:@44414.4]
  wire [7:0] RetimeWrapper_107_io_out; // @[package.scala 93:22:@44414.4]
  wire [7:0] x683_x15_1_io_a; // @[Math.scala 150:24:@44423.4]
  wire [7:0] x683_x15_1_io_b; // @[Math.scala 150:24:@44423.4]
  wire [7:0] x683_x15_1_io_result; // @[Math.scala 150:24:@44423.4]
  wire  RetimeWrapper_108_clock; // @[package.scala 93:22:@44433.4]
  wire  RetimeWrapper_108_reset; // @[package.scala 93:22:@44433.4]
  wire  RetimeWrapper_108_io_flow; // @[package.scala 93:22:@44433.4]
  wire [7:0] RetimeWrapper_108_io_in; // @[package.scala 93:22:@44433.4]
  wire [7:0] RetimeWrapper_108_io_out; // @[package.scala 93:22:@44433.4]
  wire [7:0] x684_x16_1_io_a; // @[Math.scala 150:24:@44442.4]
  wire [7:0] x684_x16_1_io_b; // @[Math.scala 150:24:@44442.4]
  wire [7:0] x684_x16_1_io_result; // @[Math.scala 150:24:@44442.4]
  wire [7:0] x685_x15_1_io_a; // @[Math.scala 150:24:@44452.4]
  wire [7:0] x685_x15_1_io_b; // @[Math.scala 150:24:@44452.4]
  wire [7:0] x685_x15_1_io_result; // @[Math.scala 150:24:@44452.4]
  wire  RetimeWrapper_109_clock; // @[package.scala 93:22:@44462.4]
  wire  RetimeWrapper_109_reset; // @[package.scala 93:22:@44462.4]
  wire  RetimeWrapper_109_io_flow; // @[package.scala 93:22:@44462.4]
  wire [7:0] RetimeWrapper_109_io_in; // @[package.scala 93:22:@44462.4]
  wire [7:0] RetimeWrapper_109_io_out; // @[package.scala 93:22:@44462.4]
  wire [7:0] x686_x16_1_io_a; // @[Math.scala 150:24:@44471.4]
  wire [7:0] x686_x16_1_io_b; // @[Math.scala 150:24:@44471.4]
  wire [7:0] x686_x16_1_io_result; // @[Math.scala 150:24:@44471.4]
  wire [7:0] x687_x15_1_io_a; // @[Math.scala 150:24:@44481.4]
  wire [7:0] x687_x15_1_io_b; // @[Math.scala 150:24:@44481.4]
  wire [7:0] x687_x15_1_io_result; // @[Math.scala 150:24:@44481.4]
  wire [7:0] x688_x16_1_io_a; // @[Math.scala 150:24:@44491.4]
  wire [7:0] x688_x16_1_io_b; // @[Math.scala 150:24:@44491.4]
  wire [7:0] x688_x16_1_io_result; // @[Math.scala 150:24:@44491.4]
  wire [7:0] x689_x15_1_io_a; // @[Math.scala 150:24:@44503.4]
  wire [7:0] x689_x15_1_io_b; // @[Math.scala 150:24:@44503.4]
  wire [7:0] x689_x15_1_io_result; // @[Math.scala 150:24:@44503.4]
  wire  RetimeWrapper_110_clock; // @[package.scala 93:22:@44513.4]
  wire  RetimeWrapper_110_reset; // @[package.scala 93:22:@44513.4]
  wire  RetimeWrapper_110_io_flow; // @[package.scala 93:22:@44513.4]
  wire [7:0] RetimeWrapper_110_io_in; // @[package.scala 93:22:@44513.4]
  wire [7:0] RetimeWrapper_110_io_out; // @[package.scala 93:22:@44513.4]
  wire  x690_sum_1_clock; // @[Math.scala 150:24:@44522.4]
  wire  x690_sum_1_reset; // @[Math.scala 150:24:@44522.4]
  wire [7:0] x690_sum_1_io_a; // @[Math.scala 150:24:@44522.4]
  wire [7:0] x690_sum_1_io_b; // @[Math.scala 150:24:@44522.4]
  wire  x690_sum_1_io_flow; // @[Math.scala 150:24:@44522.4]
  wire [7:0] x690_sum_1_io_result; // @[Math.scala 150:24:@44522.4]
  wire  RetimeWrapper_111_clock; // @[package.scala 93:22:@44541.4]
  wire  RetimeWrapper_111_reset; // @[package.scala 93:22:@44541.4]
  wire  RetimeWrapper_111_io_flow; // @[package.scala 93:22:@44541.4]
  wire [8:0] RetimeWrapper_111_io_in; // @[package.scala 93:22:@44541.4]
  wire [8:0] RetimeWrapper_111_io_out; // @[package.scala 93:22:@44541.4]
  wire  RetimeWrapper_112_clock; // @[package.scala 93:22:@44553.4]
  wire  RetimeWrapper_112_reset; // @[package.scala 93:22:@44553.4]
  wire  RetimeWrapper_112_io_flow; // @[package.scala 93:22:@44553.4]
  wire [8:0] RetimeWrapper_112_io_in; // @[package.scala 93:22:@44553.4]
  wire [8:0] RetimeWrapper_112_io_out; // @[package.scala 93:22:@44553.4]
  wire  RetimeWrapper_113_clock; // @[package.scala 93:22:@44565.4]
  wire  RetimeWrapper_113_reset; // @[package.scala 93:22:@44565.4]
  wire  RetimeWrapper_113_io_flow; // @[package.scala 93:22:@44565.4]
  wire [9:0] RetimeWrapper_113_io_in; // @[package.scala 93:22:@44565.4]
  wire [9:0] RetimeWrapper_113_io_out; // @[package.scala 93:22:@44565.4]
  wire  RetimeWrapper_114_clock; // @[package.scala 93:22:@44577.4]
  wire  RetimeWrapper_114_reset; // @[package.scala 93:22:@44577.4]
  wire  RetimeWrapper_114_io_flow; // @[package.scala 93:22:@44577.4]
  wire [8:0] RetimeWrapper_114_io_in; // @[package.scala 93:22:@44577.4]
  wire [8:0] RetimeWrapper_114_io_out; // @[package.scala 93:22:@44577.4]
  wire  RetimeWrapper_115_clock; // @[package.scala 93:22:@44589.4]
  wire  RetimeWrapper_115_reset; // @[package.scala 93:22:@44589.4]
  wire  RetimeWrapper_115_io_flow; // @[package.scala 93:22:@44589.4]
  wire [8:0] RetimeWrapper_115_io_in; // @[package.scala 93:22:@44589.4]
  wire [8:0] RetimeWrapper_115_io_out; // @[package.scala 93:22:@44589.4]
  wire  RetimeWrapper_116_clock; // @[package.scala 93:22:@44599.4]
  wire  RetimeWrapper_116_reset; // @[package.scala 93:22:@44599.4]
  wire  RetimeWrapper_116_io_flow; // @[package.scala 93:22:@44599.4]
  wire [7:0] RetimeWrapper_116_io_in; // @[package.scala 93:22:@44599.4]
  wire [7:0] RetimeWrapper_116_io_out; // @[package.scala 93:22:@44599.4]
  wire [7:0] x697_x15_1_io_a; // @[Math.scala 150:24:@44608.4]
  wire [7:0] x697_x15_1_io_b; // @[Math.scala 150:24:@44608.4]
  wire [7:0] x697_x15_1_io_result; // @[Math.scala 150:24:@44608.4]
  wire  RetimeWrapper_117_clock; // @[package.scala 93:22:@44618.4]
  wire  RetimeWrapper_117_reset; // @[package.scala 93:22:@44618.4]
  wire  RetimeWrapper_117_io_flow; // @[package.scala 93:22:@44618.4]
  wire [7:0] RetimeWrapper_117_io_in; // @[package.scala 93:22:@44618.4]
  wire [7:0] RetimeWrapper_117_io_out; // @[package.scala 93:22:@44618.4]
  wire [7:0] x698_x16_1_io_a; // @[Math.scala 150:24:@44627.4]
  wire [7:0] x698_x16_1_io_b; // @[Math.scala 150:24:@44627.4]
  wire [7:0] x698_x16_1_io_result; // @[Math.scala 150:24:@44627.4]
  wire [7:0] x699_x15_1_io_a; // @[Math.scala 150:24:@44637.4]
  wire [7:0] x699_x15_1_io_b; // @[Math.scala 150:24:@44637.4]
  wire [7:0] x699_x15_1_io_result; // @[Math.scala 150:24:@44637.4]
  wire  RetimeWrapper_118_clock; // @[package.scala 93:22:@44647.4]
  wire  RetimeWrapper_118_reset; // @[package.scala 93:22:@44647.4]
  wire  RetimeWrapper_118_io_flow; // @[package.scala 93:22:@44647.4]
  wire [7:0] RetimeWrapper_118_io_in; // @[package.scala 93:22:@44647.4]
  wire [7:0] RetimeWrapper_118_io_out; // @[package.scala 93:22:@44647.4]
  wire [7:0] x700_x16_1_io_a; // @[Math.scala 150:24:@44656.4]
  wire [7:0] x700_x16_1_io_b; // @[Math.scala 150:24:@44656.4]
  wire [7:0] x700_x16_1_io_result; // @[Math.scala 150:24:@44656.4]
  wire [7:0] x701_x15_1_io_a; // @[Math.scala 150:24:@44666.4]
  wire [7:0] x701_x15_1_io_b; // @[Math.scala 150:24:@44666.4]
  wire [7:0] x701_x15_1_io_result; // @[Math.scala 150:24:@44666.4]
  wire [7:0] x702_x16_1_io_a; // @[Math.scala 150:24:@44676.4]
  wire [7:0] x702_x16_1_io_b; // @[Math.scala 150:24:@44676.4]
  wire [7:0] x702_x16_1_io_result; // @[Math.scala 150:24:@44676.4]
  wire [7:0] x703_x15_1_io_a; // @[Math.scala 150:24:@44686.4]
  wire [7:0] x703_x15_1_io_b; // @[Math.scala 150:24:@44686.4]
  wire [7:0] x703_x15_1_io_result; // @[Math.scala 150:24:@44686.4]
  wire  RetimeWrapper_119_clock; // @[package.scala 93:22:@44696.4]
  wire  RetimeWrapper_119_reset; // @[package.scala 93:22:@44696.4]
  wire  RetimeWrapper_119_io_flow; // @[package.scala 93:22:@44696.4]
  wire [7:0] RetimeWrapper_119_io_in; // @[package.scala 93:22:@44696.4]
  wire [7:0] RetimeWrapper_119_io_out; // @[package.scala 93:22:@44696.4]
  wire  x704_sum_1_clock; // @[Math.scala 150:24:@44705.4]
  wire  x704_sum_1_reset; // @[Math.scala 150:24:@44705.4]
  wire [7:0] x704_sum_1_io_a; // @[Math.scala 150:24:@44705.4]
  wire [7:0] x704_sum_1_io_b; // @[Math.scala 150:24:@44705.4]
  wire  x704_sum_1_io_flow; // @[Math.scala 150:24:@44705.4]
  wire [7:0] x704_sum_1_io_result; // @[Math.scala 150:24:@44705.4]
  wire  RetimeWrapper_120_clock; // @[package.scala 93:22:@44724.4]
  wire  RetimeWrapper_120_reset; // @[package.scala 93:22:@44724.4]
  wire  RetimeWrapper_120_io_flow; // @[package.scala 93:22:@44724.4]
  wire [8:0] RetimeWrapper_120_io_in; // @[package.scala 93:22:@44724.4]
  wire [8:0] RetimeWrapper_120_io_out; // @[package.scala 93:22:@44724.4]
  wire  RetimeWrapper_121_clock; // @[package.scala 93:22:@44736.4]
  wire  RetimeWrapper_121_reset; // @[package.scala 93:22:@44736.4]
  wire  RetimeWrapper_121_io_flow; // @[package.scala 93:22:@44736.4]
  wire [9:0] RetimeWrapper_121_io_in; // @[package.scala 93:22:@44736.4]
  wire [9:0] RetimeWrapper_121_io_out; // @[package.scala 93:22:@44736.4]
  wire  RetimeWrapper_122_clock; // @[package.scala 93:22:@44748.4]
  wire  RetimeWrapper_122_reset; // @[package.scala 93:22:@44748.4]
  wire  RetimeWrapper_122_io_flow; // @[package.scala 93:22:@44748.4]
  wire [8:0] RetimeWrapper_122_io_in; // @[package.scala 93:22:@44748.4]
  wire [8:0] RetimeWrapper_122_io_out; // @[package.scala 93:22:@44748.4]
  wire  RetimeWrapper_123_clock; // @[package.scala 93:22:@44760.4]
  wire  RetimeWrapper_123_reset; // @[package.scala 93:22:@44760.4]
  wire  RetimeWrapper_123_io_flow; // @[package.scala 93:22:@44760.4]
  wire [8:0] RetimeWrapper_123_io_in; // @[package.scala 93:22:@44760.4]
  wire [8:0] RetimeWrapper_123_io_out; // @[package.scala 93:22:@44760.4]
  wire [7:0] x710_x15_1_io_a; // @[Math.scala 150:24:@44770.4]
  wire [7:0] x710_x15_1_io_b; // @[Math.scala 150:24:@44770.4]
  wire [7:0] x710_x15_1_io_result; // @[Math.scala 150:24:@44770.4]
  wire  RetimeWrapper_124_clock; // @[package.scala 93:22:@44780.4]
  wire  RetimeWrapper_124_reset; // @[package.scala 93:22:@44780.4]
  wire  RetimeWrapper_124_io_flow; // @[package.scala 93:22:@44780.4]
  wire [7:0] RetimeWrapper_124_io_in; // @[package.scala 93:22:@44780.4]
  wire [7:0] RetimeWrapper_124_io_out; // @[package.scala 93:22:@44780.4]
  wire [7:0] x711_x16_1_io_a; // @[Math.scala 150:24:@44789.4]
  wire [7:0] x711_x16_1_io_b; // @[Math.scala 150:24:@44789.4]
  wire [7:0] x711_x16_1_io_result; // @[Math.scala 150:24:@44789.4]
  wire [7:0] x712_x15_1_io_a; // @[Math.scala 150:24:@44799.4]
  wire [7:0] x712_x15_1_io_b; // @[Math.scala 150:24:@44799.4]
  wire [7:0] x712_x15_1_io_result; // @[Math.scala 150:24:@44799.4]
  wire [7:0] x713_x16_1_io_a; // @[Math.scala 150:24:@44809.4]
  wire [7:0] x713_x16_1_io_b; // @[Math.scala 150:24:@44809.4]
  wire [7:0] x713_x16_1_io_result; // @[Math.scala 150:24:@44809.4]
  wire [7:0] x714_x15_1_io_a; // @[Math.scala 150:24:@44819.4]
  wire [7:0] x714_x15_1_io_b; // @[Math.scala 150:24:@44819.4]
  wire [7:0] x714_x15_1_io_result; // @[Math.scala 150:24:@44819.4]
  wire [7:0] x715_x16_1_io_a; // @[Math.scala 150:24:@44829.4]
  wire [7:0] x715_x16_1_io_b; // @[Math.scala 150:24:@44829.4]
  wire [7:0] x715_x16_1_io_result; // @[Math.scala 150:24:@44829.4]
  wire [7:0] x716_x15_1_io_a; // @[Math.scala 150:24:@44839.4]
  wire [7:0] x716_x15_1_io_b; // @[Math.scala 150:24:@44839.4]
  wire [7:0] x716_x15_1_io_result; // @[Math.scala 150:24:@44839.4]
  wire  RetimeWrapper_125_clock; // @[package.scala 93:22:@44849.4]
  wire  RetimeWrapper_125_reset; // @[package.scala 93:22:@44849.4]
  wire  RetimeWrapper_125_io_flow; // @[package.scala 93:22:@44849.4]
  wire [7:0] RetimeWrapper_125_io_in; // @[package.scala 93:22:@44849.4]
  wire [7:0] RetimeWrapper_125_io_out; // @[package.scala 93:22:@44849.4]
  wire  x717_sum_1_clock; // @[Math.scala 150:24:@44858.4]
  wire  x717_sum_1_reset; // @[Math.scala 150:24:@44858.4]
  wire [7:0] x717_sum_1_io_a; // @[Math.scala 150:24:@44858.4]
  wire [7:0] x717_sum_1_io_b; // @[Math.scala 150:24:@44858.4]
  wire  x717_sum_1_io_flow; // @[Math.scala 150:24:@44858.4]
  wire [7:0] x717_sum_1_io_result; // @[Math.scala 150:24:@44858.4]
  wire  RetimeWrapper_126_clock; // @[package.scala 93:22:@44877.4]
  wire  RetimeWrapper_126_reset; // @[package.scala 93:22:@44877.4]
  wire  RetimeWrapper_126_io_flow; // @[package.scala 93:22:@44877.4]
  wire [8:0] RetimeWrapper_126_io_in; // @[package.scala 93:22:@44877.4]
  wire [8:0] RetimeWrapper_126_io_out; // @[package.scala 93:22:@44877.4]
  wire  RetimeWrapper_127_clock; // @[package.scala 93:22:@44889.4]
  wire  RetimeWrapper_127_reset; // @[package.scala 93:22:@44889.4]
  wire  RetimeWrapper_127_io_flow; // @[package.scala 93:22:@44889.4]
  wire [9:0] RetimeWrapper_127_io_in; // @[package.scala 93:22:@44889.4]
  wire [9:0] RetimeWrapper_127_io_out; // @[package.scala 93:22:@44889.4]
  wire  RetimeWrapper_128_clock; // @[package.scala 93:22:@44901.4]
  wire  RetimeWrapper_128_reset; // @[package.scala 93:22:@44901.4]
  wire  RetimeWrapper_128_io_flow; // @[package.scala 93:22:@44901.4]
  wire [8:0] RetimeWrapper_128_io_in; // @[package.scala 93:22:@44901.4]
  wire [8:0] RetimeWrapper_128_io_out; // @[package.scala 93:22:@44901.4]
  wire  RetimeWrapper_129_clock; // @[package.scala 93:22:@44913.4]
  wire  RetimeWrapper_129_reset; // @[package.scala 93:22:@44913.4]
  wire  RetimeWrapper_129_io_flow; // @[package.scala 93:22:@44913.4]
  wire [8:0] RetimeWrapper_129_io_in; // @[package.scala 93:22:@44913.4]
  wire [8:0] RetimeWrapper_129_io_out; // @[package.scala 93:22:@44913.4]
  wire [7:0] x723_x15_1_io_a; // @[Math.scala 150:24:@44923.4]
  wire [7:0] x723_x15_1_io_b; // @[Math.scala 150:24:@44923.4]
  wire [7:0] x723_x15_1_io_result; // @[Math.scala 150:24:@44923.4]
  wire  RetimeWrapper_130_clock; // @[package.scala 93:22:@44933.4]
  wire  RetimeWrapper_130_reset; // @[package.scala 93:22:@44933.4]
  wire  RetimeWrapper_130_io_flow; // @[package.scala 93:22:@44933.4]
  wire [7:0] RetimeWrapper_130_io_in; // @[package.scala 93:22:@44933.4]
  wire [7:0] RetimeWrapper_130_io_out; // @[package.scala 93:22:@44933.4]
  wire [7:0] x724_x16_1_io_a; // @[Math.scala 150:24:@44942.4]
  wire [7:0] x724_x16_1_io_b; // @[Math.scala 150:24:@44942.4]
  wire [7:0] x724_x16_1_io_result; // @[Math.scala 150:24:@44942.4]
  wire [7:0] x725_x15_1_io_a; // @[Math.scala 150:24:@44952.4]
  wire [7:0] x725_x15_1_io_b; // @[Math.scala 150:24:@44952.4]
  wire [7:0] x725_x15_1_io_result; // @[Math.scala 150:24:@44952.4]
  wire [7:0] x726_x16_1_io_a; // @[Math.scala 150:24:@44962.4]
  wire [7:0] x726_x16_1_io_b; // @[Math.scala 150:24:@44962.4]
  wire [7:0] x726_x16_1_io_result; // @[Math.scala 150:24:@44962.4]
  wire [7:0] x727_x15_1_io_a; // @[Math.scala 150:24:@44972.4]
  wire [7:0] x727_x15_1_io_b; // @[Math.scala 150:24:@44972.4]
  wire [7:0] x727_x15_1_io_result; // @[Math.scala 150:24:@44972.4]
  wire [7:0] x728_x16_1_io_a; // @[Math.scala 150:24:@44982.4]
  wire [7:0] x728_x16_1_io_b; // @[Math.scala 150:24:@44982.4]
  wire [7:0] x728_x16_1_io_result; // @[Math.scala 150:24:@44982.4]
  wire [7:0] x729_x15_1_io_a; // @[Math.scala 150:24:@44992.4]
  wire [7:0] x729_x15_1_io_b; // @[Math.scala 150:24:@44992.4]
  wire [7:0] x729_x15_1_io_result; // @[Math.scala 150:24:@44992.4]
  wire  RetimeWrapper_131_clock; // @[package.scala 93:22:@45002.4]
  wire  RetimeWrapper_131_reset; // @[package.scala 93:22:@45002.4]
  wire  RetimeWrapper_131_io_flow; // @[package.scala 93:22:@45002.4]
  wire [7:0] RetimeWrapper_131_io_in; // @[package.scala 93:22:@45002.4]
  wire [7:0] RetimeWrapper_131_io_out; // @[package.scala 93:22:@45002.4]
  wire  x730_sum_1_clock; // @[Math.scala 150:24:@45013.4]
  wire  x730_sum_1_reset; // @[Math.scala 150:24:@45013.4]
  wire [7:0] x730_sum_1_io_a; // @[Math.scala 150:24:@45013.4]
  wire [7:0] x730_sum_1_io_b; // @[Math.scala 150:24:@45013.4]
  wire  x730_sum_1_io_flow; // @[Math.scala 150:24:@45013.4]
  wire [7:0] x730_sum_1_io_result; // @[Math.scala 150:24:@45013.4]
  wire  RetimeWrapper_132_clock; // @[package.scala 93:22:@45040.4]
  wire  RetimeWrapper_132_reset; // @[package.scala 93:22:@45040.4]
  wire  RetimeWrapper_132_io_flow; // @[package.scala 93:22:@45040.4]
  wire [31:0] RetimeWrapper_132_io_in; // @[package.scala 93:22:@45040.4]
  wire [31:0] RetimeWrapper_132_io_out; // @[package.scala 93:22:@45040.4]
  wire  RetimeWrapper_133_clock; // @[package.scala 93:22:@45049.4]
  wire  RetimeWrapper_133_reset; // @[package.scala 93:22:@45049.4]
  wire  RetimeWrapper_133_io_flow; // @[package.scala 93:22:@45049.4]
  wire  RetimeWrapper_133_io_in; // @[package.scala 93:22:@45049.4]
  wire  RetimeWrapper_133_io_out; // @[package.scala 93:22:@45049.4]
  wire  RetimeWrapper_134_clock; // @[package.scala 93:22:@45058.4]
  wire  RetimeWrapper_134_reset; // @[package.scala 93:22:@45058.4]
  wire  RetimeWrapper_134_io_flow; // @[package.scala 93:22:@45058.4]
  wire  RetimeWrapper_134_io_in; // @[package.scala 93:22:@45058.4]
  wire  RetimeWrapper_134_io_out; // @[package.scala 93:22:@45058.4]
  wire  RetimeWrapper_135_clock; // @[package.scala 93:22:@45067.4]
  wire  RetimeWrapper_135_reset; // @[package.scala 93:22:@45067.4]
  wire  RetimeWrapper_135_io_flow; // @[package.scala 93:22:@45067.4]
  wire  RetimeWrapper_135_io_in; // @[package.scala 93:22:@45067.4]
  wire  RetimeWrapper_135_io_out; // @[package.scala 93:22:@45067.4]
  wire  b521; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 62:18:@42080.4]
  wire  b522; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 63:18:@42081.4]
  wire  _T_205; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 67:30:@42083.4]
  wire  _T_206; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 67:37:@42084.4]
  wire  _T_210; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 69:76:@42089.4]
  wire  _T_211; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 69:62:@42090.4]
  wire  _T_213; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 69:101:@42091.4]
  wire [31:0] x824_x523_D1_0_number; // @[package.scala 96:25:@42100.4 package.scala 96:25:@42101.4]
  wire [31:0] b519_number; // @[Math.scala 712:22:@42065.4 Math.scala 713:14:@42066.4]
  wire [31:0] _T_246; // @[Math.scala 499:52:@42265.4]
  wire  x528; // @[Math.scala 499:44:@42273.4]
  wire  x529; // @[Math.scala 499:44:@42280.4]
  wire  x530; // @[Math.scala 499:44:@42287.4]
  wire [31:0] _T_293; // @[Mux.scala 19:72:@42299.4]
  wire [31:0] _T_295; // @[Mux.scala 19:72:@42300.4]
  wire [31:0] _T_297; // @[Mux.scala 19:72:@42301.4]
  wire [31:0] _T_299; // @[Mux.scala 19:72:@42303.4]
  wire [31:0] x825_x531_D2_number; // @[package.scala 96:25:@42316.4 package.scala 96:25:@42317.4]
  wire [31:0] _T_314; // @[Math.scala 406:49:@42323.4]
  wire [31:0] _T_316; // @[Math.scala 406:56:@42325.4]
  wire [31:0] _T_317; // @[Math.scala 406:56:@42326.4]
  wire  _T_329; // @[FixedPoint.scala 50:25:@42344.4]
  wire [1:0] _T_333; // @[Bitwise.scala 72:12:@42346.4]
  wire [29:0] _T_334; // @[FixedPoint.scala 18:52:@42347.4]
  wire [31:0] x535_number; // @[Cat.scala 30:58:@42348.4]
  wire [39:0] _GEN_0; // @[Math.scala 450:32:@42353.4]
  wire [39:0] _T_339; // @[Math.scala 450:32:@42353.4]
  wire [37:0] _GEN_1; // @[Math.scala 450:32:@42358.4]
  wire [37:0] _T_343; // @[Math.scala 450:32:@42358.4]
  wire  _T_379; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 127:101:@42456.4]
  wire  _T_383; // @[package.scala 96:25:@42464.4 package.scala 96:25:@42465.4]
  wire  _T_385; // @[implicits.scala 55:10:@42466.4]
  wire  _T_386; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 127:118:@42467.4]
  wire  _T_388; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 127:207:@42469.4]
  wire  _T_389; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 127:226:@42470.4]
  wire  x830_b521_D24; // @[package.scala 96:25:@42435.4 package.scala 96:25:@42436.4]
  wire  _T_390; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 127:252:@42471.4]
  wire  x829_b522_D24; // @[package.scala 96:25:@42426.4 package.scala 96:25:@42427.4]
  wire  _T_434; // @[package.scala 96:25:@42571.4 package.scala 96:25:@42572.4]
  wire  _T_436; // @[implicits.scala 55:10:@42573.4]
  wire  _T_437; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 150:118:@42574.4]
  wire  _T_439; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 150:207:@42576.4]
  wire  _T_440; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 150:226:@42577.4]
  wire  _T_441; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 150:252:@42578.4]
  wire  _T_482; // @[package.scala 96:25:@42669.4 package.scala 96:25:@42670.4]
  wire  _T_484; // @[implicits.scala 55:10:@42671.4]
  wire  _T_485; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 171:118:@42672.4]
  wire  _T_487; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 171:207:@42674.4]
  wire  _T_488; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 171:226:@42675.4]
  wire  _T_489; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 171:252:@42676.4]
  wire  _T_532; // @[package.scala 96:25:@42769.4 package.scala 96:25:@42770.4]
  wire  _T_534; // @[implicits.scala 55:10:@42771.4]
  wire  _T_535; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 200:166:@42772.4]
  wire  _T_537; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 200:255:@42774.4]
  wire  _T_538; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 200:274:@42775.4]
  wire  _T_539; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 200:300:@42776.4]
  wire [31:0] x843_b519_D26_number; // @[package.scala 96:25:@42790.4 package.scala 96:25:@42791.4]
  wire [31:0] _T_551; // @[Math.scala 406:49:@42797.4]
  wire [31:0] _T_553; // @[Math.scala 406:56:@42799.4]
  wire [31:0] _T_554; // @[Math.scala 406:56:@42800.4]
  wire [31:0] _T_558; // @[package.scala 96:25:@42808.4]
  wire [31:0] x804_number; // @[implicits.scala 133:21:@42810.4]
  wire [31:0] x844_x552_rdcol_D26_number; // @[package.scala 96:25:@42833.4 package.scala 96:25:@42834.4]
  wire [31:0] _T_578; // @[Math.scala 465:37:@42839.4]
  wire  x845_x560_D1; // @[package.scala 96:25:@42856.4 package.scala 96:25:@42857.4]
  wire  x561; // @[package.scala 96:25:@42847.4 package.scala 96:25:@42848.4]
  wire  x562; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 215:24:@42860.4]
  wire [31:0] _T_597; // @[Math.scala 406:49:@42869.4]
  wire [31:0] _T_599; // @[Math.scala 406:56:@42871.4]
  wire [31:0] _T_600; // @[Math.scala 406:56:@42872.4]
  wire  _T_605; // @[FixedPoint.scala 50:25:@42878.4]
  wire [1:0] _T_609; // @[Bitwise.scala 72:12:@42880.4]
  wire [29:0] _T_610; // @[FixedPoint.scala 18:52:@42881.4]
  wire [31:0] x565_number; // @[Cat.scala 30:58:@42882.4]
  wire [39:0] _GEN_2; // @[Math.scala 450:32:@42887.4]
  wire [39:0] _T_615; // @[Math.scala 450:32:@42887.4]
  wire [37:0] _GEN_3; // @[Math.scala 450:32:@42892.4]
  wire [37:0] _T_619; // @[Math.scala 450:32:@42892.4]
  wire  _T_658; // @[package.scala 96:25:@42987.4 package.scala 96:25:@42988.4]
  wire  _T_660; // @[implicits.scala 55:10:@42989.4]
  wire  _T_661; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 248:194:@42990.4]
  wire  x852_x563_D20; // @[package.scala 96:25:@42975.4 package.scala 96:25:@42976.4]
  wire  _T_662; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 248:283:@42991.4]
  wire  x851_b521_D48; // @[package.scala 96:25:@42966.4 package.scala 96:25:@42967.4]
  wire  _T_663; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 248:291:@42992.4]
  wire  x848_b522_D48; // @[package.scala 96:25:@42939.4 package.scala 96:25:@42940.4]
  wire [31:0] x853_x546_rdcol_D26_number; // @[package.scala 96:25:@43008.4 package.scala 96:25:@43009.4]
  wire [31:0] _T_674; // @[Math.scala 465:37:@43014.4]
  wire  x570; // @[package.scala 96:25:@43022.4 package.scala 96:25:@43023.4]
  wire  x571; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 256:24:@43026.4]
  wire  _T_706; // @[package.scala 96:25:@43077.4 package.scala 96:25:@43078.4]
  wire  _T_708; // @[implicits.scala 55:10:@43079.4]
  wire  _T_709; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 271:194:@43080.4]
  wire  x855_x572_D20; // @[package.scala 96:25:@43056.4 package.scala 96:25:@43057.4]
  wire  _T_710; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 271:283:@43081.4]
  wire  _T_711; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 271:291:@43082.4]
  wire [31:0] x857_x540_rdcol_D26_number; // @[package.scala 96:25:@43098.4 package.scala 96:25:@43099.4]
  wire [31:0] _T_722; // @[Math.scala 465:37:@43104.4]
  wire  x576; // @[package.scala 96:25:@43112.4 package.scala 96:25:@43113.4]
  wire  x577; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 279:24:@43116.4]
  wire  _T_754; // @[package.scala 96:25:@43167.4 package.scala 96:25:@43168.4]
  wire  _T_756; // @[implicits.scala 55:10:@43169.4]
  wire  _T_757; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 300:194:@43170.4]
  wire  x860_x578_D20; // @[package.scala 96:25:@43155.4 package.scala 96:25:@43156.4]
  wire  _T_758; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 300:283:@43171.4]
  wire  _T_759; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 300:326:@43172.4]
  wire [31:0] x861_b520_D26_number; // @[package.scala 96:25:@43188.4 package.scala 96:25:@43189.4]
  wire [31:0] _T_772; // @[Math.scala 465:37:@43196.4]
  wire  x560; // @[package.scala 96:25:@42824.4 package.scala 96:25:@42825.4]
  wire  x582; // @[package.scala 96:25:@43204.4 package.scala 96:25:@43205.4]
  wire  x583; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 310:59:@43208.4]
  wire  _T_810; // @[package.scala 96:25:@43277.4 package.scala 96:25:@43278.4]
  wire  _T_812; // @[implicits.scala 55:10:@43279.4]
  wire  _T_813; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 329:194:@43280.4]
  wire  x865_x584_D21; // @[package.scala 96:25:@43256.4 package.scala 96:25:@43257.4]
  wire  _T_814; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 329:283:@43281.4]
  wire  _T_815; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 329:291:@43282.4]
  wire [31:0] x588_rdcol_number; // @[Math.scala 154:22:@43301.4 Math.scala 155:14:@43302.4]
  wire [31:0] _T_830; // @[Math.scala 465:37:@43307.4]
  wire  x589; // @[package.scala 96:25:@43315.4 package.scala 96:25:@43316.4]
  wire  x590; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 337:59:@43319.4]
  wire  _T_873; // @[package.scala 96:25:@43385.4 package.scala 96:25:@43386.4]
  wire  _T_875; // @[implicits.scala 55:10:@43387.4]
  wire  _T_876; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 354:194:@43388.4]
  wire  x867_x591_D20; // @[package.scala 96:25:@43364.4 package.scala 96:25:@43365.4]
  wire  _T_877; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 354:283:@43389.4]
  wire  _T_878; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 354:291:@43390.4]
  wire [31:0] x597_rdcol_number; // @[Math.scala 154:22:@43409.4 Math.scala 155:14:@43410.4]
  wire [31:0] _T_893; // @[Math.scala 465:37:@43415.4]
  wire  x598; // @[package.scala 96:25:@43423.4 package.scala 96:25:@43424.4]
  wire  x599; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 362:59:@43427.4]
  wire  _T_936; // @[package.scala 96:25:@43493.4 package.scala 96:25:@43494.4]
  wire  _T_938; // @[implicits.scala 55:10:@43495.4]
  wire  _T_939; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 379:194:@43496.4]
  wire  x870_x600_D20; // @[package.scala 96:25:@43481.4 package.scala 96:25:@43482.4]
  wire  _T_940; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 379:283:@43497.4]
  wire  _T_941; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 379:291:@43498.4]
  wire [31:0] x606_rdrow_number; // @[Math.scala 195:22:@43517.4 Math.scala 196:14:@43518.4]
  wire [31:0] _T_958; // @[Math.scala 406:49:@43524.4]
  wire [31:0] _T_960; // @[Math.scala 406:56:@43526.4]
  wire [31:0] _T_961; // @[Math.scala 406:56:@43527.4]
  wire [31:0] _T_965; // @[package.scala 96:25:@43535.4]
  wire [31:0] x809_number; // @[implicits.scala 133:21:@43537.4]
  wire  x608; // @[package.scala 96:25:@43551.4 package.scala 96:25:@43552.4]
  wire  x609; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 389:24:@43555.4]
  wire [31:0] _T_988; // @[Math.scala 406:49:@43564.4]
  wire [31:0] _T_990; // @[Math.scala 406:56:@43566.4]
  wire [31:0] _T_991; // @[Math.scala 406:56:@43567.4]
  wire  _T_996; // @[FixedPoint.scala 50:25:@43573.4]
  wire [1:0] _T_1000; // @[Bitwise.scala 72:12:@43575.4]
  wire [29:0] _T_1001; // @[FixedPoint.scala 18:52:@43576.4]
  wire [31:0] x612_number; // @[Cat.scala 30:58:@43577.4]
  wire [39:0] _GEN_4; // @[Math.scala 450:32:@43582.4]
  wire [39:0] _T_1006; // @[Math.scala 450:32:@43582.4]
  wire [37:0] _GEN_5; // @[Math.scala 450:32:@43587.4]
  wire [37:0] _T_1010; // @[Math.scala 450:32:@43587.4]
  wire  _T_1037; // @[package.scala 96:25:@43646.4 package.scala 96:25:@43647.4]
  wire  _T_1039; // @[implicits.scala 55:10:@43648.4]
  wire  _T_1040; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 420:194:@43649.4]
  wire  x873_x610_D20; // @[package.scala 96:25:@43634.4 package.scala 96:25:@43635.4]
  wire  _T_1041; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 420:283:@43650.4]
  wire  _T_1042; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 420:291:@43651.4]
  wire  x617; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 424:59:@43662.4]
  wire  _T_1068; // @[package.scala 96:25:@43697.4 package.scala 96:25:@43698.4]
  wire  _T_1070; // @[implicits.scala 55:10:@43699.4]
  wire  _T_1071; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 437:194:@43700.4]
  wire  x874_x618_D20; // @[package.scala 96:25:@43685.4 package.scala 96:25:@43686.4]
  wire  _T_1072; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 437:283:@43701.4]
  wire  _T_1073; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 437:291:@43702.4]
  wire  x622; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 441:59:@43713.4]
  wire  _T_1097; // @[package.scala 96:25:@43746.4 package.scala 96:25:@43747.4]
  wire  _T_1099; // @[implicits.scala 55:10:@43748.4]
  wire  _T_1100; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 452:194:@43749.4]
  wire  x875_x623_D20; // @[package.scala 96:25:@43734.4 package.scala 96:25:@43735.4]
  wire  _T_1101; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 452:283:@43750.4]
  wire  _T_1102; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 452:291:@43751.4]
  wire  x876_x582_D1; // @[package.scala 96:25:@43767.4 package.scala 96:25:@43768.4]
  wire  x627; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 458:59:@43771.4]
  wire  _T_1135; // @[package.scala 96:25:@43822.4 package.scala 96:25:@43823.4]
  wire  _T_1137; // @[implicits.scala 55:10:@43824.4]
  wire  _T_1138; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 473:194:@43825.4]
  wire  x879_x628_D20; // @[package.scala 96:25:@43810.4 package.scala 96:25:@43811.4]
  wire  _T_1139; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 473:283:@43826.4]
  wire  _T_1140; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 473:291:@43827.4]
  wire  x632; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 477:59:@43838.4]
  wire  _T_1164; // @[package.scala 96:25:@43871.4 package.scala 96:25:@43872.4]
  wire  _T_1166; // @[implicits.scala 55:10:@43873.4]
  wire  _T_1167; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 488:194:@43874.4]
  wire  x880_x633_D20; // @[package.scala 96:25:@43859.4 package.scala 96:25:@43860.4]
  wire  _T_1168; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 488:283:@43875.4]
  wire  _T_1169; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 488:291:@43876.4]
  wire  x637; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 492:59:@43887.4]
  wire  _T_1193; // @[package.scala 96:25:@43920.4 package.scala 96:25:@43921.4]
  wire  _T_1195; // @[implicits.scala 55:10:@43922.4]
  wire  _T_1196; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 503:194:@43923.4]
  wire  x881_x638_D20; // @[package.scala 96:25:@43908.4 package.scala 96:25:@43909.4]
  wire  _T_1197; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 503:283:@43924.4]
  wire  _T_1198; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 503:291:@43925.4]
  wire [31:0] x642_rdrow_number; // @[Math.scala 195:22:@43944.4 Math.scala 196:14:@43945.4]
  wire [31:0] _T_1215; // @[Math.scala 406:49:@43951.4]
  wire [31:0] _T_1217; // @[Math.scala 406:56:@43953.4]
  wire [31:0] _T_1218; // @[Math.scala 406:56:@43954.4]
  wire [31:0] _T_1222; // @[package.scala 96:25:@43962.4]
  wire [31:0] x814_number; // @[implicits.scala 133:21:@43964.4]
  wire  x644; // @[package.scala 96:25:@43978.4 package.scala 96:25:@43979.4]
  wire  x645; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 513:24:@43982.4]
  wire [31:0] _T_1245; // @[Math.scala 406:49:@43991.4]
  wire [31:0] _T_1247; // @[Math.scala 406:56:@43993.4]
  wire [31:0] _T_1248; // @[Math.scala 406:56:@43994.4]
  wire  _T_1253; // @[FixedPoint.scala 50:25:@44000.4]
  wire [1:0] _T_1257; // @[Bitwise.scala 72:12:@44002.4]
  wire [29:0] _T_1258; // @[FixedPoint.scala 18:52:@44003.4]
  wire [31:0] x648_number; // @[Cat.scala 30:58:@44004.4]
  wire [39:0] _GEN_6; // @[Math.scala 450:32:@44009.4]
  wire [39:0] _T_1263; // @[Math.scala 450:32:@44009.4]
  wire [37:0] _GEN_7; // @[Math.scala 450:32:@44014.4]
  wire [37:0] _T_1267; // @[Math.scala 450:32:@44014.4]
  wire  _T_1294; // @[package.scala 96:25:@44073.4 package.scala 96:25:@44074.4]
  wire  _T_1296; // @[implicits.scala 55:10:@44075.4]
  wire  _T_1297; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 544:194:@44076.4]
  wire  x883_x646_D20; // @[package.scala 96:25:@44052.4 package.scala 96:25:@44053.4]
  wire  _T_1298; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 544:283:@44077.4]
  wire  _T_1299; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 544:326:@44078.4]
  wire  x653; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 548:59:@44089.4]
  wire  _T_1325; // @[package.scala 96:25:@44124.4 package.scala 96:25:@44125.4]
  wire  _T_1327; // @[implicits.scala 55:10:@44126.4]
  wire  _T_1328; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 561:194:@44127.4]
  wire  x885_x654_D20; // @[package.scala 96:25:@44112.4 package.scala 96:25:@44113.4]
  wire  _T_1329; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 561:283:@44128.4]
  wire  _T_1330; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 561:291:@44129.4]
  wire  x658; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 565:59:@44140.4]
  wire  _T_1354; // @[package.scala 96:25:@44173.4 package.scala 96:25:@44174.4]
  wire  _T_1356; // @[implicits.scala 55:10:@44175.4]
  wire  _T_1357; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 576:194:@44176.4]
  wire  x886_x659_D20; // @[package.scala 96:25:@44161.4 package.scala 96:25:@44162.4]
  wire  _T_1358; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 576:283:@44177.4]
  wire  _T_1359; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 576:291:@44178.4]
  wire  x663; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 580:59:@44189.4]
  wire  _T_1389; // @[package.scala 96:25:@44240.4 package.scala 96:25:@44241.4]
  wire  _T_1391; // @[implicits.scala 55:10:@44242.4]
  wire  _T_1392; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 595:194:@44243.4]
  wire  x889_x664_D20; // @[package.scala 96:25:@44228.4 package.scala 96:25:@44229.4]
  wire  _T_1393; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 595:283:@44244.4]
  wire  _T_1394; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 595:291:@44245.4]
  wire  x668; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 599:59:@44256.4]
  wire  _T_1418; // @[package.scala 96:25:@44289.4 package.scala 96:25:@44290.4]
  wire  _T_1420; // @[implicits.scala 55:10:@44291.4]
  wire  _T_1421; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 610:194:@44292.4]
  wire  x890_x669_D20; // @[package.scala 96:25:@44277.4 package.scala 96:25:@44278.4]
  wire  _T_1422; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 610:283:@44293.4]
  wire  _T_1423; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 610:291:@44294.4]
  wire  x673; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 614:59:@44305.4]
  wire  _T_1447; // @[package.scala 96:25:@44338.4 package.scala 96:25:@44339.4]
  wire  _T_1449; // @[implicits.scala 55:10:@44340.4]
  wire  _T_1450; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 625:194:@44341.4]
  wire  x891_x674_D20; // @[package.scala 96:25:@44326.4 package.scala 96:25:@44327.4]
  wire  _T_1451; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 625:283:@44342.4]
  wire  _T_1452; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 625:291:@44343.4]
  wire [7:0] x574_rd_0_number; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 267:29:@43068.4 sm_x736_inr_Foreach_SAMPLER_BOX.scala 271:338:@43089.4]
  wire [8:0] _GEN_8; // @[Math.scala 450:32:@44355.4]
  wire [7:0] x615_rd_0_number; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 416:29:@43637.4 sm_x736_inr_Foreach_SAMPLER_BOX.scala 420:408:@43658.4]
  wire [8:0] _GEN_9; // @[Math.scala 450:32:@44367.4]
  wire [7:0] x620_rd_0_number; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 433:29:@43688.4 sm_x736_inr_Foreach_SAMPLER_BOX.scala 437:408:@43709.4]
  wire [9:0] _GEN_10; // @[Math.scala 450:32:@44379.4]
  wire [7:0] x625_rd_0_number; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 448:29:@43737.4 sm_x736_inr_Foreach_SAMPLER_BOX.scala 452:408:@43758.4]
  wire [8:0] _GEN_11; // @[Math.scala 450:32:@44391.4]
  wire [7:0] x656_rd_0_number; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 557:29:@44115.4 sm_x736_inr_Foreach_SAMPLER_BOX.scala 561:408:@44136.4]
  wire [8:0] _GEN_12; // @[Math.scala 450:32:@44403.4]
  wire [7:0] x690_sum_number; // @[Math.scala 154:22:@44528.4 Math.scala 155:14:@44529.4]
  wire [3:0] _T_1531; // @[FixedPoint.scala 18:52:@44534.4]
  wire [7:0] x580_rd_0_number; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 296:29:@43158.4 sm_x736_inr_Foreach_SAMPLER_BOX.scala 300:443:@43179.4]
  wire [8:0] _GEN_13; // @[Math.scala 450:32:@44540.4]
  wire [8:0] _GEN_14; // @[Math.scala 450:32:@44552.4]
  wire [9:0] _GEN_15; // @[Math.scala 450:32:@44564.4]
  wire [7:0] x630_rd_0_number; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 469:29:@43813.4 sm_x736_inr_Foreach_SAMPLER_BOX.scala 473:408:@43834.4]
  wire [8:0] _GEN_16; // @[Math.scala 450:32:@44576.4]
  wire [7:0] x661_rd_0_number; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 572:29:@44164.4 sm_x736_inr_Foreach_SAMPLER_BOX.scala 576:408:@44185.4]
  wire [8:0] _GEN_17; // @[Math.scala 450:32:@44588.4]
  wire [7:0] x704_sum_number; // @[Math.scala 154:22:@44711.4 Math.scala 155:14:@44712.4]
  wire [3:0] _T_1607; // @[FixedPoint.scala 18:52:@44717.4]
  wire [7:0] x586_rd_0_number; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 325:29:@43268.4 sm_x736_inr_Foreach_SAMPLER_BOX.scala 329:408:@43289.4]
  wire [8:0] _GEN_18; // @[Math.scala 450:32:@44723.4]
  wire [9:0] _GEN_19; // @[Math.scala 450:32:@44735.4]
  wire [7:0] x635_rd_0_number; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 484:29:@43862.4 sm_x736_inr_Foreach_SAMPLER_BOX.scala 488:408:@43883.4]
  wire [8:0] _GEN_20; // @[Math.scala 450:32:@44747.4]
  wire [7:0] x666_rd_0_number; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 591:29:@44231.4 sm_x736_inr_Foreach_SAMPLER_BOX.scala 595:408:@44252.4]
  wire [8:0] _GEN_21; // @[Math.scala 450:32:@44759.4]
  wire [7:0] x717_sum_number; // @[Math.scala 154:22:@44864.4 Math.scala 155:14:@44865.4]
  wire [3:0] _T_1671; // @[FixedPoint.scala 18:52:@44870.4]
  wire [7:0] x595_rd_0_number; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 350:29:@43376.4 sm_x736_inr_Foreach_SAMPLER_BOX.scala 354:408:@43397.4]
  wire [8:0] _GEN_22; // @[Math.scala 450:32:@44876.4]
  wire [9:0] _GEN_23; // @[Math.scala 450:32:@44888.4]
  wire [7:0] x640_rd_0_number; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 499:29:@43911.4 sm_x736_inr_Foreach_SAMPLER_BOX.scala 503:408:@43932.4]
  wire [8:0] _GEN_24; // @[Math.scala 450:32:@44900.4]
  wire [7:0] x671_rd_0_number; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 606:29:@44280.4 sm_x736_inr_Foreach_SAMPLER_BOX.scala 610:408:@44301.4]
  wire [8:0] _GEN_25; // @[Math.scala 450:32:@44912.4]
  wire [7:0] x730_sum_number; // @[Math.scala 154:22:@45019.4 Math.scala 155:14:@45020.4]
  wire [3:0] _T_1737; // @[FixedPoint.scala 18:52:@45025.4]
  wire [15:0] _T_1750; // @[Cat.scala 30:58:@45035.4]
  wire [15:0] _T_1751; // @[Cat.scala 30:58:@45036.4]
  wire  _T_1764; // @[package.scala 96:25:@45072.4 package.scala 96:25:@45073.4]
  wire  _T_1766; // @[implicits.scala 55:10:@45074.4]
  wire  x904_b521_D55; // @[package.scala 96:25:@45054.4 package.scala 96:25:@45055.4]
  wire  _T_1767; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 785:117:@45075.4]
  wire  x905_b522_D55; // @[package.scala 96:25:@45063.4 package.scala 96:25:@45064.4]
  wire  _T_1768; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 785:123:@45076.4]
  wire [31:0] x827_x538_sum_D3_number; // @[package.scala 96:25:@42408.4 package.scala 96:25:@42409.4]
  wire [31:0] x828_x534_D8_number; // @[package.scala 96:25:@42417.4 package.scala 96:25:@42418.4]
  wire [31:0] x831_x800_D22_number; // @[package.scala 96:25:@42444.4 package.scala 96:25:@42445.4]
  wire [31:0] x834_x542_D7_number; // @[package.scala 96:25:@42542.4 package.scala 96:25:@42543.4]
  wire [31:0] x836_x544_sum_D2_number; // @[package.scala 96:25:@42560.4 package.scala 96:25:@42561.4]
  wire [31:0] x837_x550_sum_D2_number; // @[package.scala 96:25:@42640.4 package.scala 96:25:@42641.4]
  wire [31:0] x839_x548_D7_number; // @[package.scala 96:25:@42658.4 package.scala 96:25:@42659.4]
  wire [31:0] x840_x554_D7_number; // @[package.scala 96:25:@42740.4 package.scala 96:25:@42741.4]
  wire [31:0] x842_x556_sum_D2_number; // @[package.scala 96:25:@42758.4 package.scala 96:25:@42759.4]
  wire [31:0] x567_sum_number; // @[Math.scala 154:22:@42930.4 Math.scala 155:14:@42931.4]
  wire [31:0] x849_x554_D31_number; // @[package.scala 96:25:@42948.4 package.scala 96:25:@42949.4]
  wire [31:0] x850_x805_D21_number; // @[package.scala 96:25:@42957.4 package.scala 96:25:@42958.4]
  wire [31:0] x573_sum_number; // @[Math.scala 154:22:@43047.4 Math.scala 155:14:@43048.4]
  wire [31:0] x856_x548_D31_number; // @[package.scala 96:25:@43065.4 package.scala 96:25:@43066.4]
  wire [31:0] x579_sum_number; // @[Math.scala 154:22:@43137.4 Math.scala 155:14:@43138.4]
  wire [31:0] x859_x542_D31_number; // @[package.scala 96:25:@43146.4 package.scala 96:25:@43147.4]
  wire [31:0] x864_x534_D32_number; // @[package.scala 96:25:@43247.4 package.scala 96:25:@43248.4]
  wire [31:0] x866_x585_sum_D1_number; // @[package.scala 96:25:@43265.4 package.scala 96:25:@43266.4]
  wire [31:0] x594_sum_number; // @[Math.scala 154:22:@43355.4 Math.scala 155:14:@43356.4]
  wire [31:0] x868_x592_D5_number; // @[package.scala 96:25:@43373.4 package.scala 96:25:@43374.4]
  wire [31:0] x603_sum_number; // @[Math.scala 154:22:@43463.4 Math.scala 155:14:@43464.4]
  wire [31:0] x869_x601_D5_number; // @[package.scala 96:25:@43472.4 package.scala 96:25:@43473.4]
  wire [31:0] x614_sum_number; // @[Math.scala 154:22:@43616.4 Math.scala 155:14:@43617.4]
  wire [31:0] x872_x810_D20_number; // @[package.scala 96:25:@43625.4 package.scala 96:25:@43626.4]
  wire [31:0] x619_sum_number; // @[Math.scala 154:22:@43676.4 Math.scala 155:14:@43677.4]
  wire [31:0] x624_sum_number; // @[Math.scala 154:22:@43725.4 Math.scala 155:14:@43726.4]
  wire [31:0] x878_x629_sum_D1_number; // @[package.scala 96:25:@43801.4 package.scala 96:25:@43802.4]
  wire [31:0] x634_sum_number; // @[Math.scala 154:22:@43850.4 Math.scala 155:14:@43851.4]
  wire [31:0] x639_sum_number; // @[Math.scala 154:22:@43899.4 Math.scala 155:14:@43900.4]
  wire [31:0] x650_sum_number; // @[Math.scala 154:22:@44043.4 Math.scala 155:14:@44044.4]
  wire [31:0] x884_x815_D20_number; // @[package.scala 96:25:@44061.4 package.scala 96:25:@44062.4]
  wire [31:0] x655_sum_number; // @[Math.scala 154:22:@44103.4 Math.scala 155:14:@44104.4]
  wire [31:0] x660_sum_number; // @[Math.scala 154:22:@44152.4 Math.scala 155:14:@44153.4]
  wire [31:0] x888_x665_sum_D1_number; // @[package.scala 96:25:@44219.4 package.scala 96:25:@44220.4]
  wire [31:0] x670_sum_number; // @[Math.scala 154:22:@44268.4 Math.scala 155:14:@44269.4]
  wire [31:0] x675_sum_number; // @[Math.scala 154:22:@44317.4 Math.scala 155:14:@44318.4]
  wire [8:0] _T_1460; // @[package.scala 96:25:@44361.4 package.scala 96:25:@44362.4]
  wire [8:0] _T_1466; // @[package.scala 96:25:@44373.4 package.scala 96:25:@44374.4]
  wire [9:0] _T_1472; // @[package.scala 96:25:@44385.4 package.scala 96:25:@44386.4]
  wire [8:0] _T_1478; // @[package.scala 96:25:@44397.4 package.scala 96:25:@44398.4]
  wire [8:0] _T_1484; // @[package.scala 96:25:@44409.4 package.scala 96:25:@44410.4]
  wire [8:0] _T_1538; // @[package.scala 96:25:@44546.4 package.scala 96:25:@44547.4]
  wire [8:0] _T_1544; // @[package.scala 96:25:@44558.4 package.scala 96:25:@44559.4]
  wire [9:0] _T_1550; // @[package.scala 96:25:@44570.4 package.scala 96:25:@44571.4]
  wire [8:0] _T_1556; // @[package.scala 96:25:@44582.4 package.scala 96:25:@44583.4]
  wire [8:0] _T_1562; // @[package.scala 96:25:@44594.4 package.scala 96:25:@44595.4]
  wire [8:0] _T_1614; // @[package.scala 96:25:@44729.4 package.scala 96:25:@44730.4]
  wire [9:0] _T_1620; // @[package.scala 96:25:@44741.4 package.scala 96:25:@44742.4]
  wire [8:0] _T_1626; // @[package.scala 96:25:@44753.4 package.scala 96:25:@44754.4]
  wire [8:0] _T_1632; // @[package.scala 96:25:@44765.4 package.scala 96:25:@44766.4]
  wire [8:0] _T_1678; // @[package.scala 96:25:@44882.4 package.scala 96:25:@44883.4]
  wire [9:0] _T_1684; // @[package.scala 96:25:@44894.4 package.scala 96:25:@44895.4]
  wire [8:0] _T_1690; // @[package.scala 96:25:@44906.4 package.scala 96:25:@44907.4]
  wire [8:0] _T_1696; // @[package.scala 96:25:@44918.4 package.scala 96:25:@44919.4]
  _ _ ( // @[Math.scala 709:24:@42060.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 709:24:@42072.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper ( // @[package.scala 93:22:@42095.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x525_lb_0 x525_lb_0 ( // @[m_x525_lb_0.scala 47:17:@42105.4]
    .clock(x525_lb_0_clock),
    .reset(x525_lb_0_reset),
    .io_rPort_17_banks_1(x525_lb_0_io_rPort_17_banks_1),
    .io_rPort_17_banks_0(x525_lb_0_io_rPort_17_banks_0),
    .io_rPort_17_ofs_0(x525_lb_0_io_rPort_17_ofs_0),
    .io_rPort_17_en_0(x525_lb_0_io_rPort_17_en_0),
    .io_rPort_17_backpressure(x525_lb_0_io_rPort_17_backpressure),
    .io_rPort_17_output_0(x525_lb_0_io_rPort_17_output_0),
    .io_rPort_16_banks_1(x525_lb_0_io_rPort_16_banks_1),
    .io_rPort_16_banks_0(x525_lb_0_io_rPort_16_banks_0),
    .io_rPort_16_ofs_0(x525_lb_0_io_rPort_16_ofs_0),
    .io_rPort_16_en_0(x525_lb_0_io_rPort_16_en_0),
    .io_rPort_16_backpressure(x525_lb_0_io_rPort_16_backpressure),
    .io_rPort_16_output_0(x525_lb_0_io_rPort_16_output_0),
    .io_rPort_15_banks_1(x525_lb_0_io_rPort_15_banks_1),
    .io_rPort_15_banks_0(x525_lb_0_io_rPort_15_banks_0),
    .io_rPort_15_ofs_0(x525_lb_0_io_rPort_15_ofs_0),
    .io_rPort_15_en_0(x525_lb_0_io_rPort_15_en_0),
    .io_rPort_15_backpressure(x525_lb_0_io_rPort_15_backpressure),
    .io_rPort_15_output_0(x525_lb_0_io_rPort_15_output_0),
    .io_rPort_14_banks_1(x525_lb_0_io_rPort_14_banks_1),
    .io_rPort_14_banks_0(x525_lb_0_io_rPort_14_banks_0),
    .io_rPort_14_ofs_0(x525_lb_0_io_rPort_14_ofs_0),
    .io_rPort_14_en_0(x525_lb_0_io_rPort_14_en_0),
    .io_rPort_14_backpressure(x525_lb_0_io_rPort_14_backpressure),
    .io_rPort_14_output_0(x525_lb_0_io_rPort_14_output_0),
    .io_rPort_13_banks_1(x525_lb_0_io_rPort_13_banks_1),
    .io_rPort_13_banks_0(x525_lb_0_io_rPort_13_banks_0),
    .io_rPort_13_ofs_0(x525_lb_0_io_rPort_13_ofs_0),
    .io_rPort_13_en_0(x525_lb_0_io_rPort_13_en_0),
    .io_rPort_13_backpressure(x525_lb_0_io_rPort_13_backpressure),
    .io_rPort_13_output_0(x525_lb_0_io_rPort_13_output_0),
    .io_rPort_12_banks_1(x525_lb_0_io_rPort_12_banks_1),
    .io_rPort_12_banks_0(x525_lb_0_io_rPort_12_banks_0),
    .io_rPort_12_ofs_0(x525_lb_0_io_rPort_12_ofs_0),
    .io_rPort_12_en_0(x525_lb_0_io_rPort_12_en_0),
    .io_rPort_12_backpressure(x525_lb_0_io_rPort_12_backpressure),
    .io_rPort_12_output_0(x525_lb_0_io_rPort_12_output_0),
    .io_rPort_11_banks_1(x525_lb_0_io_rPort_11_banks_1),
    .io_rPort_11_banks_0(x525_lb_0_io_rPort_11_banks_0),
    .io_rPort_11_ofs_0(x525_lb_0_io_rPort_11_ofs_0),
    .io_rPort_11_en_0(x525_lb_0_io_rPort_11_en_0),
    .io_rPort_11_backpressure(x525_lb_0_io_rPort_11_backpressure),
    .io_rPort_11_output_0(x525_lb_0_io_rPort_11_output_0),
    .io_rPort_10_banks_1(x525_lb_0_io_rPort_10_banks_1),
    .io_rPort_10_banks_0(x525_lb_0_io_rPort_10_banks_0),
    .io_rPort_10_ofs_0(x525_lb_0_io_rPort_10_ofs_0),
    .io_rPort_10_en_0(x525_lb_0_io_rPort_10_en_0),
    .io_rPort_10_backpressure(x525_lb_0_io_rPort_10_backpressure),
    .io_rPort_10_output_0(x525_lb_0_io_rPort_10_output_0),
    .io_rPort_9_banks_1(x525_lb_0_io_rPort_9_banks_1),
    .io_rPort_9_banks_0(x525_lb_0_io_rPort_9_banks_0),
    .io_rPort_9_ofs_0(x525_lb_0_io_rPort_9_ofs_0),
    .io_rPort_9_en_0(x525_lb_0_io_rPort_9_en_0),
    .io_rPort_9_backpressure(x525_lb_0_io_rPort_9_backpressure),
    .io_rPort_9_output_0(x525_lb_0_io_rPort_9_output_0),
    .io_rPort_8_banks_1(x525_lb_0_io_rPort_8_banks_1),
    .io_rPort_8_banks_0(x525_lb_0_io_rPort_8_banks_0),
    .io_rPort_8_ofs_0(x525_lb_0_io_rPort_8_ofs_0),
    .io_rPort_8_en_0(x525_lb_0_io_rPort_8_en_0),
    .io_rPort_8_backpressure(x525_lb_0_io_rPort_8_backpressure),
    .io_rPort_8_output_0(x525_lb_0_io_rPort_8_output_0),
    .io_rPort_7_banks_1(x525_lb_0_io_rPort_7_banks_1),
    .io_rPort_7_banks_0(x525_lb_0_io_rPort_7_banks_0),
    .io_rPort_7_ofs_0(x525_lb_0_io_rPort_7_ofs_0),
    .io_rPort_7_en_0(x525_lb_0_io_rPort_7_en_0),
    .io_rPort_7_backpressure(x525_lb_0_io_rPort_7_backpressure),
    .io_rPort_7_output_0(x525_lb_0_io_rPort_7_output_0),
    .io_rPort_6_banks_1(x525_lb_0_io_rPort_6_banks_1),
    .io_rPort_6_banks_0(x525_lb_0_io_rPort_6_banks_0),
    .io_rPort_6_ofs_0(x525_lb_0_io_rPort_6_ofs_0),
    .io_rPort_6_en_0(x525_lb_0_io_rPort_6_en_0),
    .io_rPort_6_backpressure(x525_lb_0_io_rPort_6_backpressure),
    .io_rPort_6_output_0(x525_lb_0_io_rPort_6_output_0),
    .io_rPort_5_banks_1(x525_lb_0_io_rPort_5_banks_1),
    .io_rPort_5_banks_0(x525_lb_0_io_rPort_5_banks_0),
    .io_rPort_5_ofs_0(x525_lb_0_io_rPort_5_ofs_0),
    .io_rPort_5_en_0(x525_lb_0_io_rPort_5_en_0),
    .io_rPort_5_backpressure(x525_lb_0_io_rPort_5_backpressure),
    .io_rPort_5_output_0(x525_lb_0_io_rPort_5_output_0),
    .io_rPort_4_banks_1(x525_lb_0_io_rPort_4_banks_1),
    .io_rPort_4_banks_0(x525_lb_0_io_rPort_4_banks_0),
    .io_rPort_4_ofs_0(x525_lb_0_io_rPort_4_ofs_0),
    .io_rPort_4_en_0(x525_lb_0_io_rPort_4_en_0),
    .io_rPort_4_backpressure(x525_lb_0_io_rPort_4_backpressure),
    .io_rPort_4_output_0(x525_lb_0_io_rPort_4_output_0),
    .io_rPort_3_banks_1(x525_lb_0_io_rPort_3_banks_1),
    .io_rPort_3_banks_0(x525_lb_0_io_rPort_3_banks_0),
    .io_rPort_3_ofs_0(x525_lb_0_io_rPort_3_ofs_0),
    .io_rPort_3_en_0(x525_lb_0_io_rPort_3_en_0),
    .io_rPort_3_backpressure(x525_lb_0_io_rPort_3_backpressure),
    .io_rPort_3_output_0(x525_lb_0_io_rPort_3_output_0),
    .io_rPort_2_banks_1(x525_lb_0_io_rPort_2_banks_1),
    .io_rPort_2_banks_0(x525_lb_0_io_rPort_2_banks_0),
    .io_rPort_2_ofs_0(x525_lb_0_io_rPort_2_ofs_0),
    .io_rPort_2_en_0(x525_lb_0_io_rPort_2_en_0),
    .io_rPort_2_backpressure(x525_lb_0_io_rPort_2_backpressure),
    .io_rPort_2_output_0(x525_lb_0_io_rPort_2_output_0),
    .io_rPort_1_banks_1(x525_lb_0_io_rPort_1_banks_1),
    .io_rPort_1_banks_0(x525_lb_0_io_rPort_1_banks_0),
    .io_rPort_1_ofs_0(x525_lb_0_io_rPort_1_ofs_0),
    .io_rPort_1_en_0(x525_lb_0_io_rPort_1_en_0),
    .io_rPort_1_backpressure(x525_lb_0_io_rPort_1_backpressure),
    .io_rPort_1_output_0(x525_lb_0_io_rPort_1_output_0),
    .io_rPort_0_banks_1(x525_lb_0_io_rPort_0_banks_1),
    .io_rPort_0_banks_0(x525_lb_0_io_rPort_0_banks_0),
    .io_rPort_0_ofs_0(x525_lb_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x525_lb_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x525_lb_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x525_lb_0_io_rPort_0_output_0),
    .io_wPort_3_banks_1(x525_lb_0_io_wPort_3_banks_1),
    .io_wPort_3_banks_0(x525_lb_0_io_wPort_3_banks_0),
    .io_wPort_3_ofs_0(x525_lb_0_io_wPort_3_ofs_0),
    .io_wPort_3_data_0(x525_lb_0_io_wPort_3_data_0),
    .io_wPort_3_en_0(x525_lb_0_io_wPort_3_en_0),
    .io_wPort_2_banks_1(x525_lb_0_io_wPort_2_banks_1),
    .io_wPort_2_banks_0(x525_lb_0_io_wPort_2_banks_0),
    .io_wPort_2_ofs_0(x525_lb_0_io_wPort_2_ofs_0),
    .io_wPort_2_data_0(x525_lb_0_io_wPort_2_data_0),
    .io_wPort_2_en_0(x525_lb_0_io_wPort_2_en_0),
    .io_wPort_1_banks_1(x525_lb_0_io_wPort_1_banks_1),
    .io_wPort_1_banks_0(x525_lb_0_io_wPort_1_banks_0),
    .io_wPort_1_ofs_0(x525_lb_0_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(x525_lb_0_io_wPort_1_data_0),
    .io_wPort_1_en_0(x525_lb_0_io_wPort_1_en_0),
    .io_wPort_0_banks_1(x525_lb_0_io_wPort_0_banks_1),
    .io_wPort_0_banks_0(x525_lb_0_io_wPort_0_banks_0),
    .io_wPort_0_ofs_0(x525_lb_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x525_lb_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x525_lb_0_io_wPort_0_en_0)
  );
  RetimeWrapper_297 RetimeWrapper_1 ( // @[package.scala 93:22:@42311.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x534 x534_1 ( // @[Math.scala 366:24:@42333.4]
    .clock(x534_1_clock),
    .reset(x534_1_reset),
    .io_a(x534_1_io_a),
    .io_flow(x534_1_io_flow),
    .io_result(x534_1_io_result)
  );
  x494_sum x803_sum_1 ( // @[Math.scala 150:24:@42362.4]
    .clock(x803_sum_1_clock),
    .reset(x803_sum_1_reset),
    .io_a(x803_sum_1_io_a),
    .io_b(x803_sum_1_io_b),
    .io_flow(x803_sum_1_io_flow),
    .io_result(x803_sum_1_io_result)
  );
  x537_div x537_div_1 ( // @[Math.scala 327:24:@42374.4]
    .clock(x537_div_1_clock),
    .reset(x537_div_1_reset),
    .io_a(x537_div_1_io_a),
    .io_flow(x537_div_1_io_flow),
    .io_result(x537_div_1_io_result)
  );
  RetimeWrapper_301 RetimeWrapper_2 ( // @[package.scala 93:22:@42384.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x494_sum x538_sum_1 ( // @[Math.scala 150:24:@42393.4]
    .clock(x538_sum_1_clock),
    .reset(x538_sum_1_reset),
    .io_a(x538_sum_1_io_a),
    .io_b(x538_sum_1_io_b),
    .io_flow(x538_sum_1_io_flow),
    .io_result(x538_sum_1_io_result)
  );
  RetimeWrapper_303 RetimeWrapper_3 ( // @[package.scala 93:22:@42403.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_304 RetimeWrapper_4 ( // @[package.scala 93:22:@42412.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_305 RetimeWrapper_5 ( // @[package.scala 93:22:@42421.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_305 RetimeWrapper_6 ( // @[package.scala 93:22:@42430.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_307 RetimeWrapper_7 ( // @[package.scala 93:22:@42439.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_308 RetimeWrapper_8 ( // @[package.scala 93:22:@42448.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_305 RetimeWrapper_9 ( // @[package.scala 93:22:@42459.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  x494_sum x540_rdcol_1 ( // @[Math.scala 150:24:@42482.4]
    .clock(x540_rdcol_1_clock),
    .reset(x540_rdcol_1_reset),
    .io_a(x540_rdcol_1_io_a),
    .io_b(x540_rdcol_1_io_b),
    .io_flow(x540_rdcol_1_io_flow),
    .io_result(x540_rdcol_1_io_result)
  );
  x534 x542_1 ( // @[Math.scala 366:24:@42496.4]
    .clock(x542_1_clock),
    .reset(x542_1_reset),
    .io_a(x542_1_io_a),
    .io_flow(x542_1_io_flow),
    .io_result(x542_1_io_result)
  );
  x537_div x543_div_1 ( // @[Math.scala 327:24:@42508.4]
    .clock(x543_div_1_clock),
    .reset(x543_div_1_reset),
    .io_a(x543_div_1_io_a),
    .io_flow(x543_div_1_io_flow),
    .io_result(x543_div_1_io_result)
  );
  RetimeWrapper_313 RetimeWrapper_10 ( // @[package.scala 93:22:@42518.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  x494_sum x544_sum_1 ( // @[Math.scala 150:24:@42527.4]
    .clock(x544_sum_1_clock),
    .reset(x544_sum_1_reset),
    .io_a(x544_sum_1_io_a),
    .io_b(x544_sum_1_io_b),
    .io_flow(x544_sum_1_io_flow),
    .io_result(x544_sum_1_io_result)
  );
  RetimeWrapper_315 RetimeWrapper_11 ( // @[package.scala 93:22:@42537.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_308 RetimeWrapper_12 ( // @[package.scala 93:22:@42546.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_297 RetimeWrapper_13 ( // @[package.scala 93:22:@42555.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_305 RetimeWrapper_14 ( // @[package.scala 93:22:@42566.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  x494_sum x546_rdcol_1 ( // @[Math.scala 150:24:@42589.4]
    .clock(x546_rdcol_1_clock),
    .reset(x546_rdcol_1_reset),
    .io_a(x546_rdcol_1_io_a),
    .io_b(x546_rdcol_1_io_b),
    .io_flow(x546_rdcol_1_io_flow),
    .io_result(x546_rdcol_1_io_result)
  );
  x534 x548_1 ( // @[Math.scala 366:24:@42603.4]
    .clock(x548_1_clock),
    .reset(x548_1_reset),
    .io_a(x548_1_io_a),
    .io_flow(x548_1_io_flow),
    .io_result(x548_1_io_result)
  );
  x537_div x549_div_1 ( // @[Math.scala 327:24:@42615.4]
    .clock(x549_div_1_clock),
    .reset(x549_div_1_reset),
    .io_a(x549_div_1_io_a),
    .io_flow(x549_div_1_io_flow),
    .io_result(x549_div_1_io_result)
  );
  x494_sum x550_sum_1 ( // @[Math.scala 150:24:@42625.4]
    .clock(x550_sum_1_clock),
    .reset(x550_sum_1_reset),
    .io_a(x550_sum_1_io_a),
    .io_b(x550_sum_1_io_b),
    .io_flow(x550_sum_1_io_flow),
    .io_result(x550_sum_1_io_result)
  );
  RetimeWrapper_297 RetimeWrapper_15 ( // @[package.scala 93:22:@42635.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_308 RetimeWrapper_16 ( // @[package.scala 93:22:@42644.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_315 RetimeWrapper_17 ( // @[package.scala 93:22:@42653.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_305 RetimeWrapper_18 ( // @[package.scala 93:22:@42664.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  x494_sum x552_rdcol_1 ( // @[Math.scala 150:24:@42687.4]
    .clock(x552_rdcol_1_clock),
    .reset(x552_rdcol_1_reset),
    .io_a(x552_rdcol_1_io_a),
    .io_b(x552_rdcol_1_io_b),
    .io_flow(x552_rdcol_1_io_flow),
    .io_result(x552_rdcol_1_io_result)
  );
  x534 x554_1 ( // @[Math.scala 366:24:@42703.4]
    .clock(x554_1_clock),
    .reset(x554_1_reset),
    .io_a(x554_1_io_a),
    .io_flow(x554_1_io_flow),
    .io_result(x554_1_io_result)
  );
  x537_div x555_div_1 ( // @[Math.scala 327:24:@42715.4]
    .clock(x555_div_1_clock),
    .reset(x555_div_1_reset),
    .io_a(x555_div_1_io_a),
    .io_flow(x555_div_1_io_flow),
    .io_result(x555_div_1_io_result)
  );
  x494_sum x556_sum_1 ( // @[Math.scala 150:24:@42725.4]
    .clock(x556_sum_1_clock),
    .reset(x556_sum_1_reset),
    .io_a(x556_sum_1_io_a),
    .io_b(x556_sum_1_io_b),
    .io_flow(x556_sum_1_io_flow),
    .io_result(x556_sum_1_io_result)
  );
  RetimeWrapper_315 RetimeWrapper_19 ( // @[package.scala 93:22:@42735.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_308 RetimeWrapper_20 ( // @[package.scala 93:22:@42744.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_297 RetimeWrapper_21 ( // @[package.scala 93:22:@42753.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_305 RetimeWrapper_22 ( // @[package.scala 93:22:@42764.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_335 RetimeWrapper_23 ( // @[package.scala 93:22:@42785.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_24 ( // @[package.scala 93:22:@42801.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper RetimeWrapper_25 ( // @[package.scala 93:22:@42819.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_335 RetimeWrapper_26 ( // @[package.scala 93:22:@42828.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper RetimeWrapper_27 ( // @[package.scala 93:22:@42842.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper RetimeWrapper_28 ( // @[package.scala 93:22:@42851.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  x494_sum x808_sum_1 ( // @[Math.scala 150:24:@42896.4]
    .clock(x808_sum_1_clock),
    .reset(x808_sum_1_reset),
    .io_a(x808_sum_1_io_a),
    .io_b(x808_sum_1_io_b),
    .io_flow(x808_sum_1_io_flow),
    .io_result(x808_sum_1_io_result)
  );
  RetimeWrapper_342 RetimeWrapper_29 ( // @[package.scala 93:22:@42906.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_335 RetimeWrapper_30 ( // @[package.scala 93:22:@42915.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  x494_sum x567_sum_1 ( // @[Math.scala 150:24:@42924.4]
    .clock(x567_sum_1_clock),
    .reset(x567_sum_1_reset),
    .io_a(x567_sum_1_io_a),
    .io_b(x567_sum_1_io_b),
    .io_flow(x567_sum_1_io_flow),
    .io_result(x567_sum_1_io_result)
  );
  RetimeWrapper_345 RetimeWrapper_31 ( // @[package.scala 93:22:@42934.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_346 RetimeWrapper_32 ( // @[package.scala 93:22:@42943.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_347 RetimeWrapper_33 ( // @[package.scala 93:22:@42952.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_345 RetimeWrapper_34 ( // @[package.scala 93:22:@42961.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_349 RetimeWrapper_35 ( // @[package.scala 93:22:@42970.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_345 RetimeWrapper_36 ( // @[package.scala 93:22:@42982.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_335 RetimeWrapper_37 ( // @[package.scala 93:22:@43003.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper RetimeWrapper_38 ( // @[package.scala 93:22:@43017.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_335 RetimeWrapper_39 ( // @[package.scala 93:22:@43032.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  x494_sum x573_sum_1 ( // @[Math.scala 150:24:@43041.4]
    .clock(x573_sum_1_clock),
    .reset(x573_sum_1_reset),
    .io_a(x573_sum_1_io_a),
    .io_b(x573_sum_1_io_b),
    .io_flow(x573_sum_1_io_flow),
    .io_result(x573_sum_1_io_result)
  );
  RetimeWrapper_349 RetimeWrapper_40 ( // @[package.scala 93:22:@43051.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper_346 RetimeWrapper_41 ( // @[package.scala 93:22:@43060.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_345 RetimeWrapper_42 ( // @[package.scala 93:22:@43072.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_335 RetimeWrapper_43 ( // @[package.scala 93:22:@43093.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper RetimeWrapper_44 ( // @[package.scala 93:22:@43107.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_335 RetimeWrapper_45 ( // @[package.scala 93:22:@43122.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  x494_sum x579_sum_1 ( // @[Math.scala 150:24:@43131.4]
    .clock(x579_sum_1_clock),
    .reset(x579_sum_1_reset),
    .io_a(x579_sum_1_io_a),
    .io_b(x579_sum_1_io_b),
    .io_flow(x579_sum_1_io_flow),
    .io_result(x579_sum_1_io_result)
  );
  RetimeWrapper_346 RetimeWrapper_46 ( // @[package.scala 93:22:@43141.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_349 RetimeWrapper_47 ( // @[package.scala 93:22:@43150.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_345 RetimeWrapper_48 ( // @[package.scala 93:22:@43162.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_335 RetimeWrapper_49 ( // @[package.scala 93:22:@43183.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper RetimeWrapper_50 ( // @[package.scala 93:22:@43199.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_313 RetimeWrapper_51 ( // @[package.scala 93:22:@43214.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_335 RetimeWrapper_52 ( // @[package.scala 93:22:@43223.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  x494_sum x585_sum_1 ( // @[Math.scala 150:24:@43232.4]
    .clock(x585_sum_1_clock),
    .reset(x585_sum_1_reset),
    .io_a(x585_sum_1_io_a),
    .io_b(x585_sum_1_io_b),
    .io_flow(x585_sum_1_io_flow),
    .io_result(x585_sum_1_io_result)
  );
  RetimeWrapper_370 RetimeWrapper_53 ( // @[package.scala 93:22:@43242.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper_371 RetimeWrapper_54 ( // @[package.scala 93:22:@43251.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_55 ( // @[package.scala 93:22:@43260.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper_345 RetimeWrapper_56 ( // @[package.scala 93:22:@43272.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  x494_sum x588_rdcol_1 ( // @[Math.scala 150:24:@43295.4]
    .clock(x588_rdcol_1_clock),
    .reset(x588_rdcol_1_reset),
    .io_a(x588_rdcol_1_io_a),
    .io_b(x588_rdcol_1_io_b),
    .io_flow(x588_rdcol_1_io_flow),
    .io_result(x588_rdcol_1_io_result)
  );
  RetimeWrapper RetimeWrapper_57 ( // @[package.scala 93:22:@43310.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  x534 x592_1 ( // @[Math.scala 366:24:@43327.4]
    .clock(x592_1_clock),
    .reset(x592_1_reset),
    .io_a(x592_1_io_a),
    .io_flow(x592_1_io_flow),
    .io_result(x592_1_io_result)
  );
  x537_div x593_div_1 ( // @[Math.scala 327:24:@43339.4]
    .clock(x593_div_1_clock),
    .reset(x593_div_1_reset),
    .io_a(x593_div_1_io_a),
    .io_flow(x593_div_1_io_flow),
    .io_result(x593_div_1_io_result)
  );
  x494_sum x594_sum_1 ( // @[Math.scala 150:24:@43349.4]
    .clock(x594_sum_1_clock),
    .reset(x594_sum_1_reset),
    .io_a(x594_sum_1_io_a),
    .io_b(x594_sum_1_io_b),
    .io_flow(x594_sum_1_io_flow),
    .io_result(x594_sum_1_io_result)
  );
  RetimeWrapper_349 RetimeWrapper_58 ( // @[package.scala 93:22:@43359.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_380 RetimeWrapper_59 ( // @[package.scala 93:22:@43368.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_345 RetimeWrapper_60 ( // @[package.scala 93:22:@43380.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  x494_sum x597_rdcol_1 ( // @[Math.scala 150:24:@43403.4]
    .clock(x597_rdcol_1_clock),
    .reset(x597_rdcol_1_reset),
    .io_a(x597_rdcol_1_io_a),
    .io_b(x597_rdcol_1_io_b),
    .io_flow(x597_rdcol_1_io_flow),
    .io_result(x597_rdcol_1_io_result)
  );
  RetimeWrapper RetimeWrapper_61 ( // @[package.scala 93:22:@43418.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  x534 x601_1 ( // @[Math.scala 366:24:@43435.4]
    .clock(x601_1_clock),
    .reset(x601_1_reset),
    .io_a(x601_1_io_a),
    .io_flow(x601_1_io_flow),
    .io_result(x601_1_io_result)
  );
  x537_div x602_div_1 ( // @[Math.scala 327:24:@43447.4]
    .clock(x602_div_1_clock),
    .reset(x602_div_1_reset),
    .io_a(x602_div_1_io_a),
    .io_flow(x602_div_1_io_flow),
    .io_result(x602_div_1_io_result)
  );
  x494_sum x603_sum_1 ( // @[Math.scala 150:24:@43457.4]
    .clock(x603_sum_1_clock),
    .reset(x603_sum_1_reset),
    .io_a(x603_sum_1_io_a),
    .io_b(x603_sum_1_io_b),
    .io_flow(x603_sum_1_io_flow),
    .io_result(x603_sum_1_io_result)
  );
  RetimeWrapper_380 RetimeWrapper_62 ( // @[package.scala 93:22:@43467.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_349 RetimeWrapper_63 ( // @[package.scala 93:22:@43476.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  RetimeWrapper_345 RetimeWrapper_64 ( // @[package.scala 93:22:@43488.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  x787_sub x606_rdrow_1 ( // @[Math.scala 191:24:@43511.4]
    .clock(x606_rdrow_1_clock),
    .reset(x606_rdrow_1_reset),
    .io_a(x606_rdrow_1_io_a),
    .io_b(x606_rdrow_1_io_b),
    .io_flow(x606_rdrow_1_io_flow),
    .io_result(x606_rdrow_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_65 ( // @[package.scala 93:22:@43528.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper RetimeWrapper_66 ( // @[package.scala 93:22:@43546.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  x494_sum x813_sum_1 ( // @[Math.scala 150:24:@43591.4]
    .clock(x813_sum_1_clock),
    .reset(x813_sum_1_reset),
    .io_a(x813_sum_1_io_a),
    .io_b(x813_sum_1_io_b),
    .io_flow(x813_sum_1_io_flow),
    .io_result(x813_sum_1_io_result)
  );
  RetimeWrapper_313 RetimeWrapper_67 ( // @[package.scala 93:22:@43601.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  x494_sum x614_sum_1 ( // @[Math.scala 150:24:@43610.4]
    .clock(x614_sum_1_clock),
    .reset(x614_sum_1_reset),
    .io_a(x614_sum_1_io_a),
    .io_b(x614_sum_1_io_b),
    .io_flow(x614_sum_1_io_flow),
    .io_result(x614_sum_1_io_result)
  );
  RetimeWrapper_300 RetimeWrapper_68 ( // @[package.scala 93:22:@43620.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_349 RetimeWrapper_69 ( // @[package.scala 93:22:@43629.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  RetimeWrapper_345 RetimeWrapper_70 ( // @[package.scala 93:22:@43641.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  x494_sum x619_sum_1 ( // @[Math.scala 150:24:@43670.4]
    .clock(x619_sum_1_clock),
    .reset(x619_sum_1_reset),
    .io_a(x619_sum_1_io_a),
    .io_b(x619_sum_1_io_b),
    .io_flow(x619_sum_1_io_flow),
    .io_result(x619_sum_1_io_result)
  );
  RetimeWrapper_349 RetimeWrapper_71 ( // @[package.scala 93:22:@43680.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  RetimeWrapper_345 RetimeWrapper_72 ( // @[package.scala 93:22:@43692.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  x494_sum x624_sum_1 ( // @[Math.scala 150:24:@43719.4]
    .clock(x624_sum_1_clock),
    .reset(x624_sum_1_reset),
    .io_a(x624_sum_1_io_a),
    .io_b(x624_sum_1_io_b),
    .io_flow(x624_sum_1_io_flow),
    .io_result(x624_sum_1_io_result)
  );
  RetimeWrapper_349 RetimeWrapper_73 ( // @[package.scala 93:22:@43729.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  RetimeWrapper_345 RetimeWrapper_74 ( // @[package.scala 93:22:@43741.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  RetimeWrapper RetimeWrapper_75 ( // @[package.scala 93:22:@43762.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_301 RetimeWrapper_76 ( // @[package.scala 93:22:@43777.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  x494_sum x629_sum_1 ( // @[Math.scala 150:24:@43786.4]
    .clock(x629_sum_1_clock),
    .reset(x629_sum_1_reset),
    .io_a(x629_sum_1_io_a),
    .io_b(x629_sum_1_io_b),
    .io_flow(x629_sum_1_io_flow),
    .io_result(x629_sum_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_77 ( // @[package.scala 93:22:@43796.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  RetimeWrapper_349 RetimeWrapper_78 ( // @[package.scala 93:22:@43805.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  RetimeWrapper_345 RetimeWrapper_79 ( // @[package.scala 93:22:@43817.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  x494_sum x634_sum_1 ( // @[Math.scala 150:24:@43844.4]
    .clock(x634_sum_1_clock),
    .reset(x634_sum_1_reset),
    .io_a(x634_sum_1_io_a),
    .io_b(x634_sum_1_io_b),
    .io_flow(x634_sum_1_io_flow),
    .io_result(x634_sum_1_io_result)
  );
  RetimeWrapper_349 RetimeWrapper_80 ( // @[package.scala 93:22:@43854.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  RetimeWrapper_345 RetimeWrapper_81 ( // @[package.scala 93:22:@43866.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  x494_sum x639_sum_1 ( // @[Math.scala 150:24:@43893.4]
    .clock(x639_sum_1_clock),
    .reset(x639_sum_1_reset),
    .io_a(x639_sum_1_io_a),
    .io_b(x639_sum_1_io_b),
    .io_flow(x639_sum_1_io_flow),
    .io_result(x639_sum_1_io_result)
  );
  RetimeWrapper_349 RetimeWrapper_82 ( // @[package.scala 93:22:@43903.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  RetimeWrapper_345 RetimeWrapper_83 ( // @[package.scala 93:22:@43915.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  x787_sub x642_rdrow_1 ( // @[Math.scala 191:24:@43938.4]
    .clock(x642_rdrow_1_clock),
    .reset(x642_rdrow_1_reset),
    .io_a(x642_rdrow_1_io_a),
    .io_b(x642_rdrow_1_io_b),
    .io_flow(x642_rdrow_1_io_flow),
    .io_result(x642_rdrow_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_84 ( // @[package.scala 93:22:@43955.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  RetimeWrapper RetimeWrapper_85 ( // @[package.scala 93:22:@43973.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  x494_sum x818_sum_1 ( // @[Math.scala 150:24:@44018.4]
    .clock(x818_sum_1_clock),
    .reset(x818_sum_1_reset),
    .io_a(x818_sum_1_io_a),
    .io_b(x818_sum_1_io_b),
    .io_flow(x818_sum_1_io_flow),
    .io_result(x818_sum_1_io_result)
  );
  RetimeWrapper_313 RetimeWrapper_86 ( // @[package.scala 93:22:@44028.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  x494_sum x650_sum_1 ( // @[Math.scala 150:24:@44037.4]
    .clock(x650_sum_1_clock),
    .reset(x650_sum_1_reset),
    .io_a(x650_sum_1_io_a),
    .io_b(x650_sum_1_io_b),
    .io_flow(x650_sum_1_io_flow),
    .io_result(x650_sum_1_io_result)
  );
  RetimeWrapper_349 RetimeWrapper_87 ( // @[package.scala 93:22:@44047.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  RetimeWrapper_300 RetimeWrapper_88 ( // @[package.scala 93:22:@44056.4]
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  RetimeWrapper_345 RetimeWrapper_89 ( // @[package.scala 93:22:@44068.4]
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  x494_sum x655_sum_1 ( // @[Math.scala 150:24:@44097.4]
    .clock(x655_sum_1_clock),
    .reset(x655_sum_1_reset),
    .io_a(x655_sum_1_io_a),
    .io_b(x655_sum_1_io_b),
    .io_flow(x655_sum_1_io_flow),
    .io_result(x655_sum_1_io_result)
  );
  RetimeWrapper_349 RetimeWrapper_90 ( // @[package.scala 93:22:@44107.4]
    .clock(RetimeWrapper_90_clock),
    .reset(RetimeWrapper_90_reset),
    .io_flow(RetimeWrapper_90_io_flow),
    .io_in(RetimeWrapper_90_io_in),
    .io_out(RetimeWrapper_90_io_out)
  );
  RetimeWrapper_345 RetimeWrapper_91 ( // @[package.scala 93:22:@44119.4]
    .clock(RetimeWrapper_91_clock),
    .reset(RetimeWrapper_91_reset),
    .io_flow(RetimeWrapper_91_io_flow),
    .io_in(RetimeWrapper_91_io_in),
    .io_out(RetimeWrapper_91_io_out)
  );
  x494_sum x660_sum_1 ( // @[Math.scala 150:24:@44146.4]
    .clock(x660_sum_1_clock),
    .reset(x660_sum_1_reset),
    .io_a(x660_sum_1_io_a),
    .io_b(x660_sum_1_io_b),
    .io_flow(x660_sum_1_io_flow),
    .io_result(x660_sum_1_io_result)
  );
  RetimeWrapper_349 RetimeWrapper_92 ( // @[package.scala 93:22:@44156.4]
    .clock(RetimeWrapper_92_clock),
    .reset(RetimeWrapper_92_reset),
    .io_flow(RetimeWrapper_92_io_flow),
    .io_in(RetimeWrapper_92_io_in),
    .io_out(RetimeWrapper_92_io_out)
  );
  RetimeWrapper_345 RetimeWrapper_93 ( // @[package.scala 93:22:@44168.4]
    .clock(RetimeWrapper_93_clock),
    .reset(RetimeWrapper_93_reset),
    .io_flow(RetimeWrapper_93_io_flow),
    .io_in(RetimeWrapper_93_io_in),
    .io_out(RetimeWrapper_93_io_out)
  );
  RetimeWrapper_301 RetimeWrapper_94 ( // @[package.scala 93:22:@44195.4]
    .clock(RetimeWrapper_94_clock),
    .reset(RetimeWrapper_94_reset),
    .io_flow(RetimeWrapper_94_io_flow),
    .io_in(RetimeWrapper_94_io_in),
    .io_out(RetimeWrapper_94_io_out)
  );
  x494_sum x665_sum_1 ( // @[Math.scala 150:24:@44204.4]
    .clock(x665_sum_1_clock),
    .reset(x665_sum_1_reset),
    .io_a(x665_sum_1_io_a),
    .io_b(x665_sum_1_io_b),
    .io_flow(x665_sum_1_io_flow),
    .io_result(x665_sum_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_95 ( // @[package.scala 93:22:@44214.4]
    .clock(RetimeWrapper_95_clock),
    .reset(RetimeWrapper_95_reset),
    .io_flow(RetimeWrapper_95_io_flow),
    .io_in(RetimeWrapper_95_io_in),
    .io_out(RetimeWrapper_95_io_out)
  );
  RetimeWrapper_349 RetimeWrapper_96 ( // @[package.scala 93:22:@44223.4]
    .clock(RetimeWrapper_96_clock),
    .reset(RetimeWrapper_96_reset),
    .io_flow(RetimeWrapper_96_io_flow),
    .io_in(RetimeWrapper_96_io_in),
    .io_out(RetimeWrapper_96_io_out)
  );
  RetimeWrapper_345 RetimeWrapper_97 ( // @[package.scala 93:22:@44235.4]
    .clock(RetimeWrapper_97_clock),
    .reset(RetimeWrapper_97_reset),
    .io_flow(RetimeWrapper_97_io_flow),
    .io_in(RetimeWrapper_97_io_in),
    .io_out(RetimeWrapper_97_io_out)
  );
  x494_sum x670_sum_1 ( // @[Math.scala 150:24:@44262.4]
    .clock(x670_sum_1_clock),
    .reset(x670_sum_1_reset),
    .io_a(x670_sum_1_io_a),
    .io_b(x670_sum_1_io_b),
    .io_flow(x670_sum_1_io_flow),
    .io_result(x670_sum_1_io_result)
  );
  RetimeWrapper_349 RetimeWrapper_98 ( // @[package.scala 93:22:@44272.4]
    .clock(RetimeWrapper_98_clock),
    .reset(RetimeWrapper_98_reset),
    .io_flow(RetimeWrapper_98_io_flow),
    .io_in(RetimeWrapper_98_io_in),
    .io_out(RetimeWrapper_98_io_out)
  );
  RetimeWrapper_345 RetimeWrapper_99 ( // @[package.scala 93:22:@44284.4]
    .clock(RetimeWrapper_99_clock),
    .reset(RetimeWrapper_99_reset),
    .io_flow(RetimeWrapper_99_io_flow),
    .io_in(RetimeWrapper_99_io_in),
    .io_out(RetimeWrapper_99_io_out)
  );
  x494_sum x675_sum_1 ( // @[Math.scala 150:24:@44311.4]
    .clock(x675_sum_1_clock),
    .reset(x675_sum_1_reset),
    .io_a(x675_sum_1_io_a),
    .io_b(x675_sum_1_io_b),
    .io_flow(x675_sum_1_io_flow),
    .io_result(x675_sum_1_io_result)
  );
  RetimeWrapper_349 RetimeWrapper_100 ( // @[package.scala 93:22:@44321.4]
    .clock(RetimeWrapper_100_clock),
    .reset(RetimeWrapper_100_reset),
    .io_flow(RetimeWrapper_100_io_flow),
    .io_in(RetimeWrapper_100_io_in),
    .io_out(RetimeWrapper_100_io_out)
  );
  RetimeWrapper_345 RetimeWrapper_101 ( // @[package.scala 93:22:@44333.4]
    .clock(RetimeWrapper_101_clock),
    .reset(RetimeWrapper_101_reset),
    .io_flow(RetimeWrapper_101_io_flow),
    .io_in(RetimeWrapper_101_io_in),
    .io_out(RetimeWrapper_101_io_out)
  );
  RetimeWrapper_57 RetimeWrapper_102 ( // @[package.scala 93:22:@44356.4]
    .clock(RetimeWrapper_102_clock),
    .reset(RetimeWrapper_102_reset),
    .io_flow(RetimeWrapper_102_io_flow),
    .io_in(RetimeWrapper_102_io_in),
    .io_out(RetimeWrapper_102_io_out)
  );
  RetimeWrapper_57 RetimeWrapper_103 ( // @[package.scala 93:22:@44368.4]
    .clock(RetimeWrapper_103_clock),
    .reset(RetimeWrapper_103_reset),
    .io_flow(RetimeWrapper_103_io_flow),
    .io_in(RetimeWrapper_103_io_in),
    .io_out(RetimeWrapper_103_io_out)
  );
  RetimeWrapper_445 RetimeWrapper_104 ( // @[package.scala 93:22:@44380.4]
    .clock(RetimeWrapper_104_clock),
    .reset(RetimeWrapper_104_reset),
    .io_flow(RetimeWrapper_104_io_flow),
    .io_in(RetimeWrapper_104_io_in),
    .io_out(RetimeWrapper_104_io_out)
  );
  RetimeWrapper_57 RetimeWrapper_105 ( // @[package.scala 93:22:@44392.4]
    .clock(RetimeWrapper_105_clock),
    .reset(RetimeWrapper_105_reset),
    .io_flow(RetimeWrapper_105_io_flow),
    .io_in(RetimeWrapper_105_io_in),
    .io_out(RetimeWrapper_105_io_out)
  );
  RetimeWrapper_57 RetimeWrapper_106 ( // @[package.scala 93:22:@44404.4]
    .clock(RetimeWrapper_106_clock),
    .reset(RetimeWrapper_106_reset),
    .io_flow(RetimeWrapper_106_io_flow),
    .io_in(RetimeWrapper_106_io_in),
    .io_out(RetimeWrapper_106_io_out)
  );
  RetimeWrapper_448 RetimeWrapper_107 ( // @[package.scala 93:22:@44414.4]
    .clock(RetimeWrapper_107_clock),
    .reset(RetimeWrapper_107_reset),
    .io_flow(RetimeWrapper_107_io_flow),
    .io_in(RetimeWrapper_107_io_in),
    .io_out(RetimeWrapper_107_io_out)
  );
  x683_x15 x683_x15_1 ( // @[Math.scala 150:24:@44423.4]
    .io_a(x683_x15_1_io_a),
    .io_b(x683_x15_1_io_b),
    .io_result(x683_x15_1_io_result)
  );
  RetimeWrapper_448 RetimeWrapper_108 ( // @[package.scala 93:22:@44433.4]
    .clock(RetimeWrapper_108_clock),
    .reset(RetimeWrapper_108_reset),
    .io_flow(RetimeWrapper_108_io_flow),
    .io_in(RetimeWrapper_108_io_in),
    .io_out(RetimeWrapper_108_io_out)
  );
  x683_x15 x684_x16_1 ( // @[Math.scala 150:24:@44442.4]
    .io_a(x684_x16_1_io_a),
    .io_b(x684_x16_1_io_b),
    .io_result(x684_x16_1_io_result)
  );
  x683_x15 x685_x15_1 ( // @[Math.scala 150:24:@44452.4]
    .io_a(x685_x15_1_io_a),
    .io_b(x685_x15_1_io_b),
    .io_result(x685_x15_1_io_result)
  );
  RetimeWrapper_448 RetimeWrapper_109 ( // @[package.scala 93:22:@44462.4]
    .clock(RetimeWrapper_109_clock),
    .reset(RetimeWrapper_109_reset),
    .io_flow(RetimeWrapper_109_io_flow),
    .io_in(RetimeWrapper_109_io_in),
    .io_out(RetimeWrapper_109_io_out)
  );
  x683_x15 x686_x16_1 ( // @[Math.scala 150:24:@44471.4]
    .io_a(x686_x16_1_io_a),
    .io_b(x686_x16_1_io_b),
    .io_result(x686_x16_1_io_result)
  );
  x683_x15 x687_x15_1 ( // @[Math.scala 150:24:@44481.4]
    .io_a(x687_x15_1_io_a),
    .io_b(x687_x15_1_io_b),
    .io_result(x687_x15_1_io_result)
  );
  x683_x15 x688_x16_1 ( // @[Math.scala 150:24:@44491.4]
    .io_a(x688_x16_1_io_a),
    .io_b(x688_x16_1_io_b),
    .io_result(x688_x16_1_io_result)
  );
  x683_x15 x689_x15_1 ( // @[Math.scala 150:24:@44503.4]
    .io_a(x689_x15_1_io_a),
    .io_b(x689_x15_1_io_b),
    .io_result(x689_x15_1_io_result)
  );
  RetimeWrapper_448 RetimeWrapper_110 ( // @[package.scala 93:22:@44513.4]
    .clock(RetimeWrapper_110_clock),
    .reset(RetimeWrapper_110_reset),
    .io_flow(RetimeWrapper_110_io_flow),
    .io_in(RetimeWrapper_110_io_in),
    .io_out(RetimeWrapper_110_io_out)
  );
  x690_sum x690_sum_1 ( // @[Math.scala 150:24:@44522.4]
    .clock(x690_sum_1_clock),
    .reset(x690_sum_1_reset),
    .io_a(x690_sum_1_io_a),
    .io_b(x690_sum_1_io_b),
    .io_flow(x690_sum_1_io_flow),
    .io_result(x690_sum_1_io_result)
  );
  RetimeWrapper_57 RetimeWrapper_111 ( // @[package.scala 93:22:@44541.4]
    .clock(RetimeWrapper_111_clock),
    .reset(RetimeWrapper_111_reset),
    .io_flow(RetimeWrapper_111_io_flow),
    .io_in(RetimeWrapper_111_io_in),
    .io_out(RetimeWrapper_111_io_out)
  );
  RetimeWrapper_57 RetimeWrapper_112 ( // @[package.scala 93:22:@44553.4]
    .clock(RetimeWrapper_112_clock),
    .reset(RetimeWrapper_112_reset),
    .io_flow(RetimeWrapper_112_io_flow),
    .io_in(RetimeWrapper_112_io_in),
    .io_out(RetimeWrapper_112_io_out)
  );
  RetimeWrapper_445 RetimeWrapper_113 ( // @[package.scala 93:22:@44565.4]
    .clock(RetimeWrapper_113_clock),
    .reset(RetimeWrapper_113_reset),
    .io_flow(RetimeWrapper_113_io_flow),
    .io_in(RetimeWrapper_113_io_in),
    .io_out(RetimeWrapper_113_io_out)
  );
  RetimeWrapper_57 RetimeWrapper_114 ( // @[package.scala 93:22:@44577.4]
    .clock(RetimeWrapper_114_clock),
    .reset(RetimeWrapper_114_reset),
    .io_flow(RetimeWrapper_114_io_flow),
    .io_in(RetimeWrapper_114_io_in),
    .io_out(RetimeWrapper_114_io_out)
  );
  RetimeWrapper_57 RetimeWrapper_115 ( // @[package.scala 93:22:@44589.4]
    .clock(RetimeWrapper_115_clock),
    .reset(RetimeWrapper_115_reset),
    .io_flow(RetimeWrapper_115_io_flow),
    .io_in(RetimeWrapper_115_io_in),
    .io_out(RetimeWrapper_115_io_out)
  );
  RetimeWrapper_448 RetimeWrapper_116 ( // @[package.scala 93:22:@44599.4]
    .clock(RetimeWrapper_116_clock),
    .reset(RetimeWrapper_116_reset),
    .io_flow(RetimeWrapper_116_io_flow),
    .io_in(RetimeWrapper_116_io_in),
    .io_out(RetimeWrapper_116_io_out)
  );
  x683_x15 x697_x15_1 ( // @[Math.scala 150:24:@44608.4]
    .io_a(x697_x15_1_io_a),
    .io_b(x697_x15_1_io_b),
    .io_result(x697_x15_1_io_result)
  );
  RetimeWrapper_448 RetimeWrapper_117 ( // @[package.scala 93:22:@44618.4]
    .clock(RetimeWrapper_117_clock),
    .reset(RetimeWrapper_117_reset),
    .io_flow(RetimeWrapper_117_io_flow),
    .io_in(RetimeWrapper_117_io_in),
    .io_out(RetimeWrapper_117_io_out)
  );
  x683_x15 x698_x16_1 ( // @[Math.scala 150:24:@44627.4]
    .io_a(x698_x16_1_io_a),
    .io_b(x698_x16_1_io_b),
    .io_result(x698_x16_1_io_result)
  );
  x683_x15 x699_x15_1 ( // @[Math.scala 150:24:@44637.4]
    .io_a(x699_x15_1_io_a),
    .io_b(x699_x15_1_io_b),
    .io_result(x699_x15_1_io_result)
  );
  RetimeWrapper_448 RetimeWrapper_118 ( // @[package.scala 93:22:@44647.4]
    .clock(RetimeWrapper_118_clock),
    .reset(RetimeWrapper_118_reset),
    .io_flow(RetimeWrapper_118_io_flow),
    .io_in(RetimeWrapper_118_io_in),
    .io_out(RetimeWrapper_118_io_out)
  );
  x683_x15 x700_x16_1 ( // @[Math.scala 150:24:@44656.4]
    .io_a(x700_x16_1_io_a),
    .io_b(x700_x16_1_io_b),
    .io_result(x700_x16_1_io_result)
  );
  x683_x15 x701_x15_1 ( // @[Math.scala 150:24:@44666.4]
    .io_a(x701_x15_1_io_a),
    .io_b(x701_x15_1_io_b),
    .io_result(x701_x15_1_io_result)
  );
  x683_x15 x702_x16_1 ( // @[Math.scala 150:24:@44676.4]
    .io_a(x702_x16_1_io_a),
    .io_b(x702_x16_1_io_b),
    .io_result(x702_x16_1_io_result)
  );
  x683_x15 x703_x15_1 ( // @[Math.scala 150:24:@44686.4]
    .io_a(x703_x15_1_io_a),
    .io_b(x703_x15_1_io_b),
    .io_result(x703_x15_1_io_result)
  );
  RetimeWrapper_448 RetimeWrapper_119 ( // @[package.scala 93:22:@44696.4]
    .clock(RetimeWrapper_119_clock),
    .reset(RetimeWrapper_119_reset),
    .io_flow(RetimeWrapper_119_io_flow),
    .io_in(RetimeWrapper_119_io_in),
    .io_out(RetimeWrapper_119_io_out)
  );
  x690_sum x704_sum_1 ( // @[Math.scala 150:24:@44705.4]
    .clock(x704_sum_1_clock),
    .reset(x704_sum_1_reset),
    .io_a(x704_sum_1_io_a),
    .io_b(x704_sum_1_io_b),
    .io_flow(x704_sum_1_io_flow),
    .io_result(x704_sum_1_io_result)
  );
  RetimeWrapper_57 RetimeWrapper_120 ( // @[package.scala 93:22:@44724.4]
    .clock(RetimeWrapper_120_clock),
    .reset(RetimeWrapper_120_reset),
    .io_flow(RetimeWrapper_120_io_flow),
    .io_in(RetimeWrapper_120_io_in),
    .io_out(RetimeWrapper_120_io_out)
  );
  RetimeWrapper_445 RetimeWrapper_121 ( // @[package.scala 93:22:@44736.4]
    .clock(RetimeWrapper_121_clock),
    .reset(RetimeWrapper_121_reset),
    .io_flow(RetimeWrapper_121_io_flow),
    .io_in(RetimeWrapper_121_io_in),
    .io_out(RetimeWrapper_121_io_out)
  );
  RetimeWrapper_57 RetimeWrapper_122 ( // @[package.scala 93:22:@44748.4]
    .clock(RetimeWrapper_122_clock),
    .reset(RetimeWrapper_122_reset),
    .io_flow(RetimeWrapper_122_io_flow),
    .io_in(RetimeWrapper_122_io_in),
    .io_out(RetimeWrapper_122_io_out)
  );
  RetimeWrapper_57 RetimeWrapper_123 ( // @[package.scala 93:22:@44760.4]
    .clock(RetimeWrapper_123_clock),
    .reset(RetimeWrapper_123_reset),
    .io_flow(RetimeWrapper_123_io_flow),
    .io_in(RetimeWrapper_123_io_in),
    .io_out(RetimeWrapper_123_io_out)
  );
  x683_x15 x710_x15_1 ( // @[Math.scala 150:24:@44770.4]
    .io_a(x710_x15_1_io_a),
    .io_b(x710_x15_1_io_b),
    .io_result(x710_x15_1_io_result)
  );
  RetimeWrapper_448 RetimeWrapper_124 ( // @[package.scala 93:22:@44780.4]
    .clock(RetimeWrapper_124_clock),
    .reset(RetimeWrapper_124_reset),
    .io_flow(RetimeWrapper_124_io_flow),
    .io_in(RetimeWrapper_124_io_in),
    .io_out(RetimeWrapper_124_io_out)
  );
  x683_x15 x711_x16_1 ( // @[Math.scala 150:24:@44789.4]
    .io_a(x711_x16_1_io_a),
    .io_b(x711_x16_1_io_b),
    .io_result(x711_x16_1_io_result)
  );
  x683_x15 x712_x15_1 ( // @[Math.scala 150:24:@44799.4]
    .io_a(x712_x15_1_io_a),
    .io_b(x712_x15_1_io_b),
    .io_result(x712_x15_1_io_result)
  );
  x683_x15 x713_x16_1 ( // @[Math.scala 150:24:@44809.4]
    .io_a(x713_x16_1_io_a),
    .io_b(x713_x16_1_io_b),
    .io_result(x713_x16_1_io_result)
  );
  x683_x15 x714_x15_1 ( // @[Math.scala 150:24:@44819.4]
    .io_a(x714_x15_1_io_a),
    .io_b(x714_x15_1_io_b),
    .io_result(x714_x15_1_io_result)
  );
  x683_x15 x715_x16_1 ( // @[Math.scala 150:24:@44829.4]
    .io_a(x715_x16_1_io_a),
    .io_b(x715_x16_1_io_b),
    .io_result(x715_x16_1_io_result)
  );
  x683_x15 x716_x15_1 ( // @[Math.scala 150:24:@44839.4]
    .io_a(x716_x15_1_io_a),
    .io_b(x716_x15_1_io_b),
    .io_result(x716_x15_1_io_result)
  );
  RetimeWrapper_448 RetimeWrapper_125 ( // @[package.scala 93:22:@44849.4]
    .clock(RetimeWrapper_125_clock),
    .reset(RetimeWrapper_125_reset),
    .io_flow(RetimeWrapper_125_io_flow),
    .io_in(RetimeWrapper_125_io_in),
    .io_out(RetimeWrapper_125_io_out)
  );
  x690_sum x717_sum_1 ( // @[Math.scala 150:24:@44858.4]
    .clock(x717_sum_1_clock),
    .reset(x717_sum_1_reset),
    .io_a(x717_sum_1_io_a),
    .io_b(x717_sum_1_io_b),
    .io_flow(x717_sum_1_io_flow),
    .io_result(x717_sum_1_io_result)
  );
  RetimeWrapper_57 RetimeWrapper_126 ( // @[package.scala 93:22:@44877.4]
    .clock(RetimeWrapper_126_clock),
    .reset(RetimeWrapper_126_reset),
    .io_flow(RetimeWrapper_126_io_flow),
    .io_in(RetimeWrapper_126_io_in),
    .io_out(RetimeWrapper_126_io_out)
  );
  RetimeWrapper_445 RetimeWrapper_127 ( // @[package.scala 93:22:@44889.4]
    .clock(RetimeWrapper_127_clock),
    .reset(RetimeWrapper_127_reset),
    .io_flow(RetimeWrapper_127_io_flow),
    .io_in(RetimeWrapper_127_io_in),
    .io_out(RetimeWrapper_127_io_out)
  );
  RetimeWrapper_57 RetimeWrapper_128 ( // @[package.scala 93:22:@44901.4]
    .clock(RetimeWrapper_128_clock),
    .reset(RetimeWrapper_128_reset),
    .io_flow(RetimeWrapper_128_io_flow),
    .io_in(RetimeWrapper_128_io_in),
    .io_out(RetimeWrapper_128_io_out)
  );
  RetimeWrapper_57 RetimeWrapper_129 ( // @[package.scala 93:22:@44913.4]
    .clock(RetimeWrapper_129_clock),
    .reset(RetimeWrapper_129_reset),
    .io_flow(RetimeWrapper_129_io_flow),
    .io_in(RetimeWrapper_129_io_in),
    .io_out(RetimeWrapper_129_io_out)
  );
  x683_x15 x723_x15_1 ( // @[Math.scala 150:24:@44923.4]
    .io_a(x723_x15_1_io_a),
    .io_b(x723_x15_1_io_b),
    .io_result(x723_x15_1_io_result)
  );
  RetimeWrapper_448 RetimeWrapper_130 ( // @[package.scala 93:22:@44933.4]
    .clock(RetimeWrapper_130_clock),
    .reset(RetimeWrapper_130_reset),
    .io_flow(RetimeWrapper_130_io_flow),
    .io_in(RetimeWrapper_130_io_in),
    .io_out(RetimeWrapper_130_io_out)
  );
  x683_x15 x724_x16_1 ( // @[Math.scala 150:24:@44942.4]
    .io_a(x724_x16_1_io_a),
    .io_b(x724_x16_1_io_b),
    .io_result(x724_x16_1_io_result)
  );
  x683_x15 x725_x15_1 ( // @[Math.scala 150:24:@44952.4]
    .io_a(x725_x15_1_io_a),
    .io_b(x725_x15_1_io_b),
    .io_result(x725_x15_1_io_result)
  );
  x683_x15 x726_x16_1 ( // @[Math.scala 150:24:@44962.4]
    .io_a(x726_x16_1_io_a),
    .io_b(x726_x16_1_io_b),
    .io_result(x726_x16_1_io_result)
  );
  x683_x15 x727_x15_1 ( // @[Math.scala 150:24:@44972.4]
    .io_a(x727_x15_1_io_a),
    .io_b(x727_x15_1_io_b),
    .io_result(x727_x15_1_io_result)
  );
  x683_x15 x728_x16_1 ( // @[Math.scala 150:24:@44982.4]
    .io_a(x728_x16_1_io_a),
    .io_b(x728_x16_1_io_b),
    .io_result(x728_x16_1_io_result)
  );
  x683_x15 x729_x15_1 ( // @[Math.scala 150:24:@44992.4]
    .io_a(x729_x15_1_io_a),
    .io_b(x729_x15_1_io_b),
    .io_result(x729_x15_1_io_result)
  );
  RetimeWrapper_448 RetimeWrapper_131 ( // @[package.scala 93:22:@45002.4]
    .clock(RetimeWrapper_131_clock),
    .reset(RetimeWrapper_131_reset),
    .io_flow(RetimeWrapper_131_io_flow),
    .io_in(RetimeWrapper_131_io_in),
    .io_out(RetimeWrapper_131_io_out)
  );
  x690_sum x730_sum_1 ( // @[Math.scala 150:24:@45013.4]
    .clock(x730_sum_1_clock),
    .reset(x730_sum_1_reset),
    .io_a(x730_sum_1_io_a),
    .io_b(x730_sum_1_io_b),
    .io_flow(x730_sum_1_io_flow),
    .io_result(x730_sum_1_io_result)
  );
  RetimeWrapper_303 RetimeWrapper_132 ( // @[package.scala 93:22:@45040.4]
    .clock(RetimeWrapper_132_clock),
    .reset(RetimeWrapper_132_reset),
    .io_flow(RetimeWrapper_132_io_flow),
    .io_in(RetimeWrapper_132_io_in),
    .io_out(RetimeWrapper_132_io_out)
  );
  RetimeWrapper_48 RetimeWrapper_133 ( // @[package.scala 93:22:@45049.4]
    .clock(RetimeWrapper_133_clock),
    .reset(RetimeWrapper_133_reset),
    .io_flow(RetimeWrapper_133_io_flow),
    .io_in(RetimeWrapper_133_io_in),
    .io_out(RetimeWrapper_133_io_out)
  );
  RetimeWrapper_48 RetimeWrapper_134 ( // @[package.scala 93:22:@45058.4]
    .clock(RetimeWrapper_134_clock),
    .reset(RetimeWrapper_134_reset),
    .io_flow(RetimeWrapper_134_io_flow),
    .io_in(RetimeWrapper_134_io_in),
    .io_out(RetimeWrapper_134_io_out)
  );
  RetimeWrapper_48 RetimeWrapper_135 ( // @[package.scala 93:22:@45067.4]
    .clock(RetimeWrapper_135_clock),
    .reset(RetimeWrapper_135_reset),
    .io_flow(RetimeWrapper_135_io_flow),
    .io_in(RetimeWrapper_135_io_in),
    .io_out(RetimeWrapper_135_io_out)
  );
  assign b521 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 62:18:@42080.4]
  assign b522 = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 63:18:@42081.4]
  assign _T_205 = b521 & b522; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 67:30:@42083.4]
  assign _T_206 = _T_205 & io_sigsIn_datapathEn; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 67:37:@42084.4]
  assign _T_210 = io_in_x480_TID == 8'h0; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 69:76:@42089.4]
  assign _T_211 = _T_206 & _T_210; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 69:62:@42090.4]
  assign _T_213 = io_in_x480_TDEST == 8'h0; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 69:101:@42091.4]
  assign x824_x523_D1_0_number = RetimeWrapper_io_out; // @[package.scala 96:25:@42100.4 package.scala 96:25:@42101.4]
  assign b519_number = __io_result; // @[Math.scala 712:22:@42065.4 Math.scala 713:14:@42066.4]
  assign _T_246 = $signed(b519_number); // @[Math.scala 499:52:@42265.4]
  assign x528 = $signed(32'sh1) == $signed(_T_246); // @[Math.scala 499:44:@42273.4]
  assign x529 = $signed(32'sh2) == $signed(_T_246); // @[Math.scala 499:44:@42280.4]
  assign x530 = $signed(32'sh3) == $signed(_T_246); // @[Math.scala 499:44:@42287.4]
  assign _T_293 = x528 ? 32'h1 : 32'h0; // @[Mux.scala 19:72:@42299.4]
  assign _T_295 = x529 ? 32'h2 : 32'h0; // @[Mux.scala 19:72:@42300.4]
  assign _T_297 = x530 ? 32'h3 : 32'h0; // @[Mux.scala 19:72:@42301.4]
  assign _T_299 = _T_293 | _T_295; // @[Mux.scala 19:72:@42303.4]
  assign x825_x531_D2_number = RetimeWrapper_1_io_out; // @[package.scala 96:25:@42316.4 package.scala 96:25:@42317.4]
  assign _T_314 = $signed(x825_x531_D2_number); // @[Math.scala 406:49:@42323.4]
  assign _T_316 = $signed(_T_314) & $signed(32'sh3); // @[Math.scala 406:56:@42325.4]
  assign _T_317 = $signed(_T_316); // @[Math.scala 406:56:@42326.4]
  assign _T_329 = x825_x531_D2_number[31]; // @[FixedPoint.scala 50:25:@42344.4]
  assign _T_333 = _T_329 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@42346.4]
  assign _T_334 = x825_x531_D2_number[31:2]; // @[FixedPoint.scala 18:52:@42347.4]
  assign x535_number = {_T_333,_T_334}; // @[Cat.scala 30:58:@42348.4]
  assign _GEN_0 = {{8'd0}, x535_number}; // @[Math.scala 450:32:@42353.4]
  assign _T_339 = _GEN_0 << 8; // @[Math.scala 450:32:@42353.4]
  assign _GEN_1 = {{6'd0}, x535_number}; // @[Math.scala 450:32:@42358.4]
  assign _T_343 = _GEN_1 << 6; // @[Math.scala 450:32:@42358.4]
  assign _T_379 = ~ io_sigsIn_break; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 127:101:@42456.4]
  assign _T_383 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@42464.4 package.scala 96:25:@42465.4]
  assign _T_385 = io_rr ? _T_383 : 1'h0; // @[implicits.scala 55:10:@42466.4]
  assign _T_386 = _T_379 & _T_385; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 127:118:@42467.4]
  assign _T_388 = _T_386 & _T_379; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 127:207:@42469.4]
  assign _T_389 = _T_388 & io_sigsIn_backpressure; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 127:226:@42470.4]
  assign x830_b521_D24 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@42435.4 package.scala 96:25:@42436.4]
  assign _T_390 = _T_389 & x830_b521_D24; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 127:252:@42471.4]
  assign x829_b522_D24 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@42426.4 package.scala 96:25:@42427.4]
  assign _T_434 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@42571.4 package.scala 96:25:@42572.4]
  assign _T_436 = io_rr ? _T_434 : 1'h0; // @[implicits.scala 55:10:@42573.4]
  assign _T_437 = _T_379 & _T_436; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 150:118:@42574.4]
  assign _T_439 = _T_437 & _T_379; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 150:207:@42576.4]
  assign _T_440 = _T_439 & io_sigsIn_backpressure; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 150:226:@42577.4]
  assign _T_441 = _T_440 & x830_b521_D24; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 150:252:@42578.4]
  assign _T_482 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@42669.4 package.scala 96:25:@42670.4]
  assign _T_484 = io_rr ? _T_482 : 1'h0; // @[implicits.scala 55:10:@42671.4]
  assign _T_485 = _T_379 & _T_484; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 171:118:@42672.4]
  assign _T_487 = _T_485 & _T_379; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 171:207:@42674.4]
  assign _T_488 = _T_487 & io_sigsIn_backpressure; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 171:226:@42675.4]
  assign _T_489 = _T_488 & x830_b521_D24; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 171:252:@42676.4]
  assign _T_532 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@42769.4 package.scala 96:25:@42770.4]
  assign _T_534 = io_rr ? _T_532 : 1'h0; // @[implicits.scala 55:10:@42771.4]
  assign _T_535 = _T_379 & _T_534; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 200:166:@42772.4]
  assign _T_537 = _T_535 & _T_379; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 200:255:@42774.4]
  assign _T_538 = _T_537 & io_sigsIn_backpressure; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 200:274:@42775.4]
  assign _T_539 = _T_538 & x830_b521_D24; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 200:300:@42776.4]
  assign x843_b519_D26_number = RetimeWrapper_23_io_out; // @[package.scala 96:25:@42790.4 package.scala 96:25:@42791.4]
  assign _T_551 = $signed(x843_b519_D26_number); // @[Math.scala 406:49:@42797.4]
  assign _T_553 = $signed(_T_551) & $signed(32'sh3); // @[Math.scala 406:56:@42799.4]
  assign _T_554 = $signed(_T_553); // @[Math.scala 406:56:@42800.4]
  assign _T_558 = $signed(RetimeWrapper_24_io_out); // @[package.scala 96:25:@42808.4]
  assign x804_number = $unsigned(_T_558); // @[implicits.scala 133:21:@42810.4]
  assign x844_x552_rdcol_D26_number = RetimeWrapper_26_io_out; // @[package.scala 96:25:@42833.4 package.scala 96:25:@42834.4]
  assign _T_578 = $signed(x844_x552_rdcol_D26_number); // @[Math.scala 465:37:@42839.4]
  assign x845_x560_D1 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@42856.4 package.scala 96:25:@42857.4]
  assign x561 = RetimeWrapper_27_io_out; // @[package.scala 96:25:@42847.4 package.scala 96:25:@42848.4]
  assign x562 = x845_x560_D1 | x561; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 215:24:@42860.4]
  assign _T_597 = $signed(x804_number); // @[Math.scala 406:49:@42869.4]
  assign _T_599 = $signed(_T_597) & $signed(32'sh3); // @[Math.scala 406:56:@42871.4]
  assign _T_600 = $signed(_T_599); // @[Math.scala 406:56:@42872.4]
  assign _T_605 = x804_number[31]; // @[FixedPoint.scala 50:25:@42878.4]
  assign _T_609 = _T_605 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@42880.4]
  assign _T_610 = x804_number[31:2]; // @[FixedPoint.scala 18:52:@42881.4]
  assign x565_number = {_T_609,_T_610}; // @[Cat.scala 30:58:@42882.4]
  assign _GEN_2 = {{8'd0}, x565_number}; // @[Math.scala 450:32:@42887.4]
  assign _T_615 = _GEN_2 << 8; // @[Math.scala 450:32:@42887.4]
  assign _GEN_3 = {{6'd0}, x565_number}; // @[Math.scala 450:32:@42892.4]
  assign _T_619 = _GEN_3 << 6; // @[Math.scala 450:32:@42892.4]
  assign _T_658 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@42987.4 package.scala 96:25:@42988.4]
  assign _T_660 = io_rr ? _T_658 : 1'h0; // @[implicits.scala 55:10:@42989.4]
  assign _T_661 = _T_379 & _T_660; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 248:194:@42990.4]
  assign x852_x563_D20 = RetimeWrapper_35_io_out; // @[package.scala 96:25:@42975.4 package.scala 96:25:@42976.4]
  assign _T_662 = _T_661 & x852_x563_D20; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 248:283:@42991.4]
  assign x851_b521_D48 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@42966.4 package.scala 96:25:@42967.4]
  assign _T_663 = _T_662 & x851_b521_D48; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 248:291:@42992.4]
  assign x848_b522_D48 = RetimeWrapper_31_io_out; // @[package.scala 96:25:@42939.4 package.scala 96:25:@42940.4]
  assign x853_x546_rdcol_D26_number = RetimeWrapper_37_io_out; // @[package.scala 96:25:@43008.4 package.scala 96:25:@43009.4]
  assign _T_674 = $signed(x853_x546_rdcol_D26_number); // @[Math.scala 465:37:@43014.4]
  assign x570 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@43022.4 package.scala 96:25:@43023.4]
  assign x571 = x845_x560_D1 | x570; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 256:24:@43026.4]
  assign _T_706 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@43077.4 package.scala 96:25:@43078.4]
  assign _T_708 = io_rr ? _T_706 : 1'h0; // @[implicits.scala 55:10:@43079.4]
  assign _T_709 = _T_379 & _T_708; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 271:194:@43080.4]
  assign x855_x572_D20 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@43056.4 package.scala 96:25:@43057.4]
  assign _T_710 = _T_709 & x855_x572_D20; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 271:283:@43081.4]
  assign _T_711 = _T_710 & x851_b521_D48; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 271:291:@43082.4]
  assign x857_x540_rdcol_D26_number = RetimeWrapper_43_io_out; // @[package.scala 96:25:@43098.4 package.scala 96:25:@43099.4]
  assign _T_722 = $signed(x857_x540_rdcol_D26_number); // @[Math.scala 465:37:@43104.4]
  assign x576 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@43112.4 package.scala 96:25:@43113.4]
  assign x577 = x845_x560_D1 | x576; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 279:24:@43116.4]
  assign _T_754 = RetimeWrapper_48_io_out; // @[package.scala 96:25:@43167.4 package.scala 96:25:@43168.4]
  assign _T_756 = io_rr ? _T_754 : 1'h0; // @[implicits.scala 55:10:@43169.4]
  assign _T_757 = _T_379 & _T_756; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 300:194:@43170.4]
  assign x860_x578_D20 = RetimeWrapper_47_io_out; // @[package.scala 96:25:@43155.4 package.scala 96:25:@43156.4]
  assign _T_758 = _T_757 & x860_x578_D20; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 300:283:@43171.4]
  assign _T_759 = _T_758 & x851_b521_D48; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 300:326:@43172.4]
  assign x861_b520_D26_number = RetimeWrapper_49_io_out; // @[package.scala 96:25:@43188.4 package.scala 96:25:@43189.4]
  assign _T_772 = $signed(x861_b520_D26_number); // @[Math.scala 465:37:@43196.4]
  assign x560 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@42824.4 package.scala 96:25:@42825.4]
  assign x582 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@43204.4 package.scala 96:25:@43205.4]
  assign x583 = x560 | x582; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 310:59:@43208.4]
  assign _T_810 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@43277.4 package.scala 96:25:@43278.4]
  assign _T_812 = io_rr ? _T_810 : 1'h0; // @[implicits.scala 55:10:@43279.4]
  assign _T_813 = _T_379 & _T_812; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 329:194:@43280.4]
  assign x865_x584_D21 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@43256.4 package.scala 96:25:@43257.4]
  assign _T_814 = _T_813 & x865_x584_D21; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 329:283:@43281.4]
  assign _T_815 = _T_814 & x851_b521_D48; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 329:291:@43282.4]
  assign x588_rdcol_number = x588_rdcol_1_io_result; // @[Math.scala 154:22:@43301.4 Math.scala 155:14:@43302.4]
  assign _T_830 = $signed(x588_rdcol_number); // @[Math.scala 465:37:@43307.4]
  assign x589 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@43315.4 package.scala 96:25:@43316.4]
  assign x590 = x845_x560_D1 | x589; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 337:59:@43319.4]
  assign _T_873 = RetimeWrapper_60_io_out; // @[package.scala 96:25:@43385.4 package.scala 96:25:@43386.4]
  assign _T_875 = io_rr ? _T_873 : 1'h0; // @[implicits.scala 55:10:@43387.4]
  assign _T_876 = _T_379 & _T_875; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 354:194:@43388.4]
  assign x867_x591_D20 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@43364.4 package.scala 96:25:@43365.4]
  assign _T_877 = _T_876 & x867_x591_D20; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 354:283:@43389.4]
  assign _T_878 = _T_877 & x851_b521_D48; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 354:291:@43390.4]
  assign x597_rdcol_number = x597_rdcol_1_io_result; // @[Math.scala 154:22:@43409.4 Math.scala 155:14:@43410.4]
  assign _T_893 = $signed(x597_rdcol_number); // @[Math.scala 465:37:@43415.4]
  assign x598 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@43423.4 package.scala 96:25:@43424.4]
  assign x599 = x845_x560_D1 | x598; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 362:59:@43427.4]
  assign _T_936 = RetimeWrapper_64_io_out; // @[package.scala 96:25:@43493.4 package.scala 96:25:@43494.4]
  assign _T_938 = io_rr ? _T_936 : 1'h0; // @[implicits.scala 55:10:@43495.4]
  assign _T_939 = _T_379 & _T_938; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 379:194:@43496.4]
  assign x870_x600_D20 = RetimeWrapper_63_io_out; // @[package.scala 96:25:@43481.4 package.scala 96:25:@43482.4]
  assign _T_940 = _T_939 & x870_x600_D20; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 379:283:@43497.4]
  assign _T_941 = _T_940 & x851_b521_D48; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 379:291:@43498.4]
  assign x606_rdrow_number = x606_rdrow_1_io_result; // @[Math.scala 195:22:@43517.4 Math.scala 196:14:@43518.4]
  assign _T_958 = $signed(x606_rdrow_number); // @[Math.scala 406:49:@43524.4]
  assign _T_960 = $signed(_T_958) & $signed(32'sh3); // @[Math.scala 406:56:@43526.4]
  assign _T_961 = $signed(_T_960); // @[Math.scala 406:56:@43527.4]
  assign _T_965 = $signed(RetimeWrapper_65_io_out); // @[package.scala 96:25:@43535.4]
  assign x809_number = $unsigned(_T_965); // @[implicits.scala 133:21:@43537.4]
  assign x608 = RetimeWrapper_66_io_out; // @[package.scala 96:25:@43551.4 package.scala 96:25:@43552.4]
  assign x609 = x608 | x561; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 389:24:@43555.4]
  assign _T_988 = $signed(x809_number); // @[Math.scala 406:49:@43564.4]
  assign _T_990 = $signed(_T_988) & $signed(32'sh3); // @[Math.scala 406:56:@43566.4]
  assign _T_991 = $signed(_T_990); // @[Math.scala 406:56:@43567.4]
  assign _T_996 = x809_number[31]; // @[FixedPoint.scala 50:25:@43573.4]
  assign _T_1000 = _T_996 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@43575.4]
  assign _T_1001 = x809_number[31:2]; // @[FixedPoint.scala 18:52:@43576.4]
  assign x612_number = {_T_1000,_T_1001}; // @[Cat.scala 30:58:@43577.4]
  assign _GEN_4 = {{8'd0}, x612_number}; // @[Math.scala 450:32:@43582.4]
  assign _T_1006 = _GEN_4 << 8; // @[Math.scala 450:32:@43582.4]
  assign _GEN_5 = {{6'd0}, x612_number}; // @[Math.scala 450:32:@43587.4]
  assign _T_1010 = _GEN_5 << 6; // @[Math.scala 450:32:@43587.4]
  assign _T_1037 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@43646.4 package.scala 96:25:@43647.4]
  assign _T_1039 = io_rr ? _T_1037 : 1'h0; // @[implicits.scala 55:10:@43648.4]
  assign _T_1040 = _T_379 & _T_1039; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 420:194:@43649.4]
  assign x873_x610_D20 = RetimeWrapper_69_io_out; // @[package.scala 96:25:@43634.4 package.scala 96:25:@43635.4]
  assign _T_1041 = _T_1040 & x873_x610_D20; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 420:283:@43650.4]
  assign _T_1042 = _T_1041 & x851_b521_D48; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 420:291:@43651.4]
  assign x617 = x608 | x570; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 424:59:@43662.4]
  assign _T_1068 = RetimeWrapper_72_io_out; // @[package.scala 96:25:@43697.4 package.scala 96:25:@43698.4]
  assign _T_1070 = io_rr ? _T_1068 : 1'h0; // @[implicits.scala 55:10:@43699.4]
  assign _T_1071 = _T_379 & _T_1070; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 437:194:@43700.4]
  assign x874_x618_D20 = RetimeWrapper_71_io_out; // @[package.scala 96:25:@43685.4 package.scala 96:25:@43686.4]
  assign _T_1072 = _T_1071 & x874_x618_D20; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 437:283:@43701.4]
  assign _T_1073 = _T_1072 & x851_b521_D48; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 437:291:@43702.4]
  assign x622 = x608 | x576; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 441:59:@43713.4]
  assign _T_1097 = RetimeWrapper_74_io_out; // @[package.scala 96:25:@43746.4 package.scala 96:25:@43747.4]
  assign _T_1099 = io_rr ? _T_1097 : 1'h0; // @[implicits.scala 55:10:@43748.4]
  assign _T_1100 = _T_379 & _T_1099; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 452:194:@43749.4]
  assign x875_x623_D20 = RetimeWrapper_73_io_out; // @[package.scala 96:25:@43734.4 package.scala 96:25:@43735.4]
  assign _T_1101 = _T_1100 & x875_x623_D20; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 452:283:@43750.4]
  assign _T_1102 = _T_1101 & x851_b521_D48; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 452:291:@43751.4]
  assign x876_x582_D1 = RetimeWrapper_75_io_out; // @[package.scala 96:25:@43767.4 package.scala 96:25:@43768.4]
  assign x627 = x608 | x876_x582_D1; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 458:59:@43771.4]
  assign _T_1135 = RetimeWrapper_79_io_out; // @[package.scala 96:25:@43822.4 package.scala 96:25:@43823.4]
  assign _T_1137 = io_rr ? _T_1135 : 1'h0; // @[implicits.scala 55:10:@43824.4]
  assign _T_1138 = _T_379 & _T_1137; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 473:194:@43825.4]
  assign x879_x628_D20 = RetimeWrapper_78_io_out; // @[package.scala 96:25:@43810.4 package.scala 96:25:@43811.4]
  assign _T_1139 = _T_1138 & x879_x628_D20; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 473:283:@43826.4]
  assign _T_1140 = _T_1139 & x851_b521_D48; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 473:291:@43827.4]
  assign x632 = x608 | x589; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 477:59:@43838.4]
  assign _T_1164 = RetimeWrapper_81_io_out; // @[package.scala 96:25:@43871.4 package.scala 96:25:@43872.4]
  assign _T_1166 = io_rr ? _T_1164 : 1'h0; // @[implicits.scala 55:10:@43873.4]
  assign _T_1167 = _T_379 & _T_1166; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 488:194:@43874.4]
  assign x880_x633_D20 = RetimeWrapper_80_io_out; // @[package.scala 96:25:@43859.4 package.scala 96:25:@43860.4]
  assign _T_1168 = _T_1167 & x880_x633_D20; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 488:283:@43875.4]
  assign _T_1169 = _T_1168 & x851_b521_D48; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 488:291:@43876.4]
  assign x637 = x608 | x598; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 492:59:@43887.4]
  assign _T_1193 = RetimeWrapper_83_io_out; // @[package.scala 96:25:@43920.4 package.scala 96:25:@43921.4]
  assign _T_1195 = io_rr ? _T_1193 : 1'h0; // @[implicits.scala 55:10:@43922.4]
  assign _T_1196 = _T_379 & _T_1195; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 503:194:@43923.4]
  assign x881_x638_D20 = RetimeWrapper_82_io_out; // @[package.scala 96:25:@43908.4 package.scala 96:25:@43909.4]
  assign _T_1197 = _T_1196 & x881_x638_D20; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 503:283:@43924.4]
  assign _T_1198 = _T_1197 & x851_b521_D48; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 503:291:@43925.4]
  assign x642_rdrow_number = x642_rdrow_1_io_result; // @[Math.scala 195:22:@43944.4 Math.scala 196:14:@43945.4]
  assign _T_1215 = $signed(x642_rdrow_number); // @[Math.scala 406:49:@43951.4]
  assign _T_1217 = $signed(_T_1215) & $signed(32'sh3); // @[Math.scala 406:56:@43953.4]
  assign _T_1218 = $signed(_T_1217); // @[Math.scala 406:56:@43954.4]
  assign _T_1222 = $signed(RetimeWrapper_84_io_out); // @[package.scala 96:25:@43962.4]
  assign x814_number = $unsigned(_T_1222); // @[implicits.scala 133:21:@43964.4]
  assign x644 = RetimeWrapper_85_io_out; // @[package.scala 96:25:@43978.4 package.scala 96:25:@43979.4]
  assign x645 = x644 | x561; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 513:24:@43982.4]
  assign _T_1245 = $signed(x814_number); // @[Math.scala 406:49:@43991.4]
  assign _T_1247 = $signed(_T_1245) & $signed(32'sh3); // @[Math.scala 406:56:@43993.4]
  assign _T_1248 = $signed(_T_1247); // @[Math.scala 406:56:@43994.4]
  assign _T_1253 = x814_number[31]; // @[FixedPoint.scala 50:25:@44000.4]
  assign _T_1257 = _T_1253 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@44002.4]
  assign _T_1258 = x814_number[31:2]; // @[FixedPoint.scala 18:52:@44003.4]
  assign x648_number = {_T_1257,_T_1258}; // @[Cat.scala 30:58:@44004.4]
  assign _GEN_6 = {{8'd0}, x648_number}; // @[Math.scala 450:32:@44009.4]
  assign _T_1263 = _GEN_6 << 8; // @[Math.scala 450:32:@44009.4]
  assign _GEN_7 = {{6'd0}, x648_number}; // @[Math.scala 450:32:@44014.4]
  assign _T_1267 = _GEN_7 << 6; // @[Math.scala 450:32:@44014.4]
  assign _T_1294 = RetimeWrapper_89_io_out; // @[package.scala 96:25:@44073.4 package.scala 96:25:@44074.4]
  assign _T_1296 = io_rr ? _T_1294 : 1'h0; // @[implicits.scala 55:10:@44075.4]
  assign _T_1297 = _T_379 & _T_1296; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 544:194:@44076.4]
  assign x883_x646_D20 = RetimeWrapper_87_io_out; // @[package.scala 96:25:@44052.4 package.scala 96:25:@44053.4]
  assign _T_1298 = _T_1297 & x883_x646_D20; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 544:283:@44077.4]
  assign _T_1299 = _T_1298 & x851_b521_D48; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 544:326:@44078.4]
  assign x653 = x644 | x570; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 548:59:@44089.4]
  assign _T_1325 = RetimeWrapper_91_io_out; // @[package.scala 96:25:@44124.4 package.scala 96:25:@44125.4]
  assign _T_1327 = io_rr ? _T_1325 : 1'h0; // @[implicits.scala 55:10:@44126.4]
  assign _T_1328 = _T_379 & _T_1327; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 561:194:@44127.4]
  assign x885_x654_D20 = RetimeWrapper_90_io_out; // @[package.scala 96:25:@44112.4 package.scala 96:25:@44113.4]
  assign _T_1329 = _T_1328 & x885_x654_D20; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 561:283:@44128.4]
  assign _T_1330 = _T_1329 & x851_b521_D48; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 561:291:@44129.4]
  assign x658 = x644 | x576; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 565:59:@44140.4]
  assign _T_1354 = RetimeWrapper_93_io_out; // @[package.scala 96:25:@44173.4 package.scala 96:25:@44174.4]
  assign _T_1356 = io_rr ? _T_1354 : 1'h0; // @[implicits.scala 55:10:@44175.4]
  assign _T_1357 = _T_379 & _T_1356; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 576:194:@44176.4]
  assign x886_x659_D20 = RetimeWrapper_92_io_out; // @[package.scala 96:25:@44161.4 package.scala 96:25:@44162.4]
  assign _T_1358 = _T_1357 & x886_x659_D20; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 576:283:@44177.4]
  assign _T_1359 = _T_1358 & x851_b521_D48; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 576:291:@44178.4]
  assign x663 = x644 | x876_x582_D1; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 580:59:@44189.4]
  assign _T_1389 = RetimeWrapper_97_io_out; // @[package.scala 96:25:@44240.4 package.scala 96:25:@44241.4]
  assign _T_1391 = io_rr ? _T_1389 : 1'h0; // @[implicits.scala 55:10:@44242.4]
  assign _T_1392 = _T_379 & _T_1391; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 595:194:@44243.4]
  assign x889_x664_D20 = RetimeWrapper_96_io_out; // @[package.scala 96:25:@44228.4 package.scala 96:25:@44229.4]
  assign _T_1393 = _T_1392 & x889_x664_D20; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 595:283:@44244.4]
  assign _T_1394 = _T_1393 & x851_b521_D48; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 595:291:@44245.4]
  assign x668 = x644 | x589; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 599:59:@44256.4]
  assign _T_1418 = RetimeWrapper_99_io_out; // @[package.scala 96:25:@44289.4 package.scala 96:25:@44290.4]
  assign _T_1420 = io_rr ? _T_1418 : 1'h0; // @[implicits.scala 55:10:@44291.4]
  assign _T_1421 = _T_379 & _T_1420; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 610:194:@44292.4]
  assign x890_x669_D20 = RetimeWrapper_98_io_out; // @[package.scala 96:25:@44277.4 package.scala 96:25:@44278.4]
  assign _T_1422 = _T_1421 & x890_x669_D20; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 610:283:@44293.4]
  assign _T_1423 = _T_1422 & x851_b521_D48; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 610:291:@44294.4]
  assign x673 = x644 | x598; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 614:59:@44305.4]
  assign _T_1447 = RetimeWrapper_101_io_out; // @[package.scala 96:25:@44338.4 package.scala 96:25:@44339.4]
  assign _T_1449 = io_rr ? _T_1447 : 1'h0; // @[implicits.scala 55:10:@44340.4]
  assign _T_1450 = _T_379 & _T_1449; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 625:194:@44341.4]
  assign x891_x674_D20 = RetimeWrapper_100_io_out; // @[package.scala 96:25:@44326.4 package.scala 96:25:@44327.4]
  assign _T_1451 = _T_1450 & x891_x674_D20; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 625:283:@44342.4]
  assign _T_1452 = _T_1451 & x851_b521_D48; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 625:291:@44343.4]
  assign x574_rd_0_number = x525_lb_0_io_rPort_2_output_0; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 267:29:@43068.4 sm_x736_inr_Foreach_SAMPLER_BOX.scala 271:338:@43089.4]
  assign _GEN_8 = {{1'd0}, x574_rd_0_number}; // @[Math.scala 450:32:@44355.4]
  assign x615_rd_0_number = x525_lb_0_io_rPort_6_output_0; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 416:29:@43637.4 sm_x736_inr_Foreach_SAMPLER_BOX.scala 420:408:@43658.4]
  assign _GEN_9 = {{1'd0}, x615_rd_0_number}; // @[Math.scala 450:32:@44367.4]
  assign x620_rd_0_number = x525_lb_0_io_rPort_15_output_0; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 433:29:@43688.4 sm_x736_inr_Foreach_SAMPLER_BOX.scala 437:408:@43709.4]
  assign _GEN_10 = {{2'd0}, x620_rd_0_number}; // @[Math.scala 450:32:@44379.4]
  assign x625_rd_0_number = x525_lb_0_io_rPort_5_output_0; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 448:29:@43737.4 sm_x736_inr_Foreach_SAMPLER_BOX.scala 452:408:@43758.4]
  assign _GEN_11 = {{1'd0}, x625_rd_0_number}; // @[Math.scala 450:32:@44391.4]
  assign x656_rd_0_number = x525_lb_0_io_rPort_11_output_0; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 557:29:@44115.4 sm_x736_inr_Foreach_SAMPLER_BOX.scala 561:408:@44136.4]
  assign _GEN_12 = {{1'd0}, x656_rd_0_number}; // @[Math.scala 450:32:@44403.4]
  assign x690_sum_number = x690_sum_1_io_result; // @[Math.scala 154:22:@44528.4 Math.scala 155:14:@44529.4]
  assign _T_1531 = x690_sum_number[7:4]; // @[FixedPoint.scala 18:52:@44534.4]
  assign x580_rd_0_number = x525_lb_0_io_rPort_9_output_0; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 296:29:@43158.4 sm_x736_inr_Foreach_SAMPLER_BOX.scala 300:443:@43179.4]
  assign _GEN_13 = {{1'd0}, x580_rd_0_number}; // @[Math.scala 450:32:@44540.4]
  assign _GEN_14 = {{1'd0}, x620_rd_0_number}; // @[Math.scala 450:32:@44552.4]
  assign _GEN_15 = {{2'd0}, x625_rd_0_number}; // @[Math.scala 450:32:@44564.4]
  assign x630_rd_0_number = x525_lb_0_io_rPort_4_output_0; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 469:29:@43813.4 sm_x736_inr_Foreach_SAMPLER_BOX.scala 473:408:@43834.4]
  assign _GEN_16 = {{1'd0}, x630_rd_0_number}; // @[Math.scala 450:32:@44576.4]
  assign x661_rd_0_number = x525_lb_0_io_rPort_3_output_0; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 572:29:@44164.4 sm_x736_inr_Foreach_SAMPLER_BOX.scala 576:408:@44185.4]
  assign _GEN_17 = {{1'd0}, x661_rd_0_number}; // @[Math.scala 450:32:@44588.4]
  assign x704_sum_number = x704_sum_1_io_result; // @[Math.scala 154:22:@44711.4 Math.scala 155:14:@44712.4]
  assign _T_1607 = x704_sum_number[7:4]; // @[FixedPoint.scala 18:52:@44717.4]
  assign x586_rd_0_number = x525_lb_0_io_rPort_7_output_0; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 325:29:@43268.4 sm_x736_inr_Foreach_SAMPLER_BOX.scala 329:408:@43289.4]
  assign _GEN_18 = {{1'd0}, x586_rd_0_number}; // @[Math.scala 450:32:@44723.4]
  assign _GEN_19 = {{2'd0}, x630_rd_0_number}; // @[Math.scala 450:32:@44735.4]
  assign x635_rd_0_number = x525_lb_0_io_rPort_16_output_0; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 484:29:@43862.4 sm_x736_inr_Foreach_SAMPLER_BOX.scala 488:408:@43883.4]
  assign _GEN_20 = {{1'd0}, x635_rd_0_number}; // @[Math.scala 450:32:@44747.4]
  assign x666_rd_0_number = x525_lb_0_io_rPort_0_output_0; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 591:29:@44231.4 sm_x736_inr_Foreach_SAMPLER_BOX.scala 595:408:@44252.4]
  assign _GEN_21 = {{1'd0}, x666_rd_0_number}; // @[Math.scala 450:32:@44759.4]
  assign x717_sum_number = x717_sum_1_io_result; // @[Math.scala 154:22:@44864.4 Math.scala 155:14:@44865.4]
  assign _T_1671 = x717_sum_number[7:4]; // @[FixedPoint.scala 18:52:@44870.4]
  assign x595_rd_0_number = x525_lb_0_io_rPort_12_output_0; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 350:29:@43376.4 sm_x736_inr_Foreach_SAMPLER_BOX.scala 354:408:@43397.4]
  assign _GEN_22 = {{1'd0}, x595_rd_0_number}; // @[Math.scala 450:32:@44876.4]
  assign _GEN_23 = {{2'd0}, x635_rd_0_number}; // @[Math.scala 450:32:@44888.4]
  assign x640_rd_0_number = x525_lb_0_io_rPort_10_output_0; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 499:29:@43911.4 sm_x736_inr_Foreach_SAMPLER_BOX.scala 503:408:@43932.4]
  assign _GEN_24 = {{1'd0}, x640_rd_0_number}; // @[Math.scala 450:32:@44900.4]
  assign x671_rd_0_number = x525_lb_0_io_rPort_13_output_0; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 606:29:@44280.4 sm_x736_inr_Foreach_SAMPLER_BOX.scala 610:408:@44301.4]
  assign _GEN_25 = {{1'd0}, x671_rd_0_number}; // @[Math.scala 450:32:@44912.4]
  assign x730_sum_number = x730_sum_1_io_result; // @[Math.scala 154:22:@45019.4 Math.scala 155:14:@45020.4]
  assign _T_1737 = x730_sum_number[7:4]; // @[FixedPoint.scala 18:52:@45025.4]
  assign _T_1750 = {4'h0,_T_1671,4'h0,_T_1737}; // @[Cat.scala 30:58:@45035.4]
  assign _T_1751 = {4'h0,_T_1531,4'h0,_T_1607}; // @[Cat.scala 30:58:@45036.4]
  assign _T_1764 = RetimeWrapper_135_io_out; // @[package.scala 96:25:@45072.4 package.scala 96:25:@45073.4]
  assign _T_1766 = io_rr ? _T_1764 : 1'h0; // @[implicits.scala 55:10:@45074.4]
  assign x904_b521_D55 = RetimeWrapper_133_io_out; // @[package.scala 96:25:@45054.4 package.scala 96:25:@45055.4]
  assign _T_1767 = _T_1766 & x904_b521_D55; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 785:117:@45075.4]
  assign x905_b522_D55 = RetimeWrapper_134_io_out; // @[package.scala 96:25:@45063.4 package.scala 96:25:@45064.4]
  assign _T_1768 = _T_1767 & x905_b522_D55; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 785:123:@45076.4]
  assign x827_x538_sum_D3_number = RetimeWrapper_3_io_out; // @[package.scala 96:25:@42408.4 package.scala 96:25:@42409.4]
  assign x828_x534_D8_number = RetimeWrapper_4_io_out; // @[package.scala 96:25:@42417.4 package.scala 96:25:@42418.4]
  assign x831_x800_D22_number = RetimeWrapper_7_io_out; // @[package.scala 96:25:@42444.4 package.scala 96:25:@42445.4]
  assign x834_x542_D7_number = RetimeWrapper_11_io_out; // @[package.scala 96:25:@42542.4 package.scala 96:25:@42543.4]
  assign x836_x544_sum_D2_number = RetimeWrapper_13_io_out; // @[package.scala 96:25:@42560.4 package.scala 96:25:@42561.4]
  assign x837_x550_sum_D2_number = RetimeWrapper_15_io_out; // @[package.scala 96:25:@42640.4 package.scala 96:25:@42641.4]
  assign x839_x548_D7_number = RetimeWrapper_17_io_out; // @[package.scala 96:25:@42658.4 package.scala 96:25:@42659.4]
  assign x840_x554_D7_number = RetimeWrapper_19_io_out; // @[package.scala 96:25:@42740.4 package.scala 96:25:@42741.4]
  assign x842_x556_sum_D2_number = RetimeWrapper_21_io_out; // @[package.scala 96:25:@42758.4 package.scala 96:25:@42759.4]
  assign x567_sum_number = x567_sum_1_io_result; // @[Math.scala 154:22:@42930.4 Math.scala 155:14:@42931.4]
  assign x849_x554_D31_number = RetimeWrapper_32_io_out; // @[package.scala 96:25:@42948.4 package.scala 96:25:@42949.4]
  assign x850_x805_D21_number = RetimeWrapper_33_io_out; // @[package.scala 96:25:@42957.4 package.scala 96:25:@42958.4]
  assign x573_sum_number = x573_sum_1_io_result; // @[Math.scala 154:22:@43047.4 Math.scala 155:14:@43048.4]
  assign x856_x548_D31_number = RetimeWrapper_41_io_out; // @[package.scala 96:25:@43065.4 package.scala 96:25:@43066.4]
  assign x579_sum_number = x579_sum_1_io_result; // @[Math.scala 154:22:@43137.4 Math.scala 155:14:@43138.4]
  assign x859_x542_D31_number = RetimeWrapper_46_io_out; // @[package.scala 96:25:@43146.4 package.scala 96:25:@43147.4]
  assign x864_x534_D32_number = RetimeWrapper_53_io_out; // @[package.scala 96:25:@43247.4 package.scala 96:25:@43248.4]
  assign x866_x585_sum_D1_number = RetimeWrapper_55_io_out; // @[package.scala 96:25:@43265.4 package.scala 96:25:@43266.4]
  assign x594_sum_number = x594_sum_1_io_result; // @[Math.scala 154:22:@43355.4 Math.scala 155:14:@43356.4]
  assign x868_x592_D5_number = RetimeWrapper_59_io_out; // @[package.scala 96:25:@43373.4 package.scala 96:25:@43374.4]
  assign x603_sum_number = x603_sum_1_io_result; // @[Math.scala 154:22:@43463.4 Math.scala 155:14:@43464.4]
  assign x869_x601_D5_number = RetimeWrapper_62_io_out; // @[package.scala 96:25:@43472.4 package.scala 96:25:@43473.4]
  assign x614_sum_number = x614_sum_1_io_result; // @[Math.scala 154:22:@43616.4 Math.scala 155:14:@43617.4]
  assign x872_x810_D20_number = RetimeWrapper_68_io_out; // @[package.scala 96:25:@43625.4 package.scala 96:25:@43626.4]
  assign x619_sum_number = x619_sum_1_io_result; // @[Math.scala 154:22:@43676.4 Math.scala 155:14:@43677.4]
  assign x624_sum_number = x624_sum_1_io_result; // @[Math.scala 154:22:@43725.4 Math.scala 155:14:@43726.4]
  assign x878_x629_sum_D1_number = RetimeWrapper_77_io_out; // @[package.scala 96:25:@43801.4 package.scala 96:25:@43802.4]
  assign x634_sum_number = x634_sum_1_io_result; // @[Math.scala 154:22:@43850.4 Math.scala 155:14:@43851.4]
  assign x639_sum_number = x639_sum_1_io_result; // @[Math.scala 154:22:@43899.4 Math.scala 155:14:@43900.4]
  assign x650_sum_number = x650_sum_1_io_result; // @[Math.scala 154:22:@44043.4 Math.scala 155:14:@44044.4]
  assign x884_x815_D20_number = RetimeWrapper_88_io_out; // @[package.scala 96:25:@44061.4 package.scala 96:25:@44062.4]
  assign x655_sum_number = x655_sum_1_io_result; // @[Math.scala 154:22:@44103.4 Math.scala 155:14:@44104.4]
  assign x660_sum_number = x660_sum_1_io_result; // @[Math.scala 154:22:@44152.4 Math.scala 155:14:@44153.4]
  assign x888_x665_sum_D1_number = RetimeWrapper_95_io_out; // @[package.scala 96:25:@44219.4 package.scala 96:25:@44220.4]
  assign x670_sum_number = x670_sum_1_io_result; // @[Math.scala 154:22:@44268.4 Math.scala 155:14:@44269.4]
  assign x675_sum_number = x675_sum_1_io_result; // @[Math.scala 154:22:@44317.4 Math.scala 155:14:@44318.4]
  assign _T_1460 = RetimeWrapper_102_io_out; // @[package.scala 96:25:@44361.4 package.scala 96:25:@44362.4]
  assign _T_1466 = RetimeWrapper_103_io_out; // @[package.scala 96:25:@44373.4 package.scala 96:25:@44374.4]
  assign _T_1472 = RetimeWrapper_104_io_out; // @[package.scala 96:25:@44385.4 package.scala 96:25:@44386.4]
  assign _T_1478 = RetimeWrapper_105_io_out; // @[package.scala 96:25:@44397.4 package.scala 96:25:@44398.4]
  assign _T_1484 = RetimeWrapper_106_io_out; // @[package.scala 96:25:@44409.4 package.scala 96:25:@44410.4]
  assign _T_1538 = RetimeWrapper_111_io_out; // @[package.scala 96:25:@44546.4 package.scala 96:25:@44547.4]
  assign _T_1544 = RetimeWrapper_112_io_out; // @[package.scala 96:25:@44558.4 package.scala 96:25:@44559.4]
  assign _T_1550 = RetimeWrapper_113_io_out; // @[package.scala 96:25:@44570.4 package.scala 96:25:@44571.4]
  assign _T_1556 = RetimeWrapper_114_io_out; // @[package.scala 96:25:@44582.4 package.scala 96:25:@44583.4]
  assign _T_1562 = RetimeWrapper_115_io_out; // @[package.scala 96:25:@44594.4 package.scala 96:25:@44595.4]
  assign _T_1614 = RetimeWrapper_120_io_out; // @[package.scala 96:25:@44729.4 package.scala 96:25:@44730.4]
  assign _T_1620 = RetimeWrapper_121_io_out; // @[package.scala 96:25:@44741.4 package.scala 96:25:@44742.4]
  assign _T_1626 = RetimeWrapper_122_io_out; // @[package.scala 96:25:@44753.4 package.scala 96:25:@44754.4]
  assign _T_1632 = RetimeWrapper_123_io_out; // @[package.scala 96:25:@44765.4 package.scala 96:25:@44766.4]
  assign _T_1678 = RetimeWrapper_126_io_out; // @[package.scala 96:25:@44882.4 package.scala 96:25:@44883.4]
  assign _T_1684 = RetimeWrapper_127_io_out; // @[package.scala 96:25:@44894.4 package.scala 96:25:@44895.4]
  assign _T_1690 = RetimeWrapper_128_io_out; // @[package.scala 96:25:@44906.4 package.scala 96:25:@44907.4]
  assign _T_1696 = RetimeWrapper_129_io_out; // @[package.scala 96:25:@44918.4 package.scala 96:25:@44919.4]
  assign io_in_x481_TVALID = _T_1768 & io_sigsIn_backpressure; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 785:22:@45078.4]
  assign io_in_x481_TDATA = {{224'd0}, RetimeWrapper_132_io_out}; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 786:24:@45079.4]
  assign io_in_x480_TREADY = _T_211 & _T_213; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 67:22:@42085.4 sm_x736_inr_Foreach_SAMPLER_BOX.scala 69:22:@42093.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 710:17:@42063.4]
  assign __1_io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_1); // @[Math.scala 710:17:@42075.4]
  assign RetimeWrapper_clock = clock; // @[:@42096.4]
  assign RetimeWrapper_reset = reset; // @[:@42097.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@42099.4]
  assign RetimeWrapper_io_in = io_in_x480_TDATA[31:0]; // @[package.scala 94:16:@42098.4]
  assign x525_lb_0_clock = clock; // @[:@42106.4]
  assign x525_lb_0_reset = reset; // @[:@42107.4]
  assign x525_lb_0_io_rPort_17_banks_1 = x869_x601_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@44346.4]
  assign x525_lb_0_io_rPort_17_banks_0 = x884_x815_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@44345.4]
  assign x525_lb_0_io_rPort_17_ofs_0 = x675_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@44347.4]
  assign x525_lb_0_io_rPort_17_en_0 = _T_1452 & x848_b522_D48; // @[MemInterfaceType.scala 110:79:@44349.4]
  assign x525_lb_0_io_rPort_17_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@44348.4]
  assign x525_lb_0_io_rPort_16_banks_1 = x868_x592_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@43879.4]
  assign x525_lb_0_io_rPort_16_banks_0 = x872_x810_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@43878.4]
  assign x525_lb_0_io_rPort_16_ofs_0 = x634_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@43880.4]
  assign x525_lb_0_io_rPort_16_en_0 = _T_1169 & x848_b522_D48; // @[MemInterfaceType.scala 110:79:@43882.4]
  assign x525_lb_0_io_rPort_16_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@43881.4]
  assign x525_lb_0_io_rPort_15_banks_1 = x856_x548_D31_number[2:0]; // @[MemInterfaceType.scala 106:58:@43705.4]
  assign x525_lb_0_io_rPort_15_banks_0 = x872_x810_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@43704.4]
  assign x525_lb_0_io_rPort_15_ofs_0 = x619_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@43706.4]
  assign x525_lb_0_io_rPort_15_en_0 = _T_1073 & x848_b522_D48; // @[MemInterfaceType.scala 110:79:@43708.4]
  assign x525_lb_0_io_rPort_15_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@43707.4]
  assign x525_lb_0_io_rPort_14_banks_1 = x849_x554_D31_number[2:0]; // @[MemInterfaceType.scala 106:58:@42995.4]
  assign x525_lb_0_io_rPort_14_banks_0 = x850_x805_D21_number[2:0]; // @[MemInterfaceType.scala 106:58:@42994.4]
  assign x525_lb_0_io_rPort_14_ofs_0 = x567_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@42996.4]
  assign x525_lb_0_io_rPort_14_en_0 = _T_663 & x848_b522_D48; // @[MemInterfaceType.scala 110:79:@42998.4]
  assign x525_lb_0_io_rPort_14_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@42997.4]
  assign x525_lb_0_io_rPort_13_banks_1 = x868_x592_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@44297.4]
  assign x525_lb_0_io_rPort_13_banks_0 = x884_x815_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@44296.4]
  assign x525_lb_0_io_rPort_13_ofs_0 = x670_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@44298.4]
  assign x525_lb_0_io_rPort_13_en_0 = _T_1423 & x848_b522_D48; // @[MemInterfaceType.scala 110:79:@44300.4]
  assign x525_lb_0_io_rPort_13_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@44299.4]
  assign x525_lb_0_io_rPort_12_banks_1 = x868_x592_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@43393.4]
  assign x525_lb_0_io_rPort_12_banks_0 = x850_x805_D21_number[2:0]; // @[MemInterfaceType.scala 106:58:@43392.4]
  assign x525_lb_0_io_rPort_12_ofs_0 = x594_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@43394.4]
  assign x525_lb_0_io_rPort_12_en_0 = _T_878 & x848_b522_D48; // @[MemInterfaceType.scala 110:79:@43396.4]
  assign x525_lb_0_io_rPort_12_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@43395.4]
  assign x525_lb_0_io_rPort_11_banks_1 = x856_x548_D31_number[2:0]; // @[MemInterfaceType.scala 106:58:@44132.4]
  assign x525_lb_0_io_rPort_11_banks_0 = x884_x815_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@44131.4]
  assign x525_lb_0_io_rPort_11_ofs_0 = x655_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@44133.4]
  assign x525_lb_0_io_rPort_11_en_0 = _T_1330 & x848_b522_D48; // @[MemInterfaceType.scala 110:79:@44135.4]
  assign x525_lb_0_io_rPort_11_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@44134.4]
  assign x525_lb_0_io_rPort_10_banks_1 = x869_x601_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@43928.4]
  assign x525_lb_0_io_rPort_10_banks_0 = x872_x810_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@43927.4]
  assign x525_lb_0_io_rPort_10_ofs_0 = x639_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@43929.4]
  assign x525_lb_0_io_rPort_10_en_0 = _T_1198 & x848_b522_D48; // @[MemInterfaceType.scala 110:79:@43931.4]
  assign x525_lb_0_io_rPort_10_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@43930.4]
  assign x525_lb_0_io_rPort_9_banks_1 = x859_x542_D31_number[2:0]; // @[MemInterfaceType.scala 106:58:@43175.4]
  assign x525_lb_0_io_rPort_9_banks_0 = x850_x805_D21_number[2:0]; // @[MemInterfaceType.scala 106:58:@43174.4]
  assign x525_lb_0_io_rPort_9_ofs_0 = x579_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@43176.4]
  assign x525_lb_0_io_rPort_9_en_0 = _T_759 & x848_b522_D48; // @[MemInterfaceType.scala 110:79:@43178.4]
  assign x525_lb_0_io_rPort_9_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@43177.4]
  assign x525_lb_0_io_rPort_8_banks_1 = x869_x601_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@43501.4]
  assign x525_lb_0_io_rPort_8_banks_0 = x850_x805_D21_number[2:0]; // @[MemInterfaceType.scala 106:58:@43500.4]
  assign x525_lb_0_io_rPort_8_ofs_0 = x603_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@43502.4]
  assign x525_lb_0_io_rPort_8_en_0 = _T_941 & x848_b522_D48; // @[MemInterfaceType.scala 110:79:@43504.4]
  assign x525_lb_0_io_rPort_8_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@43503.4]
  assign x525_lb_0_io_rPort_7_banks_1 = x864_x534_D32_number[2:0]; // @[MemInterfaceType.scala 106:58:@43285.4]
  assign x525_lb_0_io_rPort_7_banks_0 = x850_x805_D21_number[2:0]; // @[MemInterfaceType.scala 106:58:@43284.4]
  assign x525_lb_0_io_rPort_7_ofs_0 = x866_x585_sum_D1_number[8:0]; // @[MemInterfaceType.scala 107:54:@43286.4]
  assign x525_lb_0_io_rPort_7_en_0 = _T_815 & x848_b522_D48; // @[MemInterfaceType.scala 110:79:@43288.4]
  assign x525_lb_0_io_rPort_7_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@43287.4]
  assign x525_lb_0_io_rPort_6_banks_1 = x849_x554_D31_number[2:0]; // @[MemInterfaceType.scala 106:58:@43654.4]
  assign x525_lb_0_io_rPort_6_banks_0 = x872_x810_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@43653.4]
  assign x525_lb_0_io_rPort_6_ofs_0 = x614_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@43655.4]
  assign x525_lb_0_io_rPort_6_en_0 = _T_1042 & x848_b522_D48; // @[MemInterfaceType.scala 110:79:@43657.4]
  assign x525_lb_0_io_rPort_6_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@43656.4]
  assign x525_lb_0_io_rPort_5_banks_1 = x859_x542_D31_number[2:0]; // @[MemInterfaceType.scala 106:58:@43754.4]
  assign x525_lb_0_io_rPort_5_banks_0 = x872_x810_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@43753.4]
  assign x525_lb_0_io_rPort_5_ofs_0 = x624_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@43755.4]
  assign x525_lb_0_io_rPort_5_en_0 = _T_1102 & x848_b522_D48; // @[MemInterfaceType.scala 110:79:@43757.4]
  assign x525_lb_0_io_rPort_5_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@43756.4]
  assign x525_lb_0_io_rPort_4_banks_1 = x864_x534_D32_number[2:0]; // @[MemInterfaceType.scala 106:58:@43830.4]
  assign x525_lb_0_io_rPort_4_banks_0 = x872_x810_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@43829.4]
  assign x525_lb_0_io_rPort_4_ofs_0 = x878_x629_sum_D1_number[8:0]; // @[MemInterfaceType.scala 107:54:@43831.4]
  assign x525_lb_0_io_rPort_4_en_0 = _T_1140 & x848_b522_D48; // @[MemInterfaceType.scala 110:79:@43833.4]
  assign x525_lb_0_io_rPort_4_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@43832.4]
  assign x525_lb_0_io_rPort_3_banks_1 = x859_x542_D31_number[2:0]; // @[MemInterfaceType.scala 106:58:@44181.4]
  assign x525_lb_0_io_rPort_3_banks_0 = x884_x815_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@44180.4]
  assign x525_lb_0_io_rPort_3_ofs_0 = x660_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@44182.4]
  assign x525_lb_0_io_rPort_3_en_0 = _T_1359 & x848_b522_D48; // @[MemInterfaceType.scala 110:79:@44184.4]
  assign x525_lb_0_io_rPort_3_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@44183.4]
  assign x525_lb_0_io_rPort_2_banks_1 = x856_x548_D31_number[2:0]; // @[MemInterfaceType.scala 106:58:@43085.4]
  assign x525_lb_0_io_rPort_2_banks_0 = x850_x805_D21_number[2:0]; // @[MemInterfaceType.scala 106:58:@43084.4]
  assign x525_lb_0_io_rPort_2_ofs_0 = x573_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@43086.4]
  assign x525_lb_0_io_rPort_2_en_0 = _T_711 & x848_b522_D48; // @[MemInterfaceType.scala 110:79:@43088.4]
  assign x525_lb_0_io_rPort_2_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@43087.4]
  assign x525_lb_0_io_rPort_1_banks_1 = x849_x554_D31_number[2:0]; // @[MemInterfaceType.scala 106:58:@44081.4]
  assign x525_lb_0_io_rPort_1_banks_0 = x884_x815_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@44080.4]
  assign x525_lb_0_io_rPort_1_ofs_0 = x650_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@44082.4]
  assign x525_lb_0_io_rPort_1_en_0 = _T_1299 & x848_b522_D48; // @[MemInterfaceType.scala 110:79:@44084.4]
  assign x525_lb_0_io_rPort_1_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@44083.4]
  assign x525_lb_0_io_rPort_0_banks_1 = x864_x534_D32_number[2:0]; // @[MemInterfaceType.scala 106:58:@44248.4]
  assign x525_lb_0_io_rPort_0_banks_0 = x884_x815_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@44247.4]
  assign x525_lb_0_io_rPort_0_ofs_0 = x888_x665_sum_D1_number[8:0]; // @[MemInterfaceType.scala 107:54:@44249.4]
  assign x525_lb_0_io_rPort_0_en_0 = _T_1394 & x848_b522_D48; // @[MemInterfaceType.scala 110:79:@44251.4]
  assign x525_lb_0_io_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@44250.4]
  assign x525_lb_0_io_wPort_3_banks_1 = x840_x554_D7_number[2:0]; // @[MemInterfaceType.scala 88:58:@42779.4]
  assign x525_lb_0_io_wPort_3_banks_0 = x831_x800_D22_number[2:0]; // @[MemInterfaceType.scala 88:58:@42778.4]
  assign x525_lb_0_io_wPort_3_ofs_0 = x842_x556_sum_D2_number[8:0]; // @[MemInterfaceType.scala 89:54:@42780.4]
  assign x525_lb_0_io_wPort_3_data_0 = RetimeWrapper_20_io_out; // @[MemInterfaceType.scala 90:56:@42781.4]
  assign x525_lb_0_io_wPort_3_en_0 = _T_539 & x829_b522_D24; // @[MemInterfaceType.scala 93:57:@42783.4]
  assign x525_lb_0_io_wPort_2_banks_1 = x839_x548_D7_number[2:0]; // @[MemInterfaceType.scala 88:58:@42679.4]
  assign x525_lb_0_io_wPort_2_banks_0 = x831_x800_D22_number[2:0]; // @[MemInterfaceType.scala 88:58:@42678.4]
  assign x525_lb_0_io_wPort_2_ofs_0 = x837_x550_sum_D2_number[8:0]; // @[MemInterfaceType.scala 89:54:@42680.4]
  assign x525_lb_0_io_wPort_2_data_0 = RetimeWrapper_16_io_out; // @[MemInterfaceType.scala 90:56:@42681.4]
  assign x525_lb_0_io_wPort_2_en_0 = _T_489 & x829_b522_D24; // @[MemInterfaceType.scala 93:57:@42683.4]
  assign x525_lb_0_io_wPort_1_banks_1 = x834_x542_D7_number[2:0]; // @[MemInterfaceType.scala 88:58:@42581.4]
  assign x525_lb_0_io_wPort_1_banks_0 = x831_x800_D22_number[2:0]; // @[MemInterfaceType.scala 88:58:@42580.4]
  assign x525_lb_0_io_wPort_1_ofs_0 = x836_x544_sum_D2_number[8:0]; // @[MemInterfaceType.scala 89:54:@42582.4]
  assign x525_lb_0_io_wPort_1_data_0 = RetimeWrapper_12_io_out; // @[MemInterfaceType.scala 90:56:@42583.4]
  assign x525_lb_0_io_wPort_1_en_0 = _T_441 & x829_b522_D24; // @[MemInterfaceType.scala 93:57:@42585.4]
  assign x525_lb_0_io_wPort_0_banks_1 = x828_x534_D8_number[2:0]; // @[MemInterfaceType.scala 88:58:@42474.4]
  assign x525_lb_0_io_wPort_0_banks_0 = x831_x800_D22_number[2:0]; // @[MemInterfaceType.scala 88:58:@42473.4]
  assign x525_lb_0_io_wPort_0_ofs_0 = x827_x538_sum_D3_number[8:0]; // @[MemInterfaceType.scala 89:54:@42475.4]
  assign x525_lb_0_io_wPort_0_data_0 = RetimeWrapper_8_io_out; // @[MemInterfaceType.scala 90:56:@42476.4]
  assign x525_lb_0_io_wPort_0_en_0 = _T_390 & x829_b522_D24; // @[MemInterfaceType.scala 93:57:@42478.4]
  assign RetimeWrapper_1_clock = clock; // @[:@42312.4]
  assign RetimeWrapper_1_reset = reset; // @[:@42313.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@42315.4]
  assign RetimeWrapper_1_io_in = _T_299 | _T_297; // @[package.scala 94:16:@42314.4]
  assign x534_1_clock = clock; // @[:@42334.4]
  assign x534_1_reset = reset; // @[:@42335.4]
  assign x534_1_io_a = __1_io_result; // @[Math.scala 367:17:@42336.4]
  assign x534_1_io_flow = io_in_x481_TREADY; // @[Math.scala 369:20:@42338.4]
  assign x803_sum_1_clock = clock; // @[:@42363.4]
  assign x803_sum_1_reset = reset; // @[:@42364.4]
  assign x803_sum_1_io_a = _T_339[31:0]; // @[Math.scala 151:17:@42365.4]
  assign x803_sum_1_io_b = _T_343[31:0]; // @[Math.scala 152:17:@42366.4]
  assign x803_sum_1_io_flow = io_in_x481_TREADY; // @[Math.scala 153:20:@42367.4]
  assign x537_div_1_clock = clock; // @[:@42375.4]
  assign x537_div_1_reset = reset; // @[:@42376.4]
  assign x537_div_1_io_a = __1_io_result; // @[Math.scala 328:17:@42377.4]
  assign x537_div_1_io_flow = io_in_x481_TREADY; // @[Math.scala 330:20:@42379.4]
  assign RetimeWrapper_2_clock = clock; // @[:@42385.4]
  assign RetimeWrapper_2_reset = reset; // @[:@42386.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@42388.4]
  assign RetimeWrapper_2_io_in = x803_sum_1_io_result; // @[package.scala 94:16:@42387.4]
  assign x538_sum_1_clock = clock; // @[:@42394.4]
  assign x538_sum_1_reset = reset; // @[:@42395.4]
  assign x538_sum_1_io_a = RetimeWrapper_2_io_out; // @[Math.scala 151:17:@42396.4]
  assign x538_sum_1_io_b = x537_div_1_io_result; // @[Math.scala 152:17:@42397.4]
  assign x538_sum_1_io_flow = io_in_x481_TREADY; // @[Math.scala 153:20:@42398.4]
  assign RetimeWrapper_3_clock = clock; // @[:@42404.4]
  assign RetimeWrapper_3_reset = reset; // @[:@42405.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@42407.4]
  assign RetimeWrapper_3_io_in = x538_sum_1_io_result; // @[package.scala 94:16:@42406.4]
  assign RetimeWrapper_4_clock = clock; // @[:@42413.4]
  assign RetimeWrapper_4_reset = reset; // @[:@42414.4]
  assign RetimeWrapper_4_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@42416.4]
  assign RetimeWrapper_4_io_in = x534_1_io_result; // @[package.scala 94:16:@42415.4]
  assign RetimeWrapper_5_clock = clock; // @[:@42422.4]
  assign RetimeWrapper_5_reset = reset; // @[:@42423.4]
  assign RetimeWrapper_5_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@42425.4]
  assign RetimeWrapper_5_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@42424.4]
  assign RetimeWrapper_6_clock = clock; // @[:@42431.4]
  assign RetimeWrapper_6_reset = reset; // @[:@42432.4]
  assign RetimeWrapper_6_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@42434.4]
  assign RetimeWrapper_6_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@42433.4]
  assign RetimeWrapper_7_clock = clock; // @[:@42440.4]
  assign RetimeWrapper_7_reset = reset; // @[:@42441.4]
  assign RetimeWrapper_7_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@42443.4]
  assign RetimeWrapper_7_io_in = $unsigned(_T_317); // @[package.scala 94:16:@42442.4]
  assign RetimeWrapper_8_clock = clock; // @[:@42449.4]
  assign RetimeWrapper_8_reset = reset; // @[:@42450.4]
  assign RetimeWrapper_8_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@42452.4]
  assign RetimeWrapper_8_io_in = x824_x523_D1_0_number[7:0]; // @[package.scala 94:16:@42451.4]
  assign RetimeWrapper_9_clock = clock; // @[:@42460.4]
  assign RetimeWrapper_9_reset = reset; // @[:@42461.4]
  assign RetimeWrapper_9_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@42463.4]
  assign RetimeWrapper_9_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@42462.4]
  assign x540_rdcol_1_clock = clock; // @[:@42483.4]
  assign x540_rdcol_1_reset = reset; // @[:@42484.4]
  assign x540_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@42485.4]
  assign x540_rdcol_1_io_b = 32'h1; // @[Math.scala 152:17:@42486.4]
  assign x540_rdcol_1_io_flow = io_in_x481_TREADY; // @[Math.scala 153:20:@42487.4]
  assign x542_1_clock = clock; // @[:@42497.4]
  assign x542_1_reset = reset; // @[:@42498.4]
  assign x542_1_io_a = x540_rdcol_1_io_result; // @[Math.scala 367:17:@42499.4]
  assign x542_1_io_flow = io_in_x481_TREADY; // @[Math.scala 369:20:@42501.4]
  assign x543_div_1_clock = clock; // @[:@42509.4]
  assign x543_div_1_reset = reset; // @[:@42510.4]
  assign x543_div_1_io_a = x540_rdcol_1_io_result; // @[Math.scala 328:17:@42511.4]
  assign x543_div_1_io_flow = io_in_x481_TREADY; // @[Math.scala 330:20:@42513.4]
  assign RetimeWrapper_10_clock = clock; // @[:@42519.4]
  assign RetimeWrapper_10_reset = reset; // @[:@42520.4]
  assign RetimeWrapper_10_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@42522.4]
  assign RetimeWrapper_10_io_in = x803_sum_1_io_result; // @[package.scala 94:16:@42521.4]
  assign x544_sum_1_clock = clock; // @[:@42528.4]
  assign x544_sum_1_reset = reset; // @[:@42529.4]
  assign x544_sum_1_io_a = RetimeWrapper_10_io_out; // @[Math.scala 151:17:@42530.4]
  assign x544_sum_1_io_b = x543_div_1_io_result; // @[Math.scala 152:17:@42531.4]
  assign x544_sum_1_io_flow = io_in_x481_TREADY; // @[Math.scala 153:20:@42532.4]
  assign RetimeWrapper_11_clock = clock; // @[:@42538.4]
  assign RetimeWrapper_11_reset = reset; // @[:@42539.4]
  assign RetimeWrapper_11_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@42541.4]
  assign RetimeWrapper_11_io_in = x542_1_io_result; // @[package.scala 94:16:@42540.4]
  assign RetimeWrapper_12_clock = clock; // @[:@42547.4]
  assign RetimeWrapper_12_reset = reset; // @[:@42548.4]
  assign RetimeWrapper_12_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@42550.4]
  assign RetimeWrapper_12_io_in = x824_x523_D1_0_number[15:8]; // @[package.scala 94:16:@42549.4]
  assign RetimeWrapper_13_clock = clock; // @[:@42556.4]
  assign RetimeWrapper_13_reset = reset; // @[:@42557.4]
  assign RetimeWrapper_13_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@42559.4]
  assign RetimeWrapper_13_io_in = x544_sum_1_io_result; // @[package.scala 94:16:@42558.4]
  assign RetimeWrapper_14_clock = clock; // @[:@42567.4]
  assign RetimeWrapper_14_reset = reset; // @[:@42568.4]
  assign RetimeWrapper_14_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@42570.4]
  assign RetimeWrapper_14_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@42569.4]
  assign x546_rdcol_1_clock = clock; // @[:@42590.4]
  assign x546_rdcol_1_reset = reset; // @[:@42591.4]
  assign x546_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@42592.4]
  assign x546_rdcol_1_io_b = 32'h2; // @[Math.scala 152:17:@42593.4]
  assign x546_rdcol_1_io_flow = io_in_x481_TREADY; // @[Math.scala 153:20:@42594.4]
  assign x548_1_clock = clock; // @[:@42604.4]
  assign x548_1_reset = reset; // @[:@42605.4]
  assign x548_1_io_a = x546_rdcol_1_io_result; // @[Math.scala 367:17:@42606.4]
  assign x548_1_io_flow = io_in_x481_TREADY; // @[Math.scala 369:20:@42608.4]
  assign x549_div_1_clock = clock; // @[:@42616.4]
  assign x549_div_1_reset = reset; // @[:@42617.4]
  assign x549_div_1_io_a = x546_rdcol_1_io_result; // @[Math.scala 328:17:@42618.4]
  assign x549_div_1_io_flow = io_in_x481_TREADY; // @[Math.scala 330:20:@42620.4]
  assign x550_sum_1_clock = clock; // @[:@42626.4]
  assign x550_sum_1_reset = reset; // @[:@42627.4]
  assign x550_sum_1_io_a = RetimeWrapper_10_io_out; // @[Math.scala 151:17:@42628.4]
  assign x550_sum_1_io_b = x549_div_1_io_result; // @[Math.scala 152:17:@42629.4]
  assign x550_sum_1_io_flow = io_in_x481_TREADY; // @[Math.scala 153:20:@42630.4]
  assign RetimeWrapper_15_clock = clock; // @[:@42636.4]
  assign RetimeWrapper_15_reset = reset; // @[:@42637.4]
  assign RetimeWrapper_15_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@42639.4]
  assign RetimeWrapper_15_io_in = x550_sum_1_io_result; // @[package.scala 94:16:@42638.4]
  assign RetimeWrapper_16_clock = clock; // @[:@42645.4]
  assign RetimeWrapper_16_reset = reset; // @[:@42646.4]
  assign RetimeWrapper_16_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@42648.4]
  assign RetimeWrapper_16_io_in = x824_x523_D1_0_number[23:16]; // @[package.scala 94:16:@42647.4]
  assign RetimeWrapper_17_clock = clock; // @[:@42654.4]
  assign RetimeWrapper_17_reset = reset; // @[:@42655.4]
  assign RetimeWrapper_17_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@42657.4]
  assign RetimeWrapper_17_io_in = x548_1_io_result; // @[package.scala 94:16:@42656.4]
  assign RetimeWrapper_18_clock = clock; // @[:@42665.4]
  assign RetimeWrapper_18_reset = reset; // @[:@42666.4]
  assign RetimeWrapper_18_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@42668.4]
  assign RetimeWrapper_18_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@42667.4]
  assign x552_rdcol_1_clock = clock; // @[:@42688.4]
  assign x552_rdcol_1_reset = reset; // @[:@42689.4]
  assign x552_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@42690.4]
  assign x552_rdcol_1_io_b = 32'h3; // @[Math.scala 152:17:@42691.4]
  assign x552_rdcol_1_io_flow = io_in_x481_TREADY; // @[Math.scala 153:20:@42692.4]
  assign x554_1_clock = clock; // @[:@42704.4]
  assign x554_1_reset = reset; // @[:@42705.4]
  assign x554_1_io_a = x552_rdcol_1_io_result; // @[Math.scala 367:17:@42706.4]
  assign x554_1_io_flow = io_in_x481_TREADY; // @[Math.scala 369:20:@42708.4]
  assign x555_div_1_clock = clock; // @[:@42716.4]
  assign x555_div_1_reset = reset; // @[:@42717.4]
  assign x555_div_1_io_a = x552_rdcol_1_io_result; // @[Math.scala 328:17:@42718.4]
  assign x555_div_1_io_flow = io_in_x481_TREADY; // @[Math.scala 330:20:@42720.4]
  assign x556_sum_1_clock = clock; // @[:@42726.4]
  assign x556_sum_1_reset = reset; // @[:@42727.4]
  assign x556_sum_1_io_a = RetimeWrapper_10_io_out; // @[Math.scala 151:17:@42728.4]
  assign x556_sum_1_io_b = x555_div_1_io_result; // @[Math.scala 152:17:@42729.4]
  assign x556_sum_1_io_flow = io_in_x481_TREADY; // @[Math.scala 153:20:@42730.4]
  assign RetimeWrapper_19_clock = clock; // @[:@42736.4]
  assign RetimeWrapper_19_reset = reset; // @[:@42737.4]
  assign RetimeWrapper_19_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@42739.4]
  assign RetimeWrapper_19_io_in = x554_1_io_result; // @[package.scala 94:16:@42738.4]
  assign RetimeWrapper_20_clock = clock; // @[:@42745.4]
  assign RetimeWrapper_20_reset = reset; // @[:@42746.4]
  assign RetimeWrapper_20_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@42748.4]
  assign RetimeWrapper_20_io_in = x824_x523_D1_0_number[31:24]; // @[package.scala 94:16:@42747.4]
  assign RetimeWrapper_21_clock = clock; // @[:@42754.4]
  assign RetimeWrapper_21_reset = reset; // @[:@42755.4]
  assign RetimeWrapper_21_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@42757.4]
  assign RetimeWrapper_21_io_in = x556_sum_1_io_result; // @[package.scala 94:16:@42756.4]
  assign RetimeWrapper_22_clock = clock; // @[:@42765.4]
  assign RetimeWrapper_22_reset = reset; // @[:@42766.4]
  assign RetimeWrapper_22_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@42768.4]
  assign RetimeWrapper_22_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@42767.4]
  assign RetimeWrapper_23_clock = clock; // @[:@42786.4]
  assign RetimeWrapper_23_reset = reset; // @[:@42787.4]
  assign RetimeWrapper_23_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@42789.4]
  assign RetimeWrapper_23_io_in = __io_result; // @[package.scala 94:16:@42788.4]
  assign RetimeWrapper_24_clock = clock; // @[:@42802.4]
  assign RetimeWrapper_24_reset = reset; // @[:@42803.4]
  assign RetimeWrapper_24_io_flow = io_in_x481_TREADY; // @[package.scala 95:18:@42806.4]
  assign RetimeWrapper_24_io_in = $unsigned(_T_554); // @[package.scala 94:16:@42805.4]
  assign RetimeWrapper_25_clock = clock; // @[:@42820.4]
  assign RetimeWrapper_25_reset = reset; // @[:@42821.4]
  assign RetimeWrapper_25_io_flow = io_in_x481_TREADY; // @[package.scala 95:18:@42823.4]
  assign RetimeWrapper_25_io_in = $signed(_T_551) < $signed(32'sh0); // @[package.scala 94:16:@42822.4]
  assign RetimeWrapper_26_clock = clock; // @[:@42829.4]
  assign RetimeWrapper_26_reset = reset; // @[:@42830.4]
  assign RetimeWrapper_26_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@42832.4]
  assign RetimeWrapper_26_io_in = x552_rdcol_1_io_result; // @[package.scala 94:16:@42831.4]
  assign RetimeWrapper_27_clock = clock; // @[:@42843.4]
  assign RetimeWrapper_27_reset = reset; // @[:@42844.4]
  assign RetimeWrapper_27_io_flow = io_in_x481_TREADY; // @[package.scala 95:18:@42846.4]
  assign RetimeWrapper_27_io_in = $signed(_T_578) < $signed(32'sh0); // @[package.scala 94:16:@42845.4]
  assign RetimeWrapper_28_clock = clock; // @[:@42852.4]
  assign RetimeWrapper_28_reset = reset; // @[:@42853.4]
  assign RetimeWrapper_28_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@42855.4]
  assign RetimeWrapper_28_io_in = RetimeWrapper_25_io_out; // @[package.scala 94:16:@42854.4]
  assign x808_sum_1_clock = clock; // @[:@42897.4]
  assign x808_sum_1_reset = reset; // @[:@42898.4]
  assign x808_sum_1_io_a = _T_615[31:0]; // @[Math.scala 151:17:@42899.4]
  assign x808_sum_1_io_b = _T_619[31:0]; // @[Math.scala 152:17:@42900.4]
  assign x808_sum_1_io_flow = io_in_x481_TREADY; // @[Math.scala 153:20:@42901.4]
  assign RetimeWrapper_29_clock = clock; // @[:@42907.4]
  assign RetimeWrapper_29_reset = reset; // @[:@42908.4]
  assign RetimeWrapper_29_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@42910.4]
  assign RetimeWrapper_29_io_in = x808_sum_1_io_result; // @[package.scala 94:16:@42909.4]
  assign RetimeWrapper_30_clock = clock; // @[:@42916.4]
  assign RetimeWrapper_30_reset = reset; // @[:@42917.4]
  assign RetimeWrapper_30_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@42919.4]
  assign RetimeWrapper_30_io_in = x555_div_1_io_result; // @[package.scala 94:16:@42918.4]
  assign x567_sum_1_clock = clock; // @[:@42925.4]
  assign x567_sum_1_reset = reset; // @[:@42926.4]
  assign x567_sum_1_io_a = RetimeWrapper_29_io_out; // @[Math.scala 151:17:@42927.4]
  assign x567_sum_1_io_b = RetimeWrapper_30_io_out; // @[Math.scala 152:17:@42928.4]
  assign x567_sum_1_io_flow = io_in_x481_TREADY; // @[Math.scala 153:20:@42929.4]
  assign RetimeWrapper_31_clock = clock; // @[:@42935.4]
  assign RetimeWrapper_31_reset = reset; // @[:@42936.4]
  assign RetimeWrapper_31_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@42938.4]
  assign RetimeWrapper_31_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@42937.4]
  assign RetimeWrapper_32_clock = clock; // @[:@42944.4]
  assign RetimeWrapper_32_reset = reset; // @[:@42945.4]
  assign RetimeWrapper_32_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@42947.4]
  assign RetimeWrapper_32_io_in = x554_1_io_result; // @[package.scala 94:16:@42946.4]
  assign RetimeWrapper_33_clock = clock; // @[:@42953.4]
  assign RetimeWrapper_33_reset = reset; // @[:@42954.4]
  assign RetimeWrapper_33_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@42956.4]
  assign RetimeWrapper_33_io_in = $unsigned(_T_600); // @[package.scala 94:16:@42955.4]
  assign RetimeWrapper_34_clock = clock; // @[:@42962.4]
  assign RetimeWrapper_34_reset = reset; // @[:@42963.4]
  assign RetimeWrapper_34_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@42965.4]
  assign RetimeWrapper_34_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@42964.4]
  assign RetimeWrapper_35_clock = clock; // @[:@42971.4]
  assign RetimeWrapper_35_reset = reset; // @[:@42972.4]
  assign RetimeWrapper_35_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@42974.4]
  assign RetimeWrapper_35_io_in = ~ x562; // @[package.scala 94:16:@42973.4]
  assign RetimeWrapper_36_clock = clock; // @[:@42983.4]
  assign RetimeWrapper_36_reset = reset; // @[:@42984.4]
  assign RetimeWrapper_36_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@42986.4]
  assign RetimeWrapper_36_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@42985.4]
  assign RetimeWrapper_37_clock = clock; // @[:@43004.4]
  assign RetimeWrapper_37_reset = reset; // @[:@43005.4]
  assign RetimeWrapper_37_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@43007.4]
  assign RetimeWrapper_37_io_in = x546_rdcol_1_io_result; // @[package.scala 94:16:@43006.4]
  assign RetimeWrapper_38_clock = clock; // @[:@43018.4]
  assign RetimeWrapper_38_reset = reset; // @[:@43019.4]
  assign RetimeWrapper_38_io_flow = io_in_x481_TREADY; // @[package.scala 95:18:@43021.4]
  assign RetimeWrapper_38_io_in = $signed(_T_674) < $signed(32'sh0); // @[package.scala 94:16:@43020.4]
  assign RetimeWrapper_39_clock = clock; // @[:@43033.4]
  assign RetimeWrapper_39_reset = reset; // @[:@43034.4]
  assign RetimeWrapper_39_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@43036.4]
  assign RetimeWrapper_39_io_in = x549_div_1_io_result; // @[package.scala 94:16:@43035.4]
  assign x573_sum_1_clock = clock; // @[:@43042.4]
  assign x573_sum_1_reset = reset; // @[:@43043.4]
  assign x573_sum_1_io_a = RetimeWrapper_29_io_out; // @[Math.scala 151:17:@43044.4]
  assign x573_sum_1_io_b = RetimeWrapper_39_io_out; // @[Math.scala 152:17:@43045.4]
  assign x573_sum_1_io_flow = io_in_x481_TREADY; // @[Math.scala 153:20:@43046.4]
  assign RetimeWrapper_40_clock = clock; // @[:@43052.4]
  assign RetimeWrapper_40_reset = reset; // @[:@43053.4]
  assign RetimeWrapper_40_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@43055.4]
  assign RetimeWrapper_40_io_in = ~ x571; // @[package.scala 94:16:@43054.4]
  assign RetimeWrapper_41_clock = clock; // @[:@43061.4]
  assign RetimeWrapper_41_reset = reset; // @[:@43062.4]
  assign RetimeWrapper_41_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@43064.4]
  assign RetimeWrapper_41_io_in = x548_1_io_result; // @[package.scala 94:16:@43063.4]
  assign RetimeWrapper_42_clock = clock; // @[:@43073.4]
  assign RetimeWrapper_42_reset = reset; // @[:@43074.4]
  assign RetimeWrapper_42_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@43076.4]
  assign RetimeWrapper_42_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@43075.4]
  assign RetimeWrapper_43_clock = clock; // @[:@43094.4]
  assign RetimeWrapper_43_reset = reset; // @[:@43095.4]
  assign RetimeWrapper_43_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@43097.4]
  assign RetimeWrapper_43_io_in = x540_rdcol_1_io_result; // @[package.scala 94:16:@43096.4]
  assign RetimeWrapper_44_clock = clock; // @[:@43108.4]
  assign RetimeWrapper_44_reset = reset; // @[:@43109.4]
  assign RetimeWrapper_44_io_flow = io_in_x481_TREADY; // @[package.scala 95:18:@43111.4]
  assign RetimeWrapper_44_io_in = $signed(_T_722) < $signed(32'sh0); // @[package.scala 94:16:@43110.4]
  assign RetimeWrapper_45_clock = clock; // @[:@43123.4]
  assign RetimeWrapper_45_reset = reset; // @[:@43124.4]
  assign RetimeWrapper_45_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@43126.4]
  assign RetimeWrapper_45_io_in = x543_div_1_io_result; // @[package.scala 94:16:@43125.4]
  assign x579_sum_1_clock = clock; // @[:@43132.4]
  assign x579_sum_1_reset = reset; // @[:@43133.4]
  assign x579_sum_1_io_a = RetimeWrapper_29_io_out; // @[Math.scala 151:17:@43134.4]
  assign x579_sum_1_io_b = RetimeWrapper_45_io_out; // @[Math.scala 152:17:@43135.4]
  assign x579_sum_1_io_flow = io_in_x481_TREADY; // @[Math.scala 153:20:@43136.4]
  assign RetimeWrapper_46_clock = clock; // @[:@43142.4]
  assign RetimeWrapper_46_reset = reset; // @[:@43143.4]
  assign RetimeWrapper_46_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@43145.4]
  assign RetimeWrapper_46_io_in = x542_1_io_result; // @[package.scala 94:16:@43144.4]
  assign RetimeWrapper_47_clock = clock; // @[:@43151.4]
  assign RetimeWrapper_47_reset = reset; // @[:@43152.4]
  assign RetimeWrapper_47_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@43154.4]
  assign RetimeWrapper_47_io_in = ~ x577; // @[package.scala 94:16:@43153.4]
  assign RetimeWrapper_48_clock = clock; // @[:@43163.4]
  assign RetimeWrapper_48_reset = reset; // @[:@43164.4]
  assign RetimeWrapper_48_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@43166.4]
  assign RetimeWrapper_48_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@43165.4]
  assign RetimeWrapper_49_clock = clock; // @[:@43184.4]
  assign RetimeWrapper_49_reset = reset; // @[:@43185.4]
  assign RetimeWrapper_49_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@43187.4]
  assign RetimeWrapper_49_io_in = __1_io_result; // @[package.scala 94:16:@43186.4]
  assign RetimeWrapper_50_clock = clock; // @[:@43200.4]
  assign RetimeWrapper_50_reset = reset; // @[:@43201.4]
  assign RetimeWrapper_50_io_flow = io_in_x481_TREADY; // @[package.scala 95:18:@43203.4]
  assign RetimeWrapper_50_io_in = $signed(_T_772) < $signed(32'sh0); // @[package.scala 94:16:@43202.4]
  assign RetimeWrapper_51_clock = clock; // @[:@43215.4]
  assign RetimeWrapper_51_reset = reset; // @[:@43216.4]
  assign RetimeWrapper_51_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@43218.4]
  assign RetimeWrapper_51_io_in = x808_sum_1_io_result; // @[package.scala 94:16:@43217.4]
  assign RetimeWrapper_52_clock = clock; // @[:@43224.4]
  assign RetimeWrapper_52_reset = reset; // @[:@43225.4]
  assign RetimeWrapper_52_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@43227.4]
  assign RetimeWrapper_52_io_in = x537_div_1_io_result; // @[package.scala 94:16:@43226.4]
  assign x585_sum_1_clock = clock; // @[:@43233.4]
  assign x585_sum_1_reset = reset; // @[:@43234.4]
  assign x585_sum_1_io_a = RetimeWrapper_51_io_out; // @[Math.scala 151:17:@43235.4]
  assign x585_sum_1_io_b = RetimeWrapper_52_io_out; // @[Math.scala 152:17:@43236.4]
  assign x585_sum_1_io_flow = io_in_x481_TREADY; // @[Math.scala 153:20:@43237.4]
  assign RetimeWrapper_53_clock = clock; // @[:@43243.4]
  assign RetimeWrapper_53_reset = reset; // @[:@43244.4]
  assign RetimeWrapper_53_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@43246.4]
  assign RetimeWrapper_53_io_in = x534_1_io_result; // @[package.scala 94:16:@43245.4]
  assign RetimeWrapper_54_clock = clock; // @[:@43252.4]
  assign RetimeWrapper_54_reset = reset; // @[:@43253.4]
  assign RetimeWrapper_54_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@43255.4]
  assign RetimeWrapper_54_io_in = ~ x583; // @[package.scala 94:16:@43254.4]
  assign RetimeWrapper_55_clock = clock; // @[:@43261.4]
  assign RetimeWrapper_55_reset = reset; // @[:@43262.4]
  assign RetimeWrapper_55_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@43264.4]
  assign RetimeWrapper_55_io_in = x585_sum_1_io_result; // @[package.scala 94:16:@43263.4]
  assign RetimeWrapper_56_clock = clock; // @[:@43273.4]
  assign RetimeWrapper_56_reset = reset; // @[:@43274.4]
  assign RetimeWrapper_56_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@43276.4]
  assign RetimeWrapper_56_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@43275.4]
  assign x588_rdcol_1_clock = clock; // @[:@43296.4]
  assign x588_rdcol_1_reset = reset; // @[:@43297.4]
  assign x588_rdcol_1_io_a = RetimeWrapper_49_io_out; // @[Math.scala 151:17:@43298.4]
  assign x588_rdcol_1_io_b = 32'hffffffff; // @[Math.scala 152:17:@43299.4]
  assign x588_rdcol_1_io_flow = io_in_x481_TREADY; // @[Math.scala 153:20:@43300.4]
  assign RetimeWrapper_57_clock = clock; // @[:@43311.4]
  assign RetimeWrapper_57_reset = reset; // @[:@43312.4]
  assign RetimeWrapper_57_io_flow = io_in_x481_TREADY; // @[package.scala 95:18:@43314.4]
  assign RetimeWrapper_57_io_in = $signed(_T_830) < $signed(32'sh0); // @[package.scala 94:16:@43313.4]
  assign x592_1_clock = clock; // @[:@43328.4]
  assign x592_1_reset = reset; // @[:@43329.4]
  assign x592_1_io_a = x588_rdcol_1_io_result; // @[Math.scala 367:17:@43330.4]
  assign x592_1_io_flow = io_in_x481_TREADY; // @[Math.scala 369:20:@43332.4]
  assign x593_div_1_clock = clock; // @[:@43340.4]
  assign x593_div_1_reset = reset; // @[:@43341.4]
  assign x593_div_1_io_a = x588_rdcol_1_io_result; // @[Math.scala 328:17:@43342.4]
  assign x593_div_1_io_flow = io_in_x481_TREADY; // @[Math.scala 330:20:@43344.4]
  assign x594_sum_1_clock = clock; // @[:@43350.4]
  assign x594_sum_1_reset = reset; // @[:@43351.4]
  assign x594_sum_1_io_a = RetimeWrapper_29_io_out; // @[Math.scala 151:17:@43352.4]
  assign x594_sum_1_io_b = x593_div_1_io_result; // @[Math.scala 152:17:@43353.4]
  assign x594_sum_1_io_flow = io_in_x481_TREADY; // @[Math.scala 153:20:@43354.4]
  assign RetimeWrapper_58_clock = clock; // @[:@43360.4]
  assign RetimeWrapper_58_reset = reset; // @[:@43361.4]
  assign RetimeWrapper_58_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@43363.4]
  assign RetimeWrapper_58_io_in = ~ x590; // @[package.scala 94:16:@43362.4]
  assign RetimeWrapper_59_clock = clock; // @[:@43369.4]
  assign RetimeWrapper_59_reset = reset; // @[:@43370.4]
  assign RetimeWrapper_59_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@43372.4]
  assign RetimeWrapper_59_io_in = x592_1_io_result; // @[package.scala 94:16:@43371.4]
  assign RetimeWrapper_60_clock = clock; // @[:@43381.4]
  assign RetimeWrapper_60_reset = reset; // @[:@43382.4]
  assign RetimeWrapper_60_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@43384.4]
  assign RetimeWrapper_60_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@43383.4]
  assign x597_rdcol_1_clock = clock; // @[:@43404.4]
  assign x597_rdcol_1_reset = reset; // @[:@43405.4]
  assign x597_rdcol_1_io_a = RetimeWrapper_49_io_out; // @[Math.scala 151:17:@43406.4]
  assign x597_rdcol_1_io_b = 32'hfffffffe; // @[Math.scala 152:17:@43407.4]
  assign x597_rdcol_1_io_flow = io_in_x481_TREADY; // @[Math.scala 153:20:@43408.4]
  assign RetimeWrapper_61_clock = clock; // @[:@43419.4]
  assign RetimeWrapper_61_reset = reset; // @[:@43420.4]
  assign RetimeWrapper_61_io_flow = io_in_x481_TREADY; // @[package.scala 95:18:@43422.4]
  assign RetimeWrapper_61_io_in = $signed(_T_893) < $signed(32'sh0); // @[package.scala 94:16:@43421.4]
  assign x601_1_clock = clock; // @[:@43436.4]
  assign x601_1_reset = reset; // @[:@43437.4]
  assign x601_1_io_a = x597_rdcol_1_io_result; // @[Math.scala 367:17:@43438.4]
  assign x601_1_io_flow = io_in_x481_TREADY; // @[Math.scala 369:20:@43440.4]
  assign x602_div_1_clock = clock; // @[:@43448.4]
  assign x602_div_1_reset = reset; // @[:@43449.4]
  assign x602_div_1_io_a = x597_rdcol_1_io_result; // @[Math.scala 328:17:@43450.4]
  assign x602_div_1_io_flow = io_in_x481_TREADY; // @[Math.scala 330:20:@43452.4]
  assign x603_sum_1_clock = clock; // @[:@43458.4]
  assign x603_sum_1_reset = reset; // @[:@43459.4]
  assign x603_sum_1_io_a = RetimeWrapper_29_io_out; // @[Math.scala 151:17:@43460.4]
  assign x603_sum_1_io_b = x602_div_1_io_result; // @[Math.scala 152:17:@43461.4]
  assign x603_sum_1_io_flow = io_in_x481_TREADY; // @[Math.scala 153:20:@43462.4]
  assign RetimeWrapper_62_clock = clock; // @[:@43468.4]
  assign RetimeWrapper_62_reset = reset; // @[:@43469.4]
  assign RetimeWrapper_62_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@43471.4]
  assign RetimeWrapper_62_io_in = x601_1_io_result; // @[package.scala 94:16:@43470.4]
  assign RetimeWrapper_63_clock = clock; // @[:@43477.4]
  assign RetimeWrapper_63_reset = reset; // @[:@43478.4]
  assign RetimeWrapper_63_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@43480.4]
  assign RetimeWrapper_63_io_in = ~ x599; // @[package.scala 94:16:@43479.4]
  assign RetimeWrapper_64_clock = clock; // @[:@43489.4]
  assign RetimeWrapper_64_reset = reset; // @[:@43490.4]
  assign RetimeWrapper_64_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@43492.4]
  assign RetimeWrapper_64_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@43491.4]
  assign x606_rdrow_1_clock = clock; // @[:@43512.4]
  assign x606_rdrow_1_reset = reset; // @[:@43513.4]
  assign x606_rdrow_1_io_a = RetimeWrapper_23_io_out; // @[Math.scala 192:17:@43514.4]
  assign x606_rdrow_1_io_b = 32'h1; // @[Math.scala 193:17:@43515.4]
  assign x606_rdrow_1_io_flow = io_in_x481_TREADY; // @[Math.scala 194:20:@43516.4]
  assign RetimeWrapper_65_clock = clock; // @[:@43529.4]
  assign RetimeWrapper_65_reset = reset; // @[:@43530.4]
  assign RetimeWrapper_65_io_flow = io_in_x481_TREADY; // @[package.scala 95:18:@43533.4]
  assign RetimeWrapper_65_io_in = $unsigned(_T_961); // @[package.scala 94:16:@43532.4]
  assign RetimeWrapper_66_clock = clock; // @[:@43547.4]
  assign RetimeWrapper_66_reset = reset; // @[:@43548.4]
  assign RetimeWrapper_66_io_flow = io_in_x481_TREADY; // @[package.scala 95:18:@43550.4]
  assign RetimeWrapper_66_io_in = $signed(_T_958) < $signed(32'sh0); // @[package.scala 94:16:@43549.4]
  assign x813_sum_1_clock = clock; // @[:@43592.4]
  assign x813_sum_1_reset = reset; // @[:@43593.4]
  assign x813_sum_1_io_a = _T_1006[31:0]; // @[Math.scala 151:17:@43594.4]
  assign x813_sum_1_io_b = _T_1010[31:0]; // @[Math.scala 152:17:@43595.4]
  assign x813_sum_1_io_flow = io_in_x481_TREADY; // @[Math.scala 153:20:@43596.4]
  assign RetimeWrapper_67_clock = clock; // @[:@43602.4]
  assign RetimeWrapper_67_reset = reset; // @[:@43603.4]
  assign RetimeWrapper_67_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@43605.4]
  assign RetimeWrapper_67_io_in = x813_sum_1_io_result; // @[package.scala 94:16:@43604.4]
  assign x614_sum_1_clock = clock; // @[:@43611.4]
  assign x614_sum_1_reset = reset; // @[:@43612.4]
  assign x614_sum_1_io_a = RetimeWrapper_67_io_out; // @[Math.scala 151:17:@43613.4]
  assign x614_sum_1_io_b = RetimeWrapper_30_io_out; // @[Math.scala 152:17:@43614.4]
  assign x614_sum_1_io_flow = io_in_x481_TREADY; // @[Math.scala 153:20:@43615.4]
  assign RetimeWrapper_68_clock = clock; // @[:@43621.4]
  assign RetimeWrapper_68_reset = reset; // @[:@43622.4]
  assign RetimeWrapper_68_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@43624.4]
  assign RetimeWrapper_68_io_in = $unsigned(_T_991); // @[package.scala 94:16:@43623.4]
  assign RetimeWrapper_69_clock = clock; // @[:@43630.4]
  assign RetimeWrapper_69_reset = reset; // @[:@43631.4]
  assign RetimeWrapper_69_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@43633.4]
  assign RetimeWrapper_69_io_in = ~ x609; // @[package.scala 94:16:@43632.4]
  assign RetimeWrapper_70_clock = clock; // @[:@43642.4]
  assign RetimeWrapper_70_reset = reset; // @[:@43643.4]
  assign RetimeWrapper_70_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@43645.4]
  assign RetimeWrapper_70_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@43644.4]
  assign x619_sum_1_clock = clock; // @[:@43671.4]
  assign x619_sum_1_reset = reset; // @[:@43672.4]
  assign x619_sum_1_io_a = RetimeWrapper_67_io_out; // @[Math.scala 151:17:@43673.4]
  assign x619_sum_1_io_b = RetimeWrapper_39_io_out; // @[Math.scala 152:17:@43674.4]
  assign x619_sum_1_io_flow = io_in_x481_TREADY; // @[Math.scala 153:20:@43675.4]
  assign RetimeWrapper_71_clock = clock; // @[:@43681.4]
  assign RetimeWrapper_71_reset = reset; // @[:@43682.4]
  assign RetimeWrapper_71_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@43684.4]
  assign RetimeWrapper_71_io_in = ~ x617; // @[package.scala 94:16:@43683.4]
  assign RetimeWrapper_72_clock = clock; // @[:@43693.4]
  assign RetimeWrapper_72_reset = reset; // @[:@43694.4]
  assign RetimeWrapper_72_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@43696.4]
  assign RetimeWrapper_72_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@43695.4]
  assign x624_sum_1_clock = clock; // @[:@43720.4]
  assign x624_sum_1_reset = reset; // @[:@43721.4]
  assign x624_sum_1_io_a = RetimeWrapper_67_io_out; // @[Math.scala 151:17:@43722.4]
  assign x624_sum_1_io_b = RetimeWrapper_45_io_out; // @[Math.scala 152:17:@43723.4]
  assign x624_sum_1_io_flow = io_in_x481_TREADY; // @[Math.scala 153:20:@43724.4]
  assign RetimeWrapper_73_clock = clock; // @[:@43730.4]
  assign RetimeWrapper_73_reset = reset; // @[:@43731.4]
  assign RetimeWrapper_73_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@43733.4]
  assign RetimeWrapper_73_io_in = ~ x622; // @[package.scala 94:16:@43732.4]
  assign RetimeWrapper_74_clock = clock; // @[:@43742.4]
  assign RetimeWrapper_74_reset = reset; // @[:@43743.4]
  assign RetimeWrapper_74_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@43745.4]
  assign RetimeWrapper_74_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@43744.4]
  assign RetimeWrapper_75_clock = clock; // @[:@43763.4]
  assign RetimeWrapper_75_reset = reset; // @[:@43764.4]
  assign RetimeWrapper_75_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@43766.4]
  assign RetimeWrapper_75_io_in = RetimeWrapper_50_io_out; // @[package.scala 94:16:@43765.4]
  assign RetimeWrapper_76_clock = clock; // @[:@43778.4]
  assign RetimeWrapper_76_reset = reset; // @[:@43779.4]
  assign RetimeWrapper_76_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@43781.4]
  assign RetimeWrapper_76_io_in = x813_sum_1_io_result; // @[package.scala 94:16:@43780.4]
  assign x629_sum_1_clock = clock; // @[:@43787.4]
  assign x629_sum_1_reset = reset; // @[:@43788.4]
  assign x629_sum_1_io_a = RetimeWrapper_76_io_out; // @[Math.scala 151:17:@43789.4]
  assign x629_sum_1_io_b = RetimeWrapper_52_io_out; // @[Math.scala 152:17:@43790.4]
  assign x629_sum_1_io_flow = io_in_x481_TREADY; // @[Math.scala 153:20:@43791.4]
  assign RetimeWrapper_77_clock = clock; // @[:@43797.4]
  assign RetimeWrapper_77_reset = reset; // @[:@43798.4]
  assign RetimeWrapper_77_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@43800.4]
  assign RetimeWrapper_77_io_in = x629_sum_1_io_result; // @[package.scala 94:16:@43799.4]
  assign RetimeWrapper_78_clock = clock; // @[:@43806.4]
  assign RetimeWrapper_78_reset = reset; // @[:@43807.4]
  assign RetimeWrapper_78_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@43809.4]
  assign RetimeWrapper_78_io_in = ~ x627; // @[package.scala 94:16:@43808.4]
  assign RetimeWrapper_79_clock = clock; // @[:@43818.4]
  assign RetimeWrapper_79_reset = reset; // @[:@43819.4]
  assign RetimeWrapper_79_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@43821.4]
  assign RetimeWrapper_79_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@43820.4]
  assign x634_sum_1_clock = clock; // @[:@43845.4]
  assign x634_sum_1_reset = reset; // @[:@43846.4]
  assign x634_sum_1_io_a = RetimeWrapper_67_io_out; // @[Math.scala 151:17:@43847.4]
  assign x634_sum_1_io_b = x593_div_1_io_result; // @[Math.scala 152:17:@43848.4]
  assign x634_sum_1_io_flow = io_in_x481_TREADY; // @[Math.scala 153:20:@43849.4]
  assign RetimeWrapper_80_clock = clock; // @[:@43855.4]
  assign RetimeWrapper_80_reset = reset; // @[:@43856.4]
  assign RetimeWrapper_80_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@43858.4]
  assign RetimeWrapper_80_io_in = ~ x632; // @[package.scala 94:16:@43857.4]
  assign RetimeWrapper_81_clock = clock; // @[:@43867.4]
  assign RetimeWrapper_81_reset = reset; // @[:@43868.4]
  assign RetimeWrapper_81_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@43870.4]
  assign RetimeWrapper_81_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@43869.4]
  assign x639_sum_1_clock = clock; // @[:@43894.4]
  assign x639_sum_1_reset = reset; // @[:@43895.4]
  assign x639_sum_1_io_a = RetimeWrapper_67_io_out; // @[Math.scala 151:17:@43896.4]
  assign x639_sum_1_io_b = x602_div_1_io_result; // @[Math.scala 152:17:@43897.4]
  assign x639_sum_1_io_flow = io_in_x481_TREADY; // @[Math.scala 153:20:@43898.4]
  assign RetimeWrapper_82_clock = clock; // @[:@43904.4]
  assign RetimeWrapper_82_reset = reset; // @[:@43905.4]
  assign RetimeWrapper_82_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@43907.4]
  assign RetimeWrapper_82_io_in = ~ x637; // @[package.scala 94:16:@43906.4]
  assign RetimeWrapper_83_clock = clock; // @[:@43916.4]
  assign RetimeWrapper_83_reset = reset; // @[:@43917.4]
  assign RetimeWrapper_83_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@43919.4]
  assign RetimeWrapper_83_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@43918.4]
  assign x642_rdrow_1_clock = clock; // @[:@43939.4]
  assign x642_rdrow_1_reset = reset; // @[:@43940.4]
  assign x642_rdrow_1_io_a = RetimeWrapper_23_io_out; // @[Math.scala 192:17:@43941.4]
  assign x642_rdrow_1_io_b = 32'h2; // @[Math.scala 193:17:@43942.4]
  assign x642_rdrow_1_io_flow = io_in_x481_TREADY; // @[Math.scala 194:20:@43943.4]
  assign RetimeWrapper_84_clock = clock; // @[:@43956.4]
  assign RetimeWrapper_84_reset = reset; // @[:@43957.4]
  assign RetimeWrapper_84_io_flow = io_in_x481_TREADY; // @[package.scala 95:18:@43960.4]
  assign RetimeWrapper_84_io_in = $unsigned(_T_1218); // @[package.scala 94:16:@43959.4]
  assign RetimeWrapper_85_clock = clock; // @[:@43974.4]
  assign RetimeWrapper_85_reset = reset; // @[:@43975.4]
  assign RetimeWrapper_85_io_flow = io_in_x481_TREADY; // @[package.scala 95:18:@43977.4]
  assign RetimeWrapper_85_io_in = $signed(_T_1215) < $signed(32'sh0); // @[package.scala 94:16:@43976.4]
  assign x818_sum_1_clock = clock; // @[:@44019.4]
  assign x818_sum_1_reset = reset; // @[:@44020.4]
  assign x818_sum_1_io_a = _T_1263[31:0]; // @[Math.scala 151:17:@44021.4]
  assign x818_sum_1_io_b = _T_1267[31:0]; // @[Math.scala 152:17:@44022.4]
  assign x818_sum_1_io_flow = io_in_x481_TREADY; // @[Math.scala 153:20:@44023.4]
  assign RetimeWrapper_86_clock = clock; // @[:@44029.4]
  assign RetimeWrapper_86_reset = reset; // @[:@44030.4]
  assign RetimeWrapper_86_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44032.4]
  assign RetimeWrapper_86_io_in = x818_sum_1_io_result; // @[package.scala 94:16:@44031.4]
  assign x650_sum_1_clock = clock; // @[:@44038.4]
  assign x650_sum_1_reset = reset; // @[:@44039.4]
  assign x650_sum_1_io_a = RetimeWrapper_86_io_out; // @[Math.scala 151:17:@44040.4]
  assign x650_sum_1_io_b = RetimeWrapper_30_io_out; // @[Math.scala 152:17:@44041.4]
  assign x650_sum_1_io_flow = io_in_x481_TREADY; // @[Math.scala 153:20:@44042.4]
  assign RetimeWrapper_87_clock = clock; // @[:@44048.4]
  assign RetimeWrapper_87_reset = reset; // @[:@44049.4]
  assign RetimeWrapper_87_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44051.4]
  assign RetimeWrapper_87_io_in = ~ x645; // @[package.scala 94:16:@44050.4]
  assign RetimeWrapper_88_clock = clock; // @[:@44057.4]
  assign RetimeWrapper_88_reset = reset; // @[:@44058.4]
  assign RetimeWrapper_88_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44060.4]
  assign RetimeWrapper_88_io_in = $unsigned(_T_1248); // @[package.scala 94:16:@44059.4]
  assign RetimeWrapper_89_clock = clock; // @[:@44069.4]
  assign RetimeWrapper_89_reset = reset; // @[:@44070.4]
  assign RetimeWrapper_89_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44072.4]
  assign RetimeWrapper_89_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@44071.4]
  assign x655_sum_1_clock = clock; // @[:@44098.4]
  assign x655_sum_1_reset = reset; // @[:@44099.4]
  assign x655_sum_1_io_a = RetimeWrapper_86_io_out; // @[Math.scala 151:17:@44100.4]
  assign x655_sum_1_io_b = RetimeWrapper_39_io_out; // @[Math.scala 152:17:@44101.4]
  assign x655_sum_1_io_flow = io_in_x481_TREADY; // @[Math.scala 153:20:@44102.4]
  assign RetimeWrapper_90_clock = clock; // @[:@44108.4]
  assign RetimeWrapper_90_reset = reset; // @[:@44109.4]
  assign RetimeWrapper_90_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44111.4]
  assign RetimeWrapper_90_io_in = ~ x653; // @[package.scala 94:16:@44110.4]
  assign RetimeWrapper_91_clock = clock; // @[:@44120.4]
  assign RetimeWrapper_91_reset = reset; // @[:@44121.4]
  assign RetimeWrapper_91_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44123.4]
  assign RetimeWrapper_91_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@44122.4]
  assign x660_sum_1_clock = clock; // @[:@44147.4]
  assign x660_sum_1_reset = reset; // @[:@44148.4]
  assign x660_sum_1_io_a = RetimeWrapper_86_io_out; // @[Math.scala 151:17:@44149.4]
  assign x660_sum_1_io_b = RetimeWrapper_45_io_out; // @[Math.scala 152:17:@44150.4]
  assign x660_sum_1_io_flow = io_in_x481_TREADY; // @[Math.scala 153:20:@44151.4]
  assign RetimeWrapper_92_clock = clock; // @[:@44157.4]
  assign RetimeWrapper_92_reset = reset; // @[:@44158.4]
  assign RetimeWrapper_92_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44160.4]
  assign RetimeWrapper_92_io_in = ~ x658; // @[package.scala 94:16:@44159.4]
  assign RetimeWrapper_93_clock = clock; // @[:@44169.4]
  assign RetimeWrapper_93_reset = reset; // @[:@44170.4]
  assign RetimeWrapper_93_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44172.4]
  assign RetimeWrapper_93_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@44171.4]
  assign RetimeWrapper_94_clock = clock; // @[:@44196.4]
  assign RetimeWrapper_94_reset = reset; // @[:@44197.4]
  assign RetimeWrapper_94_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44199.4]
  assign RetimeWrapper_94_io_in = x818_sum_1_io_result; // @[package.scala 94:16:@44198.4]
  assign x665_sum_1_clock = clock; // @[:@44205.4]
  assign x665_sum_1_reset = reset; // @[:@44206.4]
  assign x665_sum_1_io_a = RetimeWrapper_94_io_out; // @[Math.scala 151:17:@44207.4]
  assign x665_sum_1_io_b = RetimeWrapper_52_io_out; // @[Math.scala 152:17:@44208.4]
  assign x665_sum_1_io_flow = io_in_x481_TREADY; // @[Math.scala 153:20:@44209.4]
  assign RetimeWrapper_95_clock = clock; // @[:@44215.4]
  assign RetimeWrapper_95_reset = reset; // @[:@44216.4]
  assign RetimeWrapper_95_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44218.4]
  assign RetimeWrapper_95_io_in = x665_sum_1_io_result; // @[package.scala 94:16:@44217.4]
  assign RetimeWrapper_96_clock = clock; // @[:@44224.4]
  assign RetimeWrapper_96_reset = reset; // @[:@44225.4]
  assign RetimeWrapper_96_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44227.4]
  assign RetimeWrapper_96_io_in = ~ x663; // @[package.scala 94:16:@44226.4]
  assign RetimeWrapper_97_clock = clock; // @[:@44236.4]
  assign RetimeWrapper_97_reset = reset; // @[:@44237.4]
  assign RetimeWrapper_97_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44239.4]
  assign RetimeWrapper_97_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@44238.4]
  assign x670_sum_1_clock = clock; // @[:@44263.4]
  assign x670_sum_1_reset = reset; // @[:@44264.4]
  assign x670_sum_1_io_a = RetimeWrapper_86_io_out; // @[Math.scala 151:17:@44265.4]
  assign x670_sum_1_io_b = x593_div_1_io_result; // @[Math.scala 152:17:@44266.4]
  assign x670_sum_1_io_flow = io_in_x481_TREADY; // @[Math.scala 153:20:@44267.4]
  assign RetimeWrapper_98_clock = clock; // @[:@44273.4]
  assign RetimeWrapper_98_reset = reset; // @[:@44274.4]
  assign RetimeWrapper_98_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44276.4]
  assign RetimeWrapper_98_io_in = ~ x668; // @[package.scala 94:16:@44275.4]
  assign RetimeWrapper_99_clock = clock; // @[:@44285.4]
  assign RetimeWrapper_99_reset = reset; // @[:@44286.4]
  assign RetimeWrapper_99_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44288.4]
  assign RetimeWrapper_99_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@44287.4]
  assign x675_sum_1_clock = clock; // @[:@44312.4]
  assign x675_sum_1_reset = reset; // @[:@44313.4]
  assign x675_sum_1_io_a = RetimeWrapper_86_io_out; // @[Math.scala 151:17:@44314.4]
  assign x675_sum_1_io_b = x602_div_1_io_result; // @[Math.scala 152:17:@44315.4]
  assign x675_sum_1_io_flow = io_in_x481_TREADY; // @[Math.scala 153:20:@44316.4]
  assign RetimeWrapper_100_clock = clock; // @[:@44322.4]
  assign RetimeWrapper_100_reset = reset; // @[:@44323.4]
  assign RetimeWrapper_100_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44325.4]
  assign RetimeWrapper_100_io_in = ~ x673; // @[package.scala 94:16:@44324.4]
  assign RetimeWrapper_101_clock = clock; // @[:@44334.4]
  assign RetimeWrapper_101_reset = reset; // @[:@44335.4]
  assign RetimeWrapper_101_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44337.4]
  assign RetimeWrapper_101_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@44336.4]
  assign RetimeWrapper_102_clock = clock; // @[:@44357.4]
  assign RetimeWrapper_102_reset = reset; // @[:@44358.4]
  assign RetimeWrapper_102_io_flow = io_in_x481_TREADY; // @[package.scala 95:18:@44360.4]
  assign RetimeWrapper_102_io_in = _GEN_8 << 1; // @[package.scala 94:16:@44359.4]
  assign RetimeWrapper_103_clock = clock; // @[:@44369.4]
  assign RetimeWrapper_103_reset = reset; // @[:@44370.4]
  assign RetimeWrapper_103_io_flow = io_in_x481_TREADY; // @[package.scala 95:18:@44372.4]
  assign RetimeWrapper_103_io_in = _GEN_9 << 1; // @[package.scala 94:16:@44371.4]
  assign RetimeWrapper_104_clock = clock; // @[:@44381.4]
  assign RetimeWrapper_104_reset = reset; // @[:@44382.4]
  assign RetimeWrapper_104_io_flow = io_in_x481_TREADY; // @[package.scala 95:18:@44384.4]
  assign RetimeWrapper_104_io_in = _GEN_10 << 2; // @[package.scala 94:16:@44383.4]
  assign RetimeWrapper_105_clock = clock; // @[:@44393.4]
  assign RetimeWrapper_105_reset = reset; // @[:@44394.4]
  assign RetimeWrapper_105_io_flow = io_in_x481_TREADY; // @[package.scala 95:18:@44396.4]
  assign RetimeWrapper_105_io_in = _GEN_11 << 1; // @[package.scala 94:16:@44395.4]
  assign RetimeWrapper_106_clock = clock; // @[:@44405.4]
  assign RetimeWrapper_106_reset = reset; // @[:@44406.4]
  assign RetimeWrapper_106_io_flow = io_in_x481_TREADY; // @[package.scala 95:18:@44408.4]
  assign RetimeWrapper_106_io_in = _GEN_12 << 1; // @[package.scala 94:16:@44407.4]
  assign RetimeWrapper_107_clock = clock; // @[:@44415.4]
  assign RetimeWrapper_107_reset = reset; // @[:@44416.4]
  assign RetimeWrapper_107_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44418.4]
  assign RetimeWrapper_107_io_in = x525_lb_0_io_rPort_14_output_0; // @[package.scala 94:16:@44417.4]
  assign x683_x15_1_io_a = RetimeWrapper_107_io_out; // @[Math.scala 151:17:@44426.4]
  assign x683_x15_1_io_b = _T_1460[7:0]; // @[Math.scala 152:17:@44427.4]
  assign RetimeWrapper_108_clock = clock; // @[:@44434.4]
  assign RetimeWrapper_108_reset = reset; // @[:@44435.4]
  assign RetimeWrapper_108_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44437.4]
  assign RetimeWrapper_108_io_in = x525_lb_0_io_rPort_9_output_0; // @[package.scala 94:16:@44436.4]
  assign x684_x16_1_io_a = RetimeWrapper_108_io_out; // @[Math.scala 151:17:@44445.4]
  assign x684_x16_1_io_b = _T_1466[7:0]; // @[Math.scala 152:17:@44446.4]
  assign x685_x15_1_io_a = _T_1472[7:0]; // @[Math.scala 151:17:@44455.4]
  assign x685_x15_1_io_b = _T_1478[7:0]; // @[Math.scala 152:17:@44456.4]
  assign RetimeWrapper_109_clock = clock; // @[:@44463.4]
  assign RetimeWrapper_109_reset = reset; // @[:@44464.4]
  assign RetimeWrapper_109_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44466.4]
  assign RetimeWrapper_109_io_in = x525_lb_0_io_rPort_1_output_0; // @[package.scala 94:16:@44465.4]
  assign x686_x16_1_io_a = RetimeWrapper_109_io_out; // @[Math.scala 151:17:@44474.4]
  assign x686_x16_1_io_b = _T_1484[7:0]; // @[Math.scala 152:17:@44475.4]
  assign x687_x15_1_io_a = x683_x15_1_io_result; // @[Math.scala 151:17:@44484.4]
  assign x687_x15_1_io_b = x684_x16_1_io_result; // @[Math.scala 152:17:@44485.4]
  assign x688_x16_1_io_a = x685_x15_1_io_result; // @[Math.scala 151:17:@44494.4]
  assign x688_x16_1_io_b = x686_x16_1_io_result; // @[Math.scala 152:17:@44495.4]
  assign x689_x15_1_io_a = x687_x15_1_io_result; // @[Math.scala 151:17:@44506.4]
  assign x689_x15_1_io_b = x688_x16_1_io_result; // @[Math.scala 152:17:@44507.4]
  assign RetimeWrapper_110_clock = clock; // @[:@44514.4]
  assign RetimeWrapper_110_reset = reset; // @[:@44515.4]
  assign RetimeWrapper_110_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44517.4]
  assign RetimeWrapper_110_io_in = x525_lb_0_io_rPort_3_output_0; // @[package.scala 94:16:@44516.4]
  assign x690_sum_1_clock = clock; // @[:@44523.4]
  assign x690_sum_1_reset = reset; // @[:@44524.4]
  assign x690_sum_1_io_a = x689_x15_1_io_result; // @[Math.scala 151:17:@44525.4]
  assign x690_sum_1_io_b = RetimeWrapper_110_io_out; // @[Math.scala 152:17:@44526.4]
  assign x690_sum_1_io_flow = io_in_x481_TREADY; // @[Math.scala 153:20:@44527.4]
  assign RetimeWrapper_111_clock = clock; // @[:@44542.4]
  assign RetimeWrapper_111_reset = reset; // @[:@44543.4]
  assign RetimeWrapper_111_io_flow = io_in_x481_TREADY; // @[package.scala 95:18:@44545.4]
  assign RetimeWrapper_111_io_in = _GEN_13 << 1; // @[package.scala 94:16:@44544.4]
  assign RetimeWrapper_112_clock = clock; // @[:@44554.4]
  assign RetimeWrapper_112_reset = reset; // @[:@44555.4]
  assign RetimeWrapper_112_io_flow = io_in_x481_TREADY; // @[package.scala 95:18:@44557.4]
  assign RetimeWrapper_112_io_in = _GEN_14 << 1; // @[package.scala 94:16:@44556.4]
  assign RetimeWrapper_113_clock = clock; // @[:@44566.4]
  assign RetimeWrapper_113_reset = reset; // @[:@44567.4]
  assign RetimeWrapper_113_io_flow = io_in_x481_TREADY; // @[package.scala 95:18:@44569.4]
  assign RetimeWrapper_113_io_in = _GEN_15 << 2; // @[package.scala 94:16:@44568.4]
  assign RetimeWrapper_114_clock = clock; // @[:@44578.4]
  assign RetimeWrapper_114_reset = reset; // @[:@44579.4]
  assign RetimeWrapper_114_io_flow = io_in_x481_TREADY; // @[package.scala 95:18:@44581.4]
  assign RetimeWrapper_114_io_in = _GEN_16 << 1; // @[package.scala 94:16:@44580.4]
  assign RetimeWrapper_115_clock = clock; // @[:@44590.4]
  assign RetimeWrapper_115_reset = reset; // @[:@44591.4]
  assign RetimeWrapper_115_io_flow = io_in_x481_TREADY; // @[package.scala 95:18:@44593.4]
  assign RetimeWrapper_115_io_in = _GEN_17 << 1; // @[package.scala 94:16:@44592.4]
  assign RetimeWrapper_116_clock = clock; // @[:@44600.4]
  assign RetimeWrapper_116_reset = reset; // @[:@44601.4]
  assign RetimeWrapper_116_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44603.4]
  assign RetimeWrapper_116_io_in = x525_lb_0_io_rPort_2_output_0; // @[package.scala 94:16:@44602.4]
  assign x697_x15_1_io_a = RetimeWrapper_116_io_out; // @[Math.scala 151:17:@44611.4]
  assign x697_x15_1_io_b = _T_1538[7:0]; // @[Math.scala 152:17:@44612.4]
  assign RetimeWrapper_117_clock = clock; // @[:@44619.4]
  assign RetimeWrapper_117_reset = reset; // @[:@44620.4]
  assign RetimeWrapper_117_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44622.4]
  assign RetimeWrapper_117_io_in = x525_lb_0_io_rPort_7_output_0; // @[package.scala 94:16:@44621.4]
  assign x698_x16_1_io_a = RetimeWrapper_117_io_out; // @[Math.scala 151:17:@44630.4]
  assign x698_x16_1_io_b = _T_1544[7:0]; // @[Math.scala 152:17:@44631.4]
  assign x699_x15_1_io_a = _T_1550[7:0]; // @[Math.scala 151:17:@44640.4]
  assign x699_x15_1_io_b = _T_1556[7:0]; // @[Math.scala 152:17:@44641.4]
  assign RetimeWrapper_118_clock = clock; // @[:@44648.4]
  assign RetimeWrapper_118_reset = reset; // @[:@44649.4]
  assign RetimeWrapper_118_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44651.4]
  assign RetimeWrapper_118_io_in = x525_lb_0_io_rPort_11_output_0; // @[package.scala 94:16:@44650.4]
  assign x700_x16_1_io_a = RetimeWrapper_118_io_out; // @[Math.scala 151:17:@44659.4]
  assign x700_x16_1_io_b = _T_1562[7:0]; // @[Math.scala 152:17:@44660.4]
  assign x701_x15_1_io_a = x697_x15_1_io_result; // @[Math.scala 151:17:@44669.4]
  assign x701_x15_1_io_b = x698_x16_1_io_result; // @[Math.scala 152:17:@44670.4]
  assign x702_x16_1_io_a = x699_x15_1_io_result; // @[Math.scala 151:17:@44679.4]
  assign x702_x16_1_io_b = x700_x16_1_io_result; // @[Math.scala 152:17:@44680.4]
  assign x703_x15_1_io_a = x701_x15_1_io_result; // @[Math.scala 151:17:@44689.4]
  assign x703_x15_1_io_b = x702_x16_1_io_result; // @[Math.scala 152:17:@44690.4]
  assign RetimeWrapper_119_clock = clock; // @[:@44697.4]
  assign RetimeWrapper_119_reset = reset; // @[:@44698.4]
  assign RetimeWrapper_119_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44700.4]
  assign RetimeWrapper_119_io_in = x525_lb_0_io_rPort_0_output_0; // @[package.scala 94:16:@44699.4]
  assign x704_sum_1_clock = clock; // @[:@44706.4]
  assign x704_sum_1_reset = reset; // @[:@44707.4]
  assign x704_sum_1_io_a = x703_x15_1_io_result; // @[Math.scala 151:17:@44708.4]
  assign x704_sum_1_io_b = RetimeWrapper_119_io_out; // @[Math.scala 152:17:@44709.4]
  assign x704_sum_1_io_flow = io_in_x481_TREADY; // @[Math.scala 153:20:@44710.4]
  assign RetimeWrapper_120_clock = clock; // @[:@44725.4]
  assign RetimeWrapper_120_reset = reset; // @[:@44726.4]
  assign RetimeWrapper_120_io_flow = io_in_x481_TREADY; // @[package.scala 95:18:@44728.4]
  assign RetimeWrapper_120_io_in = _GEN_18 << 1; // @[package.scala 94:16:@44727.4]
  assign RetimeWrapper_121_clock = clock; // @[:@44737.4]
  assign RetimeWrapper_121_reset = reset; // @[:@44738.4]
  assign RetimeWrapper_121_io_flow = io_in_x481_TREADY; // @[package.scala 95:18:@44740.4]
  assign RetimeWrapper_121_io_in = _GEN_19 << 2; // @[package.scala 94:16:@44739.4]
  assign RetimeWrapper_122_clock = clock; // @[:@44749.4]
  assign RetimeWrapper_122_reset = reset; // @[:@44750.4]
  assign RetimeWrapper_122_io_flow = io_in_x481_TREADY; // @[package.scala 95:18:@44752.4]
  assign RetimeWrapper_122_io_in = _GEN_20 << 1; // @[package.scala 94:16:@44751.4]
  assign RetimeWrapper_123_clock = clock; // @[:@44761.4]
  assign RetimeWrapper_123_reset = reset; // @[:@44762.4]
  assign RetimeWrapper_123_io_flow = io_in_x481_TREADY; // @[package.scala 95:18:@44764.4]
  assign RetimeWrapper_123_io_in = _GEN_21 << 1; // @[package.scala 94:16:@44763.4]
  assign x710_x15_1_io_a = RetimeWrapper_108_io_out; // @[Math.scala 151:17:@44773.4]
  assign x710_x15_1_io_b = _T_1614[7:0]; // @[Math.scala 152:17:@44774.4]
  assign RetimeWrapper_124_clock = clock; // @[:@44781.4]
  assign RetimeWrapper_124_reset = reset; // @[:@44782.4]
  assign RetimeWrapper_124_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44784.4]
  assign RetimeWrapper_124_io_in = x525_lb_0_io_rPort_12_output_0; // @[package.scala 94:16:@44783.4]
  assign x711_x16_1_io_a = RetimeWrapper_124_io_out; // @[Math.scala 151:17:@44792.4]
  assign x711_x16_1_io_b = _T_1478[7:0]; // @[Math.scala 152:17:@44793.4]
  assign x712_x15_1_io_a = _T_1620[7:0]; // @[Math.scala 151:17:@44802.4]
  assign x712_x15_1_io_b = _T_1626[7:0]; // @[Math.scala 152:17:@44803.4]
  assign x713_x16_1_io_a = RetimeWrapper_110_io_out; // @[Math.scala 151:17:@44812.4]
  assign x713_x16_1_io_b = _T_1632[7:0]; // @[Math.scala 152:17:@44813.4]
  assign x714_x15_1_io_a = x710_x15_1_io_result; // @[Math.scala 151:17:@44822.4]
  assign x714_x15_1_io_b = x711_x16_1_io_result; // @[Math.scala 152:17:@44823.4]
  assign x715_x16_1_io_a = x712_x15_1_io_result; // @[Math.scala 151:17:@44832.4]
  assign x715_x16_1_io_b = x713_x16_1_io_result; // @[Math.scala 152:17:@44833.4]
  assign x716_x15_1_io_a = x714_x15_1_io_result; // @[Math.scala 151:17:@44842.4]
  assign x716_x15_1_io_b = x715_x16_1_io_result; // @[Math.scala 152:17:@44843.4]
  assign RetimeWrapper_125_clock = clock; // @[:@44850.4]
  assign RetimeWrapper_125_reset = reset; // @[:@44851.4]
  assign RetimeWrapper_125_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44853.4]
  assign RetimeWrapper_125_io_in = x525_lb_0_io_rPort_13_output_0; // @[package.scala 94:16:@44852.4]
  assign x717_sum_1_clock = clock; // @[:@44859.4]
  assign x717_sum_1_reset = reset; // @[:@44860.4]
  assign x717_sum_1_io_a = x716_x15_1_io_result; // @[Math.scala 151:17:@44861.4]
  assign x717_sum_1_io_b = RetimeWrapper_125_io_out; // @[Math.scala 152:17:@44862.4]
  assign x717_sum_1_io_flow = io_in_x481_TREADY; // @[Math.scala 153:20:@44863.4]
  assign RetimeWrapper_126_clock = clock; // @[:@44878.4]
  assign RetimeWrapper_126_reset = reset; // @[:@44879.4]
  assign RetimeWrapper_126_io_flow = io_in_x481_TREADY; // @[package.scala 95:18:@44881.4]
  assign RetimeWrapper_126_io_in = _GEN_22 << 1; // @[package.scala 94:16:@44880.4]
  assign RetimeWrapper_127_clock = clock; // @[:@44890.4]
  assign RetimeWrapper_127_reset = reset; // @[:@44891.4]
  assign RetimeWrapper_127_io_flow = io_in_x481_TREADY; // @[package.scala 95:18:@44893.4]
  assign RetimeWrapper_127_io_in = _GEN_23 << 2; // @[package.scala 94:16:@44892.4]
  assign RetimeWrapper_128_clock = clock; // @[:@44902.4]
  assign RetimeWrapper_128_reset = reset; // @[:@44903.4]
  assign RetimeWrapper_128_io_flow = io_in_x481_TREADY; // @[package.scala 95:18:@44905.4]
  assign RetimeWrapper_128_io_in = _GEN_24 << 1; // @[package.scala 94:16:@44904.4]
  assign RetimeWrapper_129_clock = clock; // @[:@44914.4]
  assign RetimeWrapper_129_reset = reset; // @[:@44915.4]
  assign RetimeWrapper_129_io_flow = io_in_x481_TREADY; // @[package.scala 95:18:@44917.4]
  assign RetimeWrapper_129_io_in = _GEN_25 << 1; // @[package.scala 94:16:@44916.4]
  assign x723_x15_1_io_a = RetimeWrapper_117_io_out; // @[Math.scala 151:17:@44926.4]
  assign x723_x15_1_io_b = _T_1678[7:0]; // @[Math.scala 152:17:@44927.4]
  assign RetimeWrapper_130_clock = clock; // @[:@44934.4]
  assign RetimeWrapper_130_reset = reset; // @[:@44935.4]
  assign RetimeWrapper_130_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44937.4]
  assign RetimeWrapper_130_io_in = x525_lb_0_io_rPort_8_output_0; // @[package.scala 94:16:@44936.4]
  assign x724_x16_1_io_a = RetimeWrapper_130_io_out; // @[Math.scala 151:17:@44945.4]
  assign x724_x16_1_io_b = _T_1556[7:0]; // @[Math.scala 152:17:@44946.4]
  assign x725_x15_1_io_a = _T_1684[7:0]; // @[Math.scala 151:17:@44955.4]
  assign x725_x15_1_io_b = _T_1690[7:0]; // @[Math.scala 152:17:@44956.4]
  assign x726_x16_1_io_a = RetimeWrapper_119_io_out; // @[Math.scala 151:17:@44965.4]
  assign x726_x16_1_io_b = _T_1696[7:0]; // @[Math.scala 152:17:@44966.4]
  assign x727_x15_1_io_a = x723_x15_1_io_result; // @[Math.scala 151:17:@44975.4]
  assign x727_x15_1_io_b = x724_x16_1_io_result; // @[Math.scala 152:17:@44976.4]
  assign x728_x16_1_io_a = x725_x15_1_io_result; // @[Math.scala 151:17:@44985.4]
  assign x728_x16_1_io_b = x726_x16_1_io_result; // @[Math.scala 152:17:@44986.4]
  assign x729_x15_1_io_a = x727_x15_1_io_result; // @[Math.scala 151:17:@44995.4]
  assign x729_x15_1_io_b = x728_x16_1_io_result; // @[Math.scala 152:17:@44996.4]
  assign RetimeWrapper_131_clock = clock; // @[:@45003.4]
  assign RetimeWrapper_131_reset = reset; // @[:@45004.4]
  assign RetimeWrapper_131_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45006.4]
  assign RetimeWrapper_131_io_in = x525_lb_0_io_rPort_17_output_0; // @[package.scala 94:16:@45005.4]
  assign x730_sum_1_clock = clock; // @[:@45014.4]
  assign x730_sum_1_reset = reset; // @[:@45015.4]
  assign x730_sum_1_io_a = x729_x15_1_io_result; // @[Math.scala 151:17:@45016.4]
  assign x730_sum_1_io_b = RetimeWrapper_131_io_out; // @[Math.scala 152:17:@45017.4]
  assign x730_sum_1_io_flow = io_in_x481_TREADY; // @[Math.scala 153:20:@45018.4]
  assign RetimeWrapper_132_clock = clock; // @[:@45041.4]
  assign RetimeWrapper_132_reset = reset; // @[:@45042.4]
  assign RetimeWrapper_132_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45044.4]
  assign RetimeWrapper_132_io_in = {_T_1751,_T_1750}; // @[package.scala 94:16:@45043.4]
  assign RetimeWrapper_133_clock = clock; // @[:@45050.4]
  assign RetimeWrapper_133_reset = reset; // @[:@45051.4]
  assign RetimeWrapper_133_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45053.4]
  assign RetimeWrapper_133_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@45052.4]
  assign RetimeWrapper_134_clock = clock; // @[:@45059.4]
  assign RetimeWrapper_134_reset = reset; // @[:@45060.4]
  assign RetimeWrapper_134_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45062.4]
  assign RetimeWrapper_134_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@45061.4]
  assign RetimeWrapper_135_clock = clock; // @[:@45068.4]
  assign RetimeWrapper_135_reset = reset; // @[:@45069.4]
  assign RetimeWrapper_135_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45071.4]
  assign RetimeWrapper_135_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@45070.4]
endmodule
module x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1( // @[:@45089.2]
  input          clock, // @[:@45090.4]
  input          reset, // @[:@45091.4]
  output         io_in_x481_TVALID, // @[:@45092.4]
  input          io_in_x481_TREADY, // @[:@45092.4]
  output [255:0] io_in_x481_TDATA, // @[:@45092.4]
  input          io_in_x480_TVALID, // @[:@45092.4]
  output         io_in_x480_TREADY, // @[:@45092.4]
  input  [255:0] io_in_x480_TDATA, // @[:@45092.4]
  input  [7:0]   io_in_x480_TID, // @[:@45092.4]
  input  [7:0]   io_in_x480_TDEST, // @[:@45092.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@45092.4]
  input          io_sigsIn_smChildAcks_0, // @[:@45092.4]
  output         io_sigsOut_smDoneIn_0, // @[:@45092.4]
  input          io_rr // @[:@45092.4]
);
  wire  x518_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@45126.4]
  wire  x518_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@45126.4]
  wire  x518_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@45126.4]
  wire  x518_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@45126.4]
  wire [12:0] x518_ctrchain_io_output_counts_1; // @[SpatialBlocks.scala 37:22:@45126.4]
  wire [12:0] x518_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@45126.4]
  wire  x518_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@45126.4]
  wire  x518_ctrchain_io_output_oobs_1; // @[SpatialBlocks.scala 37:22:@45126.4]
  wire  x518_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@45126.4]
  wire  x736_inr_Foreach_SAMPLER_BOX_sm_clock; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 32:18:@45186.4]
  wire  x736_inr_Foreach_SAMPLER_BOX_sm_reset; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 32:18:@45186.4]
  wire  x736_inr_Foreach_SAMPLER_BOX_sm_io_enable; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 32:18:@45186.4]
  wire  x736_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 32:18:@45186.4]
  wire  x736_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 32:18:@45186.4]
  wire  x736_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 32:18:@45186.4]
  wire  x736_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 32:18:@45186.4]
  wire  x736_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 32:18:@45186.4]
  wire  x736_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 32:18:@45186.4]
  wire  x736_inr_Foreach_SAMPLER_BOX_sm_io_parentAck; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 32:18:@45186.4]
  wire  x736_inr_Foreach_SAMPLER_BOX_sm_io_backpressure; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 32:18:@45186.4]
  wire  x736_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 32:18:@45186.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@45214.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@45214.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@45214.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@45214.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@45214.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@45256.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@45256.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@45256.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@45256.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@45256.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@45264.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@45264.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@45264.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@45264.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@45264.4]
  wire  x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_clock; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 798:24:@45298.4]
  wire  x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_reset; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 798:24:@45298.4]
  wire  x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x481_TVALID; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 798:24:@45298.4]
  wire  x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x481_TREADY; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 798:24:@45298.4]
  wire [255:0] x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x481_TDATA; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 798:24:@45298.4]
  wire  x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x480_TREADY; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 798:24:@45298.4]
  wire [255:0] x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x480_TDATA; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 798:24:@45298.4]
  wire [7:0] x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x480_TID; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 798:24:@45298.4]
  wire [7:0] x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x480_TDEST; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 798:24:@45298.4]
  wire  x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 798:24:@45298.4]
  wire  x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 798:24:@45298.4]
  wire  x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 798:24:@45298.4]
  wire [31:0] x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 798:24:@45298.4]
  wire [31:0] x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 798:24:@45298.4]
  wire  x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 798:24:@45298.4]
  wire  x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 798:24:@45298.4]
  wire  x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_rr; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 798:24:@45298.4]
  wire  _T_240; // @[package.scala 96:25:@45219.4 package.scala 96:25:@45220.4]
  wire  x736_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[sm_x737_outr_UnitPipe.scala 69:66:@45225.4]
  wire  _T_253; // @[package.scala 96:25:@45261.4 package.scala 96:25:@45262.4]
  wire  _T_259; // @[package.scala 96:25:@45269.4 package.scala 96:25:@45270.4]
  wire  _T_262; // @[SpatialBlocks.scala 138:93:@45272.4]
  wire  x736_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn; // @[SpatialBlocks.scala 138:90:@45273.4]
  wire  _T_264; // @[SpatialBlocks.scala 157:36:@45281.4]
  wire  _T_265; // @[SpatialBlocks.scala 157:78:@45282.4]
  wire  _T_272; // @[SpatialBlocks.scala 159:58:@45294.4]
  x488_ctrchain x518_ctrchain ( // @[SpatialBlocks.scala 37:22:@45126.4]
    .clock(x518_ctrchain_clock),
    .reset(x518_ctrchain_reset),
    .io_input_reset(x518_ctrchain_io_input_reset),
    .io_input_enable(x518_ctrchain_io_input_enable),
    .io_output_counts_1(x518_ctrchain_io_output_counts_1),
    .io_output_counts_0(x518_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x518_ctrchain_io_output_oobs_0),
    .io_output_oobs_1(x518_ctrchain_io_output_oobs_1),
    .io_output_done(x518_ctrchain_io_output_done)
  );
  x736_inr_Foreach_SAMPLER_BOX_sm x736_inr_Foreach_SAMPLER_BOX_sm ( // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 32:18:@45186.4]
    .clock(x736_inr_Foreach_SAMPLER_BOX_sm_clock),
    .reset(x736_inr_Foreach_SAMPLER_BOX_sm_reset),
    .io_enable(x736_inr_Foreach_SAMPLER_BOX_sm_io_enable),
    .io_done(x736_inr_Foreach_SAMPLER_BOX_sm_io_done),
    .io_doneLatch(x736_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch),
    .io_ctrDone(x736_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone),
    .io_datapathEn(x736_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn),
    .io_ctrInc(x736_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc),
    .io_ctrRst(x736_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst),
    .io_parentAck(x736_inr_Foreach_SAMPLER_BOX_sm_io_parentAck),
    .io_backpressure(x736_inr_Foreach_SAMPLER_BOX_sm_io_backpressure),
    .io_break(x736_inr_Foreach_SAMPLER_BOX_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@45214.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@45256.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@45264.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1 x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1 ( // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 798:24:@45298.4]
    .clock(x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_clock),
    .reset(x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_reset),
    .io_in_x481_TVALID(x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x481_TVALID),
    .io_in_x481_TREADY(x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x481_TREADY),
    .io_in_x481_TDATA(x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x481_TDATA),
    .io_in_x480_TREADY(x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x480_TREADY),
    .io_in_x480_TDATA(x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x480_TDATA),
    .io_in_x480_TID(x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x480_TID),
    .io_in_x480_TDEST(x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x480_TDEST),
    .io_sigsIn_backpressure(x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_1(x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsIn_cchainOutputs_0_oobs_1(x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1),
    .io_rr(x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_rr)
  );
  assign _T_240 = RetimeWrapper_io_out; // @[package.scala 96:25:@45219.4 package.scala 96:25:@45220.4]
  assign x736_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure = io_in_x480_TVALID | x736_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x737_outr_UnitPipe.scala 69:66:@45225.4]
  assign _T_253 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@45261.4 package.scala 96:25:@45262.4]
  assign _T_259 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@45269.4 package.scala 96:25:@45270.4]
  assign _T_262 = ~ _T_259; // @[SpatialBlocks.scala 138:93:@45272.4]
  assign x736_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn = _T_253 & _T_262; // @[SpatialBlocks.scala 138:90:@45273.4]
  assign _T_264 = x736_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@45281.4]
  assign _T_265 = ~ x736_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@45282.4]
  assign _T_272 = x736_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[SpatialBlocks.scala 159:58:@45294.4]
  assign io_in_x481_TVALID = x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x481_TVALID; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 48:23:@45357.4]
  assign io_in_x481_TDATA = x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x481_TDATA; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 48:23:@45355.4]
  assign io_in_x480_TREADY = x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x480_TREADY; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 49:23:@45365.4]
  assign io_sigsOut_smDoneIn_0 = x736_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[SpatialBlocks.scala 156:53:@45279.4]
  assign x518_ctrchain_clock = clock; // @[:@45127.4]
  assign x518_ctrchain_reset = reset; // @[:@45128.4]
  assign x518_ctrchain_io_input_reset = x736_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@45297.4]
  assign x518_ctrchain_io_input_enable = _T_272 & x736_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 132:75:@45249.4 SpatialBlocks.scala 159:42:@45296.4]
  assign x736_inr_Foreach_SAMPLER_BOX_sm_clock = clock; // @[:@45187.4]
  assign x736_inr_Foreach_SAMPLER_BOX_sm_reset = reset; // @[:@45188.4]
  assign x736_inr_Foreach_SAMPLER_BOX_sm_io_enable = x736_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn & x736_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 140:18:@45276.4]
  assign x736_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone = io_rr ? _T_240 : 1'h0; // @[sm_x737_outr_UnitPipe.scala 67:50:@45222.4]
  assign x736_inr_Foreach_SAMPLER_BOX_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@45278.4]
  assign x736_inr_Foreach_SAMPLER_BOX_sm_io_backpressure = io_in_x481_TREADY | x736_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@45250.4]
  assign x736_inr_Foreach_SAMPLER_BOX_sm_io_break = 1'h0; // @[sm_x737_outr_UnitPipe.scala 71:48:@45228.4]
  assign RetimeWrapper_clock = clock; // @[:@45215.4]
  assign RetimeWrapper_reset = reset; // @[:@45216.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@45218.4]
  assign RetimeWrapper_io_in = x518_ctrchain_io_output_done; // @[package.scala 94:16:@45217.4]
  assign RetimeWrapper_1_clock = clock; // @[:@45257.4]
  assign RetimeWrapper_1_reset = reset; // @[:@45258.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@45260.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@45259.4]
  assign RetimeWrapper_2_clock = clock; // @[:@45265.4]
  assign RetimeWrapper_2_reset = reset; // @[:@45266.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@45268.4]
  assign RetimeWrapper_2_io_in = x736_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[package.scala 94:16:@45267.4]
  assign x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_clock = clock; // @[:@45299.4]
  assign x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_reset = reset; // @[:@45300.4]
  assign x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x481_TREADY = io_in_x481_TREADY; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 48:23:@45356.4]
  assign x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x480_TDATA = io_in_x480_TDATA; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 49:23:@45364.4]
  assign x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x480_TID = io_in_x480_TID; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 49:23:@45360.4]
  assign x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x480_TDEST = io_in_x480_TDEST; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 49:23:@45359.4]
  assign x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure = io_in_x481_TREADY | x736_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 803:22:@45383.4]
  assign x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn = _T_264 & _T_265; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 803:22:@45381.4]
  assign x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break = x736_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 803:22:@45379.4]
  assign x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1 = {{19{x518_ctrchain_io_output_counts_1[12]}},x518_ctrchain_io_output_counts_1}; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 803:22:@45374.4]
  assign x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{19{x518_ctrchain_io_output_counts_0[12]}},x518_ctrchain_io_output_counts_0}; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 803:22:@45373.4]
  assign x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x518_ctrchain_io_output_oobs_0; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 803:22:@45371.4]
  assign x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1 = x518_ctrchain_io_output_oobs_1; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 803:22:@45372.4]
  assign x736_inr_Foreach_SAMPLER_BOX_kernelx736_inr_Foreach_SAMPLER_BOX_concrete1_io_rr = io_rr; // @[sm_x736_inr_Foreach_SAMPLER_BOX.scala 802:18:@45367.4]
endmodule
module x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1( // @[:@45397.2]
  input          clock, // @[:@45398.4]
  input          reset, // @[:@45399.4]
  output         io_in_x481_TVALID, // @[:@45400.4]
  input          io_in_x481_TREADY, // @[:@45400.4]
  output [255:0] io_in_x481_TDATA, // @[:@45400.4]
  input          io_in_x480_TVALID, // @[:@45400.4]
  output         io_in_x480_TREADY, // @[:@45400.4]
  input  [255:0] io_in_x480_TDATA, // @[:@45400.4]
  input  [7:0]   io_in_x480_TID, // @[:@45400.4]
  input  [7:0]   io_in_x480_TDEST, // @[:@45400.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@45400.4]
  input          io_sigsIn_smEnableOuts_1, // @[:@45400.4]
  input          io_sigsIn_smChildAcks_0, // @[:@45400.4]
  input          io_sigsIn_smChildAcks_1, // @[:@45400.4]
  output         io_sigsOut_smDoneIn_0, // @[:@45400.4]
  output         io_sigsOut_smDoneIn_1, // @[:@45400.4]
  output         io_sigsOut_smCtrCopyDone_0, // @[:@45400.4]
  output         io_sigsOut_smCtrCopyDone_1, // @[:@45400.4]
  input          io_rr // @[:@45400.4]
);
  wire  x483_fifoinraw_0_clock; // @[m_x483_fifoinraw_0.scala 27:17:@45414.4]
  wire  x483_fifoinraw_0_reset; // @[m_x483_fifoinraw_0.scala 27:17:@45414.4]
  wire  x484_fifoinpacked_0_clock; // @[m_x484_fifoinpacked_0.scala 27:17:@45438.4]
  wire  x484_fifoinpacked_0_reset; // @[m_x484_fifoinpacked_0.scala 27:17:@45438.4]
  wire  x484_fifoinpacked_0_io_wPort_0_en_0; // @[m_x484_fifoinpacked_0.scala 27:17:@45438.4]
  wire  x484_fifoinpacked_0_io_full; // @[m_x484_fifoinpacked_0.scala 27:17:@45438.4]
  wire  x484_fifoinpacked_0_io_active_0_in; // @[m_x484_fifoinpacked_0.scala 27:17:@45438.4]
  wire  x484_fifoinpacked_0_io_active_0_out; // @[m_x484_fifoinpacked_0.scala 27:17:@45438.4]
  wire  x485_fifooutraw_0_clock; // @[m_x485_fifooutraw_0.scala 27:17:@45462.4]
  wire  x485_fifooutraw_0_reset; // @[m_x485_fifooutraw_0.scala 27:17:@45462.4]
  wire  x488_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@45486.4]
  wire  x488_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@45486.4]
  wire  x488_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@45486.4]
  wire  x488_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@45486.4]
  wire [12:0] x488_ctrchain_io_output_counts_1; // @[SpatialBlocks.scala 37:22:@45486.4]
  wire [12:0] x488_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@45486.4]
  wire  x488_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@45486.4]
  wire  x488_ctrchain_io_output_oobs_1; // @[SpatialBlocks.scala 37:22:@45486.4]
  wire  x488_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@45486.4]
  wire  x514_inr_Foreach_sm_clock; // @[sm_x514_inr_Foreach.scala 32:18:@45546.4]
  wire  x514_inr_Foreach_sm_reset; // @[sm_x514_inr_Foreach.scala 32:18:@45546.4]
  wire  x514_inr_Foreach_sm_io_enable; // @[sm_x514_inr_Foreach.scala 32:18:@45546.4]
  wire  x514_inr_Foreach_sm_io_done; // @[sm_x514_inr_Foreach.scala 32:18:@45546.4]
  wire  x514_inr_Foreach_sm_io_doneLatch; // @[sm_x514_inr_Foreach.scala 32:18:@45546.4]
  wire  x514_inr_Foreach_sm_io_ctrDone; // @[sm_x514_inr_Foreach.scala 32:18:@45546.4]
  wire  x514_inr_Foreach_sm_io_datapathEn; // @[sm_x514_inr_Foreach.scala 32:18:@45546.4]
  wire  x514_inr_Foreach_sm_io_ctrInc; // @[sm_x514_inr_Foreach.scala 32:18:@45546.4]
  wire  x514_inr_Foreach_sm_io_ctrRst; // @[sm_x514_inr_Foreach.scala 32:18:@45546.4]
  wire  x514_inr_Foreach_sm_io_parentAck; // @[sm_x514_inr_Foreach.scala 32:18:@45546.4]
  wire  x514_inr_Foreach_sm_io_backpressure; // @[sm_x514_inr_Foreach.scala 32:18:@45546.4]
  wire  x514_inr_Foreach_sm_io_break; // @[sm_x514_inr_Foreach.scala 32:18:@45546.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@45574.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@45574.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@45574.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@45574.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@45574.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@45620.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@45620.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@45620.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@45620.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@45620.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@45628.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@45628.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@45628.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@45628.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@45628.4]
  wire  x514_inr_Foreach_kernelx514_inr_Foreach_concrete1_clock; // @[sm_x514_inr_Foreach.scala 126:24:@45663.4]
  wire  x514_inr_Foreach_kernelx514_inr_Foreach_concrete1_reset; // @[sm_x514_inr_Foreach.scala 126:24:@45663.4]
  wire  x514_inr_Foreach_kernelx514_inr_Foreach_concrete1_io_in_x484_fifoinpacked_0_wPort_0_en_0; // @[sm_x514_inr_Foreach.scala 126:24:@45663.4]
  wire  x514_inr_Foreach_kernelx514_inr_Foreach_concrete1_io_in_x484_fifoinpacked_0_full; // @[sm_x514_inr_Foreach.scala 126:24:@45663.4]
  wire  x514_inr_Foreach_kernelx514_inr_Foreach_concrete1_io_in_x484_fifoinpacked_0_active_0_in; // @[sm_x514_inr_Foreach.scala 126:24:@45663.4]
  wire  x514_inr_Foreach_kernelx514_inr_Foreach_concrete1_io_in_x484_fifoinpacked_0_active_0_out; // @[sm_x514_inr_Foreach.scala 126:24:@45663.4]
  wire  x514_inr_Foreach_kernelx514_inr_Foreach_concrete1_io_sigsIn_backpressure; // @[sm_x514_inr_Foreach.scala 126:24:@45663.4]
  wire  x514_inr_Foreach_kernelx514_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x514_inr_Foreach.scala 126:24:@45663.4]
  wire  x514_inr_Foreach_kernelx514_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x514_inr_Foreach.scala 126:24:@45663.4]
  wire [31:0] x514_inr_Foreach_kernelx514_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1; // @[sm_x514_inr_Foreach.scala 126:24:@45663.4]
  wire [31:0] x514_inr_Foreach_kernelx514_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x514_inr_Foreach.scala 126:24:@45663.4]
  wire  x514_inr_Foreach_kernelx514_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x514_inr_Foreach.scala 126:24:@45663.4]
  wire  x514_inr_Foreach_kernelx514_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x514_inr_Foreach.scala 126:24:@45663.4]
  wire  x514_inr_Foreach_kernelx514_inr_Foreach_concrete1_io_rr; // @[sm_x514_inr_Foreach.scala 126:24:@45663.4]
  wire  x737_outr_UnitPipe_sm_clock; // @[sm_x737_outr_UnitPipe.scala 32:18:@45795.4]
  wire  x737_outr_UnitPipe_sm_reset; // @[sm_x737_outr_UnitPipe.scala 32:18:@45795.4]
  wire  x737_outr_UnitPipe_sm_io_enable; // @[sm_x737_outr_UnitPipe.scala 32:18:@45795.4]
  wire  x737_outr_UnitPipe_sm_io_done; // @[sm_x737_outr_UnitPipe.scala 32:18:@45795.4]
  wire  x737_outr_UnitPipe_sm_io_rst; // @[sm_x737_outr_UnitPipe.scala 32:18:@45795.4]
  wire  x737_outr_UnitPipe_sm_io_ctrDone; // @[sm_x737_outr_UnitPipe.scala 32:18:@45795.4]
  wire  x737_outr_UnitPipe_sm_io_ctrInc; // @[sm_x737_outr_UnitPipe.scala 32:18:@45795.4]
  wire  x737_outr_UnitPipe_sm_io_parentAck; // @[sm_x737_outr_UnitPipe.scala 32:18:@45795.4]
  wire  x737_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x737_outr_UnitPipe.scala 32:18:@45795.4]
  wire  x737_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x737_outr_UnitPipe.scala 32:18:@45795.4]
  wire  x737_outr_UnitPipe_sm_io_childAck_0; // @[sm_x737_outr_UnitPipe.scala 32:18:@45795.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@45852.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@45852.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@45852.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@45852.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@45852.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@45860.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@45860.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@45860.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@45860.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@45860.4]
  wire  x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1_clock; // @[sm_x737_outr_UnitPipe.scala 76:24:@45890.4]
  wire  x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1_reset; // @[sm_x737_outr_UnitPipe.scala 76:24:@45890.4]
  wire  x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1_io_in_x481_TVALID; // @[sm_x737_outr_UnitPipe.scala 76:24:@45890.4]
  wire  x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1_io_in_x481_TREADY; // @[sm_x737_outr_UnitPipe.scala 76:24:@45890.4]
  wire [255:0] x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1_io_in_x481_TDATA; // @[sm_x737_outr_UnitPipe.scala 76:24:@45890.4]
  wire  x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1_io_in_x480_TVALID; // @[sm_x737_outr_UnitPipe.scala 76:24:@45890.4]
  wire  x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1_io_in_x480_TREADY; // @[sm_x737_outr_UnitPipe.scala 76:24:@45890.4]
  wire [255:0] x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1_io_in_x480_TDATA; // @[sm_x737_outr_UnitPipe.scala 76:24:@45890.4]
  wire [7:0] x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1_io_in_x480_TID; // @[sm_x737_outr_UnitPipe.scala 76:24:@45890.4]
  wire [7:0] x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1_io_in_x480_TDEST; // @[sm_x737_outr_UnitPipe.scala 76:24:@45890.4]
  wire  x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x737_outr_UnitPipe.scala 76:24:@45890.4]
  wire  x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x737_outr_UnitPipe.scala 76:24:@45890.4]
  wire  x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x737_outr_UnitPipe.scala 76:24:@45890.4]
  wire  x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1_io_rr; // @[sm_x737_outr_UnitPipe.scala 76:24:@45890.4]
  wire  _T_254; // @[package.scala 96:25:@45579.4 package.scala 96:25:@45580.4]
  wire  _T_260; // @[implicits.scala 47:10:@45583.4]
  wire  _T_261; // @[sm_x738_outr_UnitPipe.scala 70:41:@45584.4]
  wire  _T_262; // @[sm_x738_outr_UnitPipe.scala 70:78:@45585.4]
  wire  _T_263; // @[sm_x738_outr_UnitPipe.scala 70:76:@45586.4]
  wire  _T_275; // @[package.scala 96:25:@45625.4 package.scala 96:25:@45626.4]
  wire  _T_281; // @[package.scala 96:25:@45633.4 package.scala 96:25:@45634.4]
  wire  _T_284; // @[SpatialBlocks.scala 138:93:@45636.4]
  wire  _T_286; // @[SpatialBlocks.scala 157:36:@45645.4]
  wire  _T_287; // @[SpatialBlocks.scala 157:78:@45646.4]
  wire  _T_354; // @[package.scala 100:49:@45823.4]
  reg  _T_357; // @[package.scala 48:56:@45824.4]
  reg [31:0] _RAND_0;
  wire  _T_371; // @[package.scala 96:25:@45857.4 package.scala 96:25:@45858.4]
  wire  _T_377; // @[package.scala 96:25:@45865.4 package.scala 96:25:@45866.4]
  wire  _T_380; // @[SpatialBlocks.scala 138:93:@45868.4]
  x483_fifoinraw_0 x483_fifoinraw_0 ( // @[m_x483_fifoinraw_0.scala 27:17:@45414.4]
    .clock(x483_fifoinraw_0_clock),
    .reset(x483_fifoinraw_0_reset)
  );
  x484_fifoinpacked_0 x484_fifoinpacked_0 ( // @[m_x484_fifoinpacked_0.scala 27:17:@45438.4]
    .clock(x484_fifoinpacked_0_clock),
    .reset(x484_fifoinpacked_0_reset),
    .io_wPort_0_en_0(x484_fifoinpacked_0_io_wPort_0_en_0),
    .io_full(x484_fifoinpacked_0_io_full),
    .io_active_0_in(x484_fifoinpacked_0_io_active_0_in),
    .io_active_0_out(x484_fifoinpacked_0_io_active_0_out)
  );
  x483_fifoinraw_0 x485_fifooutraw_0 ( // @[m_x485_fifooutraw_0.scala 27:17:@45462.4]
    .clock(x485_fifooutraw_0_clock),
    .reset(x485_fifooutraw_0_reset)
  );
  x488_ctrchain x488_ctrchain ( // @[SpatialBlocks.scala 37:22:@45486.4]
    .clock(x488_ctrchain_clock),
    .reset(x488_ctrchain_reset),
    .io_input_reset(x488_ctrchain_io_input_reset),
    .io_input_enable(x488_ctrchain_io_input_enable),
    .io_output_counts_1(x488_ctrchain_io_output_counts_1),
    .io_output_counts_0(x488_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x488_ctrchain_io_output_oobs_0),
    .io_output_oobs_1(x488_ctrchain_io_output_oobs_1),
    .io_output_done(x488_ctrchain_io_output_done)
  );
  x514_inr_Foreach_sm x514_inr_Foreach_sm ( // @[sm_x514_inr_Foreach.scala 32:18:@45546.4]
    .clock(x514_inr_Foreach_sm_clock),
    .reset(x514_inr_Foreach_sm_reset),
    .io_enable(x514_inr_Foreach_sm_io_enable),
    .io_done(x514_inr_Foreach_sm_io_done),
    .io_doneLatch(x514_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x514_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x514_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x514_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x514_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x514_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x514_inr_Foreach_sm_io_backpressure),
    .io_break(x514_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@45574.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@45620.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@45628.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x514_inr_Foreach_kernelx514_inr_Foreach_concrete1 x514_inr_Foreach_kernelx514_inr_Foreach_concrete1 ( // @[sm_x514_inr_Foreach.scala 126:24:@45663.4]
    .clock(x514_inr_Foreach_kernelx514_inr_Foreach_concrete1_clock),
    .reset(x514_inr_Foreach_kernelx514_inr_Foreach_concrete1_reset),
    .io_in_x484_fifoinpacked_0_wPort_0_en_0(x514_inr_Foreach_kernelx514_inr_Foreach_concrete1_io_in_x484_fifoinpacked_0_wPort_0_en_0),
    .io_in_x484_fifoinpacked_0_full(x514_inr_Foreach_kernelx514_inr_Foreach_concrete1_io_in_x484_fifoinpacked_0_full),
    .io_in_x484_fifoinpacked_0_active_0_in(x514_inr_Foreach_kernelx514_inr_Foreach_concrete1_io_in_x484_fifoinpacked_0_active_0_in),
    .io_in_x484_fifoinpacked_0_active_0_out(x514_inr_Foreach_kernelx514_inr_Foreach_concrete1_io_in_x484_fifoinpacked_0_active_0_out),
    .io_sigsIn_backpressure(x514_inr_Foreach_kernelx514_inr_Foreach_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x514_inr_Foreach_kernelx514_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x514_inr_Foreach_kernelx514_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_1(x514_inr_Foreach_kernelx514_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x514_inr_Foreach_kernelx514_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x514_inr_Foreach_kernelx514_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsIn_cchainOutputs_0_oobs_1(x514_inr_Foreach_kernelx514_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1),
    .io_rr(x514_inr_Foreach_kernelx514_inr_Foreach_concrete1_io_rr)
  );
  RootController_sm x737_outr_UnitPipe_sm ( // @[sm_x737_outr_UnitPipe.scala 32:18:@45795.4]
    .clock(x737_outr_UnitPipe_sm_clock),
    .reset(x737_outr_UnitPipe_sm_reset),
    .io_enable(x737_outr_UnitPipe_sm_io_enable),
    .io_done(x737_outr_UnitPipe_sm_io_done),
    .io_rst(x737_outr_UnitPipe_sm_io_rst),
    .io_ctrDone(x737_outr_UnitPipe_sm_io_ctrDone),
    .io_ctrInc(x737_outr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x737_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x737_outr_UnitPipe_sm_io_doneIn_0),
    .io_enableOut_0(x737_outr_UnitPipe_sm_io_enableOut_0),
    .io_childAck_0(x737_outr_UnitPipe_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@45852.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@45860.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1 x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1 ( // @[sm_x737_outr_UnitPipe.scala 76:24:@45890.4]
    .clock(x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1_clock),
    .reset(x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1_reset),
    .io_in_x481_TVALID(x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1_io_in_x481_TVALID),
    .io_in_x481_TREADY(x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1_io_in_x481_TREADY),
    .io_in_x481_TDATA(x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1_io_in_x481_TDATA),
    .io_in_x480_TVALID(x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1_io_in_x480_TVALID),
    .io_in_x480_TREADY(x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1_io_in_x480_TREADY),
    .io_in_x480_TDATA(x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1_io_in_x480_TDATA),
    .io_in_x480_TID(x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1_io_in_x480_TID),
    .io_in_x480_TDEST(x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1_io_in_x480_TDEST),
    .io_sigsIn_smEnableOuts_0(x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_254 = RetimeWrapper_io_out; // @[package.scala 96:25:@45579.4 package.scala 96:25:@45580.4]
  assign _T_260 = x484_fifoinpacked_0_io_full; // @[implicits.scala 47:10:@45583.4]
  assign _T_261 = ~ _T_260; // @[sm_x738_outr_UnitPipe.scala 70:41:@45584.4]
  assign _T_262 = ~ x484_fifoinpacked_0_io_active_0_out; // @[sm_x738_outr_UnitPipe.scala 70:78:@45585.4]
  assign _T_263 = _T_261 | _T_262; // @[sm_x738_outr_UnitPipe.scala 70:76:@45586.4]
  assign _T_275 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@45625.4 package.scala 96:25:@45626.4]
  assign _T_281 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@45633.4 package.scala 96:25:@45634.4]
  assign _T_284 = ~ _T_281; // @[SpatialBlocks.scala 138:93:@45636.4]
  assign _T_286 = x514_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@45645.4]
  assign _T_287 = ~ x514_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@45646.4]
  assign _T_354 = x737_outr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@45823.4]
  assign _T_371 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@45857.4 package.scala 96:25:@45858.4]
  assign _T_377 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@45865.4 package.scala 96:25:@45866.4]
  assign _T_380 = ~ _T_377; // @[SpatialBlocks.scala 138:93:@45868.4]
  assign io_in_x481_TVALID = x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1_io_in_x481_TVALID; // @[sm_x737_outr_UnitPipe.scala 48:23:@45947.4]
  assign io_in_x481_TDATA = x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1_io_in_x481_TDATA; // @[sm_x737_outr_UnitPipe.scala 48:23:@45945.4]
  assign io_in_x480_TREADY = x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1_io_in_x480_TREADY; // @[sm_x737_outr_UnitPipe.scala 49:23:@45955.4]
  assign io_sigsOut_smDoneIn_0 = x514_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 156:53:@45643.4]
  assign io_sigsOut_smDoneIn_1 = x737_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@45875.4]
  assign io_sigsOut_smCtrCopyDone_0 = x514_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 168:125:@45662.4]
  assign io_sigsOut_smCtrCopyDone_1 = x737_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@45889.4]
  assign x483_fifoinraw_0_clock = clock; // @[:@45415.4]
  assign x483_fifoinraw_0_reset = reset; // @[:@45416.4]
  assign x484_fifoinpacked_0_clock = clock; // @[:@45439.4]
  assign x484_fifoinpacked_0_reset = reset; // @[:@45440.4]
  assign x484_fifoinpacked_0_io_wPort_0_en_0 = x514_inr_Foreach_kernelx514_inr_Foreach_concrete1_io_in_x484_fifoinpacked_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@45723.4]
  assign x484_fifoinpacked_0_io_active_0_in = x514_inr_Foreach_kernelx514_inr_Foreach_concrete1_io_in_x484_fifoinpacked_0_active_0_in; // @[MemInterfaceType.scala 167:86:@45722.4]
  assign x485_fifooutraw_0_clock = clock; // @[:@45463.4]
  assign x485_fifooutraw_0_reset = reset; // @[:@45464.4]
  assign x488_ctrchain_clock = clock; // @[:@45487.4]
  assign x488_ctrchain_reset = reset; // @[:@45488.4]
  assign x488_ctrchain_io_input_reset = x514_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@45661.4]
  assign x488_ctrchain_io_input_enable = x514_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 132:75:@45613.4 SpatialBlocks.scala 159:42:@45660.4]
  assign x514_inr_Foreach_sm_clock = clock; // @[:@45547.4]
  assign x514_inr_Foreach_sm_reset = reset; // @[:@45548.4]
  assign x514_inr_Foreach_sm_io_enable = _T_275 & _T_284; // @[SpatialBlocks.scala 140:18:@45640.4]
  assign x514_inr_Foreach_sm_io_ctrDone = io_rr ? _T_254 : 1'h0; // @[sm_x738_outr_UnitPipe.scala 69:38:@45582.4]
  assign x514_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@45642.4]
  assign x514_inr_Foreach_sm_io_backpressure = _T_263 | x514_inr_Foreach_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@45614.4]
  assign x514_inr_Foreach_sm_io_break = 1'h0; // @[sm_x738_outr_UnitPipe.scala 73:36:@45592.4]
  assign RetimeWrapper_clock = clock; // @[:@45575.4]
  assign RetimeWrapper_reset = reset; // @[:@45576.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@45578.4]
  assign RetimeWrapper_io_in = x488_ctrchain_io_output_done; // @[package.scala 94:16:@45577.4]
  assign RetimeWrapper_1_clock = clock; // @[:@45621.4]
  assign RetimeWrapper_1_reset = reset; // @[:@45622.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@45624.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@45623.4]
  assign RetimeWrapper_2_clock = clock; // @[:@45629.4]
  assign RetimeWrapper_2_reset = reset; // @[:@45630.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@45632.4]
  assign RetimeWrapper_2_io_in = x514_inr_Foreach_sm_io_done; // @[package.scala 94:16:@45631.4]
  assign x514_inr_Foreach_kernelx514_inr_Foreach_concrete1_clock = clock; // @[:@45664.4]
  assign x514_inr_Foreach_kernelx514_inr_Foreach_concrete1_reset = reset; // @[:@45665.4]
  assign x514_inr_Foreach_kernelx514_inr_Foreach_concrete1_io_in_x484_fifoinpacked_0_full = x484_fifoinpacked_0_io_full; // @[MemInterfaceType.scala 159:15:@45717.4]
  assign x514_inr_Foreach_kernelx514_inr_Foreach_concrete1_io_in_x484_fifoinpacked_0_active_0_out = x484_fifoinpacked_0_io_active_0_out; // @[MemInterfaceType.scala 158:75:@45716.4]
  assign x514_inr_Foreach_kernelx514_inr_Foreach_concrete1_io_sigsIn_backpressure = _T_263 | x514_inr_Foreach_sm_io_doneLatch; // @[sm_x514_inr_Foreach.scala 131:22:@45746.4]
  assign x514_inr_Foreach_kernelx514_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_286 & _T_287; // @[sm_x514_inr_Foreach.scala 131:22:@45744.4]
  assign x514_inr_Foreach_kernelx514_inr_Foreach_concrete1_io_sigsIn_break = x514_inr_Foreach_sm_io_break; // @[sm_x514_inr_Foreach.scala 131:22:@45742.4]
  assign x514_inr_Foreach_kernelx514_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1 = {{19{x488_ctrchain_io_output_counts_1[12]}},x488_ctrchain_io_output_counts_1}; // @[sm_x514_inr_Foreach.scala 131:22:@45737.4]
  assign x514_inr_Foreach_kernelx514_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{19{x488_ctrchain_io_output_counts_0[12]}},x488_ctrchain_io_output_counts_0}; // @[sm_x514_inr_Foreach.scala 131:22:@45736.4]
  assign x514_inr_Foreach_kernelx514_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x488_ctrchain_io_output_oobs_0; // @[sm_x514_inr_Foreach.scala 131:22:@45734.4]
  assign x514_inr_Foreach_kernelx514_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1 = x488_ctrchain_io_output_oobs_1; // @[sm_x514_inr_Foreach.scala 131:22:@45735.4]
  assign x514_inr_Foreach_kernelx514_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x514_inr_Foreach.scala 130:18:@45730.4]
  assign x737_outr_UnitPipe_sm_clock = clock; // @[:@45796.4]
  assign x737_outr_UnitPipe_sm_reset = reset; // @[:@45797.4]
  assign x737_outr_UnitPipe_sm_io_enable = _T_371 & _T_380; // @[SpatialBlocks.scala 140:18:@45872.4]
  assign x737_outr_UnitPipe_sm_io_rst = 1'h0; // @[SpatialBlocks.scala 134:15:@45847.4]
  assign x737_outr_UnitPipe_sm_io_ctrDone = x737_outr_UnitPipe_sm_io_ctrInc & _T_357; // @[sm_x738_outr_UnitPipe.scala 78:40:@45827.4]
  assign x737_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@45874.4]
  assign x737_outr_UnitPipe_sm_io_doneIn_0 = x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@45844.4]
  assign RetimeWrapper_3_clock = clock; // @[:@45853.4]
  assign RetimeWrapper_3_reset = reset; // @[:@45854.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@45856.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@45855.4]
  assign RetimeWrapper_4_clock = clock; // @[:@45861.4]
  assign RetimeWrapper_4_reset = reset; // @[:@45862.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@45864.4]
  assign RetimeWrapper_4_io_in = x737_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@45863.4]
  assign x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1_clock = clock; // @[:@45891.4]
  assign x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1_reset = reset; // @[:@45892.4]
  assign x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1_io_in_x481_TREADY = io_in_x481_TREADY; // @[sm_x737_outr_UnitPipe.scala 48:23:@45946.4]
  assign x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1_io_in_x480_TVALID = io_in_x480_TVALID; // @[sm_x737_outr_UnitPipe.scala 49:23:@45956.4]
  assign x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1_io_in_x480_TDATA = io_in_x480_TDATA; // @[sm_x737_outr_UnitPipe.scala 49:23:@45954.4]
  assign x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1_io_in_x480_TID = io_in_x480_TID; // @[sm_x737_outr_UnitPipe.scala 49:23:@45950.4]
  assign x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1_io_in_x480_TDEST = io_in_x480_TDEST; // @[sm_x737_outr_UnitPipe.scala 49:23:@45949.4]
  assign x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x737_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x737_outr_UnitPipe.scala 81:22:@45965.4]
  assign x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x737_outr_UnitPipe_sm_io_childAck_0; // @[sm_x737_outr_UnitPipe.scala 81:22:@45963.4]
  assign x737_outr_UnitPipe_kernelx737_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x737_outr_UnitPipe.scala 80:18:@45957.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_357 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_357 <= 1'h0;
    end else begin
      _T_357 <= _T_354;
    end
  end
endmodule
module x760_outr_UnitPipe_sm( // @[:@46454.2]
  input   clock, // @[:@46455.4]
  input   reset, // @[:@46456.4]
  input   io_enable, // @[:@46457.4]
  output  io_done, // @[:@46457.4]
  input   io_parentAck, // @[:@46457.4]
  input   io_doneIn_0, // @[:@46457.4]
  input   io_doneIn_1, // @[:@46457.4]
  input   io_doneIn_2, // @[:@46457.4]
  output  io_enableOut_0, // @[:@46457.4]
  output  io_enableOut_1, // @[:@46457.4]
  output  io_enableOut_2, // @[:@46457.4]
  output  io_childAck_0, // @[:@46457.4]
  output  io_childAck_1, // @[:@46457.4]
  output  io_childAck_2, // @[:@46457.4]
  input   io_ctrCopyDone_0, // @[:@46457.4]
  input   io_ctrCopyDone_1, // @[:@46457.4]
  input   io_ctrCopyDone_2 // @[:@46457.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@46460.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@46460.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@46460.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@46460.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@46460.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@46460.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@46463.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@46463.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@46463.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@46463.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@46463.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@46463.4]
  wire  active_2_clock; // @[Controllers.scala 76:50:@46466.4]
  wire  active_2_reset; // @[Controllers.scala 76:50:@46466.4]
  wire  active_2_io_input_set; // @[Controllers.scala 76:50:@46466.4]
  wire  active_2_io_input_reset; // @[Controllers.scala 76:50:@46466.4]
  wire  active_2_io_input_asyn_reset; // @[Controllers.scala 76:50:@46466.4]
  wire  active_2_io_output; // @[Controllers.scala 76:50:@46466.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@46469.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@46469.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@46469.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@46469.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@46469.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@46469.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@46472.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@46472.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@46472.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@46472.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@46472.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@46472.4]
  wire  done_2_clock; // @[Controllers.scala 77:48:@46475.4]
  wire  done_2_reset; // @[Controllers.scala 77:48:@46475.4]
  wire  done_2_io_input_set; // @[Controllers.scala 77:48:@46475.4]
  wire  done_2_io_input_reset; // @[Controllers.scala 77:48:@46475.4]
  wire  done_2_io_input_asyn_reset; // @[Controllers.scala 77:48:@46475.4]
  wire  done_2_io_output; // @[Controllers.scala 77:48:@46475.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@46516.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@46516.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@46516.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@46516.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@46516.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@46516.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@46519.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@46519.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@46519.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@46519.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@46519.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@46519.4]
  wire  iterDone_2_clock; // @[Controllers.scala 90:52:@46522.4]
  wire  iterDone_2_reset; // @[Controllers.scala 90:52:@46522.4]
  wire  iterDone_2_io_input_set; // @[Controllers.scala 90:52:@46522.4]
  wire  iterDone_2_io_input_reset; // @[Controllers.scala 90:52:@46522.4]
  wire  iterDone_2_io_input_asyn_reset; // @[Controllers.scala 90:52:@46522.4]
  wire  iterDone_2_io_output; // @[Controllers.scala 90:52:@46522.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@46573.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@46573.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@46573.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@46573.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@46573.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@46587.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@46587.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@46587.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@46587.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@46587.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@46605.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@46605.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@46605.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@46605.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@46605.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@46642.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@46642.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@46642.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@46642.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@46642.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@46656.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@46656.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@46656.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@46656.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@46656.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@46674.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@46674.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@46674.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@46674.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@46674.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@46711.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@46711.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@46711.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@46711.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@46711.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@46725.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@46725.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@46725.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@46725.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@46725.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@46743.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@46743.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@46743.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@46743.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@46743.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@46800.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@46800.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@46800.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@46800.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@46800.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@46817.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@46817.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@46817.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@46817.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@46817.4]
  wire  _T_77; // @[Controllers.scala 80:47:@46478.4]
  wire  allDone; // @[Controllers.scala 80:47:@46479.4]
  wire  _T_151; // @[Controllers.scala 165:35:@46557.4]
  wire  _T_153; // @[Controllers.scala 165:60:@46558.4]
  wire  _T_154; // @[Controllers.scala 165:58:@46559.4]
  wire  _T_156; // @[Controllers.scala 165:76:@46560.4]
  wire  _T_157; // @[Controllers.scala 165:74:@46561.4]
  wire  _T_161; // @[Controllers.scala 165:109:@46564.4]
  wire  _T_164; // @[Controllers.scala 165:141:@46566.4]
  wire  _T_172; // @[package.scala 96:25:@46578.4 package.scala 96:25:@46579.4]
  wire  _T_176; // @[Controllers.scala 167:54:@46581.4]
  wire  _T_177; // @[Controllers.scala 167:52:@46582.4]
  wire  _T_184; // @[package.scala 96:25:@46592.4 package.scala 96:25:@46593.4]
  wire  _T_202; // @[package.scala 96:25:@46610.4 package.scala 96:25:@46611.4]
  wire  _T_206; // @[Controllers.scala 169:67:@46613.4]
  wire  _T_207; // @[Controllers.scala 169:86:@46614.4]
  wire  _T_219; // @[Controllers.scala 165:35:@46626.4]
  wire  _T_221; // @[Controllers.scala 165:60:@46627.4]
  wire  _T_222; // @[Controllers.scala 165:58:@46628.4]
  wire  _T_224; // @[Controllers.scala 165:76:@46629.4]
  wire  _T_225; // @[Controllers.scala 165:74:@46630.4]
  wire  _T_229; // @[Controllers.scala 165:109:@46633.4]
  wire  _T_232; // @[Controllers.scala 165:141:@46635.4]
  wire  _T_240; // @[package.scala 96:25:@46647.4 package.scala 96:25:@46648.4]
  wire  _T_244; // @[Controllers.scala 167:54:@46650.4]
  wire  _T_245; // @[Controllers.scala 167:52:@46651.4]
  wire  _T_252; // @[package.scala 96:25:@46661.4 package.scala 96:25:@46662.4]
  wire  _T_270; // @[package.scala 96:25:@46679.4 package.scala 96:25:@46680.4]
  wire  _T_274; // @[Controllers.scala 169:67:@46682.4]
  wire  _T_275; // @[Controllers.scala 169:86:@46683.4]
  wire  _T_287; // @[Controllers.scala 165:35:@46695.4]
  wire  _T_289; // @[Controllers.scala 165:60:@46696.4]
  wire  _T_290; // @[Controllers.scala 165:58:@46697.4]
  wire  _T_292; // @[Controllers.scala 165:76:@46698.4]
  wire  _T_293; // @[Controllers.scala 165:74:@46699.4]
  wire  _T_297; // @[Controllers.scala 165:109:@46702.4]
  wire  _T_300; // @[Controllers.scala 165:141:@46704.4]
  wire  _T_308; // @[package.scala 96:25:@46716.4 package.scala 96:25:@46717.4]
  wire  _T_312; // @[Controllers.scala 167:54:@46719.4]
  wire  _T_313; // @[Controllers.scala 167:52:@46720.4]
  wire  _T_320; // @[package.scala 96:25:@46730.4 package.scala 96:25:@46731.4]
  wire  _T_338; // @[package.scala 96:25:@46748.4 package.scala 96:25:@46749.4]
  wire  _T_342; // @[Controllers.scala 169:67:@46751.4]
  wire  _T_343; // @[Controllers.scala 169:86:@46752.4]
  wire  _T_358; // @[Controllers.scala 213:68:@46770.4]
  wire  _T_360; // @[Controllers.scala 213:90:@46772.4]
  wire  _T_362; // @[Controllers.scala 213:132:@46774.4]
  wire  _T_366; // @[Controllers.scala 213:68:@46779.4]
  wire  _T_368; // @[Controllers.scala 213:90:@46781.4]
  wire  _T_374; // @[Controllers.scala 213:68:@46787.4]
  wire  _T_376; // @[Controllers.scala 213:90:@46789.4]
  wire  _T_383; // @[package.scala 100:49:@46795.4]
  reg  _T_386; // @[package.scala 48:56:@46796.4]
  reg [31:0] _RAND_0;
  wire  _T_387; // @[package.scala 100:41:@46798.4]
  reg  _T_400; // @[package.scala 48:56:@46814.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@46460.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@46463.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF active_2 ( // @[Controllers.scala 76:50:@46466.4]
    .clock(active_2_clock),
    .reset(active_2_reset),
    .io_input_set(active_2_io_input_set),
    .io_input_reset(active_2_io_input_reset),
    .io_input_asyn_reset(active_2_io_input_asyn_reset),
    .io_output(active_2_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@46469.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@46472.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF done_2 ( // @[Controllers.scala 77:48:@46475.4]
    .clock(done_2_clock),
    .reset(done_2_reset),
    .io_input_set(done_2_io_input_set),
    .io_input_reset(done_2_io_input_reset),
    .io_input_asyn_reset(done_2_io_input_asyn_reset),
    .io_output(done_2_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@46516.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@46519.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  SRFF iterDone_2 ( // @[Controllers.scala 90:52:@46522.4]
    .clock(iterDone_2_clock),
    .reset(iterDone_2_reset),
    .io_input_set(iterDone_2_io_input_set),
    .io_input_reset(iterDone_2_io_input_reset),
    .io_input_asyn_reset(iterDone_2_io_input_asyn_reset),
    .io_output(iterDone_2_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@46573.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@46587.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@46605.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@46642.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@46656.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@46674.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@46711.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@46725.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper RetimeWrapper_8 ( // @[package.scala 93:22:@46743.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper RetimeWrapper_9 ( // @[package.scala 93:22:@46800.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper RetimeWrapper_10 ( // @[package.scala 93:22:@46817.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  assign _T_77 = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@46478.4]
  assign allDone = _T_77 & done_2_io_output; // @[Controllers.scala 80:47:@46479.4]
  assign _T_151 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@46557.4]
  assign _T_153 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@46558.4]
  assign _T_154 = _T_151 & _T_153; // @[Controllers.scala 165:58:@46559.4]
  assign _T_156 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@46560.4]
  assign _T_157 = _T_154 & _T_156; // @[Controllers.scala 165:74:@46561.4]
  assign _T_161 = _T_157 & io_enable; // @[Controllers.scala 165:109:@46564.4]
  assign _T_164 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@46566.4]
  assign _T_172 = RetimeWrapper_io_out; // @[package.scala 96:25:@46578.4 package.scala 96:25:@46579.4]
  assign _T_176 = _T_172 == 1'h0; // @[Controllers.scala 167:54:@46581.4]
  assign _T_177 = io_doneIn_0 | _T_176; // @[Controllers.scala 167:52:@46582.4]
  assign _T_184 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@46592.4 package.scala 96:25:@46593.4]
  assign _T_202 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@46610.4 package.scala 96:25:@46611.4]
  assign _T_206 = _T_202 == 1'h0; // @[Controllers.scala 169:67:@46613.4]
  assign _T_207 = _T_206 & io_enable; // @[Controllers.scala 169:86:@46614.4]
  assign _T_219 = ~ iterDone_1_io_output; // @[Controllers.scala 165:35:@46626.4]
  assign _T_221 = io_doneIn_1 == 1'h0; // @[Controllers.scala 165:60:@46627.4]
  assign _T_222 = _T_219 & _T_221; // @[Controllers.scala 165:58:@46628.4]
  assign _T_224 = done_1_io_output == 1'h0; // @[Controllers.scala 165:76:@46629.4]
  assign _T_225 = _T_222 & _T_224; // @[Controllers.scala 165:74:@46630.4]
  assign _T_229 = _T_225 & io_enable; // @[Controllers.scala 165:109:@46633.4]
  assign _T_232 = io_ctrCopyDone_1 == 1'h0; // @[Controllers.scala 165:141:@46635.4]
  assign _T_240 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@46647.4 package.scala 96:25:@46648.4]
  assign _T_244 = _T_240 == 1'h0; // @[Controllers.scala 167:54:@46650.4]
  assign _T_245 = io_doneIn_1 | _T_244; // @[Controllers.scala 167:52:@46651.4]
  assign _T_252 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@46661.4 package.scala 96:25:@46662.4]
  assign _T_270 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@46679.4 package.scala 96:25:@46680.4]
  assign _T_274 = _T_270 == 1'h0; // @[Controllers.scala 169:67:@46682.4]
  assign _T_275 = _T_274 & io_enable; // @[Controllers.scala 169:86:@46683.4]
  assign _T_287 = ~ iterDone_2_io_output; // @[Controllers.scala 165:35:@46695.4]
  assign _T_289 = io_doneIn_2 == 1'h0; // @[Controllers.scala 165:60:@46696.4]
  assign _T_290 = _T_287 & _T_289; // @[Controllers.scala 165:58:@46697.4]
  assign _T_292 = done_2_io_output == 1'h0; // @[Controllers.scala 165:76:@46698.4]
  assign _T_293 = _T_290 & _T_292; // @[Controllers.scala 165:74:@46699.4]
  assign _T_297 = _T_293 & io_enable; // @[Controllers.scala 165:109:@46702.4]
  assign _T_300 = io_ctrCopyDone_2 == 1'h0; // @[Controllers.scala 165:141:@46704.4]
  assign _T_308 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@46716.4 package.scala 96:25:@46717.4]
  assign _T_312 = _T_308 == 1'h0; // @[Controllers.scala 167:54:@46719.4]
  assign _T_313 = io_doneIn_2 | _T_312; // @[Controllers.scala 167:52:@46720.4]
  assign _T_320 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@46730.4 package.scala 96:25:@46731.4]
  assign _T_338 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@46748.4 package.scala 96:25:@46749.4]
  assign _T_342 = _T_338 == 1'h0; // @[Controllers.scala 169:67:@46751.4]
  assign _T_343 = _T_342 & io_enable; // @[Controllers.scala 169:86:@46752.4]
  assign _T_358 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@46770.4]
  assign _T_360 = _T_358 & _T_151; // @[Controllers.scala 213:90:@46772.4]
  assign _T_362 = ~ allDone; // @[Controllers.scala 213:132:@46774.4]
  assign _T_366 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@46779.4]
  assign _T_368 = _T_366 & _T_219; // @[Controllers.scala 213:90:@46781.4]
  assign _T_374 = io_enable & active_2_io_output; // @[Controllers.scala 213:68:@46787.4]
  assign _T_376 = _T_374 & _T_287; // @[Controllers.scala 213:90:@46789.4]
  assign _T_383 = allDone == 1'h0; // @[package.scala 100:49:@46795.4]
  assign _T_387 = allDone & _T_386; // @[package.scala 100:41:@46798.4]
  assign io_done = RetimeWrapper_10_io_out; // @[Controllers.scala 245:13:@46824.4]
  assign io_enableOut_0 = _T_360 & _T_362; // @[Controllers.scala 213:55:@46778.4]
  assign io_enableOut_1 = _T_368 & _T_362; // @[Controllers.scala 213:55:@46786.4]
  assign io_enableOut_2 = _T_376 & _T_362; // @[Controllers.scala 213:55:@46794.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@46765.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@46767.4]
  assign io_childAck_2 = iterDone_2_io_output; // @[Controllers.scala 212:58:@46769.4]
  assign active_0_clock = clock; // @[:@46461.4]
  assign active_0_reset = reset; // @[:@46462.4]
  assign active_0_io_input_set = _T_161 & _T_164; // @[Controllers.scala 165:32:@46568.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@46572.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@46482.4]
  assign active_1_clock = clock; // @[:@46464.4]
  assign active_1_reset = reset; // @[:@46465.4]
  assign active_1_io_input_set = _T_229 & _T_232; // @[Controllers.scala 165:32:@46637.4]
  assign active_1_io_input_reset = io_ctrCopyDone_1 | io_parentAck; // @[Controllers.scala 166:34:@46641.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@46483.4]
  assign active_2_clock = clock; // @[:@46467.4]
  assign active_2_reset = reset; // @[:@46468.4]
  assign active_2_io_input_set = _T_297 & _T_300; // @[Controllers.scala 165:32:@46706.4]
  assign active_2_io_input_reset = io_ctrCopyDone_2 | io_parentAck; // @[Controllers.scala 166:34:@46710.4]
  assign active_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@46484.4]
  assign done_0_clock = clock; // @[:@46470.4]
  assign done_0_reset = reset; // @[:@46471.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_207; // @[Controllers.scala 169:30:@46618.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@46496.4 Controllers.scala 170:32:@46625.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@46485.4]
  assign done_1_clock = clock; // @[:@46473.4]
  assign done_1_reset = reset; // @[:@46474.4]
  assign done_1_io_input_set = io_ctrCopyDone_1 | _T_275; // @[Controllers.scala 169:30:@46687.4]
  assign done_1_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@46505.4 Controllers.scala 170:32:@46694.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@46486.4]
  assign done_2_clock = clock; // @[:@46476.4]
  assign done_2_reset = reset; // @[:@46477.4]
  assign done_2_io_input_set = io_ctrCopyDone_2 | _T_343; // @[Controllers.scala 169:30:@46756.4]
  assign done_2_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@46514.4 Controllers.scala 170:32:@46763.4]
  assign done_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@46487.4]
  assign iterDone_0_clock = clock; // @[:@46517.4]
  assign iterDone_0_reset = reset; // @[:@46518.4]
  assign iterDone_0_io_input_set = _T_177 & io_enable; // @[Controllers.scala 167:34:@46586.4]
  assign iterDone_0_io_input_reset = _T_184 | io_parentAck; // @[Controllers.scala 92:37:@46536.4 Controllers.scala 168:36:@46602.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@46525.4]
  assign iterDone_1_clock = clock; // @[:@46520.4]
  assign iterDone_1_reset = reset; // @[:@46521.4]
  assign iterDone_1_io_input_set = _T_245 & io_enable; // @[Controllers.scala 167:34:@46655.4]
  assign iterDone_1_io_input_reset = _T_252 | io_parentAck; // @[Controllers.scala 92:37:@46545.4 Controllers.scala 168:36:@46671.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@46526.4]
  assign iterDone_2_clock = clock; // @[:@46523.4]
  assign iterDone_2_reset = reset; // @[:@46524.4]
  assign iterDone_2_io_input_set = _T_313 & io_enable; // @[Controllers.scala 167:34:@46724.4]
  assign iterDone_2_io_input_reset = _T_320 | io_parentAck; // @[Controllers.scala 92:37:@46554.4 Controllers.scala 168:36:@46740.4]
  assign iterDone_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@46527.4]
  assign RetimeWrapper_clock = clock; // @[:@46574.4]
  assign RetimeWrapper_reset = reset; // @[:@46575.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@46577.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@46576.4]
  assign RetimeWrapper_1_clock = clock; // @[:@46588.4]
  assign RetimeWrapper_1_reset = reset; // @[:@46589.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@46591.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@46590.4]
  assign RetimeWrapper_2_clock = clock; // @[:@46606.4]
  assign RetimeWrapper_2_reset = reset; // @[:@46607.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@46609.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@46608.4]
  assign RetimeWrapper_3_clock = clock; // @[:@46643.4]
  assign RetimeWrapper_3_reset = reset; // @[:@46644.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@46646.4]
  assign RetimeWrapper_3_io_in = 1'h1; // @[package.scala 94:16:@46645.4]
  assign RetimeWrapper_4_clock = clock; // @[:@46657.4]
  assign RetimeWrapper_4_reset = reset; // @[:@46658.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@46660.4]
  assign RetimeWrapper_4_io_in = io_doneIn_1; // @[package.scala 94:16:@46659.4]
  assign RetimeWrapper_5_clock = clock; // @[:@46675.4]
  assign RetimeWrapper_5_reset = reset; // @[:@46676.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@46678.4]
  assign RetimeWrapper_5_io_in = 1'h1; // @[package.scala 94:16:@46677.4]
  assign RetimeWrapper_6_clock = clock; // @[:@46712.4]
  assign RetimeWrapper_6_reset = reset; // @[:@46713.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@46715.4]
  assign RetimeWrapper_6_io_in = 1'h1; // @[package.scala 94:16:@46714.4]
  assign RetimeWrapper_7_clock = clock; // @[:@46726.4]
  assign RetimeWrapper_7_reset = reset; // @[:@46727.4]
  assign RetimeWrapper_7_io_flow = 1'h1; // @[package.scala 95:18:@46729.4]
  assign RetimeWrapper_7_io_in = io_doneIn_2; // @[package.scala 94:16:@46728.4]
  assign RetimeWrapper_8_clock = clock; // @[:@46744.4]
  assign RetimeWrapper_8_reset = reset; // @[:@46745.4]
  assign RetimeWrapper_8_io_flow = 1'h1; // @[package.scala 95:18:@46747.4]
  assign RetimeWrapper_8_io_in = 1'h1; // @[package.scala 94:16:@46746.4]
  assign RetimeWrapper_9_clock = clock; // @[:@46801.4]
  assign RetimeWrapper_9_reset = reset; // @[:@46802.4]
  assign RetimeWrapper_9_io_flow = 1'h1; // @[package.scala 95:18:@46804.4]
  assign RetimeWrapper_9_io_in = _T_387 | io_parentAck; // @[package.scala 94:16:@46803.4]
  assign RetimeWrapper_10_clock = clock; // @[:@46818.4]
  assign RetimeWrapper_10_reset = reset; // @[:@46819.4]
  assign RetimeWrapper_10_io_flow = io_enable; // @[package.scala 95:18:@46821.4]
  assign RetimeWrapper_10_io_in = allDone & _T_400; // @[package.scala 94:16:@46820.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_386 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_400 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_386 <= 1'h0;
    end else begin
      _T_386 <= _T_383;
    end
    if (reset) begin
      _T_400 <= 1'h0;
    end else begin
      _T_400 <= _T_383;
    end
  end
endmodule
module x746_inr_UnitPipe_sm( // @[:@46997.2]
  input   clock, // @[:@46998.4]
  input   reset, // @[:@46999.4]
  input   io_enable, // @[:@47000.4]
  output  io_done, // @[:@47000.4]
  output  io_doneLatch, // @[:@47000.4]
  input   io_ctrDone, // @[:@47000.4]
  output  io_datapathEn, // @[:@47000.4]
  output  io_ctrInc, // @[:@47000.4]
  input   io_parentAck, // @[:@47000.4]
  input   io_backpressure // @[:@47000.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@47002.4]
  wire  active_reset; // @[Controllers.scala 261:22:@47002.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@47002.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@47002.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@47002.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@47002.4]
  wire  done_clock; // @[Controllers.scala 262:20:@47005.4]
  wire  done_reset; // @[Controllers.scala 262:20:@47005.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@47005.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@47005.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@47005.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@47005.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@47059.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@47059.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@47059.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@47059.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@47059.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@47067.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@47067.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@47067.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@47067.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@47067.4]
  wire  _T_80; // @[Controllers.scala 264:48:@47010.4]
  wire  _T_81; // @[Controllers.scala 264:46:@47011.4]
  wire  _T_82; // @[Controllers.scala 264:62:@47012.4]
  wire  _T_83; // @[Controllers.scala 264:60:@47013.4]
  wire  _T_100; // @[package.scala 100:49:@47030.4]
  reg  _T_103; // @[package.scala 48:56:@47031.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 100:49:@47039.4]
  wire  _T_116; // @[Controllers.scala 283:41:@47047.4]
  wire  _T_117; // @[Controllers.scala 283:59:@47048.4]
  wire  _T_119; // @[Controllers.scala 284:37:@47051.4]
  reg  _T_125; // @[package.scala 48:56:@47055.4]
  reg [31:0] _RAND_1;
  reg  _T_142; // @[Controllers.scala 291:31:@47077.4]
  reg [31:0] _RAND_2;
  reg  _T_149; // @[package.scala 48:56:@47080.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:41:@47082.4]
  wire  _T_152; // @[Controllers.scala 292:61:@47083.4]
  wire  _T_153; // @[Controllers.scala 292:24:@47084.4]
  SRFF active ( // @[Controllers.scala 261:22:@47002.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@47005.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@47059.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@47067.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@47010.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@47011.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@47012.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@47013.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@47030.4]
  assign _T_108 = done_io_output == 1'h0; // @[package.scala 100:49:@47039.4]
  assign _T_116 = active_io_output & _T_82; // @[Controllers.scala 283:41:@47047.4]
  assign _T_117 = _T_116 & io_enable; // @[Controllers.scala 283:59:@47048.4]
  assign _T_119 = active_io_output & io_enable; // @[Controllers.scala 284:37:@47051.4]
  assign _T_150 = done_io_output & _T_149; // @[package.scala 100:41:@47082.4]
  assign _T_152 = _T_150 ? 1'h1 : _T_142; // @[Controllers.scala 292:61:@47083.4]
  assign _T_153 = io_parentAck ? 1'h0 : _T_152; // @[Controllers.scala 292:24:@47084.4]
  assign io_done = done_io_output & _T_125; // @[Controllers.scala 287:13:@47058.4]
  assign io_doneLatch = _T_142; // @[Controllers.scala 293:18:@47086.4]
  assign io_datapathEn = _T_117 & io_backpressure; // @[Controllers.scala 283:21:@47050.4]
  assign io_ctrInc = _T_119 & io_backpressure; // @[Controllers.scala 284:17:@47053.4]
  assign active_clock = clock; // @[:@47003.4]
  assign active_reset = reset; // @[:@47004.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@47015.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@47019.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@47020.4]
  assign done_clock = clock; // @[:@47006.4]
  assign done_reset = reset; // @[:@47007.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@47035.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@47028.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@47029.4]
  assign RetimeWrapper_clock = clock; // @[:@47060.4]
  assign RetimeWrapper_reset = reset; // @[:@47061.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@47063.4]
  assign RetimeWrapper_io_in = 1'h0; // @[package.scala 94:16:@47062.4]
  assign RetimeWrapper_1_clock = clock; // @[:@47068.4]
  assign RetimeWrapper_1_reset = reset; // @[:@47069.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@47071.4]
  assign RetimeWrapper_1_io_in = io_ctrDone; // @[package.scala 94:16:@47070.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_125 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_142 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_149 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_125 <= 1'h0;
    end else begin
      _T_125 <= _T_108;
    end
    if (reset) begin
      _T_142 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_142 <= 1'h0;
      end else begin
        if (_T_150) begin
          _T_142 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_149 <= 1'h0;
    end else begin
      _T_149 <= _T_108;
    end
  end
endmodule
module x746_inr_UnitPipe_kernelx746_inr_UnitPipe_concrete1( // @[:@47161.2]
  output        io_in_x739_valid, // @[:@47164.4]
  output [63:0] io_in_x739_bits_addr, // @[:@47164.4]
  output [31:0] io_in_x739_bits_size, // @[:@47164.4]
  input  [63:0] io_in_x478_outdram_number, // @[:@47164.4]
  input         io_sigsIn_backpressure, // @[:@47164.4]
  input         io_sigsIn_datapathEn, // @[:@47164.4]
  input         io_rr // @[:@47164.4]
);
  wire [96:0] x743_tuple; // @[Cat.scala 30:58:@47178.4]
  wire  _T_135; // @[implicits.scala 55:10:@47181.4]
  assign x743_tuple = {33'h1fa400,io_in_x478_outdram_number}; // @[Cat.scala 30:58:@47178.4]
  assign _T_135 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 55:10:@47181.4]
  assign io_in_x739_valid = _T_135 & io_sigsIn_backpressure; // @[sm_x746_inr_UnitPipe.scala 65:18:@47184.4]
  assign io_in_x739_bits_addr = x743_tuple[63:0]; // @[sm_x746_inr_UnitPipe.scala 66:22:@47186.4]
  assign io_in_x739_bits_size = x743_tuple[95:64]; // @[sm_x746_inr_UnitPipe.scala 67:22:@47188.4]
endmodule
module FF_13( // @[:@47190.2]
  input         clock, // @[:@47191.4]
  input         reset, // @[:@47192.4]
  output [22:0] io_rPort_0_output_0, // @[:@47193.4]
  input  [22:0] io_wPort_0_data_0, // @[:@47193.4]
  input         io_wPort_0_reset, // @[:@47193.4]
  input         io_wPort_0_en_0 // @[:@47193.4]
);
  reg [22:0] ff; // @[MemPrimitives.scala 311:19:@47208.4]
  reg [31:0] _RAND_0;
  wire [22:0] _T_68; // @[MemPrimitives.scala 315:32:@47210.4]
  wire [22:0] _T_69; // @[MemPrimitives.scala 315:12:@47211.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 315:32:@47210.4]
  assign _T_69 = io_wPort_0_reset ? 23'h0 : _T_68; // @[MemPrimitives.scala 315:12:@47211.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 316:34:@47213.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[22:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 23'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 23'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SingleCounter_5( // @[:@47228.2]
  input         clock, // @[:@47229.4]
  input         reset, // @[:@47230.4]
  input         io_input_reset, // @[:@47231.4]
  input         io_input_enable, // @[:@47231.4]
  output [22:0] io_output_count_0, // @[:@47231.4]
  output        io_output_oobs_0, // @[:@47231.4]
  output        io_output_done // @[:@47231.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@47244.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@47244.4]
  wire [22:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@47244.4]
  wire [22:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@47244.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@47244.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@47244.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@47260.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@47260.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@47260.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@47260.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@47260.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@47260.4]
  wire  _T_36; // @[Counter.scala 264:45:@47263.4]
  wire [22:0] _T_48; // @[Counter.scala 287:52:@47288.4]
  wire [23:0] _T_50; // @[Counter.scala 291:33:@47289.4]
  wire [22:0] _T_51; // @[Counter.scala 291:33:@47290.4]
  wire [22:0] _T_52; // @[Counter.scala 291:33:@47291.4]
  wire  _T_57; // @[Counter.scala 293:18:@47293.4]
  wire [22:0] _T_68; // @[Counter.scala 299:115:@47301.4]
  wire [22:0] _T_71; // @[Counter.scala 299:152:@47304.4]
  wire [22:0] _T_72; // @[Counter.scala 299:74:@47305.4]
  wire  _T_75; // @[Counter.scala 322:102:@47309.4]
  wire  _T_77; // @[Counter.scala 322:130:@47310.4]
  FF_13 bases_0 ( // @[Counter.scala 261:53:@47244.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@47260.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@47263.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@47288.4]
  assign _T_50 = $signed(_T_48) + $signed(23'sh1); // @[Counter.scala 291:33:@47289.4]
  assign _T_51 = $signed(_T_48) + $signed(23'sh1); // @[Counter.scala 291:33:@47290.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@47291.4]
  assign _T_57 = $signed(_T_52) >= $signed(23'sh1fa400); // @[Counter.scala 293:18:@47293.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@47301.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@47304.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 299:74:@47305.4]
  assign _T_75 = $signed(_T_48) < $signed(23'sh0); // @[Counter.scala 322:102:@47309.4]
  assign _T_77 = $signed(_T_48) >= $signed(23'sh1fa400); // @[Counter.scala 322:130:@47310.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@47308.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@47312.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@47314.4]
  assign bases_0_clock = clock; // @[:@47245.4]
  assign bases_0_reset = reset; // @[:@47246.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 23'h0 : _T_72; // @[Counter.scala 299:31:@47307.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@47286.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@47287.4]
  assign SRFF_clock = clock; // @[:@47261.4]
  assign SRFF_reset = reset; // @[:@47262.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@47265.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@47267.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@47268.4]
endmodule
module x748_ctrchain( // @[:@47319.2]
  input         clock, // @[:@47320.4]
  input         reset, // @[:@47321.4]
  input         io_input_reset, // @[:@47322.4]
  input         io_input_enable, // @[:@47322.4]
  output [22:0] io_output_counts_0, // @[:@47322.4]
  output        io_output_oobs_0, // @[:@47322.4]
  output        io_output_done // @[:@47322.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 513:46:@47324.4]
  wire  ctrs_0_reset; // @[Counter.scala 513:46:@47324.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 513:46:@47324.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 513:46:@47324.4]
  wire [22:0] ctrs_0_io_output_count_0; // @[Counter.scala 513:46:@47324.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 513:46:@47324.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 513:46:@47324.4]
  reg  wasDone; // @[Counter.scala 542:24:@47333.4]
  reg [31:0] _RAND_0;
  wire  _T_45; // @[Counter.scala 546:69:@47339.4]
  wire  _T_47; // @[Counter.scala 546:80:@47340.4]
  reg  doneLatch; // @[Counter.scala 550:26:@47345.4]
  reg [31:0] _RAND_1;
  wire  _T_54; // @[Counter.scala 551:48:@47346.4]
  wire  _T_55; // @[Counter.scala 551:19:@47347.4]
  SingleCounter_5 ctrs_0 ( // @[Counter.scala 513:46:@47324.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done)
  );
  assign _T_45 = io_input_enable & ctrs_0_io_output_done; // @[Counter.scala 546:69:@47339.4]
  assign _T_47 = wasDone == 1'h0; // @[Counter.scala 546:80:@47340.4]
  assign _T_54 = ctrs_0_io_output_done ? 1'h1 : doneLatch; // @[Counter.scala 551:48:@47346.4]
  assign _T_55 = io_input_reset ? 1'h0 : _T_54; // @[Counter.scala 551:19:@47347.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 557:32:@47349.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@47351.4]
  assign io_output_done = _T_45 & _T_47; // @[Counter.scala 546:18:@47342.4]
  assign ctrs_0_clock = clock; // @[:@47325.4]
  assign ctrs_0_reset = reset; // @[:@47326.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@47330.4]
  assign ctrs_0_io_input_enable = io_input_enable; // @[Counter.scala 524:33:@47331.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= ctrs_0_io_output_done;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (ctrs_0_io_output_done) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module x755_inr_Foreach_sm( // @[:@47539.2]
  input   clock, // @[:@47540.4]
  input   reset, // @[:@47541.4]
  input   io_enable, // @[:@47542.4]
  output  io_done, // @[:@47542.4]
  output  io_doneLatch, // @[:@47542.4]
  input   io_ctrDone, // @[:@47542.4]
  output  io_datapathEn, // @[:@47542.4]
  output  io_ctrInc, // @[:@47542.4]
  output  io_ctrRst, // @[:@47542.4]
  input   io_parentAck, // @[:@47542.4]
  input   io_backpressure, // @[:@47542.4]
  input   io_break // @[:@47542.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@47544.4]
  wire  active_reset; // @[Controllers.scala 261:22:@47544.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@47544.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@47544.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@47544.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@47544.4]
  wire  done_clock; // @[Controllers.scala 262:20:@47547.4]
  wire  done_reset; // @[Controllers.scala 262:20:@47547.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@47547.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@47547.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@47547.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@47547.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@47581.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@47581.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@47581.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@47581.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@47581.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@47603.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@47603.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@47603.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@47603.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@47603.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@47615.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@47615.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@47615.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@47615.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@47615.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@47623.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@47623.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@47623.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@47623.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@47623.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@47639.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@47639.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@47639.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@47639.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@47639.4]
  wire  _T_80; // @[Controllers.scala 264:48:@47552.4]
  wire  _T_81; // @[Controllers.scala 264:46:@47553.4]
  wire  _T_82; // @[Controllers.scala 264:62:@47554.4]
  wire  _T_83; // @[Controllers.scala 264:60:@47555.4]
  wire  _T_100; // @[package.scala 100:49:@47572.4]
  reg  _T_103; // @[package.scala 48:56:@47573.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@47586.4 package.scala 96:25:@47587.4]
  wire  _T_110; // @[package.scala 100:49:@47588.4]
  reg  _T_113; // @[package.scala 48:56:@47589.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@47591.4]
  wire  _T_118; // @[Controllers.scala 283:41:@47596.4]
  wire  _T_119; // @[Controllers.scala 283:59:@47597.4]
  wire  _T_121; // @[Controllers.scala 284:37:@47600.4]
  wire  _T_124; // @[package.scala 96:25:@47608.4 package.scala 96:25:@47609.4]
  wire  _T_126; // @[package.scala 100:49:@47610.4]
  reg  _T_129; // @[package.scala 48:56:@47611.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@47633.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@47635.4]
  reg  _T_153; // @[package.scala 48:56:@47636.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@47644.4 package.scala 96:25:@47645.4]
  wire  _T_158; // @[Controllers.scala 292:61:@47646.4]
  wire  _T_159; // @[Controllers.scala 292:24:@47647.4]
  SRFF active ( // @[Controllers.scala 261:22:@47544.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@47547.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@47581.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@47603.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@47615.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@47623.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@47639.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@47552.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@47553.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@47554.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@47555.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@47572.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@47586.4 package.scala 96:25:@47587.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@47588.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@47591.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@47596.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@47597.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@47600.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@47608.4 package.scala 96:25:@47609.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@47610.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@47635.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@47644.4 package.scala 96:25:@47645.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@47646.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@47647.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@47614.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@47649.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@47599.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@47602.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@47594.4]
  assign active_clock = clock; // @[:@47545.4]
  assign active_reset = reset; // @[:@47546.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@47557.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@47561.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@47562.4]
  assign done_clock = clock; // @[:@47548.4]
  assign done_reset = reset; // @[:@47549.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@47577.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@47570.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@47571.4]
  assign RetimeWrapper_clock = clock; // @[:@47582.4]
  assign RetimeWrapper_reset = reset; // @[:@47583.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@47585.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@47584.4]
  assign RetimeWrapper_1_clock = clock; // @[:@47604.4]
  assign RetimeWrapper_1_reset = reset; // @[:@47605.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@47607.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@47606.4]
  assign RetimeWrapper_2_clock = clock; // @[:@47616.4]
  assign RetimeWrapper_2_reset = reset; // @[:@47617.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@47619.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@47618.4]
  assign RetimeWrapper_3_clock = clock; // @[:@47624.4]
  assign RetimeWrapper_3_reset = reset; // @[:@47625.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@47627.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@47626.4]
  assign RetimeWrapper_4_clock = clock; // @[:@47640.4]
  assign RetimeWrapper_4_reset = reset; // @[:@47641.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@47643.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@47642.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x755_inr_Foreach_kernelx755_inr_Foreach_concrete1( // @[:@47861.2]
  input         clock, // @[:@47862.4]
  input         reset, // @[:@47863.4]
  output [20:0] io_in_x482_outbuf_0_rPort_0_ofs_0, // @[:@47864.4]
  output        io_in_x482_outbuf_0_rPort_0_en_0, // @[:@47864.4]
  output        io_in_x482_outbuf_0_rPort_0_backpressure, // @[:@47864.4]
  input  [7:0]  io_in_x482_outbuf_0_rPort_0_output_0, // @[:@47864.4]
  output        io_in_x740_valid, // @[:@47864.4]
  output [7:0]  io_in_x740_bits_wdata_0, // @[:@47864.4]
  output        io_in_x740_bits_wstrb, // @[:@47864.4]
  input         io_sigsIn_backpressure, // @[:@47864.4]
  input         io_sigsIn_datapathEn, // @[:@47864.4]
  input         io_sigsIn_break, // @[:@47864.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@47864.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@47864.4]
  input         io_rr // @[:@47864.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@47891.4]
  wire [31:0] __io_result; // @[Math.scala 709:24:@47891.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@47920.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@47920.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@47920.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@47920.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@47920.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@47929.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@47929.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@47929.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@47929.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@47929.4]
  wire  b750; // @[sm_x755_inr_Foreach.scala 62:18:@47899.4]
  wire  _T_274; // @[sm_x755_inr_Foreach.scala 67:129:@47903.4]
  wire  _T_278; // @[implicits.scala 55:10:@47906.4]
  wire  _T_279; // @[sm_x755_inr_Foreach.scala 67:146:@47907.4]
  wire [8:0] x753_tuple; // @[Cat.scala 30:58:@47917.4]
  wire  _T_290; // @[package.scala 96:25:@47934.4 package.scala 96:25:@47935.4]
  wire  _T_292; // @[implicits.scala 55:10:@47936.4]
  wire  x906_b750_D2; // @[package.scala 96:25:@47925.4 package.scala 96:25:@47926.4]
  wire  _T_293; // @[sm_x755_inr_Foreach.scala 74:112:@47937.4]
  wire [31:0] b749_number; // @[Math.scala 712:22:@47896.4 Math.scala 713:14:@47897.4]
  _ _ ( // @[Math.scala 709:24:@47891.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@47920.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@47929.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign b750 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x755_inr_Foreach.scala 62:18:@47899.4]
  assign _T_274 = ~ io_sigsIn_break; // @[sm_x755_inr_Foreach.scala 67:129:@47903.4]
  assign _T_278 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 55:10:@47906.4]
  assign _T_279 = _T_274 & _T_278; // @[sm_x755_inr_Foreach.scala 67:146:@47907.4]
  assign x753_tuple = {1'h1,io_in_x482_outbuf_0_rPort_0_output_0}; // @[Cat.scala 30:58:@47917.4]
  assign _T_290 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@47934.4 package.scala 96:25:@47935.4]
  assign _T_292 = io_rr ? _T_290 : 1'h0; // @[implicits.scala 55:10:@47936.4]
  assign x906_b750_D2 = RetimeWrapper_io_out; // @[package.scala 96:25:@47925.4 package.scala 96:25:@47926.4]
  assign _T_293 = _T_292 & x906_b750_D2; // @[sm_x755_inr_Foreach.scala 74:112:@47937.4]
  assign b749_number = __io_result; // @[Math.scala 712:22:@47896.4 Math.scala 713:14:@47897.4]
  assign io_in_x482_outbuf_0_rPort_0_ofs_0 = b749_number[20:0]; // @[MemInterfaceType.scala 107:54:@47910.4]
  assign io_in_x482_outbuf_0_rPort_0_en_0 = _T_279 & b750; // @[MemInterfaceType.scala 110:79:@47912.4]
  assign io_in_x482_outbuf_0_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@47911.4]
  assign io_in_x740_valid = _T_293 & io_sigsIn_backpressure; // @[sm_x755_inr_Foreach.scala 74:18:@47939.4]
  assign io_in_x740_bits_wdata_0 = x753_tuple[7:0]; // @[sm_x755_inr_Foreach.scala 75:26:@47941.4]
  assign io_in_x740_bits_wstrb = x753_tuple[8]; // @[sm_x755_inr_Foreach.scala 76:23:@47943.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 710:17:@47894.4]
  assign RetimeWrapper_clock = clock; // @[:@47921.4]
  assign RetimeWrapper_reset = reset; // @[:@47922.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47924.4]
  assign RetimeWrapper_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@47923.4]
  assign RetimeWrapper_1_clock = clock; // @[:@47930.4]
  assign RetimeWrapper_1_reset = reset; // @[:@47931.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47933.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@47932.4]
endmodule
module x759_inr_UnitPipe_sm( // @[:@48099.2]
  input   clock, // @[:@48100.4]
  input   reset, // @[:@48101.4]
  input   io_enable, // @[:@48102.4]
  output  io_done, // @[:@48102.4]
  output  io_doneLatch, // @[:@48102.4]
  input   io_ctrDone, // @[:@48102.4]
  output  io_datapathEn, // @[:@48102.4]
  output  io_ctrInc, // @[:@48102.4]
  input   io_parentAck // @[:@48102.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@48104.4]
  wire  active_reset; // @[Controllers.scala 261:22:@48104.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@48104.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@48104.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@48104.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@48104.4]
  wire  done_clock; // @[Controllers.scala 262:20:@48107.4]
  wire  done_reset; // @[Controllers.scala 262:20:@48107.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@48107.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@48107.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@48107.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@48107.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@48141.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@48141.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@48141.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@48141.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@48141.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@48163.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@48163.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@48163.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@48163.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@48163.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@48175.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@48175.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@48175.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@48175.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@48175.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@48183.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@48183.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@48183.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@48183.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@48183.4]
  wire  _T_80; // @[Controllers.scala 264:48:@48112.4]
  wire  _T_81; // @[Controllers.scala 264:46:@48113.4]
  wire  _T_82; // @[Controllers.scala 264:62:@48114.4]
  wire  _T_100; // @[package.scala 100:49:@48132.4]
  reg  _T_103; // @[package.scala 48:56:@48133.4]
  reg [31:0] _RAND_0;
  wire  _T_118; // @[Controllers.scala 283:41:@48156.4]
  wire  _T_124; // @[package.scala 96:25:@48168.4 package.scala 96:25:@48169.4]
  wire  _T_126; // @[package.scala 100:49:@48170.4]
  reg  _T_129; // @[package.scala 48:56:@48171.4]
  reg [31:0] _RAND_1;
  reg  _T_146; // @[Controllers.scala 291:31:@48193.4]
  reg [31:0] _RAND_2;
  wire  _T_150; // @[package.scala 100:49:@48195.4]
  reg  _T_153; // @[package.scala 48:56:@48196.4]
  reg [31:0] _RAND_3;
  wire  _T_154; // @[package.scala 100:41:@48198.4]
  wire  _T_156; // @[Controllers.scala 292:61:@48199.4]
  wire  _T_157; // @[Controllers.scala 292:24:@48200.4]
  SRFF active ( // @[Controllers.scala 261:22:@48104.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@48107.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@48141.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@48163.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@48175.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@48183.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@48112.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@48113.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@48114.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@48132.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@48156.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@48168.4 package.scala 96:25:@48169.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@48170.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@48195.4]
  assign _T_154 = done_io_output & _T_153; // @[package.scala 100:41:@48198.4]
  assign _T_156 = _T_154 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@48199.4]
  assign _T_157 = io_parentAck ? 1'h0 : _T_156; // @[Controllers.scala 292:24:@48200.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@48174.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@48202.4]
  assign io_datapathEn = _T_118 & io_enable; // @[Controllers.scala 283:21:@48159.4]
  assign io_ctrInc = active_io_output & io_enable; // @[Controllers.scala 284:17:@48162.4]
  assign active_clock = clock; // @[:@48105.4]
  assign active_reset = reset; // @[:@48106.4]
  assign active_io_input_set = _T_81 & _T_82; // @[Controllers.scala 264:23:@48117.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@48121.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@48122.4]
  assign done_clock = clock; // @[:@48108.4]
  assign done_reset = reset; // @[:@48109.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@48137.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@48130.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@48131.4]
  assign RetimeWrapper_clock = clock; // @[:@48142.4]
  assign RetimeWrapper_reset = reset; // @[:@48143.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@48145.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@48144.4]
  assign RetimeWrapper_1_clock = clock; // @[:@48164.4]
  assign RetimeWrapper_1_reset = reset; // @[:@48165.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@48167.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@48166.4]
  assign RetimeWrapper_2_clock = clock; // @[:@48176.4]
  assign RetimeWrapper_2_reset = reset; // @[:@48177.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@48179.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@48178.4]
  assign RetimeWrapper_3_clock = clock; // @[:@48184.4]
  assign RetimeWrapper_3_reset = reset; // @[:@48185.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@48187.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@48186.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_129 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_146 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_153 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_154) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x759_inr_UnitPipe_kernelx759_inr_UnitPipe_concrete1( // @[:@48277.2]
  output  io_in_x741_ready, // @[:@48280.4]
  input   io_sigsIn_datapathEn // @[:@48280.4]
);
  assign io_in_x741_ready = io_sigsIn_datapathEn; // @[sm_x759_inr_UnitPipe.scala 57:18:@48292.4]
endmodule
module x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1( // @[:@48295.2]
  input         clock, // @[:@48296.4]
  input         reset, // @[:@48297.4]
  output        io_in_x741_ready, // @[:@48298.4]
  input         io_in_x741_valid, // @[:@48298.4]
  input         io_in_x739_ready, // @[:@48298.4]
  output        io_in_x739_valid, // @[:@48298.4]
  output [63:0] io_in_x739_bits_addr, // @[:@48298.4]
  output [31:0] io_in_x739_bits_size, // @[:@48298.4]
  output [20:0] io_in_x482_outbuf_0_rPort_0_ofs_0, // @[:@48298.4]
  output        io_in_x482_outbuf_0_rPort_0_en_0, // @[:@48298.4]
  output        io_in_x482_outbuf_0_rPort_0_backpressure, // @[:@48298.4]
  input  [7:0]  io_in_x482_outbuf_0_rPort_0_output_0, // @[:@48298.4]
  input  [63:0] io_in_x478_outdram_number, // @[:@48298.4]
  input         io_in_x740_ready, // @[:@48298.4]
  output        io_in_x740_valid, // @[:@48298.4]
  output [7:0]  io_in_x740_bits_wdata_0, // @[:@48298.4]
  output        io_in_x740_bits_wstrb, // @[:@48298.4]
  input         io_sigsIn_smEnableOuts_0, // @[:@48298.4]
  input         io_sigsIn_smEnableOuts_1, // @[:@48298.4]
  input         io_sigsIn_smEnableOuts_2, // @[:@48298.4]
  input         io_sigsIn_smChildAcks_0, // @[:@48298.4]
  input         io_sigsIn_smChildAcks_1, // @[:@48298.4]
  input         io_sigsIn_smChildAcks_2, // @[:@48298.4]
  output        io_sigsOut_smDoneIn_0, // @[:@48298.4]
  output        io_sigsOut_smDoneIn_1, // @[:@48298.4]
  output        io_sigsOut_smDoneIn_2, // @[:@48298.4]
  output        io_sigsOut_smCtrCopyDone_0, // @[:@48298.4]
  output        io_sigsOut_smCtrCopyDone_1, // @[:@48298.4]
  output        io_sigsOut_smCtrCopyDone_2, // @[:@48298.4]
  input         io_rr // @[:@48298.4]
);
  wire  x746_inr_UnitPipe_sm_clock; // @[sm_x746_inr_UnitPipe.scala 33:18:@48365.4]
  wire  x746_inr_UnitPipe_sm_reset; // @[sm_x746_inr_UnitPipe.scala 33:18:@48365.4]
  wire  x746_inr_UnitPipe_sm_io_enable; // @[sm_x746_inr_UnitPipe.scala 33:18:@48365.4]
  wire  x746_inr_UnitPipe_sm_io_done; // @[sm_x746_inr_UnitPipe.scala 33:18:@48365.4]
  wire  x746_inr_UnitPipe_sm_io_doneLatch; // @[sm_x746_inr_UnitPipe.scala 33:18:@48365.4]
  wire  x746_inr_UnitPipe_sm_io_ctrDone; // @[sm_x746_inr_UnitPipe.scala 33:18:@48365.4]
  wire  x746_inr_UnitPipe_sm_io_datapathEn; // @[sm_x746_inr_UnitPipe.scala 33:18:@48365.4]
  wire  x746_inr_UnitPipe_sm_io_ctrInc; // @[sm_x746_inr_UnitPipe.scala 33:18:@48365.4]
  wire  x746_inr_UnitPipe_sm_io_parentAck; // @[sm_x746_inr_UnitPipe.scala 33:18:@48365.4]
  wire  x746_inr_UnitPipe_sm_io_backpressure; // @[sm_x746_inr_UnitPipe.scala 33:18:@48365.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@48422.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@48422.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@48422.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@48422.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@48422.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@48430.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@48430.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@48430.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@48430.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@48430.4]
  wire  x746_inr_UnitPipe_kernelx746_inr_UnitPipe_concrete1_io_in_x739_valid; // @[sm_x746_inr_UnitPipe.scala 69:24:@48460.4]
  wire [63:0] x746_inr_UnitPipe_kernelx746_inr_UnitPipe_concrete1_io_in_x739_bits_addr; // @[sm_x746_inr_UnitPipe.scala 69:24:@48460.4]
  wire [31:0] x746_inr_UnitPipe_kernelx746_inr_UnitPipe_concrete1_io_in_x739_bits_size; // @[sm_x746_inr_UnitPipe.scala 69:24:@48460.4]
  wire [63:0] x746_inr_UnitPipe_kernelx746_inr_UnitPipe_concrete1_io_in_x478_outdram_number; // @[sm_x746_inr_UnitPipe.scala 69:24:@48460.4]
  wire  x746_inr_UnitPipe_kernelx746_inr_UnitPipe_concrete1_io_sigsIn_backpressure; // @[sm_x746_inr_UnitPipe.scala 69:24:@48460.4]
  wire  x746_inr_UnitPipe_kernelx746_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x746_inr_UnitPipe.scala 69:24:@48460.4]
  wire  x746_inr_UnitPipe_kernelx746_inr_UnitPipe_concrete1_io_rr; // @[sm_x746_inr_UnitPipe.scala 69:24:@48460.4]
  wire  x748_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@48528.4]
  wire  x748_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@48528.4]
  wire  x748_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@48528.4]
  wire  x748_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@48528.4]
  wire [22:0] x748_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@48528.4]
  wire  x748_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@48528.4]
  wire  x748_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@48528.4]
  wire  x755_inr_Foreach_sm_clock; // @[sm_x755_inr_Foreach.scala 33:18:@48581.4]
  wire  x755_inr_Foreach_sm_reset; // @[sm_x755_inr_Foreach.scala 33:18:@48581.4]
  wire  x755_inr_Foreach_sm_io_enable; // @[sm_x755_inr_Foreach.scala 33:18:@48581.4]
  wire  x755_inr_Foreach_sm_io_done; // @[sm_x755_inr_Foreach.scala 33:18:@48581.4]
  wire  x755_inr_Foreach_sm_io_doneLatch; // @[sm_x755_inr_Foreach.scala 33:18:@48581.4]
  wire  x755_inr_Foreach_sm_io_ctrDone; // @[sm_x755_inr_Foreach.scala 33:18:@48581.4]
  wire  x755_inr_Foreach_sm_io_datapathEn; // @[sm_x755_inr_Foreach.scala 33:18:@48581.4]
  wire  x755_inr_Foreach_sm_io_ctrInc; // @[sm_x755_inr_Foreach.scala 33:18:@48581.4]
  wire  x755_inr_Foreach_sm_io_ctrRst; // @[sm_x755_inr_Foreach.scala 33:18:@48581.4]
  wire  x755_inr_Foreach_sm_io_parentAck; // @[sm_x755_inr_Foreach.scala 33:18:@48581.4]
  wire  x755_inr_Foreach_sm_io_backpressure; // @[sm_x755_inr_Foreach.scala 33:18:@48581.4]
  wire  x755_inr_Foreach_sm_io_break; // @[sm_x755_inr_Foreach.scala 33:18:@48581.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@48609.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@48609.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@48609.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@48609.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@48609.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@48649.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@48649.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@48649.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@48649.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@48649.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@48657.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@48657.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@48657.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@48657.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@48657.4]
  wire  x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_clock; // @[sm_x755_inr_Foreach.scala 78:24:@48692.4]
  wire  x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_reset; // @[sm_x755_inr_Foreach.scala 78:24:@48692.4]
  wire [20:0] x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_io_in_x482_outbuf_0_rPort_0_ofs_0; // @[sm_x755_inr_Foreach.scala 78:24:@48692.4]
  wire  x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_io_in_x482_outbuf_0_rPort_0_en_0; // @[sm_x755_inr_Foreach.scala 78:24:@48692.4]
  wire  x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_io_in_x482_outbuf_0_rPort_0_backpressure; // @[sm_x755_inr_Foreach.scala 78:24:@48692.4]
  wire [7:0] x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_io_in_x482_outbuf_0_rPort_0_output_0; // @[sm_x755_inr_Foreach.scala 78:24:@48692.4]
  wire  x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_io_in_x740_valid; // @[sm_x755_inr_Foreach.scala 78:24:@48692.4]
  wire [7:0] x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_io_in_x740_bits_wdata_0; // @[sm_x755_inr_Foreach.scala 78:24:@48692.4]
  wire  x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_io_in_x740_bits_wstrb; // @[sm_x755_inr_Foreach.scala 78:24:@48692.4]
  wire  x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_io_sigsIn_backpressure; // @[sm_x755_inr_Foreach.scala 78:24:@48692.4]
  wire  x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x755_inr_Foreach.scala 78:24:@48692.4]
  wire  x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x755_inr_Foreach.scala 78:24:@48692.4]
  wire [31:0] x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x755_inr_Foreach.scala 78:24:@48692.4]
  wire  x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x755_inr_Foreach.scala 78:24:@48692.4]
  wire  x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_io_rr; // @[sm_x755_inr_Foreach.scala 78:24:@48692.4]
  wire  x759_inr_UnitPipe_sm_clock; // @[sm_x759_inr_UnitPipe.scala 32:18:@48812.4]
  wire  x759_inr_UnitPipe_sm_reset; // @[sm_x759_inr_UnitPipe.scala 32:18:@48812.4]
  wire  x759_inr_UnitPipe_sm_io_enable; // @[sm_x759_inr_UnitPipe.scala 32:18:@48812.4]
  wire  x759_inr_UnitPipe_sm_io_done; // @[sm_x759_inr_UnitPipe.scala 32:18:@48812.4]
  wire  x759_inr_UnitPipe_sm_io_doneLatch; // @[sm_x759_inr_UnitPipe.scala 32:18:@48812.4]
  wire  x759_inr_UnitPipe_sm_io_ctrDone; // @[sm_x759_inr_UnitPipe.scala 32:18:@48812.4]
  wire  x759_inr_UnitPipe_sm_io_datapathEn; // @[sm_x759_inr_UnitPipe.scala 32:18:@48812.4]
  wire  x759_inr_UnitPipe_sm_io_ctrInc; // @[sm_x759_inr_UnitPipe.scala 32:18:@48812.4]
  wire  x759_inr_UnitPipe_sm_io_parentAck; // @[sm_x759_inr_UnitPipe.scala 32:18:@48812.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@48869.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@48869.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@48869.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@48869.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@48869.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@48877.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@48877.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@48877.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@48877.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@48877.4]
  wire  x759_inr_UnitPipe_kernelx759_inr_UnitPipe_concrete1_io_in_x741_ready; // @[sm_x759_inr_UnitPipe.scala 60:24:@48907.4]
  wire  x759_inr_UnitPipe_kernelx759_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x759_inr_UnitPipe.scala 60:24:@48907.4]
  wire  _T_359; // @[package.scala 100:49:@48393.4]
  reg  _T_362; // @[package.scala 48:56:@48394.4]
  reg [31:0] _RAND_0;
  wire  _T_375; // @[package.scala 96:25:@48427.4 package.scala 96:25:@48428.4]
  wire  _T_381; // @[package.scala 96:25:@48435.4 package.scala 96:25:@48436.4]
  wire  _T_384; // @[SpatialBlocks.scala 138:93:@48438.4]
  wire  _T_454; // @[package.scala 96:25:@48614.4 package.scala 96:25:@48615.4]
  wire  _T_468; // @[package.scala 96:25:@48654.4 package.scala 96:25:@48655.4]
  wire  _T_474; // @[package.scala 96:25:@48662.4 package.scala 96:25:@48663.4]
  wire  _T_477; // @[SpatialBlocks.scala 138:93:@48665.4]
  wire  _T_479; // @[SpatialBlocks.scala 157:36:@48674.4]
  wire  _T_480; // @[SpatialBlocks.scala 157:78:@48675.4]
  wire  _T_547; // @[package.scala 100:49:@48840.4]
  reg  _T_550; // @[package.scala 48:56:@48841.4]
  reg [31:0] _RAND_1;
  wire  x759_inr_UnitPipe_sigsIn_forwardpressure; // @[sm_x760_outr_UnitPipe.scala 101:55:@48847.4]
  wire  _T_563; // @[package.scala 96:25:@48874.4 package.scala 96:25:@48875.4]
  wire  _T_569; // @[package.scala 96:25:@48882.4 package.scala 96:25:@48883.4]
  wire  _T_572; // @[SpatialBlocks.scala 138:93:@48885.4]
  wire  x759_inr_UnitPipe_sigsIn_baseEn; // @[SpatialBlocks.scala 138:90:@48886.4]
  x746_inr_UnitPipe_sm x746_inr_UnitPipe_sm ( // @[sm_x746_inr_UnitPipe.scala 33:18:@48365.4]
    .clock(x746_inr_UnitPipe_sm_clock),
    .reset(x746_inr_UnitPipe_sm_reset),
    .io_enable(x746_inr_UnitPipe_sm_io_enable),
    .io_done(x746_inr_UnitPipe_sm_io_done),
    .io_doneLatch(x746_inr_UnitPipe_sm_io_doneLatch),
    .io_ctrDone(x746_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x746_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x746_inr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x746_inr_UnitPipe_sm_io_parentAck),
    .io_backpressure(x746_inr_UnitPipe_sm_io_backpressure)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@48422.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@48430.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x746_inr_UnitPipe_kernelx746_inr_UnitPipe_concrete1 x746_inr_UnitPipe_kernelx746_inr_UnitPipe_concrete1 ( // @[sm_x746_inr_UnitPipe.scala 69:24:@48460.4]
    .io_in_x739_valid(x746_inr_UnitPipe_kernelx746_inr_UnitPipe_concrete1_io_in_x739_valid),
    .io_in_x739_bits_addr(x746_inr_UnitPipe_kernelx746_inr_UnitPipe_concrete1_io_in_x739_bits_addr),
    .io_in_x739_bits_size(x746_inr_UnitPipe_kernelx746_inr_UnitPipe_concrete1_io_in_x739_bits_size),
    .io_in_x478_outdram_number(x746_inr_UnitPipe_kernelx746_inr_UnitPipe_concrete1_io_in_x478_outdram_number),
    .io_sigsIn_backpressure(x746_inr_UnitPipe_kernelx746_inr_UnitPipe_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x746_inr_UnitPipe_kernelx746_inr_UnitPipe_concrete1_io_sigsIn_datapathEn),
    .io_rr(x746_inr_UnitPipe_kernelx746_inr_UnitPipe_concrete1_io_rr)
  );
  x748_ctrchain x748_ctrchain ( // @[SpatialBlocks.scala 37:22:@48528.4]
    .clock(x748_ctrchain_clock),
    .reset(x748_ctrchain_reset),
    .io_input_reset(x748_ctrchain_io_input_reset),
    .io_input_enable(x748_ctrchain_io_input_enable),
    .io_output_counts_0(x748_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x748_ctrchain_io_output_oobs_0),
    .io_output_done(x748_ctrchain_io_output_done)
  );
  x755_inr_Foreach_sm x755_inr_Foreach_sm ( // @[sm_x755_inr_Foreach.scala 33:18:@48581.4]
    .clock(x755_inr_Foreach_sm_clock),
    .reset(x755_inr_Foreach_sm_reset),
    .io_enable(x755_inr_Foreach_sm_io_enable),
    .io_done(x755_inr_Foreach_sm_io_done),
    .io_doneLatch(x755_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x755_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x755_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x755_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x755_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x755_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x755_inr_Foreach_sm_io_backpressure),
    .io_break(x755_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@48609.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@48649.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@48657.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x755_inr_Foreach_kernelx755_inr_Foreach_concrete1 x755_inr_Foreach_kernelx755_inr_Foreach_concrete1 ( // @[sm_x755_inr_Foreach.scala 78:24:@48692.4]
    .clock(x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_clock),
    .reset(x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_reset),
    .io_in_x482_outbuf_0_rPort_0_ofs_0(x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_io_in_x482_outbuf_0_rPort_0_ofs_0),
    .io_in_x482_outbuf_0_rPort_0_en_0(x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_io_in_x482_outbuf_0_rPort_0_en_0),
    .io_in_x482_outbuf_0_rPort_0_backpressure(x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_io_in_x482_outbuf_0_rPort_0_backpressure),
    .io_in_x482_outbuf_0_rPort_0_output_0(x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_io_in_x482_outbuf_0_rPort_0_output_0),
    .io_in_x740_valid(x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_io_in_x740_valid),
    .io_in_x740_bits_wdata_0(x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_io_in_x740_bits_wdata_0),
    .io_in_x740_bits_wstrb(x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_io_in_x740_bits_wstrb),
    .io_sigsIn_backpressure(x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_0(x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_rr(x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_io_rr)
  );
  x759_inr_UnitPipe_sm x759_inr_UnitPipe_sm ( // @[sm_x759_inr_UnitPipe.scala 32:18:@48812.4]
    .clock(x759_inr_UnitPipe_sm_clock),
    .reset(x759_inr_UnitPipe_sm_reset),
    .io_enable(x759_inr_UnitPipe_sm_io_enable),
    .io_done(x759_inr_UnitPipe_sm_io_done),
    .io_doneLatch(x759_inr_UnitPipe_sm_io_doneLatch),
    .io_ctrDone(x759_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x759_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x759_inr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x759_inr_UnitPipe_sm_io_parentAck)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@48869.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@48877.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  x759_inr_UnitPipe_kernelx759_inr_UnitPipe_concrete1 x759_inr_UnitPipe_kernelx759_inr_UnitPipe_concrete1 ( // @[sm_x759_inr_UnitPipe.scala 60:24:@48907.4]
    .io_in_x741_ready(x759_inr_UnitPipe_kernelx759_inr_UnitPipe_concrete1_io_in_x741_ready),
    .io_sigsIn_datapathEn(x759_inr_UnitPipe_kernelx759_inr_UnitPipe_concrete1_io_sigsIn_datapathEn)
  );
  assign _T_359 = x746_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@48393.4]
  assign _T_375 = RetimeWrapper_io_out; // @[package.scala 96:25:@48427.4 package.scala 96:25:@48428.4]
  assign _T_381 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@48435.4 package.scala 96:25:@48436.4]
  assign _T_384 = ~ _T_381; // @[SpatialBlocks.scala 138:93:@48438.4]
  assign _T_454 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@48614.4 package.scala 96:25:@48615.4]
  assign _T_468 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@48654.4 package.scala 96:25:@48655.4]
  assign _T_474 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@48662.4 package.scala 96:25:@48663.4]
  assign _T_477 = ~ _T_474; // @[SpatialBlocks.scala 138:93:@48665.4]
  assign _T_479 = x755_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@48674.4]
  assign _T_480 = ~ x755_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@48675.4]
  assign _T_547 = x759_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@48840.4]
  assign x759_inr_UnitPipe_sigsIn_forwardpressure = io_in_x741_valid | x759_inr_UnitPipe_sm_io_doneLatch; // @[sm_x760_outr_UnitPipe.scala 101:55:@48847.4]
  assign _T_563 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@48874.4 package.scala 96:25:@48875.4]
  assign _T_569 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@48882.4 package.scala 96:25:@48883.4]
  assign _T_572 = ~ _T_569; // @[SpatialBlocks.scala 138:93:@48885.4]
  assign x759_inr_UnitPipe_sigsIn_baseEn = _T_563 & _T_572; // @[SpatialBlocks.scala 138:90:@48886.4]
  assign io_in_x741_ready = x759_inr_UnitPipe_kernelx759_inr_UnitPipe_concrete1_io_in_x741_ready; // @[sm_x759_inr_UnitPipe.scala 46:23:@48943.4]
  assign io_in_x739_valid = x746_inr_UnitPipe_kernelx746_inr_UnitPipe_concrete1_io_in_x739_valid; // @[sm_x746_inr_UnitPipe.scala 49:23:@48498.4]
  assign io_in_x739_bits_addr = x746_inr_UnitPipe_kernelx746_inr_UnitPipe_concrete1_io_in_x739_bits_addr; // @[sm_x746_inr_UnitPipe.scala 49:23:@48497.4]
  assign io_in_x739_bits_size = x746_inr_UnitPipe_kernelx746_inr_UnitPipe_concrete1_io_in_x739_bits_size; // @[sm_x746_inr_UnitPipe.scala 49:23:@48496.4]
  assign io_in_x482_outbuf_0_rPort_0_ofs_0 = x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_io_in_x482_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@48743.4]
  assign io_in_x482_outbuf_0_rPort_0_en_0 = x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_io_in_x482_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@48742.4]
  assign io_in_x482_outbuf_0_rPort_0_backpressure = x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_io_in_x482_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@48741.4]
  assign io_in_x740_valid = x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_io_in_x740_valid; // @[sm_x755_inr_Foreach.scala 50:23:@48747.4]
  assign io_in_x740_bits_wdata_0 = x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_io_in_x740_bits_wdata_0; // @[sm_x755_inr_Foreach.scala 50:23:@48746.4]
  assign io_in_x740_bits_wstrb = x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_io_in_x740_bits_wstrb; // @[sm_x755_inr_Foreach.scala 50:23:@48745.4]
  assign io_sigsOut_smDoneIn_0 = x746_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@48445.4]
  assign io_sigsOut_smDoneIn_1 = x755_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 156:53:@48672.4]
  assign io_sigsOut_smDoneIn_2 = x759_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@48892.4]
  assign io_sigsOut_smCtrCopyDone_0 = x746_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@48459.4]
  assign io_sigsOut_smCtrCopyDone_1 = x755_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 168:125:@48691.4]
  assign io_sigsOut_smCtrCopyDone_2 = x759_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@48906.4]
  assign x746_inr_UnitPipe_sm_clock = clock; // @[:@48366.4]
  assign x746_inr_UnitPipe_sm_reset = reset; // @[:@48367.4]
  assign x746_inr_UnitPipe_sm_io_enable = _T_375 & _T_384; // @[SpatialBlocks.scala 140:18:@48442.4]
  assign x746_inr_UnitPipe_sm_io_ctrDone = x746_inr_UnitPipe_sm_io_ctrInc & _T_362; // @[sm_x760_outr_UnitPipe.scala 77:39:@48397.4]
  assign x746_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@48444.4]
  assign x746_inr_UnitPipe_sm_io_backpressure = io_in_x739_ready | x746_inr_UnitPipe_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@48416.4]
  assign RetimeWrapper_clock = clock; // @[:@48423.4]
  assign RetimeWrapper_reset = reset; // @[:@48424.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@48426.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@48425.4]
  assign RetimeWrapper_1_clock = clock; // @[:@48431.4]
  assign RetimeWrapper_1_reset = reset; // @[:@48432.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@48434.4]
  assign RetimeWrapper_1_io_in = x746_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@48433.4]
  assign x746_inr_UnitPipe_kernelx746_inr_UnitPipe_concrete1_io_in_x478_outdram_number = io_in_x478_outdram_number; // @[sm_x746_inr_UnitPipe.scala 50:31:@48500.4]
  assign x746_inr_UnitPipe_kernelx746_inr_UnitPipe_concrete1_io_sigsIn_backpressure = io_in_x739_ready | x746_inr_UnitPipe_sm_io_doneLatch; // @[sm_x746_inr_UnitPipe.scala 74:22:@48515.4]
  assign x746_inr_UnitPipe_kernelx746_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x746_inr_UnitPipe_sm_io_datapathEn; // @[sm_x746_inr_UnitPipe.scala 74:22:@48513.4]
  assign x746_inr_UnitPipe_kernelx746_inr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x746_inr_UnitPipe.scala 73:18:@48501.4]
  assign x748_ctrchain_clock = clock; // @[:@48529.4]
  assign x748_ctrchain_reset = reset; // @[:@48530.4]
  assign x748_ctrchain_io_input_reset = x755_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@48690.4]
  assign x748_ctrchain_io_input_enable = x755_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 132:75:@48642.4 SpatialBlocks.scala 159:42:@48689.4]
  assign x755_inr_Foreach_sm_clock = clock; // @[:@48582.4]
  assign x755_inr_Foreach_sm_reset = reset; // @[:@48583.4]
  assign x755_inr_Foreach_sm_io_enable = _T_468 & _T_477; // @[SpatialBlocks.scala 140:18:@48669.4]
  assign x755_inr_Foreach_sm_io_ctrDone = io_rr ? _T_454 : 1'h0; // @[sm_x760_outr_UnitPipe.scala 90:38:@48617.4]
  assign x755_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@48671.4]
  assign x755_inr_Foreach_sm_io_backpressure = io_in_x740_ready | x755_inr_Foreach_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@48643.4]
  assign x755_inr_Foreach_sm_io_break = 1'h0; // @[sm_x760_outr_UnitPipe.scala 94:36:@48623.4]
  assign RetimeWrapper_2_clock = clock; // @[:@48610.4]
  assign RetimeWrapper_2_reset = reset; // @[:@48611.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@48613.4]
  assign RetimeWrapper_2_io_in = x748_ctrchain_io_output_done; // @[package.scala 94:16:@48612.4]
  assign RetimeWrapper_3_clock = clock; // @[:@48650.4]
  assign RetimeWrapper_3_reset = reset; // @[:@48651.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@48653.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@48652.4]
  assign RetimeWrapper_4_clock = clock; // @[:@48658.4]
  assign RetimeWrapper_4_reset = reset; // @[:@48659.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@48661.4]
  assign RetimeWrapper_4_io_in = x755_inr_Foreach_sm_io_done; // @[package.scala 94:16:@48660.4]
  assign x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_clock = clock; // @[:@48693.4]
  assign x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_reset = reset; // @[:@48694.4]
  assign x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_io_in_x482_outbuf_0_rPort_0_output_0 = io_in_x482_outbuf_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@48740.4]
  assign x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_io_sigsIn_backpressure = io_in_x740_ready | x755_inr_Foreach_sm_io_doneLatch; // @[sm_x755_inr_Foreach.scala 83:22:@48763.4]
  assign x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_479 & _T_480; // @[sm_x755_inr_Foreach.scala 83:22:@48761.4]
  assign x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_io_sigsIn_break = x755_inr_Foreach_sm_io_break; // @[sm_x755_inr_Foreach.scala 83:22:@48759.4]
  assign x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{9{x748_ctrchain_io_output_counts_0[22]}},x748_ctrchain_io_output_counts_0}; // @[sm_x755_inr_Foreach.scala 83:22:@48754.4]
  assign x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x748_ctrchain_io_output_oobs_0; // @[sm_x755_inr_Foreach.scala 83:22:@48753.4]
  assign x755_inr_Foreach_kernelx755_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x755_inr_Foreach.scala 82:18:@48749.4]
  assign x759_inr_UnitPipe_sm_clock = clock; // @[:@48813.4]
  assign x759_inr_UnitPipe_sm_reset = reset; // @[:@48814.4]
  assign x759_inr_UnitPipe_sm_io_enable = x759_inr_UnitPipe_sigsIn_baseEn & x759_inr_UnitPipe_sigsIn_forwardpressure; // @[SpatialBlocks.scala 140:18:@48889.4]
  assign x759_inr_UnitPipe_sm_io_ctrDone = x759_inr_UnitPipe_sm_io_ctrInc & _T_550; // @[sm_x760_outr_UnitPipe.scala 99:39:@48844.4]
  assign x759_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_2; // @[SpatialBlocks.scala 142:21:@48891.4]
  assign RetimeWrapper_5_clock = clock; // @[:@48870.4]
  assign RetimeWrapper_5_reset = reset; // @[:@48871.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@48873.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_smEnableOuts_2; // @[package.scala 94:16:@48872.4]
  assign RetimeWrapper_6_clock = clock; // @[:@48878.4]
  assign RetimeWrapper_6_reset = reset; // @[:@48879.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@48881.4]
  assign RetimeWrapper_6_io_in = x759_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@48880.4]
  assign x759_inr_UnitPipe_kernelx759_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x759_inr_UnitPipe_sm_io_datapathEn; // @[sm_x759_inr_UnitPipe.scala 65:22:@48956.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_362 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_550 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_362 <= 1'h0;
    end else begin
      _T_362 <= _T_359;
    end
    if (reset) begin
      _T_550 <= 1'h0;
    end else begin
      _T_550 <= _T_547;
    end
  end
endmodule
module x819_kernelx819_concrete1( // @[:@48972.2]
  input          clock, // @[:@48973.4]
  input          reset, // @[:@48974.4]
  output         io_in_x481_TVALID, // @[:@48975.4]
  input          io_in_x481_TREADY, // @[:@48975.4]
  output [255:0] io_in_x481_TDATA, // @[:@48975.4]
  output         io_in_x741_ready, // @[:@48975.4]
  input          io_in_x741_valid, // @[:@48975.4]
  input          io_in_x480_TVALID, // @[:@48975.4]
  output         io_in_x480_TREADY, // @[:@48975.4]
  input  [255:0] io_in_x480_TDATA, // @[:@48975.4]
  input  [7:0]   io_in_x480_TID, // @[:@48975.4]
  input  [7:0]   io_in_x480_TDEST, // @[:@48975.4]
  input          io_in_x739_ready, // @[:@48975.4]
  output         io_in_x739_valid, // @[:@48975.4]
  output [63:0]  io_in_x739_bits_addr, // @[:@48975.4]
  output [31:0]  io_in_x739_bits_size, // @[:@48975.4]
  output [20:0]  io_in_x482_outbuf_0_rPort_0_ofs_0, // @[:@48975.4]
  output         io_in_x482_outbuf_0_rPort_0_en_0, // @[:@48975.4]
  output         io_in_x482_outbuf_0_rPort_0_backpressure, // @[:@48975.4]
  input  [7:0]   io_in_x482_outbuf_0_rPort_0_output_0, // @[:@48975.4]
  input  [63:0]  io_in_x478_outdram_number, // @[:@48975.4]
  input          io_in_x740_ready, // @[:@48975.4]
  output         io_in_x740_valid, // @[:@48975.4]
  output [7:0]   io_in_x740_bits_wdata_0, // @[:@48975.4]
  output         io_in_x740_bits_wstrb, // @[:@48975.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@48975.4]
  input          io_sigsIn_smEnableOuts_1, // @[:@48975.4]
  input          io_sigsIn_smChildAcks_0, // @[:@48975.4]
  input          io_sigsIn_smChildAcks_1, // @[:@48975.4]
  output         io_sigsOut_smDoneIn_0, // @[:@48975.4]
  output         io_sigsOut_smDoneIn_1, // @[:@48975.4]
  input          io_rr // @[:@48975.4]
);
  wire  x738_outr_UnitPipe_sm_clock; // @[sm_x738_outr_UnitPipe.scala 32:18:@49048.4]
  wire  x738_outr_UnitPipe_sm_reset; // @[sm_x738_outr_UnitPipe.scala 32:18:@49048.4]
  wire  x738_outr_UnitPipe_sm_io_enable; // @[sm_x738_outr_UnitPipe.scala 32:18:@49048.4]
  wire  x738_outr_UnitPipe_sm_io_done; // @[sm_x738_outr_UnitPipe.scala 32:18:@49048.4]
  wire  x738_outr_UnitPipe_sm_io_parentAck; // @[sm_x738_outr_UnitPipe.scala 32:18:@49048.4]
  wire  x738_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x738_outr_UnitPipe.scala 32:18:@49048.4]
  wire  x738_outr_UnitPipe_sm_io_doneIn_1; // @[sm_x738_outr_UnitPipe.scala 32:18:@49048.4]
  wire  x738_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x738_outr_UnitPipe.scala 32:18:@49048.4]
  wire  x738_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x738_outr_UnitPipe.scala 32:18:@49048.4]
  wire  x738_outr_UnitPipe_sm_io_childAck_0; // @[sm_x738_outr_UnitPipe.scala 32:18:@49048.4]
  wire  x738_outr_UnitPipe_sm_io_childAck_1; // @[sm_x738_outr_UnitPipe.scala 32:18:@49048.4]
  wire  x738_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x738_outr_UnitPipe.scala 32:18:@49048.4]
  wire  x738_outr_UnitPipe_sm_io_ctrCopyDone_1; // @[sm_x738_outr_UnitPipe.scala 32:18:@49048.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@49110.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@49110.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@49110.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@49110.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@49110.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@49118.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@49118.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@49118.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@49118.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@49118.4]
  wire  x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_clock; // @[sm_x738_outr_UnitPipe.scala 87:24:@49149.4]
  wire  x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_reset; // @[sm_x738_outr_UnitPipe.scala 87:24:@49149.4]
  wire  x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_in_x481_TVALID; // @[sm_x738_outr_UnitPipe.scala 87:24:@49149.4]
  wire  x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_in_x481_TREADY; // @[sm_x738_outr_UnitPipe.scala 87:24:@49149.4]
  wire [255:0] x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_in_x481_TDATA; // @[sm_x738_outr_UnitPipe.scala 87:24:@49149.4]
  wire  x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_in_x480_TVALID; // @[sm_x738_outr_UnitPipe.scala 87:24:@49149.4]
  wire  x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_in_x480_TREADY; // @[sm_x738_outr_UnitPipe.scala 87:24:@49149.4]
  wire [255:0] x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_in_x480_TDATA; // @[sm_x738_outr_UnitPipe.scala 87:24:@49149.4]
  wire [7:0] x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_in_x480_TID; // @[sm_x738_outr_UnitPipe.scala 87:24:@49149.4]
  wire [7:0] x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_in_x480_TDEST; // @[sm_x738_outr_UnitPipe.scala 87:24:@49149.4]
  wire  x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x738_outr_UnitPipe.scala 87:24:@49149.4]
  wire  x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x738_outr_UnitPipe.scala 87:24:@49149.4]
  wire  x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x738_outr_UnitPipe.scala 87:24:@49149.4]
  wire  x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x738_outr_UnitPipe.scala 87:24:@49149.4]
  wire  x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x738_outr_UnitPipe.scala 87:24:@49149.4]
  wire  x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x738_outr_UnitPipe.scala 87:24:@49149.4]
  wire  x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x738_outr_UnitPipe.scala 87:24:@49149.4]
  wire  x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[sm_x738_outr_UnitPipe.scala 87:24:@49149.4]
  wire  x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_rr; // @[sm_x738_outr_UnitPipe.scala 87:24:@49149.4]
  wire  x760_outr_UnitPipe_sm_clock; // @[sm_x760_outr_UnitPipe.scala 36:18:@49327.4]
  wire  x760_outr_UnitPipe_sm_reset; // @[sm_x760_outr_UnitPipe.scala 36:18:@49327.4]
  wire  x760_outr_UnitPipe_sm_io_enable; // @[sm_x760_outr_UnitPipe.scala 36:18:@49327.4]
  wire  x760_outr_UnitPipe_sm_io_done; // @[sm_x760_outr_UnitPipe.scala 36:18:@49327.4]
  wire  x760_outr_UnitPipe_sm_io_parentAck; // @[sm_x760_outr_UnitPipe.scala 36:18:@49327.4]
  wire  x760_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x760_outr_UnitPipe.scala 36:18:@49327.4]
  wire  x760_outr_UnitPipe_sm_io_doneIn_1; // @[sm_x760_outr_UnitPipe.scala 36:18:@49327.4]
  wire  x760_outr_UnitPipe_sm_io_doneIn_2; // @[sm_x760_outr_UnitPipe.scala 36:18:@49327.4]
  wire  x760_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x760_outr_UnitPipe.scala 36:18:@49327.4]
  wire  x760_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x760_outr_UnitPipe.scala 36:18:@49327.4]
  wire  x760_outr_UnitPipe_sm_io_enableOut_2; // @[sm_x760_outr_UnitPipe.scala 36:18:@49327.4]
  wire  x760_outr_UnitPipe_sm_io_childAck_0; // @[sm_x760_outr_UnitPipe.scala 36:18:@49327.4]
  wire  x760_outr_UnitPipe_sm_io_childAck_1; // @[sm_x760_outr_UnitPipe.scala 36:18:@49327.4]
  wire  x760_outr_UnitPipe_sm_io_childAck_2; // @[sm_x760_outr_UnitPipe.scala 36:18:@49327.4]
  wire  x760_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x760_outr_UnitPipe.scala 36:18:@49327.4]
  wire  x760_outr_UnitPipe_sm_io_ctrCopyDone_1; // @[sm_x760_outr_UnitPipe.scala 36:18:@49327.4]
  wire  x760_outr_UnitPipe_sm_io_ctrCopyDone_2; // @[sm_x760_outr_UnitPipe.scala 36:18:@49327.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@49399.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@49399.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@49399.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@49399.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@49399.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@49407.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@49407.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@49407.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@49407.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@49407.4]
  wire  x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_clock; // @[sm_x760_outr_UnitPipe.scala 108:24:@49439.4]
  wire  x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_reset; // @[sm_x760_outr_UnitPipe.scala 108:24:@49439.4]
  wire  x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x741_ready; // @[sm_x760_outr_UnitPipe.scala 108:24:@49439.4]
  wire  x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x741_valid; // @[sm_x760_outr_UnitPipe.scala 108:24:@49439.4]
  wire  x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x739_ready; // @[sm_x760_outr_UnitPipe.scala 108:24:@49439.4]
  wire  x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x739_valid; // @[sm_x760_outr_UnitPipe.scala 108:24:@49439.4]
  wire [63:0] x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x739_bits_addr; // @[sm_x760_outr_UnitPipe.scala 108:24:@49439.4]
  wire [31:0] x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x739_bits_size; // @[sm_x760_outr_UnitPipe.scala 108:24:@49439.4]
  wire [20:0] x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x482_outbuf_0_rPort_0_ofs_0; // @[sm_x760_outr_UnitPipe.scala 108:24:@49439.4]
  wire  x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x482_outbuf_0_rPort_0_en_0; // @[sm_x760_outr_UnitPipe.scala 108:24:@49439.4]
  wire  x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x482_outbuf_0_rPort_0_backpressure; // @[sm_x760_outr_UnitPipe.scala 108:24:@49439.4]
  wire [7:0] x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x482_outbuf_0_rPort_0_output_0; // @[sm_x760_outr_UnitPipe.scala 108:24:@49439.4]
  wire [63:0] x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x478_outdram_number; // @[sm_x760_outr_UnitPipe.scala 108:24:@49439.4]
  wire  x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x740_ready; // @[sm_x760_outr_UnitPipe.scala 108:24:@49439.4]
  wire  x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x740_valid; // @[sm_x760_outr_UnitPipe.scala 108:24:@49439.4]
  wire [7:0] x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x740_bits_wdata_0; // @[sm_x760_outr_UnitPipe.scala 108:24:@49439.4]
  wire  x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x740_bits_wstrb; // @[sm_x760_outr_UnitPipe.scala 108:24:@49439.4]
  wire  x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x760_outr_UnitPipe.scala 108:24:@49439.4]
  wire  x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x760_outr_UnitPipe.scala 108:24:@49439.4]
  wire  x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2; // @[sm_x760_outr_UnitPipe.scala 108:24:@49439.4]
  wire  x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x760_outr_UnitPipe.scala 108:24:@49439.4]
  wire  x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x760_outr_UnitPipe.scala 108:24:@49439.4]
  wire  x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2; // @[sm_x760_outr_UnitPipe.scala 108:24:@49439.4]
  wire  x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x760_outr_UnitPipe.scala 108:24:@49439.4]
  wire  x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x760_outr_UnitPipe.scala 108:24:@49439.4]
  wire  x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2; // @[sm_x760_outr_UnitPipe.scala 108:24:@49439.4]
  wire  x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x760_outr_UnitPipe.scala 108:24:@49439.4]
  wire  x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[sm_x760_outr_UnitPipe.scala 108:24:@49439.4]
  wire  x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2; // @[sm_x760_outr_UnitPipe.scala 108:24:@49439.4]
  wire  x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_rr; // @[sm_x760_outr_UnitPipe.scala 108:24:@49439.4]
  wire  _T_408; // @[package.scala 96:25:@49115.4 package.scala 96:25:@49116.4]
  wire  _T_414; // @[package.scala 96:25:@49123.4 package.scala 96:25:@49124.4]
  wire  _T_417; // @[SpatialBlocks.scala 138:93:@49126.4]
  wire  _T_508; // @[package.scala 96:25:@49404.4 package.scala 96:25:@49405.4]
  wire  _T_514; // @[package.scala 96:25:@49412.4 package.scala 96:25:@49413.4]
  wire  _T_517; // @[SpatialBlocks.scala 138:93:@49415.4]
  x738_outr_UnitPipe_sm x738_outr_UnitPipe_sm ( // @[sm_x738_outr_UnitPipe.scala 32:18:@49048.4]
    .clock(x738_outr_UnitPipe_sm_clock),
    .reset(x738_outr_UnitPipe_sm_reset),
    .io_enable(x738_outr_UnitPipe_sm_io_enable),
    .io_done(x738_outr_UnitPipe_sm_io_done),
    .io_parentAck(x738_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x738_outr_UnitPipe_sm_io_doneIn_0),
    .io_doneIn_1(x738_outr_UnitPipe_sm_io_doneIn_1),
    .io_enableOut_0(x738_outr_UnitPipe_sm_io_enableOut_0),
    .io_enableOut_1(x738_outr_UnitPipe_sm_io_enableOut_1),
    .io_childAck_0(x738_outr_UnitPipe_sm_io_childAck_0),
    .io_childAck_1(x738_outr_UnitPipe_sm_io_childAck_1),
    .io_ctrCopyDone_0(x738_outr_UnitPipe_sm_io_ctrCopyDone_0),
    .io_ctrCopyDone_1(x738_outr_UnitPipe_sm_io_ctrCopyDone_1)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@49110.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@49118.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1 x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1 ( // @[sm_x738_outr_UnitPipe.scala 87:24:@49149.4]
    .clock(x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_clock),
    .reset(x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_reset),
    .io_in_x481_TVALID(x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_in_x481_TVALID),
    .io_in_x481_TREADY(x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_in_x481_TREADY),
    .io_in_x481_TDATA(x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_in_x481_TDATA),
    .io_in_x480_TVALID(x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_in_x480_TVALID),
    .io_in_x480_TREADY(x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_in_x480_TREADY),
    .io_in_x480_TDATA(x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_in_x480_TDATA),
    .io_in_x480_TID(x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_in_x480_TID),
    .io_in_x480_TDEST(x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_in_x480_TDEST),
    .io_sigsIn_smEnableOuts_0(x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsOut_smDoneIn_0(x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smCtrCopyDone_0(x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_sigsOut_smCtrCopyDone_1(x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1),
    .io_rr(x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_rr)
  );
  x760_outr_UnitPipe_sm x760_outr_UnitPipe_sm ( // @[sm_x760_outr_UnitPipe.scala 36:18:@49327.4]
    .clock(x760_outr_UnitPipe_sm_clock),
    .reset(x760_outr_UnitPipe_sm_reset),
    .io_enable(x760_outr_UnitPipe_sm_io_enable),
    .io_done(x760_outr_UnitPipe_sm_io_done),
    .io_parentAck(x760_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x760_outr_UnitPipe_sm_io_doneIn_0),
    .io_doneIn_1(x760_outr_UnitPipe_sm_io_doneIn_1),
    .io_doneIn_2(x760_outr_UnitPipe_sm_io_doneIn_2),
    .io_enableOut_0(x760_outr_UnitPipe_sm_io_enableOut_0),
    .io_enableOut_1(x760_outr_UnitPipe_sm_io_enableOut_1),
    .io_enableOut_2(x760_outr_UnitPipe_sm_io_enableOut_2),
    .io_childAck_0(x760_outr_UnitPipe_sm_io_childAck_0),
    .io_childAck_1(x760_outr_UnitPipe_sm_io_childAck_1),
    .io_childAck_2(x760_outr_UnitPipe_sm_io_childAck_2),
    .io_ctrCopyDone_0(x760_outr_UnitPipe_sm_io_ctrCopyDone_0),
    .io_ctrCopyDone_1(x760_outr_UnitPipe_sm_io_ctrCopyDone_1),
    .io_ctrCopyDone_2(x760_outr_UnitPipe_sm_io_ctrCopyDone_2)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@49399.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@49407.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1 x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1 ( // @[sm_x760_outr_UnitPipe.scala 108:24:@49439.4]
    .clock(x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_clock),
    .reset(x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_reset),
    .io_in_x741_ready(x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x741_ready),
    .io_in_x741_valid(x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x741_valid),
    .io_in_x739_ready(x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x739_ready),
    .io_in_x739_valid(x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x739_valid),
    .io_in_x739_bits_addr(x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x739_bits_addr),
    .io_in_x739_bits_size(x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x739_bits_size),
    .io_in_x482_outbuf_0_rPort_0_ofs_0(x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x482_outbuf_0_rPort_0_ofs_0),
    .io_in_x482_outbuf_0_rPort_0_en_0(x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x482_outbuf_0_rPort_0_en_0),
    .io_in_x482_outbuf_0_rPort_0_backpressure(x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x482_outbuf_0_rPort_0_backpressure),
    .io_in_x482_outbuf_0_rPort_0_output_0(x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x482_outbuf_0_rPort_0_output_0),
    .io_in_x478_outdram_number(x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x478_outdram_number),
    .io_in_x740_ready(x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x740_ready),
    .io_in_x740_valid(x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x740_valid),
    .io_in_x740_bits_wdata_0(x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x740_bits_wdata_0),
    .io_in_x740_bits_wstrb(x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x740_bits_wstrb),
    .io_sigsIn_smEnableOuts_0(x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smEnableOuts_2(x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2),
    .io_sigsIn_smChildAcks_0(x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsIn_smChildAcks_2(x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2),
    .io_sigsOut_smDoneIn_0(x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smDoneIn_2(x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2),
    .io_sigsOut_smCtrCopyDone_0(x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_sigsOut_smCtrCopyDone_1(x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1),
    .io_sigsOut_smCtrCopyDone_2(x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2),
    .io_rr(x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_408 = RetimeWrapper_io_out; // @[package.scala 96:25:@49115.4 package.scala 96:25:@49116.4]
  assign _T_414 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@49123.4 package.scala 96:25:@49124.4]
  assign _T_417 = ~ _T_414; // @[SpatialBlocks.scala 138:93:@49126.4]
  assign _T_508 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@49404.4 package.scala 96:25:@49405.4]
  assign _T_514 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@49412.4 package.scala 96:25:@49413.4]
  assign _T_517 = ~ _T_514; // @[SpatialBlocks.scala 138:93:@49415.4]
  assign io_in_x481_TVALID = x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_in_x481_TVALID; // @[sm_x738_outr_UnitPipe.scala 48:23:@49218.4]
  assign io_in_x481_TDATA = x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_in_x481_TDATA; // @[sm_x738_outr_UnitPipe.scala 48:23:@49216.4]
  assign io_in_x741_ready = x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x741_ready; // @[sm_x760_outr_UnitPipe.scala 58:23:@49521.4]
  assign io_in_x480_TREADY = x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_in_x480_TREADY; // @[sm_x738_outr_UnitPipe.scala 49:23:@49226.4]
  assign io_in_x739_valid = x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x739_valid; // @[sm_x760_outr_UnitPipe.scala 59:23:@49524.4]
  assign io_in_x739_bits_addr = x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x739_bits_addr; // @[sm_x760_outr_UnitPipe.scala 59:23:@49523.4]
  assign io_in_x739_bits_size = x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x739_bits_size; // @[sm_x760_outr_UnitPipe.scala 59:23:@49522.4]
  assign io_in_x482_outbuf_0_rPort_0_ofs_0 = x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x482_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@49529.4]
  assign io_in_x482_outbuf_0_rPort_0_en_0 = x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x482_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@49528.4]
  assign io_in_x482_outbuf_0_rPort_0_backpressure = x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x482_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@49527.4]
  assign io_in_x740_valid = x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x740_valid; // @[sm_x760_outr_UnitPipe.scala 62:23:@49534.4]
  assign io_in_x740_bits_wdata_0 = x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x740_bits_wdata_0; // @[sm_x760_outr_UnitPipe.scala 62:23:@49533.4]
  assign io_in_x740_bits_wstrb = x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x740_bits_wstrb; // @[sm_x760_outr_UnitPipe.scala 62:23:@49532.4]
  assign io_sigsOut_smDoneIn_0 = x738_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@49133.4]
  assign io_sigsOut_smDoneIn_1 = x760_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@49422.4]
  assign x738_outr_UnitPipe_sm_clock = clock; // @[:@49049.4]
  assign x738_outr_UnitPipe_sm_reset = reset; // @[:@49050.4]
  assign x738_outr_UnitPipe_sm_io_enable = _T_408 & _T_417; // @[SpatialBlocks.scala 140:18:@49130.4]
  assign x738_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@49132.4]
  assign x738_outr_UnitPipe_sm_io_doneIn_0 = x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@49100.4]
  assign x738_outr_UnitPipe_sm_io_doneIn_1 = x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@49101.4]
  assign x738_outr_UnitPipe_sm_io_ctrCopyDone_0 = x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 161:90:@49147.4]
  assign x738_outr_UnitPipe_sm_io_ctrCopyDone_1 = x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[SpatialBlocks.scala 161:90:@49148.4]
  assign RetimeWrapper_clock = clock; // @[:@49111.4]
  assign RetimeWrapper_reset = reset; // @[:@49112.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@49114.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@49113.4]
  assign RetimeWrapper_1_clock = clock; // @[:@49119.4]
  assign RetimeWrapper_1_reset = reset; // @[:@49120.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@49122.4]
  assign RetimeWrapper_1_io_in = x738_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@49121.4]
  assign x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_clock = clock; // @[:@49150.4]
  assign x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_reset = reset; // @[:@49151.4]
  assign x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_in_x481_TREADY = io_in_x481_TREADY; // @[sm_x738_outr_UnitPipe.scala 48:23:@49217.4]
  assign x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_in_x480_TVALID = io_in_x480_TVALID; // @[sm_x738_outr_UnitPipe.scala 49:23:@49227.4]
  assign x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_in_x480_TDATA = io_in_x480_TDATA; // @[sm_x738_outr_UnitPipe.scala 49:23:@49225.4]
  assign x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_in_x480_TID = io_in_x480_TID; // @[sm_x738_outr_UnitPipe.scala 49:23:@49221.4]
  assign x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_in_x480_TDEST = io_in_x480_TDEST; // @[sm_x738_outr_UnitPipe.scala 49:23:@49220.4]
  assign x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x738_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x738_outr_UnitPipe.scala 92:22:@49243.4]
  assign x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1 = x738_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x738_outr_UnitPipe.scala 92:22:@49244.4]
  assign x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x738_outr_UnitPipe_sm_io_childAck_0; // @[sm_x738_outr_UnitPipe.scala 92:22:@49239.4]
  assign x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1 = x738_outr_UnitPipe_sm_io_childAck_1; // @[sm_x738_outr_UnitPipe.scala 92:22:@49240.4]
  assign x738_outr_UnitPipe_kernelx738_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x738_outr_UnitPipe.scala 91:18:@49228.4]
  assign x760_outr_UnitPipe_sm_clock = clock; // @[:@49328.4]
  assign x760_outr_UnitPipe_sm_reset = reset; // @[:@49329.4]
  assign x760_outr_UnitPipe_sm_io_enable = _T_508 & _T_517; // @[SpatialBlocks.scala 140:18:@49419.4]
  assign x760_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@49421.4]
  assign x760_outr_UnitPipe_sm_io_doneIn_0 = x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@49387.4]
  assign x760_outr_UnitPipe_sm_io_doneIn_1 = x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@49388.4]
  assign x760_outr_UnitPipe_sm_io_doneIn_2 = x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2; // @[SpatialBlocks.scala 130:67:@49389.4]
  assign x760_outr_UnitPipe_sm_io_ctrCopyDone_0 = x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 161:90:@49436.4]
  assign x760_outr_UnitPipe_sm_io_ctrCopyDone_1 = x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[SpatialBlocks.scala 161:90:@49437.4]
  assign x760_outr_UnitPipe_sm_io_ctrCopyDone_2 = x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2; // @[SpatialBlocks.scala 161:90:@49438.4]
  assign RetimeWrapper_2_clock = clock; // @[:@49400.4]
  assign RetimeWrapper_2_reset = reset; // @[:@49401.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@49403.4]
  assign RetimeWrapper_2_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@49402.4]
  assign RetimeWrapper_3_clock = clock; // @[:@49408.4]
  assign RetimeWrapper_3_reset = reset; // @[:@49409.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@49411.4]
  assign RetimeWrapper_3_io_in = x760_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@49410.4]
  assign x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_clock = clock; // @[:@49440.4]
  assign x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_reset = reset; // @[:@49441.4]
  assign x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x741_valid = io_in_x741_valid; // @[sm_x760_outr_UnitPipe.scala 58:23:@49520.4]
  assign x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x739_ready = io_in_x739_ready; // @[sm_x760_outr_UnitPipe.scala 59:23:@49525.4]
  assign x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x482_outbuf_0_rPort_0_output_0 = io_in_x482_outbuf_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@49526.4]
  assign x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x478_outdram_number = io_in_x478_outdram_number; // @[sm_x760_outr_UnitPipe.scala 61:31:@49531.4]
  assign x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_in_x740_ready = io_in_x740_ready; // @[sm_x760_outr_UnitPipe.scala 62:23:@49535.4]
  assign x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x760_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x760_outr_UnitPipe.scala 113:22:@49558.4]
  assign x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1 = x760_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x760_outr_UnitPipe.scala 113:22:@49559.4]
  assign x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2 = x760_outr_UnitPipe_sm_io_enableOut_2; // @[sm_x760_outr_UnitPipe.scala 113:22:@49560.4]
  assign x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x760_outr_UnitPipe_sm_io_childAck_0; // @[sm_x760_outr_UnitPipe.scala 113:22:@49552.4]
  assign x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1 = x760_outr_UnitPipe_sm_io_childAck_1; // @[sm_x760_outr_UnitPipe.scala 113:22:@49553.4]
  assign x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2 = x760_outr_UnitPipe_sm_io_childAck_2; // @[sm_x760_outr_UnitPipe.scala 113:22:@49554.4]
  assign x760_outr_UnitPipe_kernelx760_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x760_outr_UnitPipe.scala 112:18:@49536.4]
endmodule
module RootController_kernelRootController_concrete1( // @[:@49588.2]
  input          clock, // @[:@49589.4]
  input          reset, // @[:@49590.4]
  output         io_in_x481_TVALID, // @[:@49591.4]
  input          io_in_x481_TREADY, // @[:@49591.4]
  output [255:0] io_in_x481_TDATA, // @[:@49591.4]
  output         io_in_x741_ready, // @[:@49591.4]
  input          io_in_x741_valid, // @[:@49591.4]
  input          io_in_x480_TVALID, // @[:@49591.4]
  output         io_in_x480_TREADY, // @[:@49591.4]
  input  [255:0] io_in_x480_TDATA, // @[:@49591.4]
  input  [7:0]   io_in_x480_TID, // @[:@49591.4]
  input  [7:0]   io_in_x480_TDEST, // @[:@49591.4]
  input          io_in_x739_ready, // @[:@49591.4]
  output         io_in_x739_valid, // @[:@49591.4]
  output [63:0]  io_in_x739_bits_addr, // @[:@49591.4]
  output [31:0]  io_in_x739_bits_size, // @[:@49591.4]
  input  [63:0]  io_in_x478_outdram_number, // @[:@49591.4]
  input          io_in_x740_ready, // @[:@49591.4]
  output         io_in_x740_valid, // @[:@49591.4]
  output [7:0]   io_in_x740_bits_wdata_0, // @[:@49591.4]
  output         io_in_x740_bits_wstrb, // @[:@49591.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@49591.4]
  input          io_sigsIn_smChildAcks_0, // @[:@49591.4]
  output         io_sigsOut_smDoneIn_0, // @[:@49591.4]
  input          io_rr // @[:@49591.4]
);
  wire  x482_outbuf_0_clock; // @[m_x482_outbuf_0.scala 27:17:@49601.4]
  wire  x482_outbuf_0_reset; // @[m_x482_outbuf_0.scala 27:17:@49601.4]
  wire [20:0] x482_outbuf_0_io_rPort_0_ofs_0; // @[m_x482_outbuf_0.scala 27:17:@49601.4]
  wire  x482_outbuf_0_io_rPort_0_en_0; // @[m_x482_outbuf_0.scala 27:17:@49601.4]
  wire  x482_outbuf_0_io_rPort_0_backpressure; // @[m_x482_outbuf_0.scala 27:17:@49601.4]
  wire [7:0] x482_outbuf_0_io_rPort_0_output_0; // @[m_x482_outbuf_0.scala 27:17:@49601.4]
  wire  x819_sm_clock; // @[sm_x819.scala 37:18:@49659.4]
  wire  x819_sm_reset; // @[sm_x819.scala 37:18:@49659.4]
  wire  x819_sm_io_enable; // @[sm_x819.scala 37:18:@49659.4]
  wire  x819_sm_io_done; // @[sm_x819.scala 37:18:@49659.4]
  wire  x819_sm_io_ctrDone; // @[sm_x819.scala 37:18:@49659.4]
  wire  x819_sm_io_ctrInc; // @[sm_x819.scala 37:18:@49659.4]
  wire  x819_sm_io_parentAck; // @[sm_x819.scala 37:18:@49659.4]
  wire  x819_sm_io_doneIn_0; // @[sm_x819.scala 37:18:@49659.4]
  wire  x819_sm_io_doneIn_1; // @[sm_x819.scala 37:18:@49659.4]
  wire  x819_sm_io_enableOut_0; // @[sm_x819.scala 37:18:@49659.4]
  wire  x819_sm_io_enableOut_1; // @[sm_x819.scala 37:18:@49659.4]
  wire  x819_sm_io_childAck_0; // @[sm_x819.scala 37:18:@49659.4]
  wire  x819_sm_io_childAck_1; // @[sm_x819.scala 37:18:@49659.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@49726.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@49726.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@49726.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@49726.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@49726.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@49734.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@49734.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@49734.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@49734.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@49734.4]
  wire  x819_kernelx819_concrete1_clock; // @[sm_x819.scala 102:24:@49763.4]
  wire  x819_kernelx819_concrete1_reset; // @[sm_x819.scala 102:24:@49763.4]
  wire  x819_kernelx819_concrete1_io_in_x481_TVALID; // @[sm_x819.scala 102:24:@49763.4]
  wire  x819_kernelx819_concrete1_io_in_x481_TREADY; // @[sm_x819.scala 102:24:@49763.4]
  wire [255:0] x819_kernelx819_concrete1_io_in_x481_TDATA; // @[sm_x819.scala 102:24:@49763.4]
  wire  x819_kernelx819_concrete1_io_in_x741_ready; // @[sm_x819.scala 102:24:@49763.4]
  wire  x819_kernelx819_concrete1_io_in_x741_valid; // @[sm_x819.scala 102:24:@49763.4]
  wire  x819_kernelx819_concrete1_io_in_x480_TVALID; // @[sm_x819.scala 102:24:@49763.4]
  wire  x819_kernelx819_concrete1_io_in_x480_TREADY; // @[sm_x819.scala 102:24:@49763.4]
  wire [255:0] x819_kernelx819_concrete1_io_in_x480_TDATA; // @[sm_x819.scala 102:24:@49763.4]
  wire [7:0] x819_kernelx819_concrete1_io_in_x480_TID; // @[sm_x819.scala 102:24:@49763.4]
  wire [7:0] x819_kernelx819_concrete1_io_in_x480_TDEST; // @[sm_x819.scala 102:24:@49763.4]
  wire  x819_kernelx819_concrete1_io_in_x739_ready; // @[sm_x819.scala 102:24:@49763.4]
  wire  x819_kernelx819_concrete1_io_in_x739_valid; // @[sm_x819.scala 102:24:@49763.4]
  wire [63:0] x819_kernelx819_concrete1_io_in_x739_bits_addr; // @[sm_x819.scala 102:24:@49763.4]
  wire [31:0] x819_kernelx819_concrete1_io_in_x739_bits_size; // @[sm_x819.scala 102:24:@49763.4]
  wire [20:0] x819_kernelx819_concrete1_io_in_x482_outbuf_0_rPort_0_ofs_0; // @[sm_x819.scala 102:24:@49763.4]
  wire  x819_kernelx819_concrete1_io_in_x482_outbuf_0_rPort_0_en_0; // @[sm_x819.scala 102:24:@49763.4]
  wire  x819_kernelx819_concrete1_io_in_x482_outbuf_0_rPort_0_backpressure; // @[sm_x819.scala 102:24:@49763.4]
  wire [7:0] x819_kernelx819_concrete1_io_in_x482_outbuf_0_rPort_0_output_0; // @[sm_x819.scala 102:24:@49763.4]
  wire [63:0] x819_kernelx819_concrete1_io_in_x478_outdram_number; // @[sm_x819.scala 102:24:@49763.4]
  wire  x819_kernelx819_concrete1_io_in_x740_ready; // @[sm_x819.scala 102:24:@49763.4]
  wire  x819_kernelx819_concrete1_io_in_x740_valid; // @[sm_x819.scala 102:24:@49763.4]
  wire [7:0] x819_kernelx819_concrete1_io_in_x740_bits_wdata_0; // @[sm_x819.scala 102:24:@49763.4]
  wire  x819_kernelx819_concrete1_io_in_x740_bits_wstrb; // @[sm_x819.scala 102:24:@49763.4]
  wire  x819_kernelx819_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x819.scala 102:24:@49763.4]
  wire  x819_kernelx819_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x819.scala 102:24:@49763.4]
  wire  x819_kernelx819_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x819.scala 102:24:@49763.4]
  wire  x819_kernelx819_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x819.scala 102:24:@49763.4]
  wire  x819_kernelx819_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x819.scala 102:24:@49763.4]
  wire  x819_kernelx819_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x819.scala 102:24:@49763.4]
  wire  x819_kernelx819_concrete1_io_rr; // @[sm_x819.scala 102:24:@49763.4]
  wire  _T_266; // @[package.scala 100:49:@49692.4]
  reg  _T_269; // @[package.scala 48:56:@49693.4]
  reg [31:0] _RAND_0;
  wire  _T_283; // @[package.scala 96:25:@49731.4 package.scala 96:25:@49732.4]
  wire  _T_289; // @[package.scala 96:25:@49739.4 package.scala 96:25:@49740.4]
  wire  _T_292; // @[SpatialBlocks.scala 138:93:@49742.4]
  x482_outbuf_0 x482_outbuf_0 ( // @[m_x482_outbuf_0.scala 27:17:@49601.4]
    .clock(x482_outbuf_0_clock),
    .reset(x482_outbuf_0_reset),
    .io_rPort_0_ofs_0(x482_outbuf_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x482_outbuf_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x482_outbuf_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x482_outbuf_0_io_rPort_0_output_0)
  );
  x819_sm x819_sm ( // @[sm_x819.scala 37:18:@49659.4]
    .clock(x819_sm_clock),
    .reset(x819_sm_reset),
    .io_enable(x819_sm_io_enable),
    .io_done(x819_sm_io_done),
    .io_ctrDone(x819_sm_io_ctrDone),
    .io_ctrInc(x819_sm_io_ctrInc),
    .io_parentAck(x819_sm_io_parentAck),
    .io_doneIn_0(x819_sm_io_doneIn_0),
    .io_doneIn_1(x819_sm_io_doneIn_1),
    .io_enableOut_0(x819_sm_io_enableOut_0),
    .io_enableOut_1(x819_sm_io_enableOut_1),
    .io_childAck_0(x819_sm_io_childAck_0),
    .io_childAck_1(x819_sm_io_childAck_1)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@49726.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@49734.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x819_kernelx819_concrete1 x819_kernelx819_concrete1 ( // @[sm_x819.scala 102:24:@49763.4]
    .clock(x819_kernelx819_concrete1_clock),
    .reset(x819_kernelx819_concrete1_reset),
    .io_in_x481_TVALID(x819_kernelx819_concrete1_io_in_x481_TVALID),
    .io_in_x481_TREADY(x819_kernelx819_concrete1_io_in_x481_TREADY),
    .io_in_x481_TDATA(x819_kernelx819_concrete1_io_in_x481_TDATA),
    .io_in_x741_ready(x819_kernelx819_concrete1_io_in_x741_ready),
    .io_in_x741_valid(x819_kernelx819_concrete1_io_in_x741_valid),
    .io_in_x480_TVALID(x819_kernelx819_concrete1_io_in_x480_TVALID),
    .io_in_x480_TREADY(x819_kernelx819_concrete1_io_in_x480_TREADY),
    .io_in_x480_TDATA(x819_kernelx819_concrete1_io_in_x480_TDATA),
    .io_in_x480_TID(x819_kernelx819_concrete1_io_in_x480_TID),
    .io_in_x480_TDEST(x819_kernelx819_concrete1_io_in_x480_TDEST),
    .io_in_x739_ready(x819_kernelx819_concrete1_io_in_x739_ready),
    .io_in_x739_valid(x819_kernelx819_concrete1_io_in_x739_valid),
    .io_in_x739_bits_addr(x819_kernelx819_concrete1_io_in_x739_bits_addr),
    .io_in_x739_bits_size(x819_kernelx819_concrete1_io_in_x739_bits_size),
    .io_in_x482_outbuf_0_rPort_0_ofs_0(x819_kernelx819_concrete1_io_in_x482_outbuf_0_rPort_0_ofs_0),
    .io_in_x482_outbuf_0_rPort_0_en_0(x819_kernelx819_concrete1_io_in_x482_outbuf_0_rPort_0_en_0),
    .io_in_x482_outbuf_0_rPort_0_backpressure(x819_kernelx819_concrete1_io_in_x482_outbuf_0_rPort_0_backpressure),
    .io_in_x482_outbuf_0_rPort_0_output_0(x819_kernelx819_concrete1_io_in_x482_outbuf_0_rPort_0_output_0),
    .io_in_x478_outdram_number(x819_kernelx819_concrete1_io_in_x478_outdram_number),
    .io_in_x740_ready(x819_kernelx819_concrete1_io_in_x740_ready),
    .io_in_x740_valid(x819_kernelx819_concrete1_io_in_x740_valid),
    .io_in_x740_bits_wdata_0(x819_kernelx819_concrete1_io_in_x740_bits_wdata_0),
    .io_in_x740_bits_wstrb(x819_kernelx819_concrete1_io_in_x740_bits_wstrb),
    .io_sigsIn_smEnableOuts_0(x819_kernelx819_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x819_kernelx819_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(x819_kernelx819_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x819_kernelx819_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsOut_smDoneIn_0(x819_kernelx819_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x819_kernelx819_concrete1_io_sigsOut_smDoneIn_1),
    .io_rr(x819_kernelx819_concrete1_io_rr)
  );
  assign _T_266 = x819_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@49692.4]
  assign _T_283 = RetimeWrapper_io_out; // @[package.scala 96:25:@49731.4 package.scala 96:25:@49732.4]
  assign _T_289 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@49739.4 package.scala 96:25:@49740.4]
  assign _T_292 = ~ _T_289; // @[SpatialBlocks.scala 138:93:@49742.4]
  assign io_in_x481_TVALID = x819_kernelx819_concrete1_io_in_x481_TVALID; // @[sm_x819.scala 63:23:@49850.4]
  assign io_in_x481_TDATA = x819_kernelx819_concrete1_io_in_x481_TDATA; // @[sm_x819.scala 63:23:@49848.4]
  assign io_in_x741_ready = x819_kernelx819_concrete1_io_in_x741_ready; // @[sm_x819.scala 64:23:@49853.4]
  assign io_in_x480_TREADY = x819_kernelx819_concrete1_io_in_x480_TREADY; // @[sm_x819.scala 65:23:@49861.4]
  assign io_in_x739_valid = x819_kernelx819_concrete1_io_in_x739_valid; // @[sm_x819.scala 66:23:@49865.4]
  assign io_in_x739_bits_addr = x819_kernelx819_concrete1_io_in_x739_bits_addr; // @[sm_x819.scala 66:23:@49864.4]
  assign io_in_x739_bits_size = x819_kernelx819_concrete1_io_in_x739_bits_size; // @[sm_x819.scala 66:23:@49863.4]
  assign io_in_x740_valid = x819_kernelx819_concrete1_io_in_x740_valid; // @[sm_x819.scala 69:23:@49875.4]
  assign io_in_x740_bits_wdata_0 = x819_kernelx819_concrete1_io_in_x740_bits_wdata_0; // @[sm_x819.scala 69:23:@49874.4]
  assign io_in_x740_bits_wstrb = x819_kernelx819_concrete1_io_in_x740_bits_wstrb; // @[sm_x819.scala 69:23:@49873.4]
  assign io_sigsOut_smDoneIn_0 = x819_sm_io_done; // @[SpatialBlocks.scala 156:53:@49749.4]
  assign x482_outbuf_0_clock = clock; // @[:@49602.4]
  assign x482_outbuf_0_reset = reset; // @[:@49603.4]
  assign x482_outbuf_0_io_rPort_0_ofs_0 = x819_kernelx819_concrete1_io_in_x482_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@49870.4]
  assign x482_outbuf_0_io_rPort_0_en_0 = x819_kernelx819_concrete1_io_in_x482_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@49869.4]
  assign x482_outbuf_0_io_rPort_0_backpressure = x819_kernelx819_concrete1_io_in_x482_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@49868.4]
  assign x819_sm_clock = clock; // @[:@49660.4]
  assign x819_sm_reset = reset; // @[:@49661.4]
  assign x819_sm_io_enable = _T_283 & _T_292; // @[SpatialBlocks.scala 140:18:@49746.4]
  assign x819_sm_io_ctrDone = x819_sm_io_ctrInc & _T_269; // @[sm_RootController.scala 82:26:@49696.4]
  assign x819_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@49748.4]
  assign x819_sm_io_doneIn_0 = x819_kernelx819_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@49716.4]
  assign x819_sm_io_doneIn_1 = x819_kernelx819_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@49717.4]
  assign RetimeWrapper_clock = clock; // @[:@49727.4]
  assign RetimeWrapper_reset = reset; // @[:@49728.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@49730.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@49729.4]
  assign RetimeWrapper_1_clock = clock; // @[:@49735.4]
  assign RetimeWrapper_1_reset = reset; // @[:@49736.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@49738.4]
  assign RetimeWrapper_1_io_in = x819_sm_io_done; // @[package.scala 94:16:@49737.4]
  assign x819_kernelx819_concrete1_clock = clock; // @[:@49764.4]
  assign x819_kernelx819_concrete1_reset = reset; // @[:@49765.4]
  assign x819_kernelx819_concrete1_io_in_x481_TREADY = io_in_x481_TREADY; // @[sm_x819.scala 63:23:@49849.4]
  assign x819_kernelx819_concrete1_io_in_x741_valid = io_in_x741_valid; // @[sm_x819.scala 64:23:@49852.4]
  assign x819_kernelx819_concrete1_io_in_x480_TVALID = io_in_x480_TVALID; // @[sm_x819.scala 65:23:@49862.4]
  assign x819_kernelx819_concrete1_io_in_x480_TDATA = io_in_x480_TDATA; // @[sm_x819.scala 65:23:@49860.4]
  assign x819_kernelx819_concrete1_io_in_x480_TID = io_in_x480_TID; // @[sm_x819.scala 65:23:@49856.4]
  assign x819_kernelx819_concrete1_io_in_x480_TDEST = io_in_x480_TDEST; // @[sm_x819.scala 65:23:@49855.4]
  assign x819_kernelx819_concrete1_io_in_x739_ready = io_in_x739_ready; // @[sm_x819.scala 66:23:@49866.4]
  assign x819_kernelx819_concrete1_io_in_x482_outbuf_0_rPort_0_output_0 = x482_outbuf_0_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@49867.4]
  assign x819_kernelx819_concrete1_io_in_x478_outdram_number = io_in_x478_outdram_number; // @[sm_x819.scala 68:31:@49872.4]
  assign x819_kernelx819_concrete1_io_in_x740_ready = io_in_x740_ready; // @[sm_x819.scala 69:23:@49876.4]
  assign x819_kernelx819_concrete1_io_sigsIn_smEnableOuts_0 = x819_sm_io_enableOut_0; // @[sm_x819.scala 107:22:@49887.4]
  assign x819_kernelx819_concrete1_io_sigsIn_smEnableOuts_1 = x819_sm_io_enableOut_1; // @[sm_x819.scala 107:22:@49888.4]
  assign x819_kernelx819_concrete1_io_sigsIn_smChildAcks_0 = x819_sm_io_childAck_0; // @[sm_x819.scala 107:22:@49883.4]
  assign x819_kernelx819_concrete1_io_sigsIn_smChildAcks_1 = x819_sm_io_childAck_1; // @[sm_x819.scala 107:22:@49884.4]
  assign x819_kernelx819_concrete1_io_rr = io_rr; // @[sm_x819.scala 106:18:@49877.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_269 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_269 <= 1'h0;
    end else begin
      _T_269 <= _T_266;
    end
  end
endmodule
module AccelUnit( // @[:@49910.2]
  input          clock, // @[:@49911.4]
  input          reset, // @[:@49912.4]
  input          io_enable, // @[:@49913.4]
  output         io_done, // @[:@49913.4]
  input          io_reset, // @[:@49913.4]
  input          io_memStreams_loads_0_cmd_ready, // @[:@49913.4]
  output         io_memStreams_loads_0_cmd_valid, // @[:@49913.4]
  output [63:0]  io_memStreams_loads_0_cmd_bits_addr, // @[:@49913.4]
  output [31:0]  io_memStreams_loads_0_cmd_bits_size, // @[:@49913.4]
  output         io_memStreams_loads_0_data_ready, // @[:@49913.4]
  input          io_memStreams_loads_0_data_valid, // @[:@49913.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_0, // @[:@49913.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_1, // @[:@49913.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_2, // @[:@49913.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_3, // @[:@49913.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_4, // @[:@49913.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_5, // @[:@49913.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_6, // @[:@49913.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_7, // @[:@49913.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_8, // @[:@49913.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_9, // @[:@49913.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_10, // @[:@49913.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_11, // @[:@49913.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_12, // @[:@49913.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_13, // @[:@49913.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_14, // @[:@49913.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_15, // @[:@49913.4]
  input          io_memStreams_stores_0_cmd_ready, // @[:@49913.4]
  output         io_memStreams_stores_0_cmd_valid, // @[:@49913.4]
  output [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@49913.4]
  output [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@49913.4]
  input          io_memStreams_stores_0_data_ready, // @[:@49913.4]
  output         io_memStreams_stores_0_data_valid, // @[:@49913.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_0, // @[:@49913.4]
  output         io_memStreams_stores_0_data_bits_wstrb, // @[:@49913.4]
  output         io_memStreams_stores_0_wresp_ready, // @[:@49913.4]
  input          io_memStreams_stores_0_wresp_valid, // @[:@49913.4]
  input          io_memStreams_stores_0_wresp_bits, // @[:@49913.4]
  input          io_memStreams_gathers_0_cmd_ready, // @[:@49913.4]
  output         io_memStreams_gathers_0_cmd_valid, // @[:@49913.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_0, // @[:@49913.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_1, // @[:@49913.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_2, // @[:@49913.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_3, // @[:@49913.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_4, // @[:@49913.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_5, // @[:@49913.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_6, // @[:@49913.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_7, // @[:@49913.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_8, // @[:@49913.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_9, // @[:@49913.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_10, // @[:@49913.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_11, // @[:@49913.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_12, // @[:@49913.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_13, // @[:@49913.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_14, // @[:@49913.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_15, // @[:@49913.4]
  output         io_memStreams_gathers_0_data_ready, // @[:@49913.4]
  input          io_memStreams_gathers_0_data_valid, // @[:@49913.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_0, // @[:@49913.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_1, // @[:@49913.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_2, // @[:@49913.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_3, // @[:@49913.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_4, // @[:@49913.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_5, // @[:@49913.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_6, // @[:@49913.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_7, // @[:@49913.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_8, // @[:@49913.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_9, // @[:@49913.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_10, // @[:@49913.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_11, // @[:@49913.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_12, // @[:@49913.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_13, // @[:@49913.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_14, // @[:@49913.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_15, // @[:@49913.4]
  input          io_memStreams_scatters_0_cmd_ready, // @[:@49913.4]
  output         io_memStreams_scatters_0_cmd_valid, // @[:@49913.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_0, // @[:@49913.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_1, // @[:@49913.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_2, // @[:@49913.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_3, // @[:@49913.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_4, // @[:@49913.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_5, // @[:@49913.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_6, // @[:@49913.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_7, // @[:@49913.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_8, // @[:@49913.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_9, // @[:@49913.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_10, // @[:@49913.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_11, // @[:@49913.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_12, // @[:@49913.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_13, // @[:@49913.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_14, // @[:@49913.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_15, // @[:@49913.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_0, // @[:@49913.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_1, // @[:@49913.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_2, // @[:@49913.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_3, // @[:@49913.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_4, // @[:@49913.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_5, // @[:@49913.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_6, // @[:@49913.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_7, // @[:@49913.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_8, // @[:@49913.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_9, // @[:@49913.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_10, // @[:@49913.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_11, // @[:@49913.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_12, // @[:@49913.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_13, // @[:@49913.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_14, // @[:@49913.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_15, // @[:@49913.4]
  output         io_memStreams_scatters_0_wresp_ready, // @[:@49913.4]
  input          io_memStreams_scatters_0_wresp_valid, // @[:@49913.4]
  input          io_memStreams_scatters_0_wresp_bits, // @[:@49913.4]
  input          io_axiStreamsIn_0_TVALID, // @[:@49913.4]
  output         io_axiStreamsIn_0_TREADY, // @[:@49913.4]
  input  [255:0] io_axiStreamsIn_0_TDATA, // @[:@49913.4]
  input  [31:0]  io_axiStreamsIn_0_TSTRB, // @[:@49913.4]
  input  [31:0]  io_axiStreamsIn_0_TKEEP, // @[:@49913.4]
  input          io_axiStreamsIn_0_TLAST, // @[:@49913.4]
  input  [7:0]   io_axiStreamsIn_0_TID, // @[:@49913.4]
  input  [7:0]   io_axiStreamsIn_0_TDEST, // @[:@49913.4]
  input  [31:0]  io_axiStreamsIn_0_TUSER, // @[:@49913.4]
  output         io_axiStreamsOut_0_TVALID, // @[:@49913.4]
  input          io_axiStreamsOut_0_TREADY, // @[:@49913.4]
  output [255:0] io_axiStreamsOut_0_TDATA, // @[:@49913.4]
  output [31:0]  io_axiStreamsOut_0_TSTRB, // @[:@49913.4]
  output [31:0]  io_axiStreamsOut_0_TKEEP, // @[:@49913.4]
  output         io_axiStreamsOut_0_TLAST, // @[:@49913.4]
  output [7:0]   io_axiStreamsOut_0_TID, // @[:@49913.4]
  output [7:0]   io_axiStreamsOut_0_TDEST, // @[:@49913.4]
  output [31:0]  io_axiStreamsOut_0_TUSER, // @[:@49913.4]
  output         io_heap_0_req_valid, // @[:@49913.4]
  output         io_heap_0_req_bits_allocDealloc, // @[:@49913.4]
  output [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@49913.4]
  input          io_heap_0_resp_valid, // @[:@49913.4]
  input          io_heap_0_resp_bits_allocDealloc, // @[:@49913.4]
  input  [63:0]  io_heap_0_resp_bits_sizeAddr, // @[:@49913.4]
  input  [63:0]  io_argIns_0, // @[:@49913.4]
  input  [63:0]  io_argIns_1, // @[:@49913.4]
  input          io_argOuts_0_port_ready, // @[:@49913.4]
  output         io_argOuts_0_port_valid, // @[:@49913.4]
  output [63:0]  io_argOuts_0_port_bits, // @[:@49913.4]
  input  [63:0]  io_argOuts_0_echo // @[:@49913.4]
);
  wire  SingleCounter_clock; // @[Main.scala 40:32:@50061.4]
  wire  SingleCounter_reset; // @[Main.scala 40:32:@50061.4]
  wire  SingleCounter_io_input_reset; // @[Main.scala 40:32:@50061.4]
  wire  SingleCounter_io_output_done; // @[Main.scala 40:32:@50061.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@50079.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@50079.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@50079.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@50079.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@50079.4]
  wire  SRFF_clock; // @[Main.scala 44:28:@50088.4]
  wire  SRFF_reset; // @[Main.scala 44:28:@50088.4]
  wire  SRFF_io_input_set; // @[Main.scala 44:28:@50088.4]
  wire  SRFF_io_input_reset; // @[Main.scala 44:28:@50088.4]
  wire  SRFF_io_input_asyn_reset; // @[Main.scala 44:28:@50088.4]
  wire  SRFF_io_output; // @[Main.scala 44:28:@50088.4]
  wire  RootController_sm_clock; // @[sm_RootController.scala 36:18:@50127.4]
  wire  RootController_sm_reset; // @[sm_RootController.scala 36:18:@50127.4]
  wire  RootController_sm_io_enable; // @[sm_RootController.scala 36:18:@50127.4]
  wire  RootController_sm_io_done; // @[sm_RootController.scala 36:18:@50127.4]
  wire  RootController_sm_io_rst; // @[sm_RootController.scala 36:18:@50127.4]
  wire  RootController_sm_io_ctrDone; // @[sm_RootController.scala 36:18:@50127.4]
  wire  RootController_sm_io_ctrInc; // @[sm_RootController.scala 36:18:@50127.4]
  wire  RootController_sm_io_parentAck; // @[sm_RootController.scala 36:18:@50127.4]
  wire  RootController_sm_io_doneIn_0; // @[sm_RootController.scala 36:18:@50127.4]
  wire  RootController_sm_io_enableOut_0; // @[sm_RootController.scala 36:18:@50127.4]
  wire  RootController_sm_io_childAck_0; // @[sm_RootController.scala 36:18:@50127.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@50159.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@50159.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@50159.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@50159.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@50159.4]
  wire  RootController_kernelRootController_concrete1_clock; // @[sm_RootController.scala 91:24:@50221.4]
  wire  RootController_kernelRootController_concrete1_reset; // @[sm_RootController.scala 91:24:@50221.4]
  wire  RootController_kernelRootController_concrete1_io_in_x481_TVALID; // @[sm_RootController.scala 91:24:@50221.4]
  wire  RootController_kernelRootController_concrete1_io_in_x481_TREADY; // @[sm_RootController.scala 91:24:@50221.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x481_TDATA; // @[sm_RootController.scala 91:24:@50221.4]
  wire  RootController_kernelRootController_concrete1_io_in_x741_ready; // @[sm_RootController.scala 91:24:@50221.4]
  wire  RootController_kernelRootController_concrete1_io_in_x741_valid; // @[sm_RootController.scala 91:24:@50221.4]
  wire  RootController_kernelRootController_concrete1_io_in_x480_TVALID; // @[sm_RootController.scala 91:24:@50221.4]
  wire  RootController_kernelRootController_concrete1_io_in_x480_TREADY; // @[sm_RootController.scala 91:24:@50221.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x480_TDATA; // @[sm_RootController.scala 91:24:@50221.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x480_TID; // @[sm_RootController.scala 91:24:@50221.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x480_TDEST; // @[sm_RootController.scala 91:24:@50221.4]
  wire  RootController_kernelRootController_concrete1_io_in_x739_ready; // @[sm_RootController.scala 91:24:@50221.4]
  wire  RootController_kernelRootController_concrete1_io_in_x739_valid; // @[sm_RootController.scala 91:24:@50221.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x739_bits_addr; // @[sm_RootController.scala 91:24:@50221.4]
  wire [31:0] RootController_kernelRootController_concrete1_io_in_x739_bits_size; // @[sm_RootController.scala 91:24:@50221.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x478_outdram_number; // @[sm_RootController.scala 91:24:@50221.4]
  wire  RootController_kernelRootController_concrete1_io_in_x740_ready; // @[sm_RootController.scala 91:24:@50221.4]
  wire  RootController_kernelRootController_concrete1_io_in_x740_valid; // @[sm_RootController.scala 91:24:@50221.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x740_bits_wdata_0; // @[sm_RootController.scala 91:24:@50221.4]
  wire  RootController_kernelRootController_concrete1_io_in_x740_bits_wstrb; // @[sm_RootController.scala 91:24:@50221.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_RootController.scala 91:24:@50221.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0; // @[sm_RootController.scala 91:24:@50221.4]
  wire  RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[sm_RootController.scala 91:24:@50221.4]
  wire  RootController_kernelRootController_concrete1_io_rr; // @[sm_RootController.scala 91:24:@50221.4]
  wire  _T_599; // @[package.scala 96:25:@50084.4 package.scala 96:25:@50085.4]
  wire  _T_664; // @[Main.scala 46:50:@50155.4]
  wire  _T_665; // @[Main.scala 46:59:@50156.4]
  wire  _T_677; // @[package.scala 100:49:@50176.4]
  reg  _T_680; // @[package.scala 48:56:@50177.4]
  reg [31:0] _RAND_0;
  SingleCounter SingleCounter ( // @[Main.scala 40:32:@50061.4]
    .clock(SingleCounter_clock),
    .reset(SingleCounter_reset),
    .io_input_reset(SingleCounter_io_input_reset),
    .io_output_done(SingleCounter_io_output_done)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@50079.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  SRFF SRFF ( // @[Main.scala 44:28:@50088.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  RootController_sm RootController_sm ( // @[sm_RootController.scala 36:18:@50127.4]
    .clock(RootController_sm_clock),
    .reset(RootController_sm_reset),
    .io_enable(RootController_sm_io_enable),
    .io_done(RootController_sm_io_done),
    .io_rst(RootController_sm_io_rst),
    .io_ctrDone(RootController_sm_io_ctrDone),
    .io_ctrInc(RootController_sm_io_ctrInc),
    .io_parentAck(RootController_sm_io_parentAck),
    .io_doneIn_0(RootController_sm_io_doneIn_0),
    .io_enableOut_0(RootController_sm_io_enableOut_0),
    .io_childAck_0(RootController_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@50159.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RootController_kernelRootController_concrete1 RootController_kernelRootController_concrete1 ( // @[sm_RootController.scala 91:24:@50221.4]
    .clock(RootController_kernelRootController_concrete1_clock),
    .reset(RootController_kernelRootController_concrete1_reset),
    .io_in_x481_TVALID(RootController_kernelRootController_concrete1_io_in_x481_TVALID),
    .io_in_x481_TREADY(RootController_kernelRootController_concrete1_io_in_x481_TREADY),
    .io_in_x481_TDATA(RootController_kernelRootController_concrete1_io_in_x481_TDATA),
    .io_in_x741_ready(RootController_kernelRootController_concrete1_io_in_x741_ready),
    .io_in_x741_valid(RootController_kernelRootController_concrete1_io_in_x741_valid),
    .io_in_x480_TVALID(RootController_kernelRootController_concrete1_io_in_x480_TVALID),
    .io_in_x480_TREADY(RootController_kernelRootController_concrete1_io_in_x480_TREADY),
    .io_in_x480_TDATA(RootController_kernelRootController_concrete1_io_in_x480_TDATA),
    .io_in_x480_TID(RootController_kernelRootController_concrete1_io_in_x480_TID),
    .io_in_x480_TDEST(RootController_kernelRootController_concrete1_io_in_x480_TDEST),
    .io_in_x739_ready(RootController_kernelRootController_concrete1_io_in_x739_ready),
    .io_in_x739_valid(RootController_kernelRootController_concrete1_io_in_x739_valid),
    .io_in_x739_bits_addr(RootController_kernelRootController_concrete1_io_in_x739_bits_addr),
    .io_in_x739_bits_size(RootController_kernelRootController_concrete1_io_in_x739_bits_size),
    .io_in_x478_outdram_number(RootController_kernelRootController_concrete1_io_in_x478_outdram_number),
    .io_in_x740_ready(RootController_kernelRootController_concrete1_io_in_x740_ready),
    .io_in_x740_valid(RootController_kernelRootController_concrete1_io_in_x740_valid),
    .io_in_x740_bits_wdata_0(RootController_kernelRootController_concrete1_io_in_x740_bits_wdata_0),
    .io_in_x740_bits_wstrb(RootController_kernelRootController_concrete1_io_in_x740_bits_wstrb),
    .io_sigsIn_smEnableOuts_0(RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(RootController_kernelRootController_concrete1_io_rr)
  );
  assign _T_599 = RetimeWrapper_io_out; // @[package.scala 96:25:@50084.4 package.scala 96:25:@50085.4]
  assign _T_664 = io_enable & _T_599; // @[Main.scala 46:50:@50155.4]
  assign _T_665 = ~ SRFF_io_output; // @[Main.scala 46:59:@50156.4]
  assign _T_677 = RootController_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@50176.4]
  assign io_done = SRFF_io_output; // @[Main.scala 53:23:@50175.4]
  assign io_memStreams_loads_0_cmd_valid = 1'h0;
  assign io_memStreams_loads_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_loads_0_cmd_bits_size = 32'h0;
  assign io_memStreams_loads_0_data_ready = 1'h0;
  assign io_memStreams_stores_0_cmd_valid = RootController_kernelRootController_concrete1_io_in_x739_valid; // @[sm_RootController.scala 63:23:@50305.4]
  assign io_memStreams_stores_0_cmd_bits_addr = RootController_kernelRootController_concrete1_io_in_x739_bits_addr; // @[sm_RootController.scala 63:23:@50304.4]
  assign io_memStreams_stores_0_cmd_bits_size = RootController_kernelRootController_concrete1_io_in_x739_bits_size; // @[sm_RootController.scala 63:23:@50303.4]
  assign io_memStreams_stores_0_data_valid = RootController_kernelRootController_concrete1_io_in_x740_valid; // @[sm_RootController.scala 65:23:@50310.4]
  assign io_memStreams_stores_0_data_bits_wdata_0 = RootController_kernelRootController_concrete1_io_in_x740_bits_wdata_0; // @[sm_RootController.scala 65:23:@50309.4]
  assign io_memStreams_stores_0_data_bits_wstrb = RootController_kernelRootController_concrete1_io_in_x740_bits_wstrb; // @[sm_RootController.scala 65:23:@50308.4]
  assign io_memStreams_stores_0_wresp_ready = RootController_kernelRootController_concrete1_io_in_x741_ready; // @[sm_RootController.scala 61:23:@50293.4]
  assign io_memStreams_gathers_0_cmd_valid = 1'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_0 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_1 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_2 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_3 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_4 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_5 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_6 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_7 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_8 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_9 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_10 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_11 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_12 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_13 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_14 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_15 = 64'h0;
  assign io_memStreams_gathers_0_data_ready = 1'h0;
  assign io_memStreams_scatters_0_cmd_valid = 1'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_0 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_1 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_2 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_3 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_4 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_5 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_6 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_7 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_8 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_9 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_10 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_11 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_12 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_13 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_14 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_15 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_0 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_1 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_2 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_3 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_4 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_5 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_6 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_7 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_8 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_9 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_10 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_11 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_12 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_13 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_14 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_15 = 32'h0;
  assign io_memStreams_scatters_0_wresp_ready = 1'h0;
  assign io_axiStreamsIn_0_TREADY = RootController_kernelRootController_concrete1_io_in_x480_TREADY; // @[sm_RootController.scala 62:23:@50301.4]
  assign io_axiStreamsOut_0_TVALID = RootController_kernelRootController_concrete1_io_in_x481_TVALID; // @[sm_RootController.scala 60:23:@50290.4]
  assign io_axiStreamsOut_0_TDATA = RootController_kernelRootController_concrete1_io_in_x481_TDATA; // @[sm_RootController.scala 60:23:@50288.4]
  assign io_axiStreamsOut_0_TSTRB = 32'hffffffff; // @[sm_RootController.scala 60:23:@50287.4]
  assign io_axiStreamsOut_0_TKEEP = 32'hffffffff; // @[sm_RootController.scala 60:23:@50286.4]
  assign io_axiStreamsOut_0_TLAST = 1'h0; // @[sm_RootController.scala 60:23:@50285.4]
  assign io_axiStreamsOut_0_TID = 8'h0; // @[sm_RootController.scala 60:23:@50284.4]
  assign io_axiStreamsOut_0_TDEST = 8'h0; // @[sm_RootController.scala 60:23:@50283.4]
  assign io_axiStreamsOut_0_TUSER = 32'h4; // @[sm_RootController.scala 60:23:@50282.4]
  assign io_heap_0_req_valid = 1'h0;
  assign io_heap_0_req_bits_allocDealloc = 1'h0;
  assign io_heap_0_req_bits_sizeAddr = 64'h0;
  assign io_argOuts_0_port_valid = 1'h0;
  assign io_argOuts_0_port_bits = 64'h0;
  assign SingleCounter_clock = clock; // @[:@50062.4]
  assign SingleCounter_reset = reset; // @[:@50063.4]
  assign SingleCounter_io_input_reset = reset; // @[Main.scala 41:79:@50077.4]
  assign RetimeWrapper_clock = clock; // @[:@50080.4]
  assign RetimeWrapper_reset = reset; // @[:@50081.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@50083.4]
  assign RetimeWrapper_io_in = SingleCounter_io_output_done; // @[package.scala 94:16:@50082.4]
  assign SRFF_clock = clock; // @[:@50089.4]
  assign SRFF_reset = reset; // @[:@50090.4]
  assign SRFF_io_input_set = RootController_sm_io_done; // @[Main.scala 62:29:@50339.4]
  assign SRFF_io_input_reset = RetimeWrapper_1_io_out; // @[Main.scala 51:31:@50173.4]
  assign SRFF_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[Main.scala 52:36:@50174.4]
  assign RootController_sm_clock = clock; // @[:@50128.4]
  assign RootController_sm_reset = reset; // @[:@50129.4]
  assign RootController_sm_io_enable = _T_664 & _T_665; // @[Main.scala 50:33:@50172.4 SpatialBlocks.scala 140:18:@50206.4]
  assign RootController_sm_io_rst = RetimeWrapper_1_io_out; // @[SpatialBlocks.scala 134:15:@50200.4]
  assign RootController_sm_io_ctrDone = RootController_sm_io_ctrInc & _T_680; // @[Main.scala 54:34:@50180.4]
  assign RootController_sm_io_parentAck = 1'h0; // @[Main.scala 49:36:@50168.4 SpatialBlocks.scala 142:21:@50208.4]
  assign RootController_sm_io_doneIn_0 = RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@50197.4]
  assign RetimeWrapper_1_clock = clock; // @[:@50160.4]
  assign RetimeWrapper_1_reset = reset; // @[:@50161.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@50163.4]
  assign RetimeWrapper_1_io_in = reset | io_reset; // @[package.scala 94:16:@50162.4]
  assign RootController_kernelRootController_concrete1_clock = clock; // @[:@50222.4]
  assign RootController_kernelRootController_concrete1_reset = reset; // @[:@50223.4]
  assign RootController_kernelRootController_concrete1_io_in_x481_TREADY = io_axiStreamsOut_0_TREADY; // @[sm_RootController.scala 60:23:@50289.4]
  assign RootController_kernelRootController_concrete1_io_in_x741_valid = io_memStreams_stores_0_wresp_valid; // @[sm_RootController.scala 61:23:@50292.4]
  assign RootController_kernelRootController_concrete1_io_in_x480_TVALID = io_axiStreamsIn_0_TVALID; // @[sm_RootController.scala 62:23:@50302.4]
  assign RootController_kernelRootController_concrete1_io_in_x480_TDATA = io_axiStreamsIn_0_TDATA; // @[sm_RootController.scala 62:23:@50300.4]
  assign RootController_kernelRootController_concrete1_io_in_x480_TID = io_axiStreamsIn_0_TID; // @[sm_RootController.scala 62:23:@50296.4]
  assign RootController_kernelRootController_concrete1_io_in_x480_TDEST = io_axiStreamsIn_0_TDEST; // @[sm_RootController.scala 62:23:@50295.4]
  assign RootController_kernelRootController_concrete1_io_in_x739_ready = io_memStreams_stores_0_cmd_ready; // @[sm_RootController.scala 63:23:@50306.4]
  assign RootController_kernelRootController_concrete1_io_in_x478_outdram_number = io_argIns_1; // @[sm_RootController.scala 64:31:@50307.4]
  assign RootController_kernelRootController_concrete1_io_in_x740_ready = io_memStreams_stores_0_data_ready; // @[sm_RootController.scala 65:23:@50311.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0 = RootController_sm_io_enableOut_0; // @[sm_RootController.scala 96:22:@50320.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0 = RootController_sm_io_childAck_0; // @[sm_RootController.scala 96:22:@50318.4]
  assign RootController_kernelRootController_concrete1_io_rr = RetimeWrapper_io_out; // @[sm_RootController.scala 95:18:@50312.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_680 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_680 <= 1'h0;
    end else begin
      _T_680 <= _T_677;
    end
  end
endmodule
module SpatialIP( // @[:@50341.2]
  input         clock, // @[:@50342.4]
  input         reset, // @[:@50343.4]
  input  [31:0] io_raddr, // @[:@50344.4]
  input         io_wen, // @[:@50344.4]
  input  [31:0] io_waddr, // @[:@50344.4]
  input  [63:0] io_wdata, // @[:@50344.4]
  output [63:0] io_rdata // @[:@50344.4]
);
  wire  accel_clock; // @[Instantiator.scala 53:44:@50346.4]
  wire  accel_reset; // @[Instantiator.scala 53:44:@50346.4]
  wire  accel_io_enable; // @[Instantiator.scala 53:44:@50346.4]
  wire  accel_io_done; // @[Instantiator.scala 53:44:@50346.4]
  wire  accel_io_reset; // @[Instantiator.scala 53:44:@50346.4]
  wire  accel_io_memStreams_loads_0_cmd_ready; // @[Instantiator.scala 53:44:@50346.4]
  wire  accel_io_memStreams_loads_0_cmd_valid; // @[Instantiator.scala 53:44:@50346.4]
  wire [63:0] accel_io_memStreams_loads_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_loads_0_cmd_bits_size; // @[Instantiator.scala 53:44:@50346.4]
  wire  accel_io_memStreams_loads_0_data_ready; // @[Instantiator.scala 53:44:@50346.4]
  wire  accel_io_memStreams_loads_0_data_valid; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_0; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_1; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_2; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_3; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_4; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_5; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_6; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_7; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_8; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_9; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_10; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_11; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_12; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_13; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_14; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_15; // @[Instantiator.scala 53:44:@50346.4]
  wire  accel_io_memStreams_stores_0_cmd_ready; // @[Instantiator.scala 53:44:@50346.4]
  wire  accel_io_memStreams_stores_0_cmd_valid; // @[Instantiator.scala 53:44:@50346.4]
  wire [63:0] accel_io_memStreams_stores_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_stores_0_cmd_bits_size; // @[Instantiator.scala 53:44:@50346.4]
  wire  accel_io_memStreams_stores_0_data_ready; // @[Instantiator.scala 53:44:@50346.4]
  wire  accel_io_memStreams_stores_0_data_valid; // @[Instantiator.scala 53:44:@50346.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Instantiator.scala 53:44:@50346.4]
  wire  accel_io_memStreams_stores_0_data_bits_wstrb; // @[Instantiator.scala 53:44:@50346.4]
  wire  accel_io_memStreams_stores_0_wresp_ready; // @[Instantiator.scala 53:44:@50346.4]
  wire  accel_io_memStreams_stores_0_wresp_valid; // @[Instantiator.scala 53:44:@50346.4]
  wire  accel_io_memStreams_stores_0_wresp_bits; // @[Instantiator.scala 53:44:@50346.4]
  wire  accel_io_memStreams_gathers_0_cmd_ready; // @[Instantiator.scala 53:44:@50346.4]
  wire  accel_io_memStreams_gathers_0_cmd_valid; // @[Instantiator.scala 53:44:@50346.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_0; // @[Instantiator.scala 53:44:@50346.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_1; // @[Instantiator.scala 53:44:@50346.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_2; // @[Instantiator.scala 53:44:@50346.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_3; // @[Instantiator.scala 53:44:@50346.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_4; // @[Instantiator.scala 53:44:@50346.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_5; // @[Instantiator.scala 53:44:@50346.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_6; // @[Instantiator.scala 53:44:@50346.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_7; // @[Instantiator.scala 53:44:@50346.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_8; // @[Instantiator.scala 53:44:@50346.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_9; // @[Instantiator.scala 53:44:@50346.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_10; // @[Instantiator.scala 53:44:@50346.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_11; // @[Instantiator.scala 53:44:@50346.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_12; // @[Instantiator.scala 53:44:@50346.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_13; // @[Instantiator.scala 53:44:@50346.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_14; // @[Instantiator.scala 53:44:@50346.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_15; // @[Instantiator.scala 53:44:@50346.4]
  wire  accel_io_memStreams_gathers_0_data_ready; // @[Instantiator.scala 53:44:@50346.4]
  wire  accel_io_memStreams_gathers_0_data_valid; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_0; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_1; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_2; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_3; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_4; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_5; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_6; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_7; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_8; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_9; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_10; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_11; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_12; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_13; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_14; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_15; // @[Instantiator.scala 53:44:@50346.4]
  wire  accel_io_memStreams_scatters_0_cmd_ready; // @[Instantiator.scala 53:44:@50346.4]
  wire  accel_io_memStreams_scatters_0_cmd_valid; // @[Instantiator.scala 53:44:@50346.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0; // @[Instantiator.scala 53:44:@50346.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1; // @[Instantiator.scala 53:44:@50346.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2; // @[Instantiator.scala 53:44:@50346.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3; // @[Instantiator.scala 53:44:@50346.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4; // @[Instantiator.scala 53:44:@50346.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5; // @[Instantiator.scala 53:44:@50346.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6; // @[Instantiator.scala 53:44:@50346.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7; // @[Instantiator.scala 53:44:@50346.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8; // @[Instantiator.scala 53:44:@50346.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9; // @[Instantiator.scala 53:44:@50346.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10; // @[Instantiator.scala 53:44:@50346.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11; // @[Instantiator.scala 53:44:@50346.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12; // @[Instantiator.scala 53:44:@50346.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13; // @[Instantiator.scala 53:44:@50346.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14; // @[Instantiator.scala 53:44:@50346.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_0; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_1; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_2; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_3; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_4; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_5; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_6; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_7; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_8; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_9; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_10; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_11; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_12; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_13; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_14; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_15; // @[Instantiator.scala 53:44:@50346.4]
  wire  accel_io_memStreams_scatters_0_wresp_ready; // @[Instantiator.scala 53:44:@50346.4]
  wire  accel_io_memStreams_scatters_0_wresp_valid; // @[Instantiator.scala 53:44:@50346.4]
  wire  accel_io_memStreams_scatters_0_wresp_bits; // @[Instantiator.scala 53:44:@50346.4]
  wire  accel_io_axiStreamsIn_0_TVALID; // @[Instantiator.scala 53:44:@50346.4]
  wire  accel_io_axiStreamsIn_0_TREADY; // @[Instantiator.scala 53:44:@50346.4]
  wire [255:0] accel_io_axiStreamsIn_0_TDATA; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_axiStreamsIn_0_TSTRB; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_axiStreamsIn_0_TKEEP; // @[Instantiator.scala 53:44:@50346.4]
  wire  accel_io_axiStreamsIn_0_TLAST; // @[Instantiator.scala 53:44:@50346.4]
  wire [7:0] accel_io_axiStreamsIn_0_TID; // @[Instantiator.scala 53:44:@50346.4]
  wire [7:0] accel_io_axiStreamsIn_0_TDEST; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_axiStreamsIn_0_TUSER; // @[Instantiator.scala 53:44:@50346.4]
  wire  accel_io_axiStreamsOut_0_TVALID; // @[Instantiator.scala 53:44:@50346.4]
  wire  accel_io_axiStreamsOut_0_TREADY; // @[Instantiator.scala 53:44:@50346.4]
  wire [255:0] accel_io_axiStreamsOut_0_TDATA; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_axiStreamsOut_0_TSTRB; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_axiStreamsOut_0_TKEEP; // @[Instantiator.scala 53:44:@50346.4]
  wire  accel_io_axiStreamsOut_0_TLAST; // @[Instantiator.scala 53:44:@50346.4]
  wire [7:0] accel_io_axiStreamsOut_0_TID; // @[Instantiator.scala 53:44:@50346.4]
  wire [7:0] accel_io_axiStreamsOut_0_TDEST; // @[Instantiator.scala 53:44:@50346.4]
  wire [31:0] accel_io_axiStreamsOut_0_TUSER; // @[Instantiator.scala 53:44:@50346.4]
  wire  accel_io_heap_0_req_valid; // @[Instantiator.scala 53:44:@50346.4]
  wire  accel_io_heap_0_req_bits_allocDealloc; // @[Instantiator.scala 53:44:@50346.4]
  wire [63:0] accel_io_heap_0_req_bits_sizeAddr; // @[Instantiator.scala 53:44:@50346.4]
  wire  accel_io_heap_0_resp_valid; // @[Instantiator.scala 53:44:@50346.4]
  wire  accel_io_heap_0_resp_bits_allocDealloc; // @[Instantiator.scala 53:44:@50346.4]
  wire [63:0] accel_io_heap_0_resp_bits_sizeAddr; // @[Instantiator.scala 53:44:@50346.4]
  wire [63:0] accel_io_argIns_0; // @[Instantiator.scala 53:44:@50346.4]
  wire [63:0] accel_io_argIns_1; // @[Instantiator.scala 53:44:@50346.4]
  wire  accel_io_argOuts_0_port_ready; // @[Instantiator.scala 53:44:@50346.4]
  wire  accel_io_argOuts_0_port_valid; // @[Instantiator.scala 53:44:@50346.4]
  wire [63:0] accel_io_argOuts_0_port_bits; // @[Instantiator.scala 53:44:@50346.4]
  wire [63:0] accel_io_argOuts_0_echo; // @[Instantiator.scala 53:44:@50346.4]
  AccelUnit accel ( // @[Instantiator.scala 53:44:@50346.4]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_enable(accel_io_enable),
    .io_done(accel_io_done),
    .io_reset(accel_io_reset),
    .io_memStreams_loads_0_cmd_ready(accel_io_memStreams_loads_0_cmd_ready),
    .io_memStreams_loads_0_cmd_valid(accel_io_memStreams_loads_0_cmd_valid),
    .io_memStreams_loads_0_cmd_bits_addr(accel_io_memStreams_loads_0_cmd_bits_addr),
    .io_memStreams_loads_0_cmd_bits_size(accel_io_memStreams_loads_0_cmd_bits_size),
    .io_memStreams_loads_0_data_ready(accel_io_memStreams_loads_0_data_ready),
    .io_memStreams_loads_0_data_valid(accel_io_memStreams_loads_0_data_valid),
    .io_memStreams_loads_0_data_bits_rdata_0(accel_io_memStreams_loads_0_data_bits_rdata_0),
    .io_memStreams_loads_0_data_bits_rdata_1(accel_io_memStreams_loads_0_data_bits_rdata_1),
    .io_memStreams_loads_0_data_bits_rdata_2(accel_io_memStreams_loads_0_data_bits_rdata_2),
    .io_memStreams_loads_0_data_bits_rdata_3(accel_io_memStreams_loads_0_data_bits_rdata_3),
    .io_memStreams_loads_0_data_bits_rdata_4(accel_io_memStreams_loads_0_data_bits_rdata_4),
    .io_memStreams_loads_0_data_bits_rdata_5(accel_io_memStreams_loads_0_data_bits_rdata_5),
    .io_memStreams_loads_0_data_bits_rdata_6(accel_io_memStreams_loads_0_data_bits_rdata_6),
    .io_memStreams_loads_0_data_bits_rdata_7(accel_io_memStreams_loads_0_data_bits_rdata_7),
    .io_memStreams_loads_0_data_bits_rdata_8(accel_io_memStreams_loads_0_data_bits_rdata_8),
    .io_memStreams_loads_0_data_bits_rdata_9(accel_io_memStreams_loads_0_data_bits_rdata_9),
    .io_memStreams_loads_0_data_bits_rdata_10(accel_io_memStreams_loads_0_data_bits_rdata_10),
    .io_memStreams_loads_0_data_bits_rdata_11(accel_io_memStreams_loads_0_data_bits_rdata_11),
    .io_memStreams_loads_0_data_bits_rdata_12(accel_io_memStreams_loads_0_data_bits_rdata_12),
    .io_memStreams_loads_0_data_bits_rdata_13(accel_io_memStreams_loads_0_data_bits_rdata_13),
    .io_memStreams_loads_0_data_bits_rdata_14(accel_io_memStreams_loads_0_data_bits_rdata_14),
    .io_memStreams_loads_0_data_bits_rdata_15(accel_io_memStreams_loads_0_data_bits_rdata_15),
    .io_memStreams_stores_0_cmd_ready(accel_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(accel_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(accel_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(accel_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(accel_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(accel_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(accel_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(accel_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(accel_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(accel_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(accel_io_memStreams_stores_0_wresp_bits),
    .io_memStreams_gathers_0_cmd_ready(accel_io_memStreams_gathers_0_cmd_ready),
    .io_memStreams_gathers_0_cmd_valid(accel_io_memStreams_gathers_0_cmd_valid),
    .io_memStreams_gathers_0_cmd_bits_addr_0(accel_io_memStreams_gathers_0_cmd_bits_addr_0),
    .io_memStreams_gathers_0_cmd_bits_addr_1(accel_io_memStreams_gathers_0_cmd_bits_addr_1),
    .io_memStreams_gathers_0_cmd_bits_addr_2(accel_io_memStreams_gathers_0_cmd_bits_addr_2),
    .io_memStreams_gathers_0_cmd_bits_addr_3(accel_io_memStreams_gathers_0_cmd_bits_addr_3),
    .io_memStreams_gathers_0_cmd_bits_addr_4(accel_io_memStreams_gathers_0_cmd_bits_addr_4),
    .io_memStreams_gathers_0_cmd_bits_addr_5(accel_io_memStreams_gathers_0_cmd_bits_addr_5),
    .io_memStreams_gathers_0_cmd_bits_addr_6(accel_io_memStreams_gathers_0_cmd_bits_addr_6),
    .io_memStreams_gathers_0_cmd_bits_addr_7(accel_io_memStreams_gathers_0_cmd_bits_addr_7),
    .io_memStreams_gathers_0_cmd_bits_addr_8(accel_io_memStreams_gathers_0_cmd_bits_addr_8),
    .io_memStreams_gathers_0_cmd_bits_addr_9(accel_io_memStreams_gathers_0_cmd_bits_addr_9),
    .io_memStreams_gathers_0_cmd_bits_addr_10(accel_io_memStreams_gathers_0_cmd_bits_addr_10),
    .io_memStreams_gathers_0_cmd_bits_addr_11(accel_io_memStreams_gathers_0_cmd_bits_addr_11),
    .io_memStreams_gathers_0_cmd_bits_addr_12(accel_io_memStreams_gathers_0_cmd_bits_addr_12),
    .io_memStreams_gathers_0_cmd_bits_addr_13(accel_io_memStreams_gathers_0_cmd_bits_addr_13),
    .io_memStreams_gathers_0_cmd_bits_addr_14(accel_io_memStreams_gathers_0_cmd_bits_addr_14),
    .io_memStreams_gathers_0_cmd_bits_addr_15(accel_io_memStreams_gathers_0_cmd_bits_addr_15),
    .io_memStreams_gathers_0_data_ready(accel_io_memStreams_gathers_0_data_ready),
    .io_memStreams_gathers_0_data_valid(accel_io_memStreams_gathers_0_data_valid),
    .io_memStreams_gathers_0_data_bits_0(accel_io_memStreams_gathers_0_data_bits_0),
    .io_memStreams_gathers_0_data_bits_1(accel_io_memStreams_gathers_0_data_bits_1),
    .io_memStreams_gathers_0_data_bits_2(accel_io_memStreams_gathers_0_data_bits_2),
    .io_memStreams_gathers_0_data_bits_3(accel_io_memStreams_gathers_0_data_bits_3),
    .io_memStreams_gathers_0_data_bits_4(accel_io_memStreams_gathers_0_data_bits_4),
    .io_memStreams_gathers_0_data_bits_5(accel_io_memStreams_gathers_0_data_bits_5),
    .io_memStreams_gathers_0_data_bits_6(accel_io_memStreams_gathers_0_data_bits_6),
    .io_memStreams_gathers_0_data_bits_7(accel_io_memStreams_gathers_0_data_bits_7),
    .io_memStreams_gathers_0_data_bits_8(accel_io_memStreams_gathers_0_data_bits_8),
    .io_memStreams_gathers_0_data_bits_9(accel_io_memStreams_gathers_0_data_bits_9),
    .io_memStreams_gathers_0_data_bits_10(accel_io_memStreams_gathers_0_data_bits_10),
    .io_memStreams_gathers_0_data_bits_11(accel_io_memStreams_gathers_0_data_bits_11),
    .io_memStreams_gathers_0_data_bits_12(accel_io_memStreams_gathers_0_data_bits_12),
    .io_memStreams_gathers_0_data_bits_13(accel_io_memStreams_gathers_0_data_bits_13),
    .io_memStreams_gathers_0_data_bits_14(accel_io_memStreams_gathers_0_data_bits_14),
    .io_memStreams_gathers_0_data_bits_15(accel_io_memStreams_gathers_0_data_bits_15),
    .io_memStreams_scatters_0_cmd_ready(accel_io_memStreams_scatters_0_cmd_ready),
    .io_memStreams_scatters_0_cmd_valid(accel_io_memStreams_scatters_0_cmd_valid),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_0(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_1(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_2(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_3(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_4(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_5(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_6(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_7(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_8(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_9(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_10(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_11(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_12(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_13(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_14(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_15(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15),
    .io_memStreams_scatters_0_cmd_bits_wdata_0(accel_io_memStreams_scatters_0_cmd_bits_wdata_0),
    .io_memStreams_scatters_0_cmd_bits_wdata_1(accel_io_memStreams_scatters_0_cmd_bits_wdata_1),
    .io_memStreams_scatters_0_cmd_bits_wdata_2(accel_io_memStreams_scatters_0_cmd_bits_wdata_2),
    .io_memStreams_scatters_0_cmd_bits_wdata_3(accel_io_memStreams_scatters_0_cmd_bits_wdata_3),
    .io_memStreams_scatters_0_cmd_bits_wdata_4(accel_io_memStreams_scatters_0_cmd_bits_wdata_4),
    .io_memStreams_scatters_0_cmd_bits_wdata_5(accel_io_memStreams_scatters_0_cmd_bits_wdata_5),
    .io_memStreams_scatters_0_cmd_bits_wdata_6(accel_io_memStreams_scatters_0_cmd_bits_wdata_6),
    .io_memStreams_scatters_0_cmd_bits_wdata_7(accel_io_memStreams_scatters_0_cmd_bits_wdata_7),
    .io_memStreams_scatters_0_cmd_bits_wdata_8(accel_io_memStreams_scatters_0_cmd_bits_wdata_8),
    .io_memStreams_scatters_0_cmd_bits_wdata_9(accel_io_memStreams_scatters_0_cmd_bits_wdata_9),
    .io_memStreams_scatters_0_cmd_bits_wdata_10(accel_io_memStreams_scatters_0_cmd_bits_wdata_10),
    .io_memStreams_scatters_0_cmd_bits_wdata_11(accel_io_memStreams_scatters_0_cmd_bits_wdata_11),
    .io_memStreams_scatters_0_cmd_bits_wdata_12(accel_io_memStreams_scatters_0_cmd_bits_wdata_12),
    .io_memStreams_scatters_0_cmd_bits_wdata_13(accel_io_memStreams_scatters_0_cmd_bits_wdata_13),
    .io_memStreams_scatters_0_cmd_bits_wdata_14(accel_io_memStreams_scatters_0_cmd_bits_wdata_14),
    .io_memStreams_scatters_0_cmd_bits_wdata_15(accel_io_memStreams_scatters_0_cmd_bits_wdata_15),
    .io_memStreams_scatters_0_wresp_ready(accel_io_memStreams_scatters_0_wresp_ready),
    .io_memStreams_scatters_0_wresp_valid(accel_io_memStreams_scatters_0_wresp_valid),
    .io_memStreams_scatters_0_wresp_bits(accel_io_memStreams_scatters_0_wresp_bits),
    .io_axiStreamsIn_0_TVALID(accel_io_axiStreamsIn_0_TVALID),
    .io_axiStreamsIn_0_TREADY(accel_io_axiStreamsIn_0_TREADY),
    .io_axiStreamsIn_0_TDATA(accel_io_axiStreamsIn_0_TDATA),
    .io_axiStreamsIn_0_TSTRB(accel_io_axiStreamsIn_0_TSTRB),
    .io_axiStreamsIn_0_TKEEP(accel_io_axiStreamsIn_0_TKEEP),
    .io_axiStreamsIn_0_TLAST(accel_io_axiStreamsIn_0_TLAST),
    .io_axiStreamsIn_0_TID(accel_io_axiStreamsIn_0_TID),
    .io_axiStreamsIn_0_TDEST(accel_io_axiStreamsIn_0_TDEST),
    .io_axiStreamsIn_0_TUSER(accel_io_axiStreamsIn_0_TUSER),
    .io_axiStreamsOut_0_TVALID(accel_io_axiStreamsOut_0_TVALID),
    .io_axiStreamsOut_0_TREADY(accel_io_axiStreamsOut_0_TREADY),
    .io_axiStreamsOut_0_TDATA(accel_io_axiStreamsOut_0_TDATA),
    .io_axiStreamsOut_0_TSTRB(accel_io_axiStreamsOut_0_TSTRB),
    .io_axiStreamsOut_0_TKEEP(accel_io_axiStreamsOut_0_TKEEP),
    .io_axiStreamsOut_0_TLAST(accel_io_axiStreamsOut_0_TLAST),
    .io_axiStreamsOut_0_TID(accel_io_axiStreamsOut_0_TID),
    .io_axiStreamsOut_0_TDEST(accel_io_axiStreamsOut_0_TDEST),
    .io_axiStreamsOut_0_TUSER(accel_io_axiStreamsOut_0_TUSER),
    .io_heap_0_req_valid(accel_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(accel_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(accel_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(accel_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(accel_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(accel_io_heap_0_resp_bits_sizeAddr),
    .io_argIns_0(accel_io_argIns_0),
    .io_argIns_1(accel_io_argIns_1),
    .io_argOuts_0_port_ready(accel_io_argOuts_0_port_ready),
    .io_argOuts_0_port_valid(accel_io_argOuts_0_port_valid),
    .io_argOuts_0_port_bits(accel_io_argOuts_0_port_bits),
    .io_argOuts_0_echo(accel_io_argOuts_0_echo)
  );
  assign io_rdata = 64'h0;
  assign accel_clock = clock; // @[:@50347.4]
  assign accel_reset = reset; // @[:@50348.4]
  assign accel_io_enable = 1'h0;
  assign accel_io_reset = 1'h0;
  assign accel_io_memStreams_loads_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_loads_0_data_valid = 1'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_0 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_1 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_2 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_3 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_4 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_5 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_6 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_7 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_8 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_9 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_10 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_11 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_12 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_13 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_14 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_15 = 32'h0;
  assign accel_io_memStreams_stores_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_stores_0_data_ready = 1'h0;
  assign accel_io_memStreams_stores_0_wresp_valid = 1'h0;
  assign accel_io_memStreams_stores_0_wresp_bits = 1'h0;
  assign accel_io_memStreams_gathers_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_gathers_0_data_valid = 1'h0;
  assign accel_io_memStreams_gathers_0_data_bits_0 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_1 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_2 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_3 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_4 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_5 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_6 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_7 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_8 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_9 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_10 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_11 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_12 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_13 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_14 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_15 = 32'h0;
  assign accel_io_memStreams_scatters_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_scatters_0_wresp_valid = 1'h0;
  assign accel_io_memStreams_scatters_0_wresp_bits = 1'h0;
  assign accel_io_axiStreamsIn_0_TVALID = 1'h0;
  assign accel_io_axiStreamsIn_0_TDATA = 256'h0;
  assign accel_io_axiStreamsIn_0_TSTRB = 32'h0;
  assign accel_io_axiStreamsIn_0_TKEEP = 32'h0;
  assign accel_io_axiStreamsIn_0_TLAST = 1'h0;
  assign accel_io_axiStreamsIn_0_TID = 8'h0;
  assign accel_io_axiStreamsIn_0_TDEST = 8'h0;
  assign accel_io_axiStreamsIn_0_TUSER = 32'h0;
  assign accel_io_axiStreamsOut_0_TREADY = 1'h0;
  assign accel_io_heap_0_resp_valid = 1'h0;
  assign accel_io_heap_0_resp_bits_allocDealloc = 1'h0;
  assign accel_io_heap_0_resp_bits_sizeAddr = 64'h0;
  assign accel_io_argIns_0 = 64'h0;
  assign accel_io_argIns_1 = 64'h0;
  assign accel_io_argOuts_0_port_ready = 1'h0;
  assign accel_io_argOuts_0_echo = 64'h0;
endmodule
